//Latest Update Date: 11th Nov, 2025
//Owner: B Nithin Reddy


//Multiplier Design

module mul(
  input [3:0] a,b,
  output [7:0] y
);
  
  assign y = a * b;
  
endmodule
