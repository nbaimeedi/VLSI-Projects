module cve2_core (crash_dump_o_64_,
    data_addr_o_0_,
    data_addr_o_1_,
    instr_addr_o_0_,
    instr_addr_o_1_,
    boot_addr_i_0_,
    boot_addr_i_10_,
    boot_addr_i_11_,
    boot_addr_i_12_,
    boot_addr_i_13_,
    boot_addr_i_14_,
    boot_addr_i_15_,
    boot_addr_i_16_,
    boot_addr_i_17_,
    boot_addr_i_18_,
    boot_addr_i_19_,
    boot_addr_i_1_,
    boot_addr_i_20_,
    boot_addr_i_21_,
    boot_addr_i_22_,
    boot_addr_i_23_,
    boot_addr_i_24_,
    boot_addr_i_25_,
    boot_addr_i_26_,
    boot_addr_i_27_,
    boot_addr_i_28_,
    boot_addr_i_29_,
    boot_addr_i_2_,
    boot_addr_i_30_,
    boot_addr_i_31_,
    boot_addr_i_3_,
    boot_addr_i_4_,
    boot_addr_i_5_,
    boot_addr_i_6_,
    boot_addr_i_7_,
    boot_addr_i_8_,
    boot_addr_i_9_,
    clk_i,
    core_busy_o,
    crash_dump_o_0_,
    crash_dump_o_100_,
    crash_dump_o_101_,
    crash_dump_o_102_,
    crash_dump_o_103_,
    crash_dump_o_104_,
    crash_dump_o_105_,
    crash_dump_o_106_,
    crash_dump_o_107_,
    crash_dump_o_108_,
    crash_dump_o_109_,
    crash_dump_o_10_,
    crash_dump_o_110_,
    crash_dump_o_111_,
    crash_dump_o_112_,
    crash_dump_o_113_,
    crash_dump_o_114_,
    crash_dump_o_115_,
    crash_dump_o_116_,
    crash_dump_o_117_,
    crash_dump_o_118_,
    crash_dump_o_119_,
    crash_dump_o_11_,
    crash_dump_o_120_,
    crash_dump_o_121_,
    crash_dump_o_122_,
    crash_dump_o_123_,
    crash_dump_o_124_,
    crash_dump_o_125_,
    crash_dump_o_126_,
    crash_dump_o_127_,
    crash_dump_o_12_,
    crash_dump_o_13_,
    crash_dump_o_14_,
    crash_dump_o_15_,
    crash_dump_o_16_,
    crash_dump_o_17_,
    crash_dump_o_18_,
    crash_dump_o_19_,
    crash_dump_o_1_,
    crash_dump_o_20_,
    crash_dump_o_21_,
    crash_dump_o_22_,
    crash_dump_o_23_,
    crash_dump_o_24_,
    crash_dump_o_25_,
    crash_dump_o_26_,
    crash_dump_o_27_,
    crash_dump_o_28_,
    crash_dump_o_29_,
    crash_dump_o_2_,
    crash_dump_o_30_,
    crash_dump_o_31_,
    crash_dump_o_32_,
    crash_dump_o_33_,
    crash_dump_o_34_,
    crash_dump_o_35_,
    crash_dump_o_36_,
    crash_dump_o_37_,
    crash_dump_o_38_,
    crash_dump_o_39_,
    crash_dump_o_3_,
    crash_dump_o_40_,
    crash_dump_o_41_,
    crash_dump_o_42_,
    crash_dump_o_43_,
    crash_dump_o_44_,
    crash_dump_o_45_,
    crash_dump_o_46_,
    crash_dump_o_47_,
    crash_dump_o_48_,
    crash_dump_o_49_,
    crash_dump_o_4_,
    crash_dump_o_50_,
    crash_dump_o_51_,
    crash_dump_o_52_,
    crash_dump_o_53_,
    crash_dump_o_54_,
    crash_dump_o_55_,
    crash_dump_o_56_,
    crash_dump_o_57_,
    crash_dump_o_58_,
    crash_dump_o_59_,
    crash_dump_o_5_,
    crash_dump_o_60_,
    crash_dump_o_61_,
    crash_dump_o_62_,
    crash_dump_o_63_,
    crash_dump_o_65_,
    crash_dump_o_66_,
    crash_dump_o_67_,
    crash_dump_o_68_,
    crash_dump_o_69_,
    crash_dump_o_6_,
    crash_dump_o_70_,
    crash_dump_o_71_,
    crash_dump_o_72_,
    crash_dump_o_73_,
    crash_dump_o_74_,
    crash_dump_o_75_,
    crash_dump_o_76_,
    crash_dump_o_77_,
    crash_dump_o_78_,
    crash_dump_o_79_,
    crash_dump_o_7_,
    crash_dump_o_80_,
    crash_dump_o_81_,
    crash_dump_o_82_,
    crash_dump_o_83_,
    crash_dump_o_84_,
    crash_dump_o_85_,
    crash_dump_o_86_,
    crash_dump_o_87_,
    crash_dump_o_88_,
    crash_dump_o_89_,
    crash_dump_o_8_,
    crash_dump_o_90_,
    crash_dump_o_91_,
    crash_dump_o_92_,
    crash_dump_o_93_,
    crash_dump_o_94_,
    crash_dump_o_95_,
    crash_dump_o_96_,
    crash_dump_o_97_,
    crash_dump_o_98_,
    crash_dump_o_99_,
    crash_dump_o_9_,
    data_addr_o_10_,
    data_addr_o_11_,
    data_addr_o_12_,
    data_addr_o_13_,
    data_addr_o_14_,
    data_addr_o_15_,
    data_addr_o_16_,
    data_addr_o_17_,
    data_addr_o_18_,
    data_addr_o_19_,
    data_addr_o_20_,
    data_addr_o_21_,
    data_addr_o_22_,
    data_addr_o_23_,
    data_addr_o_24_,
    data_addr_o_25_,
    data_addr_o_26_,
    data_addr_o_27_,
    data_addr_o_28_,
    data_addr_o_29_,
    data_addr_o_2_,
    data_addr_o_30_,
    data_addr_o_31_,
    data_addr_o_3_,
    data_addr_o_4_,
    data_addr_o_5_,
    data_addr_o_6_,
    data_addr_o_7_,
    data_addr_o_8_,
    data_addr_o_9_,
    data_be_o_0_,
    data_be_o_1_,
    data_be_o_2_,
    data_be_o_3_,
    data_err_i,
    data_gnt_i,
    data_rdata_i_0_,
    data_rdata_i_10_,
    data_rdata_i_11_,
    data_rdata_i_12_,
    data_rdata_i_13_,
    data_rdata_i_14_,
    data_rdata_i_15_,
    data_rdata_i_16_,
    data_rdata_i_17_,
    data_rdata_i_18_,
    data_rdata_i_19_,
    data_rdata_i_1_,
    data_rdata_i_20_,
    data_rdata_i_21_,
    data_rdata_i_22_,
    data_rdata_i_23_,
    data_rdata_i_24_,
    data_rdata_i_25_,
    data_rdata_i_26_,
    data_rdata_i_27_,
    data_rdata_i_28_,
    data_rdata_i_29_,
    data_rdata_i_2_,
    data_rdata_i_30_,
    data_rdata_i_31_,
    data_rdata_i_3_,
    data_rdata_i_4_,
    data_rdata_i_5_,
    data_rdata_i_6_,
    data_rdata_i_7_,
    data_rdata_i_8_,
    data_rdata_i_9_,
    data_req_o,
    data_rvalid_i,
    data_wdata_o_0_,
    data_wdata_o_10_,
    data_wdata_o_11_,
    data_wdata_o_12_,
    data_wdata_o_13_,
    data_wdata_o_14_,
    data_wdata_o_15_,
    data_wdata_o_16_,
    data_wdata_o_17_,
    data_wdata_o_18_,
    data_wdata_o_19_,
    data_wdata_o_1_,
    data_wdata_o_20_,
    data_wdata_o_21_,
    data_wdata_o_22_,
    data_wdata_o_23_,
    data_wdata_o_24_,
    data_wdata_o_25_,
    data_wdata_o_26_,
    data_wdata_o_27_,
    data_wdata_o_28_,
    data_wdata_o_29_,
    data_wdata_o_2_,
    data_wdata_o_30_,
    data_wdata_o_31_,
    data_wdata_o_3_,
    data_wdata_o_4_,
    data_wdata_o_5_,
    data_wdata_o_6_,
    data_wdata_o_7_,
    data_wdata_o_8_,
    data_wdata_o_9_,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    hart_id_i_0_,
    hart_id_i_10_,
    hart_id_i_11_,
    hart_id_i_12_,
    hart_id_i_13_,
    hart_id_i_14_,
    hart_id_i_15_,
    hart_id_i_16_,
    hart_id_i_17_,
    hart_id_i_18_,
    hart_id_i_19_,
    hart_id_i_1_,
    hart_id_i_20_,
    hart_id_i_21_,
    hart_id_i_22_,
    hart_id_i_23_,
    hart_id_i_24_,
    hart_id_i_25_,
    hart_id_i_26_,
    hart_id_i_27_,
    hart_id_i_28_,
    hart_id_i_29_,
    hart_id_i_2_,
    hart_id_i_30_,
    hart_id_i_31_,
    hart_id_i_3_,
    hart_id_i_4_,
    hart_id_i_5_,
    hart_id_i_6_,
    hart_id_i_7_,
    hart_id_i_8_,
    hart_id_i_9_,
    instr_addr_o_10_,
    instr_addr_o_11_,
    instr_addr_o_12_,
    instr_addr_o_13_,
    instr_addr_o_14_,
    instr_addr_o_15_,
    instr_addr_o_16_,
    instr_addr_o_17_,
    instr_addr_o_18_,
    instr_addr_o_19_,
    instr_addr_o_20_,
    instr_addr_o_21_,
    instr_addr_o_22_,
    instr_addr_o_23_,
    instr_addr_o_24_,
    instr_addr_o_25_,
    instr_addr_o_26_,
    instr_addr_o_27_,
    instr_addr_o_28_,
    instr_addr_o_29_,
    instr_addr_o_2_,
    instr_addr_o_30_,
    instr_addr_o_31_,
    instr_addr_o_3_,
    instr_addr_o_4_,
    instr_addr_o_5_,
    instr_addr_o_6_,
    instr_addr_o_7_,
    instr_addr_o_8_,
    instr_addr_o_9_,
    instr_err_i,
    instr_gnt_i,
    instr_rdata_i_0_,
    instr_rdata_i_10_,
    instr_rdata_i_11_,
    instr_rdata_i_12_,
    instr_rdata_i_13_,
    instr_rdata_i_14_,
    instr_rdata_i_15_,
    instr_rdata_i_16_,
    instr_rdata_i_17_,
    instr_rdata_i_18_,
    instr_rdata_i_19_,
    instr_rdata_i_1_,
    instr_rdata_i_20_,
    instr_rdata_i_21_,
    instr_rdata_i_22_,
    instr_rdata_i_23_,
    instr_rdata_i_24_,
    instr_rdata_i_25_,
    instr_rdata_i_26_,
    instr_rdata_i_27_,
    instr_rdata_i_28_,
    instr_rdata_i_29_,
    instr_rdata_i_2_,
    instr_rdata_i_30_,
    instr_rdata_i_31_,
    instr_rdata_i_3_,
    instr_rdata_i_4_,
    instr_rdata_i_5_,
    instr_rdata_i_6_,
    instr_rdata_i_7_,
    instr_rdata_i_8_,
    instr_rdata_i_9_,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_fast_i_0_,
    irq_fast_i_10_,
    irq_fast_i_11_,
    irq_fast_i_12_,
    irq_fast_i_13_,
    irq_fast_i_14_,
    irq_fast_i_15_,
    irq_fast_i_1_,
    irq_fast_i_2_,
    irq_fast_i_3_,
    irq_fast_i_4_,
    irq_fast_i_5_,
    irq_fast_i_6_,
    irq_fast_i_7_,
    irq_fast_i_8_,
    irq_fast_i_9_,
    irq_nm_i,
    irq_pending_o,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i);
 output crash_dump_o_64_;
 output data_addr_o_0_;
 output data_addr_o_1_;
 output instr_addr_o_0_;
 output instr_addr_o_1_;
 input boot_addr_i_0_;
 input boot_addr_i_10_;
 input boot_addr_i_11_;
 input boot_addr_i_12_;
 input boot_addr_i_13_;
 input boot_addr_i_14_;
 input boot_addr_i_15_;
 input boot_addr_i_16_;
 input boot_addr_i_17_;
 input boot_addr_i_18_;
 input boot_addr_i_19_;
 input boot_addr_i_1_;
 input boot_addr_i_20_;
 input boot_addr_i_21_;
 input boot_addr_i_22_;
 input boot_addr_i_23_;
 input boot_addr_i_24_;
 input boot_addr_i_25_;
 input boot_addr_i_26_;
 input boot_addr_i_27_;
 input boot_addr_i_28_;
 input boot_addr_i_29_;
 input boot_addr_i_2_;
 input boot_addr_i_30_;
 input boot_addr_i_31_;
 input boot_addr_i_3_;
 input boot_addr_i_4_;
 input boot_addr_i_5_;
 input boot_addr_i_6_;
 input boot_addr_i_7_;
 input boot_addr_i_8_;
 input boot_addr_i_9_;
 input clk_i;
 output core_busy_o;
 output crash_dump_o_0_;
 output crash_dump_o_100_;
 output crash_dump_o_101_;
 output crash_dump_o_102_;
 output crash_dump_o_103_;
 output crash_dump_o_104_;
 output crash_dump_o_105_;
 output crash_dump_o_106_;
 output crash_dump_o_107_;
 output crash_dump_o_108_;
 output crash_dump_o_109_;
 output crash_dump_o_10_;
 output crash_dump_o_110_;
 output crash_dump_o_111_;
 output crash_dump_o_112_;
 output crash_dump_o_113_;
 output crash_dump_o_114_;
 output crash_dump_o_115_;
 output crash_dump_o_116_;
 output crash_dump_o_117_;
 output crash_dump_o_118_;
 output crash_dump_o_119_;
 output crash_dump_o_11_;
 output crash_dump_o_120_;
 output crash_dump_o_121_;
 output crash_dump_o_122_;
 output crash_dump_o_123_;
 output crash_dump_o_124_;
 output crash_dump_o_125_;
 output crash_dump_o_126_;
 output crash_dump_o_127_;
 output crash_dump_o_12_;
 output crash_dump_o_13_;
 output crash_dump_o_14_;
 output crash_dump_o_15_;
 output crash_dump_o_16_;
 output crash_dump_o_17_;
 output crash_dump_o_18_;
 output crash_dump_o_19_;
 output crash_dump_o_1_;
 output crash_dump_o_20_;
 output crash_dump_o_21_;
 output crash_dump_o_22_;
 output crash_dump_o_23_;
 output crash_dump_o_24_;
 output crash_dump_o_25_;
 output crash_dump_o_26_;
 output crash_dump_o_27_;
 output crash_dump_o_28_;
 output crash_dump_o_29_;
 output crash_dump_o_2_;
 output crash_dump_o_30_;
 output crash_dump_o_31_;
 output crash_dump_o_32_;
 output crash_dump_o_33_;
 output crash_dump_o_34_;
 output crash_dump_o_35_;
 output crash_dump_o_36_;
 output crash_dump_o_37_;
 output crash_dump_o_38_;
 output crash_dump_o_39_;
 output crash_dump_o_3_;
 output crash_dump_o_40_;
 output crash_dump_o_41_;
 output crash_dump_o_42_;
 output crash_dump_o_43_;
 output crash_dump_o_44_;
 output crash_dump_o_45_;
 output crash_dump_o_46_;
 output crash_dump_o_47_;
 output crash_dump_o_48_;
 output crash_dump_o_49_;
 output crash_dump_o_4_;
 output crash_dump_o_50_;
 output crash_dump_o_51_;
 output crash_dump_o_52_;
 output crash_dump_o_53_;
 output crash_dump_o_54_;
 output crash_dump_o_55_;
 output crash_dump_o_56_;
 output crash_dump_o_57_;
 output crash_dump_o_58_;
 output crash_dump_o_59_;
 output crash_dump_o_5_;
 output crash_dump_o_60_;
 output crash_dump_o_61_;
 output crash_dump_o_62_;
 output crash_dump_o_63_;
 output crash_dump_o_65_;
 output crash_dump_o_66_;
 output crash_dump_o_67_;
 output crash_dump_o_68_;
 output crash_dump_o_69_;
 output crash_dump_o_6_;
 output crash_dump_o_70_;
 output crash_dump_o_71_;
 output crash_dump_o_72_;
 output crash_dump_o_73_;
 output crash_dump_o_74_;
 output crash_dump_o_75_;
 output crash_dump_o_76_;
 output crash_dump_o_77_;
 output crash_dump_o_78_;
 output crash_dump_o_79_;
 output crash_dump_o_7_;
 output crash_dump_o_80_;
 output crash_dump_o_81_;
 output crash_dump_o_82_;
 output crash_dump_o_83_;
 output crash_dump_o_84_;
 output crash_dump_o_85_;
 output crash_dump_o_86_;
 output crash_dump_o_87_;
 output crash_dump_o_88_;
 output crash_dump_o_89_;
 output crash_dump_o_8_;
 output crash_dump_o_90_;
 output crash_dump_o_91_;
 output crash_dump_o_92_;
 output crash_dump_o_93_;
 output crash_dump_o_94_;
 output crash_dump_o_95_;
 output crash_dump_o_96_;
 output crash_dump_o_97_;
 output crash_dump_o_98_;
 output crash_dump_o_99_;
 output crash_dump_o_9_;
 output data_addr_o_10_;
 output data_addr_o_11_;
 output data_addr_o_12_;
 output data_addr_o_13_;
 output data_addr_o_14_;
 output data_addr_o_15_;
 output data_addr_o_16_;
 output data_addr_o_17_;
 output data_addr_o_18_;
 output data_addr_o_19_;
 output data_addr_o_20_;
 output data_addr_o_21_;
 output data_addr_o_22_;
 output data_addr_o_23_;
 output data_addr_o_24_;
 output data_addr_o_25_;
 output data_addr_o_26_;
 output data_addr_o_27_;
 output data_addr_o_28_;
 output data_addr_o_29_;
 output data_addr_o_2_;
 output data_addr_o_30_;
 output data_addr_o_31_;
 output data_addr_o_3_;
 output data_addr_o_4_;
 output data_addr_o_5_;
 output data_addr_o_6_;
 output data_addr_o_7_;
 output data_addr_o_8_;
 output data_addr_o_9_;
 output data_be_o_0_;
 output data_be_o_1_;
 output data_be_o_2_;
 output data_be_o_3_;
 input data_err_i;
 input data_gnt_i;
 input data_rdata_i_0_;
 input data_rdata_i_10_;
 input data_rdata_i_11_;
 input data_rdata_i_12_;
 input data_rdata_i_13_;
 input data_rdata_i_14_;
 input data_rdata_i_15_;
 input data_rdata_i_16_;
 input data_rdata_i_17_;
 input data_rdata_i_18_;
 input data_rdata_i_19_;
 input data_rdata_i_1_;
 input data_rdata_i_20_;
 input data_rdata_i_21_;
 input data_rdata_i_22_;
 input data_rdata_i_23_;
 input data_rdata_i_24_;
 input data_rdata_i_25_;
 input data_rdata_i_26_;
 input data_rdata_i_27_;
 input data_rdata_i_28_;
 input data_rdata_i_29_;
 input data_rdata_i_2_;
 input data_rdata_i_30_;
 input data_rdata_i_31_;
 input data_rdata_i_3_;
 input data_rdata_i_4_;
 input data_rdata_i_5_;
 input data_rdata_i_6_;
 input data_rdata_i_7_;
 input data_rdata_i_8_;
 input data_rdata_i_9_;
 output data_req_o;
 input data_rvalid_i;
 output data_wdata_o_0_;
 output data_wdata_o_10_;
 output data_wdata_o_11_;
 output data_wdata_o_12_;
 output data_wdata_o_13_;
 output data_wdata_o_14_;
 output data_wdata_o_15_;
 output data_wdata_o_16_;
 output data_wdata_o_17_;
 output data_wdata_o_18_;
 output data_wdata_o_19_;
 output data_wdata_o_1_;
 output data_wdata_o_20_;
 output data_wdata_o_21_;
 output data_wdata_o_22_;
 output data_wdata_o_23_;
 output data_wdata_o_24_;
 output data_wdata_o_25_;
 output data_wdata_o_26_;
 output data_wdata_o_27_;
 output data_wdata_o_28_;
 output data_wdata_o_29_;
 output data_wdata_o_2_;
 output data_wdata_o_30_;
 output data_wdata_o_31_;
 output data_wdata_o_3_;
 output data_wdata_o_4_;
 output data_wdata_o_5_;
 output data_wdata_o_6_;
 output data_wdata_o_7_;
 output data_wdata_o_8_;
 output data_wdata_o_9_;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input hart_id_i_0_;
 input hart_id_i_10_;
 input hart_id_i_11_;
 input hart_id_i_12_;
 input hart_id_i_13_;
 input hart_id_i_14_;
 input hart_id_i_15_;
 input hart_id_i_16_;
 input hart_id_i_17_;
 input hart_id_i_18_;
 input hart_id_i_19_;
 input hart_id_i_1_;
 input hart_id_i_20_;
 input hart_id_i_21_;
 input hart_id_i_22_;
 input hart_id_i_23_;
 input hart_id_i_24_;
 input hart_id_i_25_;
 input hart_id_i_26_;
 input hart_id_i_27_;
 input hart_id_i_28_;
 input hart_id_i_29_;
 input hart_id_i_2_;
 input hart_id_i_30_;
 input hart_id_i_31_;
 input hart_id_i_3_;
 input hart_id_i_4_;
 input hart_id_i_5_;
 input hart_id_i_6_;
 input hart_id_i_7_;
 input hart_id_i_8_;
 input hart_id_i_9_;
 output instr_addr_o_10_;
 output instr_addr_o_11_;
 output instr_addr_o_12_;
 output instr_addr_o_13_;
 output instr_addr_o_14_;
 output instr_addr_o_15_;
 output instr_addr_o_16_;
 output instr_addr_o_17_;
 output instr_addr_o_18_;
 output instr_addr_o_19_;
 output instr_addr_o_20_;
 output instr_addr_o_21_;
 output instr_addr_o_22_;
 output instr_addr_o_23_;
 output instr_addr_o_24_;
 output instr_addr_o_25_;
 output instr_addr_o_26_;
 output instr_addr_o_27_;
 output instr_addr_o_28_;
 output instr_addr_o_29_;
 output instr_addr_o_2_;
 output instr_addr_o_30_;
 output instr_addr_o_31_;
 output instr_addr_o_3_;
 output instr_addr_o_4_;
 output instr_addr_o_5_;
 output instr_addr_o_6_;
 output instr_addr_o_7_;
 output instr_addr_o_8_;
 output instr_addr_o_9_;
 input instr_err_i;
 input instr_gnt_i;
 input instr_rdata_i_0_;
 input instr_rdata_i_10_;
 input instr_rdata_i_11_;
 input instr_rdata_i_12_;
 input instr_rdata_i_13_;
 input instr_rdata_i_14_;
 input instr_rdata_i_15_;
 input instr_rdata_i_16_;
 input instr_rdata_i_17_;
 input instr_rdata_i_18_;
 input instr_rdata_i_19_;
 input instr_rdata_i_1_;
 input instr_rdata_i_20_;
 input instr_rdata_i_21_;
 input instr_rdata_i_22_;
 input instr_rdata_i_23_;
 input instr_rdata_i_24_;
 input instr_rdata_i_25_;
 input instr_rdata_i_26_;
 input instr_rdata_i_27_;
 input instr_rdata_i_28_;
 input instr_rdata_i_29_;
 input instr_rdata_i_2_;
 input instr_rdata_i_30_;
 input instr_rdata_i_31_;
 input instr_rdata_i_3_;
 input instr_rdata_i_4_;
 input instr_rdata_i_5_;
 input instr_rdata_i_6_;
 input instr_rdata_i_7_;
 input instr_rdata_i_8_;
 input instr_rdata_i_9_;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_fast_i_0_;
 input irq_fast_i_10_;
 input irq_fast_i_11_;
 input irq_fast_i_12_;
 input irq_fast_i_13_;
 input irq_fast_i_14_;
 input irq_fast_i_15_;
 input irq_fast_i_1_;
 input irq_fast_i_2_;
 input irq_fast_i_3_;
 input irq_fast_i_4_;
 input irq_fast_i_5_;
 input irq_fast_i_6_;
 input irq_fast_i_7_;
 input irq_fast_i_8_;
 input irq_fast_i_9_;
 input irq_nm_i;
 output irq_pending_o;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire net668;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire net667;
 wire net666;
 wire net665;
 wire net664;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire net663;
 wire _00585_;
 wire _00586_;
 wire net662;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire net661;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire net660;
 wire _00611_;
 wire _00612_;
 wire net659;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire net1333;
 wire net1332;
 wire _01130_;
 wire net1331;
 wire net1330;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire net1329;
 wire net1328;
 wire net1327;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire net1326;
 wire net1325;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire net1324;
 wire net1323;
 wire net1322;
 wire net1321;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire net1320;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire net1319;
 wire net1318;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire net1317;
 wire net1316;
 wire _01181_;
 wire _01182_;
 wire net1315;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire net1314;
 wire net1313;
 wire net1312;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire net1311;
 wire _01202_;
 wire net1310;
 wire net1309;
 wire _01205_;
 wire _01206_;
 wire net1308;
 wire net1307;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire net1303;
 wire net1302;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire net1301;
 wire _01236_;
 wire _01237_;
 wire net1300;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire net1298;
 wire _01270_;
 wire _01271_;
 wire net1297;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire net1293;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire net1292;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire net1288;
 wire net1287;
 wire _01329_;
 wire net1286;
 wire net1285;
 wire net1284;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire net1283;
 wire _01348_;
 wire net1282;
 wire net1281;
 wire net1280;
 wire net1279;
 wire net1278;
 wire _01354_;
 wire _01355_;
 wire net1277;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire net1276;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire net1275;
 wire net1274;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire net1273;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire net1272;
 wire net1271;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire net1270;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire net1269;
 wire net1268;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire net1267;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire net1266;
 wire _01471_;
 wire _01472_;
 wire net1265;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire net1264;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire net1263;
 wire net1262;
 wire net1261;
 wire net1260;
 wire net1259;
 wire net1258;
 wire _01506_;
 wire net1257;
 wire _01508_;
 wire _01509_;
 wire net1256;
 wire net1255;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire net1254;
 wire net1253;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire net1252;
 wire _01533_;
 wire net1251;
 wire _01535_;
 wire _01536_;
 wire net1250;
 wire net1249;
 wire net1248;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire net1247;
 wire net1246;
 wire net1245;
 wire net1244;
 wire net1243;
 wire net1242;
 wire net1241;
 wire net1240;
 wire net1239;
 wire _01552_;
 wire _01553_;
 wire net1238;
 wire net1237;
 wire net1236;
 wire net1235;
 wire net1234;
 wire net1233;
 wire net1232;
 wire _01561_;
 wire net1231;
 wire net1230;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire net1229;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire net1228;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire net1227;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire net1226;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire net1225;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire net1224;
 wire net1223;
 wire net1222;
 wire net1221;
 wire net1220;
 wire net1219;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire net1218;
 wire net1217;
 wire net1216;
 wire net1215;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire net1214;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire net1213;
 wire net1212;
 wire net1211;
 wire net1210;
 wire net1209;
 wire net1208;
 wire net1207;
 wire net1206;
 wire _01823_;
 wire _01824_;
 wire net1205;
 wire _01826_;
 wire net1204;
 wire net1203;
 wire net1202;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire net1201;
 wire net1200;
 wire net1199;
 wire net1198;
 wire net1197;
 wire net1196;
 wire _01839_;
 wire _01840_;
 wire net1195;
 wire net1194;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire net1193;
 wire _01848_;
 wire net1192;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire net1191;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire net1190;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire net1189;
 wire net1188;
 wire _01880_;
 wire net1187;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire net1186;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire net1185;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire net1184;
 wire net1183;
 wire net1182;
 wire net1181;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire net1180;
 wire net1179;
 wire net1178;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire net1177;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire net1176;
 wire net1175;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire net1174;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire net1173;
 wire _01953_;
 wire _01954_;
 wire net1172;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire net1171;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire net1170;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire net1169;
 wire net1168;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire net1167;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire net1166;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire net1165;
 wire _02006_;
 wire net1164;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire net1163;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire net1162;
 wire net1161;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire net1160;
 wire _02055_;
 wire _02056_;
 wire net1159;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire net1158;
 wire net1157;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire net1156;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire net1155;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire net1154;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire net1153;
 wire _02127_;
 wire _02128_;
 wire net1152;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire net1151;
 wire _02142_;
 wire _02143_;
 wire net1150;
 wire _02145_;
 wire _02146_;
 wire net1149;
 wire _02148_;
 wire net1148;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire net1147;
 wire _02159_;
 wire _02160_;
 wire net1146;
 wire net1145;
 wire net1144;
 wire _02164_;
 wire net1143;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire net1142;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire net1141;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire net1140;
 wire net1139;
 wire net1138;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire net1137;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire net1136;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire net1135;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire net1134;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire net1133;
 wire net1132;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire net1131;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire net1130;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire net1129;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire net1128;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire net1127;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire net1126;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire net1125;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire net1124;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire net1123;
 wire net1122;
 wire net1121;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire net1120;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire net1119;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire net1118;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire net1117;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire net1116;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire net1115;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire net1114;
 wire net1113;
 wire _02685_;
 wire _02686_;
 wire net1112;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire net1111;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire net1110;
 wire _02773_;
 wire _02774_;
 wire net1109;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire net1108;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire net1087;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire net1107;
 wire net1106;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire net1105;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire net1104;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire net1103;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire net1102;
 wire net1101;
 wire net1100;
 wire _03200_;
 wire net1099;
 wire net1098;
 wire net1097;
 wire _03204_;
 wire _03205_;
 wire net1096;
 wire _03207_;
 wire _03208_;
 wire net1095;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire net1094;
 wire _03214_;
 wire net1093;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire net1092;
 wire net1091;
 wire net1090;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire net1089;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire net1088;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire net1086;
 wire net1085;
 wire net1084;
 wire net1083;
 wire net1082;
 wire net1081;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire net1080;
 wire _03298_;
 wire _03299_;
 wire net1079;
 wire net1078;
 wire net1077;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire net1076;
 wire net1075;
 wire net1074;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire net1073;
 wire net1072;
 wire net1071;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire net1070;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire net1069;
 wire _03370_;
 wire net1068;
 wire net1067;
 wire net1066;
 wire net1065;
 wire _03375_;
 wire _03376_;
 wire net1064;
 wire net1063;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire net1062;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire net1061;
 wire _03423_;
 wire _03424_;
 wire net1060;
 wire _03426_;
 wire net1059;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire net1058;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire net1057;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire net1056;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire net1055;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire net1054;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire net1053;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire net1052;
 wire net1051;
 wire net1050;
 wire net1049;
 wire net1048;
 wire net1047;
 wire net1046;
 wire net1045;
 wire net1044;
 wire net1043;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire net1042;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire net1041;
 wire _03700_;
 wire _03701_;
 wire net1040;
 wire net1039;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire net1038;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire net1037;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire net1036;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire net1035;
 wire net1034;
 wire _03866_;
 wire net1033;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire net1032;
 wire _03881_;
 wire _03882_;
 wire net1031;
 wire _03884_;
 wire _03885_;
 wire net1030;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire net1029;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire net1028;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire net1027;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire net1026;
 wire net1025;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire net1024;
 wire net1023;
 wire net1022;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire net1021;
 wire net1020;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire net1019;
 wire _03974_;
 wire net1018;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire net1017;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire net1016;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire net1015;
 wire net1014;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire net1013;
 wire net1012;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire net1011;
 wire net1010;
 wire net1009;
 wire _04050_;
 wire _04051_;
 wire net1008;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire net1007;
 wire net1006;
 wire net1005;
 wire net1004;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire net1003;
 wire net1002;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire net1001;
 wire net1000;
 wire net999;
 wire _04081_;
 wire net998;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire net997;
 wire _04087_;
 wire net996;
 wire net995;
 wire _04090_;
 wire _04091_;
 wire net994;
 wire net993;
 wire net992;
 wire net991;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire net990;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire net989;
 wire net988;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire net987;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire net986;
 wire _04146_;
 wire _04147_;
 wire net985;
 wire net984;
 wire net983;
 wire _04151_;
 wire net982;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire net981;
 wire _04160_;
 wire _04161_;
 wire net980;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire net979;
 wire net978;
 wire _04169_;
 wire _04170_;
 wire net977;
 wire net976;
 wire _04173_;
 wire _04174_;
 wire net975;
 wire _04176_;
 wire _04177_;
 wire net974;
 wire net973;
 wire net972;
 wire net971;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire net970;
 wire net969;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire net968;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire net967;
 wire net966;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire net965;
 wire net964;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire net963;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire net962;
 wire net961;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire net960;
 wire net959;
 wire net958;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire net957;
 wire net956;
 wire net955;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire net954;
 wire net953;
 wire net952;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire net951;
 wire net950;
 wire net949;
 wire _04293_;
 wire _04294_;
 wire net948;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire net947;
 wire net946;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire net945;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire net944;
 wire net943;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire net942;
 wire _04347_;
 wire net941;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire net940;
 wire net939;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire net938;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire net937;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire net936;
 wire _04401_;
 wire net935;
 wire net934;
 wire net933;
 wire net932;
 wire net931;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire net930;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire net929;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire net928;
 wire net927;
 wire net926;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire net925;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire net924;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire net923;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire net922;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire net921;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire net920;
 wire net919;
 wire _04526_;
 wire _04527_;
 wire net918;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire net917;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire net916;
 wire net915;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire net914;
 wire net913;
 wire _04592_;
 wire _04593_;
 wire net912;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire net911;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire net910;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire net909;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire net908;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire net907;
 wire _04661_;
 wire net906;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire net905;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire net904;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire net903;
 wire net902;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire net901;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire net900;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire net899;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire net898;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire net897;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire net896;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire net895;
 wire net894;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire net893;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire net892;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire net891;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire net890;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire net889;
 wire _05086_;
 wire net888;
 wire net887;
 wire net886;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire net885;
 wire _05155_;
 wire net884;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire net883;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire net882;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire net881;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire net880;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire net879;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire net878;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire net877;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire net876;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire net875;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire net874;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire net873;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire net872;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire net871;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire net870;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire net869;
 wire _05806_;
 wire net868;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire net867;
 wire net866;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire net865;
 wire _05847_;
 wire net864;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire net863;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire net862;
 wire _05958_;
 wire net861;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire net860;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire net859;
 wire _06181_;
 wire net858;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire net857;
 wire net856;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire net855;
 wire net854;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire net853;
 wire net852;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire net851;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire net850;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire net849;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire net848;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire net847;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire net846;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire net845;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire net844;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire net843;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire net842;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire net841;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire net840;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire net839;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire net838;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire net837;
 wire net836;
 wire _07265_;
 wire net835;
 wire net834;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire net833;
 wire net832;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire net831;
 wire net830;
 wire _07279_;
 wire _07280_;
 wire net829;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire net828;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire net827;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire net826;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire net825;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire net824;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire net823;
 wire net822;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire net821;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire net820;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire net819;
 wire net818;
 wire net817;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire net816;
 wire net815;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire net814;
 wire net813;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire net812;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire net811;
 wire _07516_;
 wire _07517_;
 wire net810;
 wire _07519_;
 wire net809;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire net808;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire net807;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire net806;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire net805;
 wire _07537_;
 wire net804;
 wire net803;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire net802;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire net801;
 wire net800;
 wire net799;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire net798;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire net797;
 wire net796;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire net795;
 wire net794;
 wire _07571_;
 wire _07572_;
 wire net793;
 wire net792;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire net791;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire net790;
 wire net789;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire net788;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire net787;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire net786;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire net785;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire net784;
 wire _07621_;
 wire _07622_;
 wire net783;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire net782;
 wire _07639_;
 wire _07640_;
 wire net781;
 wire net780;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire net779;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire net778;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire net777;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire net776;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire net775;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire net774;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire net773;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire net772;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire net771;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire net770;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire net769;
 wire net768;
 wire net767;
 wire _08241_;
 wire _08242_;
 wire net766;
 wire _08244_;
 wire _08245_;
 wire net765;
 wire net764;
 wire net763;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire net762;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire net761;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire net760;
 wire _08277_;
 wire net759;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire net758;
 wire _08289_;
 wire net757;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire net756;
 wire net755;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire net754;
 wire _08312_;
 wire net753;
 wire net752;
 wire net751;
 wire net750;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire net749;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire net748;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire net747;
 wire net746;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire net745;
 wire _08386_;
 wire net744;
 wire _08388_;
 wire net743;
 wire _08390_;
 wire net742;
 wire _08392_;
 wire net741;
 wire net740;
 wire _08395_;
 wire net739;
 wire net738;
 wire _08398_;
 wire net737;
 wire net736;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire net735;
 wire net734;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire net733;
 wire net732;
 wire _08428_;
 wire _08429_;
 wire net731;
 wire net730;
 wire net729;
 wire _08433_;
 wire _08434_;
 wire net728;
 wire net727;
 wire net726;
 wire _08438_;
 wire _08439_;
 wire net725;
 wire net724;
 wire _08442_;
 wire _08443_;
 wire net723;
 wire net722;
 wire net721;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire net720;
 wire _08451_;
 wire _08452_;
 wire net719;
 wire net718;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire net717;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire net716;
 wire net715;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire net714;
 wire net713;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire net712;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire net711;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire net710;
 wire net709;
 wire _08518_;
 wire _08519_;
 wire net708;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire net707;
 wire net706;
 wire _08526_;
 wire net705;
 wire net704;
 wire net703;
 wire net702;
 wire net701;
 wire net700;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire net699;
 wire net698;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire net697;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire net696;
 wire net695;
 wire net694;
 wire net693;
 wire net692;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire net691;
 wire net690;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire net689;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire net688;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire net687;
 wire net686;
 wire _08605_;
 wire _08606_;
 wire net685;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire net684;
 wire _08622_;
 wire net683;
 wire net682;
 wire _08625_;
 wire _08626_;
 wire net681;
 wire net680;
 wire net679;
 wire net678;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire net677;
 wire _08636_;
 wire _08637_;
 wire net676;
 wire _08639_;
 wire _08640_;
 wire net675;
 wire net674;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire net673;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire net672;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire net671;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire net670;
 wire _08703_;
 wire net669;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire net7;
 wire alu_operand_a_ex_0_;
 wire net1306;
 wire net1305;
 wire net1304;
 wire alu_operand_a_ex_13_;
 wire alu_operand_a_ex_14_;
 wire alu_operand_a_ex_15_;
 wire alu_operand_a_ex_16_;
 wire alu_operand_a_ex_17_;
 wire alu_operand_a_ex_18_;
 wire net1299;
 wire alu_operand_a_ex_1_;
 wire alu_operand_a_ex_20_;
 wire alu_operand_a_ex_21_;
 wire alu_operand_a_ex_22_;
 wire alu_operand_a_ex_23_;
 wire alu_operand_a_ex_24_;
 wire alu_operand_a_ex_25_;
 wire alu_operand_a_ex_26_;
 wire net1296;
 wire net1295;
 wire net1294;
 wire alu_operand_a_ex_2_;
 wire alu_operand_a_ex_30_;
 wire alu_operand_a_ex_31_;
 wire alu_operand_a_ex_3_;
 wire net1291;
 wire alu_operand_a_ex_5_;
 wire net1290;
 wire alu_operand_a_ex_7_;
 wire alu_operand_a_ex_8_;
 wire net1289;
 wire csr_access;
 wire csr_addr_0_;
 wire csr_addr_10_;
 wire csr_addr_11_;
 wire csr_addr_1_;
 wire csr_addr_2_;
 wire csr_addr_3_;
 wire csr_addr_4_;
 wire csr_addr_5_;
 wire csr_addr_6_;
 wire csr_addr_7_;
 wire csr_addr_8_;
 wire csr_addr_9_;
 wire csr_depc_0_;
 wire csr_depc_10_;
 wire csr_depc_11_;
 wire csr_depc_12_;
 wire csr_depc_13_;
 wire csr_depc_14_;
 wire csr_depc_15_;
 wire csr_depc_16_;
 wire csr_depc_17_;
 wire csr_depc_18_;
 wire csr_depc_19_;
 wire csr_depc_1_;
 wire csr_depc_20_;
 wire csr_depc_21_;
 wire csr_depc_22_;
 wire csr_depc_23_;
 wire csr_depc_24_;
 wire csr_depc_25_;
 wire csr_depc_26_;
 wire csr_depc_27_;
 wire csr_depc_28_;
 wire csr_depc_29_;
 wire csr_depc_2_;
 wire csr_depc_30_;
 wire csr_depc_31_;
 wire csr_depc_3_;
 wire csr_depc_4_;
 wire csr_depc_5_;
 wire csr_depc_6_;
 wire csr_depc_7_;
 wire csr_depc_8_;
 wire csr_depc_9_;
 wire csr_mstatus_mie;
 wire csr_mstatus_tw;
 wire csr_mtval_0_;
 wire csr_mtval_10_;
 wire csr_mtval_11_;
 wire csr_mtval_12_;
 wire csr_mtval_13_;
 wire csr_mtval_14_;
 wire csr_mtval_15_;
 wire csr_mtval_16_;
 wire csr_mtval_17_;
 wire csr_mtval_18_;
 wire csr_mtval_19_;
 wire csr_mtval_1_;
 wire \csr_mtval_1__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_MUX__Y_B ;
 wire csr_mtval_20_;
 wire csr_mtval_21_;
 wire csr_mtval_22_;
 wire csr_mtval_23_;
 wire csr_mtval_24_;
 wire csr_mtval_25_;
 wire csr_mtval_26_;
 wire csr_mtval_27_;
 wire csr_mtval_28_;
 wire csr_mtval_29_;
 wire csr_mtval_2_;
 wire csr_mtval_30_;
 wire csr_mtval_31_;
 wire csr_mtval_3_;
 wire csr_mtval_4_;
 wire csr_mtval_5_;
 wire csr_mtval_6_;
 wire csr_mtval_7_;
 wire csr_mtval_8_;
 wire csr_mtval_9_;
 wire csr_mtvec_0_;
 wire csr_mtvec_10_;
 wire csr_mtvec_11_;
 wire csr_mtvec_12_;
 wire csr_mtvec_13_;
 wire csr_mtvec_14_;
 wire csr_mtvec_15_;
 wire csr_mtvec_16_;
 wire csr_mtvec_17_;
 wire csr_mtvec_18_;
 wire csr_mtvec_19_;
 wire csr_mtvec_1_;
 wire csr_mtvec_20_;
 wire csr_mtvec_21_;
 wire csr_mtvec_22_;
 wire csr_mtvec_23_;
 wire csr_mtvec_24_;
 wire csr_mtvec_25_;
 wire csr_mtvec_26_;
 wire csr_mtvec_27_;
 wire csr_mtvec_28_;
 wire csr_mtvec_29_;
 wire csr_mtvec_2_;
 wire csr_mtvec_30_;
 wire csr_mtvec_31_;
 wire csr_mtvec_3_;
 wire csr_mtvec_4_;
 wire csr_mtvec_5_;
 wire csr_mtvec_6_;
 wire csr_mtvec_7_;
 wire csr_mtvec_8_;
 wire csr_mtvec_9_;
 wire csr_mtvec_init;
 wire csr_op_0_;
 wire csr_op_1_;
 wire csr_op_en;
 wire csr_pmp_addr_0_;
 wire csr_pmp_addr_100_;
 wire csr_pmp_addr_101_;
 wire csr_pmp_addr_102_;
 wire csr_pmp_addr_103_;
 wire csr_pmp_addr_104_;
 wire csr_pmp_addr_105_;
 wire csr_pmp_addr_106_;
 wire csr_pmp_addr_107_;
 wire csr_pmp_addr_108_;
 wire csr_pmp_addr_109_;
 wire csr_pmp_addr_10_;
 wire csr_pmp_addr_110_;
 wire csr_pmp_addr_111_;
 wire csr_pmp_addr_112_;
 wire csr_pmp_addr_113_;
 wire csr_pmp_addr_114_;
 wire csr_pmp_addr_115_;
 wire csr_pmp_addr_116_;
 wire csr_pmp_addr_117_;
 wire csr_pmp_addr_118_;
 wire csr_pmp_addr_119_;
 wire csr_pmp_addr_11_;
 wire csr_pmp_addr_120_;
 wire csr_pmp_addr_121_;
 wire csr_pmp_addr_122_;
 wire csr_pmp_addr_123_;
 wire csr_pmp_addr_124_;
 wire csr_pmp_addr_125_;
 wire csr_pmp_addr_126_;
 wire csr_pmp_addr_127_;
 wire csr_pmp_addr_128_;
 wire csr_pmp_addr_129_;
 wire csr_pmp_addr_12_;
 wire csr_pmp_addr_130_;
 wire csr_pmp_addr_131_;
 wire csr_pmp_addr_132_;
 wire csr_pmp_addr_133_;
 wire csr_pmp_addr_134_;
 wire csr_pmp_addr_135_;
 wire csr_pmp_addr_13_;
 wire csr_pmp_addr_14_;
 wire csr_pmp_addr_15_;
 wire csr_pmp_addr_16_;
 wire csr_pmp_addr_17_;
 wire csr_pmp_addr_18_;
 wire csr_pmp_addr_19_;
 wire csr_pmp_addr_1_;
 wire csr_pmp_addr_20_;
 wire csr_pmp_addr_21_;
 wire csr_pmp_addr_22_;
 wire csr_pmp_addr_23_;
 wire csr_pmp_addr_24_;
 wire csr_pmp_addr_25_;
 wire csr_pmp_addr_26_;
 wire csr_pmp_addr_27_;
 wire csr_pmp_addr_28_;
 wire csr_pmp_addr_29_;
 wire csr_pmp_addr_2_;
 wire csr_pmp_addr_30_;
 wire csr_pmp_addr_31_;
 wire csr_pmp_addr_32_;
 wire csr_pmp_addr_33_;
 wire csr_pmp_addr_34_;
 wire csr_pmp_addr_35_;
 wire csr_pmp_addr_36_;
 wire csr_pmp_addr_37_;
 wire csr_pmp_addr_38_;
 wire csr_pmp_addr_39_;
 wire csr_pmp_addr_3_;
 wire csr_pmp_addr_40_;
 wire csr_pmp_addr_41_;
 wire csr_pmp_addr_42_;
 wire csr_pmp_addr_43_;
 wire csr_pmp_addr_44_;
 wire csr_pmp_addr_45_;
 wire csr_pmp_addr_46_;
 wire csr_pmp_addr_47_;
 wire csr_pmp_addr_48_;
 wire csr_pmp_addr_49_;
 wire csr_pmp_addr_4_;
 wire csr_pmp_addr_50_;
 wire csr_pmp_addr_51_;
 wire csr_pmp_addr_52_;
 wire csr_pmp_addr_53_;
 wire csr_pmp_addr_54_;
 wire csr_pmp_addr_55_;
 wire csr_pmp_addr_56_;
 wire csr_pmp_addr_57_;
 wire csr_pmp_addr_58_;
 wire csr_pmp_addr_59_;
 wire csr_pmp_addr_5_;
 wire csr_pmp_addr_60_;
 wire csr_pmp_addr_61_;
 wire csr_pmp_addr_62_;
 wire csr_pmp_addr_63_;
 wire csr_pmp_addr_64_;
 wire csr_pmp_addr_65_;
 wire csr_pmp_addr_66_;
 wire csr_pmp_addr_67_;
 wire csr_pmp_addr_68_;
 wire csr_pmp_addr_69_;
 wire csr_pmp_addr_6_;
 wire csr_pmp_addr_70_;
 wire csr_pmp_addr_71_;
 wire csr_pmp_addr_72_;
 wire csr_pmp_addr_73_;
 wire csr_pmp_addr_74_;
 wire csr_pmp_addr_75_;
 wire csr_pmp_addr_76_;
 wire csr_pmp_addr_77_;
 wire csr_pmp_addr_78_;
 wire csr_pmp_addr_79_;
 wire csr_pmp_addr_7_;
 wire csr_pmp_addr_80_;
 wire csr_pmp_addr_81_;
 wire csr_pmp_addr_82_;
 wire csr_pmp_addr_83_;
 wire csr_pmp_addr_84_;
 wire csr_pmp_addr_85_;
 wire csr_pmp_addr_86_;
 wire csr_pmp_addr_87_;
 wire csr_pmp_addr_88_;
 wire csr_pmp_addr_89_;
 wire csr_pmp_addr_8_;
 wire csr_pmp_addr_90_;
 wire csr_pmp_addr_91_;
 wire csr_pmp_addr_92_;
 wire csr_pmp_addr_93_;
 wire csr_pmp_addr_94_;
 wire csr_pmp_addr_95_;
 wire csr_pmp_addr_96_;
 wire csr_pmp_addr_97_;
 wire csr_pmp_addr_98_;
 wire csr_pmp_addr_99_;
 wire csr_pmp_addr_9_;
 wire csr_pmp_cfg_0_;
 wire csr_pmp_cfg_10_;
 wire csr_pmp_cfg_11_;
 wire csr_pmp_cfg_12_;
 wire csr_pmp_cfg_13_;
 wire csr_pmp_cfg_14_;
 wire csr_pmp_cfg_15_;
 wire csr_pmp_cfg_16_;
 wire csr_pmp_cfg_17_;
 wire csr_pmp_cfg_18_;
 wire csr_pmp_cfg_19_;
 wire csr_pmp_cfg_1_;
 wire csr_pmp_cfg_20_;
 wire csr_pmp_cfg_21_;
 wire csr_pmp_cfg_22_;
 wire csr_pmp_cfg_23_;
 wire csr_pmp_cfg_2_;
 wire csr_pmp_cfg_3_;
 wire csr_pmp_cfg_4_;
 wire csr_pmp_cfg_5_;
 wire csr_pmp_cfg_6_;
 wire csr_pmp_cfg_7_;
 wire csr_pmp_cfg_8_;
 wire csr_pmp_cfg_9_;
 wire csr_pmp_mseccfg_0_;
 wire csr_pmp_mseccfg_1_;
 wire csr_pmp_mseccfg_2_;
 wire csr_rdata_0_;
 wire csr_rdata_10_;
 wire csr_rdata_11_;
 wire csr_rdata_12_;
 wire csr_rdata_13_;
 wire csr_rdata_14_;
 wire csr_rdata_15_;
 wire csr_rdata_16_;
 wire csr_rdata_17_;
 wire csr_rdata_18_;
 wire csr_rdata_19_;
 wire csr_rdata_1_;
 wire csr_rdata_20_;
 wire csr_rdata_21_;
 wire csr_rdata_22_;
 wire csr_rdata_23_;
 wire csr_rdata_24_;
 wire csr_rdata_25_;
 wire csr_rdata_26_;
 wire csr_rdata_27_;
 wire csr_rdata_28_;
 wire csr_rdata_29_;
 wire csr_rdata_2_;
 wire csr_rdata_30_;
 wire csr_rdata_31_;
 wire csr_rdata_3_;
 wire csr_rdata_4_;
 wire csr_rdata_5_;
 wire csr_rdata_6_;
 wire csr_rdata_7_;
 wire csr_rdata_8_;
 wire csr_rdata_9_;
 wire csr_restore_dret_id;
 wire csr_restore_mret_id;
 wire csr_save_cause;
 wire csr_save_id;
 wire \csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A ;
 wire \csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_B ;
 wire csr_save_if;
 wire \data_be_o_$_MUX__Y_A ;
 wire debug_cause_0_;
 wire debug_cause_1_;
 wire debug_cause_2_;
 wire debug_csr_save;
 wire debug_ebreakm;
 wire debug_ebreaku;
 wire debug_mode;
 wire debug_single_step;
 wire \debug_single_step_$_AND__B_A ;
 wire \div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ;
 wire \div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ;
 wire \div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ;
 wire \div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ;
 wire \ex_block_i.alu_i.imd_val_q_i_0_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_0__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_10_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_10__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_11_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_11__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_12_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_12__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_13_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_13__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_14_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_14__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_15_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_15__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_16_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_16__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_17_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_17__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_18_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_18__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_19_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_19__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_1_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_1__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_20_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_20__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_21_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_21__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_22_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_22__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_23_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_23__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_24_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_24__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_25_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_25__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_26_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_26__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_27_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_27__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_28_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_28__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_29_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_29__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_2_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_2__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_30_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_30__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_31_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_31__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_32_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_33_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_34_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_35_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_36_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_37_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_38_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_39_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_3_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_3__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_40_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_41_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_42_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_43_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_44_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_45_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_46_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_47_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_48_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_49_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_4_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_4__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_50_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_51_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_52_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_53_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_54_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_55_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_56_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_57_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_58_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_59_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_5_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_5__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_60_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_61_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_62_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_63_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_6_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_6__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_7_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_7__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_8_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_8__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.imd_val_q_i_9_ ;
 wire \ex_block_i.alu_i.imd_val_q_i_9__$_NOT__A_Y ;
 wire \ex_block_i.alu_i.instr_first_cycle_i_$_AND__Y_B ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_10__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_11__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_12__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_13__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_14__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_15__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_16__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_17__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_18__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_19__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_1__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_20__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_21__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_22__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_23__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_24__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_25__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_26__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_27__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_28__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_29__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_30__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_31__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_32__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_3__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_4__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_5__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_6__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_7__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_8__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.alu_i.multdiv_operand_b_i_9__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_change_sign_$_AND__Y_B ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_B_$_OR__Y_B_$_AND__Y_A ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_3_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_28_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_10_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_15_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_16_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_18_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_21_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_22_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_23_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_25_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_26_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_27_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_31_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_3_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_5_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_6_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_7_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_9_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_10_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_11_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_12_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_13_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_14_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_15_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_16_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_17_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_18_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_19_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_20_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_21_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_22_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_23_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_24_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_25_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_26_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_27_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_28_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_29_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_30_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_3_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_4_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_5_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_6_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_7_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_8_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_9_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_0_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_10_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_11_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_12_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_13_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_14_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_15_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_16_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_17_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_18_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_19_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_1_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_20_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_21_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_22_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_23_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_24_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_25_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_26_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_27_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_28_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_29_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_2_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_30_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_31_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_3_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_4_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_5_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_6_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_7_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_8_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_9_ ;
 wire \ex_block_i.gen_multdiv_fast.multdiv_i.operator_i_0__$_MUX__Y_A_$_MUX__Y_S_$_OR__Y_B ;
 wire exc_cause_0_;
 wire exc_cause_1_;
 wire exc_cause_2_;
 wire exc_cause_3_;
 wire exc_cause_4_;
 wire exc_cause_5_;
 wire exc_cause_6_;
 wire \g_no_pmp.unused_priv_lvl_ls_0_ ;
 wire \g_no_pmp.unused_priv_lvl_ls_1_ ;
 wire \id_in_ready_$_AND__Y_A_$_AND__Y_A_$_AND__A_Y_$_AND__A_B ;
 wire \id_stage_i.alu_op_b_mux_sel_dec_$_MUX__Y_B_$_OR__Y_A_$_AND__Y_A ;
 wire \id_stage_i.branch_jump_set_done_d ;
 wire \id_stage_i.branch_jump_set_done_q ;
 wire \id_stage_i.branch_set_$_AND__Y_B ;
 wire \id_stage_i.branch_set_raw ;
 wire \id_stage_i.branch_set_raw_d ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__B_A ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ;
 wire \id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs_0_ ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs_1_ ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs_2_ ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs_2__$_NOT__A_Y ;
 wire \id_stage_i.controller_i.ctrl_fsm_cs_3_ ;
 wire \id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ;
 wire \id_stage_i.controller_i.do_single_step_d ;
 wire \id_stage_i.controller_i.do_single_step_q ;
 wire \id_stage_i.controller_i.enter_debug_mode_prio_d ;
 wire \id_stage_i.controller_i.enter_debug_mode_prio_q ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.exc_req_q ;
 wire \id_stage_i.controller_i.handle_irq_$_AND__Y_A_$_AND__Y_B ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.illegal_insn_q ;
 wire \id_stage_i.controller_i.instr_compressed_i_0_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_10_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_11_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_12_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_13_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_14_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_15_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_1_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_2_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_3_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_4_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_5_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_6_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_7_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_8_ ;
 wire \id_stage_i.controller_i.instr_compressed_i_9_ ;
 wire \id_stage_i.controller_i.instr_fetch_err_i ;
 wire \id_stage_i.controller_i.instr_fetch_err_plus2_i ;
 wire \id_stage_i.controller_i.instr_i_0_ ;
 wire \id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ;
 wire \id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ;
 wire \id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ;
 wire \id_stage_i.controller_i.instr_i_10_ ;
 wire \id_stage_i.controller_i.instr_i_11_ ;
 wire \id_stage_i.controller_i.instr_i_12_ ;
 wire \id_stage_i.controller_i.instr_i_13_ ;
 wire \id_stage_i.controller_i.instr_i_14_ ;
 wire \id_stage_i.controller_i.instr_i_15_ ;
 wire \id_stage_i.controller_i.instr_i_16_ ;
 wire \id_stage_i.controller_i.instr_i_17_ ;
 wire \id_stage_i.controller_i.instr_i_18_ ;
 wire \id_stage_i.controller_i.instr_i_19_ ;
 wire \id_stage_i.controller_i.instr_i_1_ ;
 wire \id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ;
 wire \id_stage_i.controller_i.instr_i_20_ ;
 wire \id_stage_i.controller_i.instr_i_21_ ;
 wire \id_stage_i.controller_i.instr_i_22_ ;
 wire \id_stage_i.controller_i.instr_i_23_ ;
 wire \id_stage_i.controller_i.instr_i_24_ ;
 wire \id_stage_i.controller_i.instr_i_25_ ;
 wire \id_stage_i.controller_i.instr_i_26_ ;
 wire \id_stage_i.controller_i.instr_i_27_ ;
 wire \id_stage_i.controller_i.instr_i_28_ ;
 wire \id_stage_i.controller_i.instr_i_29_ ;
 wire \id_stage_i.controller_i.instr_i_2_ ;
 wire \id_stage_i.controller_i.instr_i_30_ ;
 wire \id_stage_i.controller_i.instr_i_31_ ;
 wire \id_stage_i.controller_i.instr_i_3_ ;
 wire \id_stage_i.controller_i.instr_i_4_ ;
 wire \id_stage_i.controller_i.instr_i_5_ ;
 wire \id_stage_i.controller_i.instr_i_6_ ;
 wire \id_stage_i.controller_i.instr_i_7_ ;
 wire \id_stage_i.controller_i.instr_i_8_ ;
 wire \id_stage_i.controller_i.instr_i_9_ ;
 wire \id_stage_i.controller_i.instr_is_compressed_i ;
 wire \id_stage_i.controller_i.instr_valid_i ;
 wire \id_stage_i.controller_i.irqs_i_0_ ;
 wire \id_stage_i.controller_i.irqs_i_10_ ;
 wire \id_stage_i.controller_i.irqs_i_11_ ;
 wire \id_stage_i.controller_i.irqs_i_12_ ;
 wire \id_stage_i.controller_i.irqs_i_13_ ;
 wire \id_stage_i.controller_i.irqs_i_14_ ;
 wire \id_stage_i.controller_i.irqs_i_15_ ;
 wire \id_stage_i.controller_i.irqs_i_16_ ;
 wire \id_stage_i.controller_i.irqs_i_17_ ;
 wire \id_stage_i.controller_i.irqs_i_18_ ;
 wire \id_stage_i.controller_i.irqs_i_1_ ;
 wire \id_stage_i.controller_i.irqs_i_2_ ;
 wire \id_stage_i.controller_i.irqs_i_3_ ;
 wire \id_stage_i.controller_i.irqs_i_4_ ;
 wire \id_stage_i.controller_i.irqs_i_5_ ;
 wire \id_stage_i.controller_i.irqs_i_6_ ;
 wire \id_stage_i.controller_i.irqs_i_7_ ;
 wire \id_stage_i.controller_i.irqs_i_8_ ;
 wire \id_stage_i.controller_i.irqs_i_9_ ;
 wire \id_stage_i.controller_i.load_err_i ;
 wire \id_stage_i.controller_i.load_err_q ;
 wire \id_stage_i.controller_i.nmi_mode_o ;
 wire \id_stage_i.controller_i.perf_jump_o ;
 wire \id_stage_i.controller_i.perf_tbranch_o ;
 wire \id_stage_i.controller_i.priv_mode_i_0_ ;
 wire \id_stage_i.controller_i.priv_mode_i_1_ ;
 wire \id_stage_i.controller_i.store_err_i ;
 wire \id_stage_i.controller_i.store_err_q ;
 wire net1334;
 wire \id_stage_i.controller_i.wfi_insn_i ;
 wire \id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ;
 wire \id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ;
 wire \id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ;
 wire \id_stage_i.decoder_i.illegal_c_insn_i ;
 wire \id_stage_i.id_fsm_q ;
 wire \id_stage_i.illegal_csr_insn_i ;
 wire \id_stage_i.imm_b_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ;
 wire \id_stage_i.instr_perf_count_id_o_$_AND__Y_B ;
 wire \id_stage_i.perf_branch_o ;
 wire \id_stage_i.perf_div_wait_o ;
 wire \id_stage_i.perf_dside_wait_o ;
 wire \if_stage_i.instr_valid_id_d ;
 wire \if_stage_i.prefetch_buffer_i.branch_discard_q_0_ ;
 wire \if_stage_i.prefetch_buffer_i.branch_discard_q_1_ ;
 wire \if_stage_i.prefetch_buffer_i.branch_discard_s_0_ ;
 wire \if_stage_i.prefetch_buffer_i.branch_discard_s_1_ ;
 wire \if_stage_i.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.prefetch_buffer_i.discard_req_q ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_10_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_11_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_12_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_15_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_16_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_17_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_18_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_19_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_20_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_21_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_23_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_24_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_25_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_27_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_28_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_29_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_30_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_31_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_5_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_6_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_7_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_8_ ;
 wire \if_stage_i.prefetch_buffer_i.fetch_addr_q_9_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_busy_0_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_busy_1_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.err_plus2_$_AND__Y_B ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.err_q_2_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.in_valid_i_$_AND__Y_B ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_0_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_1__$_AND__Y_A ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_2__$_AND__Y_A ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_10_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_11_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_12_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_13_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_14_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_15_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_18_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_19_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_20_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_21_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_22_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_24_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_25_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_26_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_27_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_28_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_29_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_2_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_30_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_31_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_32_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_33_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_34_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_35_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_36_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_37_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_38_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_39_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_3_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_40_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_41_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_42_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_43_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_44_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_45_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_46_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_47_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_48_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_49_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_4_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_50_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_51_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_52_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_53_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_54_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_55_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_56_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_57_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_58_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_59_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_5_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_60_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_61_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_62_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_63_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_64_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_65_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_66_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_67_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_68_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_69_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_6_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_70_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_71_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_72_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_73_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_74_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_75_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_76_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_77_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_78_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_79_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_7_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_80_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_81_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_82_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_83_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_84_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_85_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_86_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_87_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_88_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_89_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_8_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_90_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_91_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_92_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_93_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_94_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_95_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_9_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.valid_d_0_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.valid_d_1_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.valid_d_2_ ;
 wire \if_stage_i.prefetch_buffer_i.fifo_i.valid_q_0_ ;
 wire \if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ;
 wire \if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ;
 wire \if_stage_i.prefetch_buffer_i.rdata_outstanding_s_0_ ;
 wire \if_stage_i.prefetch_buffer_i.rdata_outstanding_s_1_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_10_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_11_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_12_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_13_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_14_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_15_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_16_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_17_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_18_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_19_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_20_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_21_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_22_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_23_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_24_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_25_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_26_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_27_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_28_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_29_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_2_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_30_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_31_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_3_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_4_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_5_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_6_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_7_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_8_ ;
 wire \if_stage_i.prefetch_buffer_i.stored_addr_q_9_ ;
 wire \if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__A_B ;
 wire \if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__Y_B ;
 wire \if_stage_i.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.prefetch_buffer_i.valid_req_q ;
 wire \load_store_unit_i.busy_o_$_OR__Y_A_$_OR__A_B ;
 wire \load_store_unit_i.data_sign_ext_q ;
 wire \load_store_unit_i.data_type_q_0_ ;
 wire \load_store_unit_i.data_type_q_0__$_NOT__A_Y ;
 wire \load_store_unit_i.data_type_q_1_ ;
 wire \load_store_unit_i.data_type_q_1__$_NOT__A_Y ;
 wire \load_store_unit_i.data_we_q ;
 wire \load_store_unit_i.handle_misaligned_q ;
 wire \load_store_unit_i.ls_fsm_cs_0_ ;
 wire \load_store_unit_i.ls_fsm_cs_0__$_NOT__A_Y ;
 wire \load_store_unit_i.ls_fsm_cs_1_ ;
 wire \load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ;
 wire \load_store_unit_i.ls_fsm_cs_2_ ;
 wire \load_store_unit_i.lsu_err_q ;
 wire \load_store_unit_i.lsu_err_q_$_NOT__A_Y ;
 wire \load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ;
 wire \load_store_unit_i.perf_load_o ;
 wire \load_store_unit_i.perf_store_o ;
 wire \load_store_unit_i.pmp_err_q ;
 wire \load_store_unit_i.rdata_offset_q_0_ ;
 wire \load_store_unit_i.rdata_offset_q_0__$_NOT__A_Y ;
 wire \load_store_unit_i.rdata_offset_q_1_ ;
 wire \load_store_unit_i.rdata_offset_q_1__$_NOT__A_Y ;
 wire \load_store_unit_i.rdata_q_0_ ;
 wire \load_store_unit_i.rdata_q_10_ ;
 wire \load_store_unit_i.rdata_q_11_ ;
 wire \load_store_unit_i.rdata_q_12_ ;
 wire \load_store_unit_i.rdata_q_13_ ;
 wire \load_store_unit_i.rdata_q_14_ ;
 wire \load_store_unit_i.rdata_q_15_ ;
 wire \load_store_unit_i.rdata_q_16_ ;
 wire \load_store_unit_i.rdata_q_17_ ;
 wire \load_store_unit_i.rdata_q_18_ ;
 wire \load_store_unit_i.rdata_q_19_ ;
 wire \load_store_unit_i.rdata_q_1_ ;
 wire \load_store_unit_i.rdata_q_20_ ;
 wire \load_store_unit_i.rdata_q_21_ ;
 wire \load_store_unit_i.rdata_q_22_ ;
 wire \load_store_unit_i.rdata_q_23_ ;
 wire \load_store_unit_i.rdata_q_2_ ;
 wire \load_store_unit_i.rdata_q_3_ ;
 wire \load_store_unit_i.rdata_q_4_ ;
 wire \load_store_unit_i.rdata_q_5_ ;
 wire \load_store_unit_i.rdata_q_6_ ;
 wire \load_store_unit_i.rdata_q_7_ ;
 wire \load_store_unit_i.rdata_q_8_ ;
 wire \load_store_unit_i.rdata_q_9_ ;
 wire perf_instr_ret_compressed_wb;
 wire perf_instr_ret_wb;
 wire perf_iside_wait;
 wire rf_wdata_wb_0_;
 wire rf_wdata_wb_10_;
 wire rf_wdata_wb_11_;
 wire rf_wdata_wb_12_;
 wire rf_wdata_wb_13_;
 wire rf_wdata_wb_14_;
 wire rf_wdata_wb_15_;
 wire rf_wdata_wb_16_;
 wire rf_wdata_wb_17_;
 wire rf_wdata_wb_18_;
 wire rf_wdata_wb_19_;
 wire rf_wdata_wb_1_;
 wire rf_wdata_wb_20_;
 wire rf_wdata_wb_21_;
 wire rf_wdata_wb_22_;
 wire rf_wdata_wb_23_;
 wire rf_wdata_wb_24_;
 wire rf_wdata_wb_25_;
 wire rf_wdata_wb_26_;
 wire rf_wdata_wb_27_;
 wire rf_wdata_wb_28_;
 wire rf_wdata_wb_29_;
 wire rf_wdata_wb_2_;
 wire rf_wdata_wb_30_;
 wire rf_wdata_wb_31_;
 wire rf_wdata_wb_3_;
 wire rf_wdata_wb_4_;
 wire rf_wdata_wb_5_;
 wire rf_wdata_wb_6_;
 wire rf_wdata_wb_7_;
 wire rf_wdata_wb_8_;
 wire rf_wdata_wb_9_;
 wire rf_we_wb;
 wire \cs_registers_i/_0000_ ;
 wire \cs_registers_i/_0001_ ;
 wire \cs_registers_i/_0002_ ;
 wire \cs_registers_i/_0003_ ;
 wire \cs_registers_i/_0004_ ;
 wire \cs_registers_i/_0005_ ;
 wire \cs_registers_i/_0006_ ;
 wire \cs_registers_i/_0007_ ;
 wire \cs_registers_i/_0008_ ;
 wire \cs_registers_i/_0009_ ;
 wire \cs_registers_i/_0010_ ;
 wire \cs_registers_i/_0011_ ;
 wire \cs_registers_i/_0012_ ;
 wire \cs_registers_i/_0013_ ;
 wire \cs_registers_i/_0014_ ;
 wire \cs_registers_i/_0015_ ;
 wire \cs_registers_i/_0016_ ;
 wire \cs_registers_i/_0017_ ;
 wire \cs_registers_i/_0018_ ;
 wire \cs_registers_i/_0019_ ;
 wire \cs_registers_i/_0020_ ;
 wire \cs_registers_i/_0021_ ;
 wire \cs_registers_i/_0022_ ;
 wire \cs_registers_i/_0023_ ;
 wire \cs_registers_i/_0024_ ;
 wire \cs_registers_i/_0025_ ;
 wire \cs_registers_i/_0026_ ;
 wire \cs_registers_i/_0027_ ;
 wire \cs_registers_i/_0028_ ;
 wire \cs_registers_i/_0029_ ;
 wire \cs_registers_i/_0030_ ;
 wire \cs_registers_i/_0031_ ;
 wire \cs_registers_i/_0032_ ;
 wire \cs_registers_i/_0033_ ;
 wire \cs_registers_i/_0034_ ;
 wire \cs_registers_i/_0035_ ;
 wire \cs_registers_i/_0036_ ;
 wire \cs_registers_i/_0037_ ;
 wire \cs_registers_i/_0038_ ;
 wire \cs_registers_i/_0039_ ;
 wire \cs_registers_i/_0040_ ;
 wire \cs_registers_i/_0041_ ;
 wire \cs_registers_i/_0042_ ;
 wire \cs_registers_i/_0043_ ;
 wire \cs_registers_i/_0044_ ;
 wire \cs_registers_i/_0045_ ;
 wire \cs_registers_i/_0046_ ;
 wire \cs_registers_i/_0047_ ;
 wire \cs_registers_i/_0048_ ;
 wire \cs_registers_i/_0049_ ;
 wire \cs_registers_i/_0050_ ;
 wire \cs_registers_i/_0051_ ;
 wire \cs_registers_i/_0052_ ;
 wire \cs_registers_i/_0053_ ;
 wire \cs_registers_i/_0054_ ;
 wire \cs_registers_i/_0055_ ;
 wire \cs_registers_i/_0056_ ;
 wire \cs_registers_i/_0057_ ;
 wire \cs_registers_i/_0058_ ;
 wire \cs_registers_i/_0059_ ;
 wire \cs_registers_i/_0060_ ;
 wire \cs_registers_i/_0061_ ;
 wire \cs_registers_i/_0062_ ;
 wire \cs_registers_i/_0063_ ;
 wire \cs_registers_i/_0064_ ;
 wire \cs_registers_i/_0065_ ;
 wire \cs_registers_i/_0066_ ;
 wire \cs_registers_i/_0067_ ;
 wire \cs_registers_i/_0068_ ;
 wire \cs_registers_i/_0069_ ;
 wire \cs_registers_i/_0070_ ;
 wire \cs_registers_i/_0071_ ;
 wire \cs_registers_i/_0072_ ;
 wire \cs_registers_i/_0073_ ;
 wire \cs_registers_i/_0074_ ;
 wire \cs_registers_i/_0075_ ;
 wire \cs_registers_i/_0076_ ;
 wire \cs_registers_i/_0077_ ;
 wire \cs_registers_i/_0078_ ;
 wire \cs_registers_i/_0079_ ;
 wire \cs_registers_i/_0080_ ;
 wire \cs_registers_i/_0081_ ;
 wire \cs_registers_i/_0082_ ;
 wire \cs_registers_i/_0083_ ;
 wire \cs_registers_i/_0084_ ;
 wire \cs_registers_i/_0085_ ;
 wire \cs_registers_i/_0086_ ;
 wire \cs_registers_i/_0087_ ;
 wire \cs_registers_i/_0088_ ;
 wire \cs_registers_i/_0089_ ;
 wire \cs_registers_i/_0090_ ;
 wire \cs_registers_i/_0091_ ;
 wire \cs_registers_i/_0092_ ;
 wire \cs_registers_i/_0093_ ;
 wire \cs_registers_i/_0094_ ;
 wire \cs_registers_i/_0095_ ;
 wire \cs_registers_i/_0096_ ;
 wire \cs_registers_i/_0097_ ;
 wire \cs_registers_i/_0098_ ;
 wire \cs_registers_i/_0099_ ;
 wire \cs_registers_i/_0100_ ;
 wire \cs_registers_i/_0101_ ;
 wire \cs_registers_i/_0102_ ;
 wire \cs_registers_i/_0103_ ;
 wire \cs_registers_i/_0104_ ;
 wire \cs_registers_i/_0105_ ;
 wire \cs_registers_i/_0106_ ;
 wire \cs_registers_i/_0107_ ;
 wire \cs_registers_i/_0108_ ;
 wire \cs_registers_i/_0109_ ;
 wire \cs_registers_i/_0110_ ;
 wire \cs_registers_i/_0111_ ;
 wire \cs_registers_i/_0112_ ;
 wire \cs_registers_i/_0113_ ;
 wire \cs_registers_i/_0114_ ;
 wire \cs_registers_i/_0115_ ;
 wire \cs_registers_i/_0116_ ;
 wire \cs_registers_i/_0117_ ;
 wire \cs_registers_i/_0118_ ;
 wire \cs_registers_i/_0119_ ;
 wire \cs_registers_i/_0120_ ;
 wire \cs_registers_i/_0121_ ;
 wire \cs_registers_i/_0122_ ;
 wire \cs_registers_i/_0123_ ;
 wire \cs_registers_i/_0124_ ;
 wire \cs_registers_i/_0125_ ;
 wire \cs_registers_i/_0126_ ;
 wire \cs_registers_i/_0127_ ;
 wire \cs_registers_i/_0128_ ;
 wire \cs_registers_i/_0129_ ;
 wire \cs_registers_i/_0130_ ;
 wire \cs_registers_i/_0131_ ;
 wire \cs_registers_i/_0132_ ;
 wire \cs_registers_i/_0133_ ;
 wire \cs_registers_i/_0134_ ;
 wire \cs_registers_i/_0135_ ;
 wire \cs_registers_i/_0136_ ;
 wire \cs_registers_i/_0137_ ;
 wire \cs_registers_i/_0138_ ;
 wire \cs_registers_i/_0139_ ;
 wire \cs_registers_i/_0140_ ;
 wire \cs_registers_i/_0141_ ;
 wire \cs_registers_i/_0142_ ;
 wire \cs_registers_i/_0143_ ;
 wire \cs_registers_i/_0144_ ;
 wire \cs_registers_i/_0145_ ;
 wire \cs_registers_i/_0146_ ;
 wire \cs_registers_i/_0147_ ;
 wire \cs_registers_i/_0148_ ;
 wire \cs_registers_i/_0149_ ;
 wire \cs_registers_i/_0150_ ;
 wire \cs_registers_i/_0151_ ;
 wire \cs_registers_i/_0152_ ;
 wire \cs_registers_i/_0153_ ;
 wire \cs_registers_i/_0154_ ;
 wire \cs_registers_i/_0155_ ;
 wire \cs_registers_i/_0156_ ;
 wire \cs_registers_i/_0157_ ;
 wire \cs_registers_i/_0158_ ;
 wire \cs_registers_i/_0159_ ;
 wire \cs_registers_i/_0160_ ;
 wire \cs_registers_i/_0161_ ;
 wire \cs_registers_i/_0162_ ;
 wire \cs_registers_i/_0163_ ;
 wire \cs_registers_i/_0164_ ;
 wire \cs_registers_i/_0165_ ;
 wire \cs_registers_i/_0166_ ;
 wire \cs_registers_i/_0167_ ;
 wire \cs_registers_i/_0168_ ;
 wire \cs_registers_i/_0169_ ;
 wire \cs_registers_i/_0170_ ;
 wire \cs_registers_i/_0171_ ;
 wire \cs_registers_i/_0172_ ;
 wire \cs_registers_i/_0173_ ;
 wire \cs_registers_i/_0174_ ;
 wire \cs_registers_i/_0175_ ;
 wire \cs_registers_i/_0176_ ;
 wire \cs_registers_i/_0177_ ;
 wire \cs_registers_i/_0178_ ;
 wire \cs_registers_i/_0179_ ;
 wire \cs_registers_i/_0180_ ;
 wire \cs_registers_i/_0181_ ;
 wire \cs_registers_i/_0182_ ;
 wire \cs_registers_i/_0183_ ;
 wire \cs_registers_i/_0184_ ;
 wire \cs_registers_i/_0185_ ;
 wire \cs_registers_i/_0186_ ;
 wire \cs_registers_i/_0187_ ;
 wire \cs_registers_i/_0188_ ;
 wire \cs_registers_i/_0189_ ;
 wire \cs_registers_i/_0190_ ;
 wire \cs_registers_i/_0191_ ;
 wire \cs_registers_i/_0192_ ;
 wire \cs_registers_i/_0193_ ;
 wire \cs_registers_i/_0194_ ;
 wire \cs_registers_i/_0195_ ;
 wire \cs_registers_i/_0196_ ;
 wire \cs_registers_i/_0197_ ;
 wire \cs_registers_i/_0198_ ;
 wire \cs_registers_i/_0199_ ;
 wire \cs_registers_i/_0200_ ;
 wire \cs_registers_i/_0201_ ;
 wire \cs_registers_i/_0202_ ;
 wire \cs_registers_i/_0203_ ;
 wire \cs_registers_i/_0204_ ;
 wire \cs_registers_i/_0205_ ;
 wire \cs_registers_i/_0206_ ;
 wire \cs_registers_i/_0207_ ;
 wire \cs_registers_i/_0208_ ;
 wire \cs_registers_i/_0209_ ;
 wire \cs_registers_i/_0210_ ;
 wire \cs_registers_i/_0211_ ;
 wire \cs_registers_i/_0212_ ;
 wire \cs_registers_i/_0213_ ;
 wire \cs_registers_i/_0214_ ;
 wire \cs_registers_i/_0215_ ;
 wire \cs_registers_i/_0216_ ;
 wire \cs_registers_i/_0217_ ;
 wire \cs_registers_i/_0218_ ;
 wire \cs_registers_i/_0219_ ;
 wire \cs_registers_i/_0220_ ;
 wire \cs_registers_i/_0221_ ;
 wire \cs_registers_i/_0222_ ;
 wire \cs_registers_i/_0223_ ;
 wire \cs_registers_i/_0224_ ;
 wire \cs_registers_i/_0225_ ;
 wire \cs_registers_i/_0226_ ;
 wire \cs_registers_i/_0227_ ;
 wire \cs_registers_i/_0228_ ;
 wire \cs_registers_i/_0229_ ;
 wire \cs_registers_i/_0230_ ;
 wire \cs_registers_i/_0231_ ;
 wire \cs_registers_i/_0232_ ;
 wire \cs_registers_i/_0233_ ;
 wire \cs_registers_i/_0234_ ;
 wire \cs_registers_i/_0235_ ;
 wire \cs_registers_i/_0236_ ;
 wire \cs_registers_i/_0237_ ;
 wire \cs_registers_i/_0238_ ;
 wire \cs_registers_i/_0239_ ;
 wire \cs_registers_i/_0240_ ;
 wire \cs_registers_i/_0241_ ;
 wire \cs_registers_i/_0242_ ;
 wire \cs_registers_i/_0243_ ;
 wire \cs_registers_i/_0244_ ;
 wire \cs_registers_i/_0245_ ;
 wire \cs_registers_i/_0246_ ;
 wire \cs_registers_i/_0247_ ;
 wire \cs_registers_i/_0248_ ;
 wire \cs_registers_i/_0249_ ;
 wire \cs_registers_i/_0250_ ;
 wire \cs_registers_i/_0251_ ;
 wire \cs_registers_i/_0252_ ;
 wire \cs_registers_i/_0253_ ;
 wire \cs_registers_i/_0254_ ;
 wire \cs_registers_i/_0255_ ;
 wire \cs_registers_i/_0256_ ;
 wire \cs_registers_i/_0257_ ;
 wire \cs_registers_i/_0258_ ;
 wire \cs_registers_i/_0259_ ;
 wire \cs_registers_i/_0260_ ;
 wire \cs_registers_i/_0261_ ;
 wire \cs_registers_i/_0262_ ;
 wire \cs_registers_i/_0263_ ;
 wire \cs_registers_i/_0264_ ;
 wire \cs_registers_i/_0265_ ;
 wire \cs_registers_i/_0266_ ;
 wire \cs_registers_i/_0267_ ;
 wire \cs_registers_i/_0268_ ;
 wire \cs_registers_i/_0269_ ;
 wire \cs_registers_i/_0270_ ;
 wire \cs_registers_i/_0271_ ;
 wire \cs_registers_i/_0272_ ;
 wire \cs_registers_i/_0273_ ;
 wire \cs_registers_i/_0274_ ;
 wire \cs_registers_i/_0275_ ;
 wire \cs_registers_i/_0276_ ;
 wire \cs_registers_i/_0277_ ;
 wire \cs_registers_i/_0278_ ;
 wire \cs_registers_i/_0279_ ;
 wire \cs_registers_i/_0280_ ;
 wire \cs_registers_i/_0281_ ;
 wire \cs_registers_i/_0282_ ;
 wire \cs_registers_i/_0283_ ;
 wire \cs_registers_i/_0284_ ;
 wire \cs_registers_i/_0285_ ;
 wire \cs_registers_i/_0286_ ;
 wire \cs_registers_i/_0287_ ;
 wire \cs_registers_i/_0288_ ;
 wire \cs_registers_i/_0289_ ;
 wire \cs_registers_i/_0290_ ;
 wire \cs_registers_i/_0291_ ;
 wire \cs_registers_i/_0292_ ;
 wire \cs_registers_i/_0293_ ;
 wire \cs_registers_i/_0294_ ;
 wire \cs_registers_i/_0295_ ;
 wire \cs_registers_i/_0296_ ;
 wire \cs_registers_i/_0297_ ;
 wire \cs_registers_i/_0298_ ;
 wire \cs_registers_i/_0299_ ;
 wire \cs_registers_i/_0300_ ;
 wire \cs_registers_i/_0301_ ;
 wire \cs_registers_i/_0302_ ;
 wire \cs_registers_i/_0303_ ;
 wire \cs_registers_i/_0304_ ;
 wire \cs_registers_i/_0305_ ;
 wire \cs_registers_i/_0306_ ;
 wire \cs_registers_i/_0307_ ;
 wire \cs_registers_i/_0308_ ;
 wire \cs_registers_i/_0309_ ;
 wire \cs_registers_i/_0310_ ;
 wire \cs_registers_i/_0311_ ;
 wire \cs_registers_i/_0312_ ;
 wire \cs_registers_i/_0313_ ;
 wire \cs_registers_i/_0314_ ;
 wire \cs_registers_i/_0315_ ;
 wire \cs_registers_i/_0316_ ;
 wire \cs_registers_i/_0317_ ;
 wire \cs_registers_i/_0318_ ;
 wire \cs_registers_i/_0319_ ;
 wire \cs_registers_i/_0320_ ;
 wire \cs_registers_i/_0321_ ;
 wire \cs_registers_i/_0322_ ;
 wire \cs_registers_i/_0323_ ;
 wire \cs_registers_i/_0324_ ;
 wire \cs_registers_i/_0325_ ;
 wire \cs_registers_i/_0326_ ;
 wire \cs_registers_i/_0327_ ;
 wire \cs_registers_i/_0328_ ;
 wire \cs_registers_i/_0329_ ;
 wire \cs_registers_i/_0330_ ;
 wire \cs_registers_i/_0331_ ;
 wire \cs_registers_i/_0332_ ;
 wire \cs_registers_i/_0333_ ;
 wire \cs_registers_i/_0334_ ;
 wire \cs_registers_i/_0335_ ;
 wire \cs_registers_i/_0336_ ;
 wire \cs_registers_i/_0337_ ;
 wire \cs_registers_i/_0338_ ;
 wire \cs_registers_i/_0339_ ;
 wire \cs_registers_i/_0340_ ;
 wire \cs_registers_i/_0341_ ;
 wire \cs_registers_i/_0342_ ;
 wire \cs_registers_i/_0343_ ;
 wire \cs_registers_i/_0344_ ;
 wire \cs_registers_i/_0345_ ;
 wire \cs_registers_i/_0346_ ;
 wire \cs_registers_i/_0347_ ;
 wire \cs_registers_i/_0348_ ;
 wire \cs_registers_i/_0349_ ;
 wire \cs_registers_i/_0350_ ;
 wire \cs_registers_i/_0351_ ;
 wire \cs_registers_i/_0352_ ;
 wire \cs_registers_i/_0353_ ;
 wire \cs_registers_i/_0354_ ;
 wire \cs_registers_i/_0355_ ;
 wire \cs_registers_i/_0356_ ;
 wire \cs_registers_i/_0357_ ;
 wire \cs_registers_i/_0358_ ;
 wire \cs_registers_i/_0359_ ;
 wire \cs_registers_i/_0360_ ;
 wire \cs_registers_i/_0361_ ;
 wire \cs_registers_i/_0362_ ;
 wire \cs_registers_i/_0363_ ;
 wire \cs_registers_i/_0364_ ;
 wire \cs_registers_i/_0365_ ;
 wire \cs_registers_i/_0366_ ;
 wire \cs_registers_i/_0367_ ;
 wire \cs_registers_i/_0368_ ;
 wire \cs_registers_i/_0369_ ;
 wire \cs_registers_i/_0370_ ;
 wire \cs_registers_i/_0371_ ;
 wire \cs_registers_i/_0372_ ;
 wire \cs_registers_i/_0373_ ;
 wire \cs_registers_i/_0374_ ;
 wire \cs_registers_i/_0375_ ;
 wire \cs_registers_i/_0376_ ;
 wire \cs_registers_i/_0377_ ;
 wire \cs_registers_i/_0378_ ;
 wire \cs_registers_i/_0379_ ;
 wire \cs_registers_i/_0380_ ;
 wire \cs_registers_i/_0381_ ;
 wire \cs_registers_i/_0382_ ;
 wire \cs_registers_i/_0383_ ;
 wire \cs_registers_i/_0384_ ;
 wire \cs_registers_i/_0385_ ;
 wire \cs_registers_i/_0386_ ;
 wire \cs_registers_i/_0387_ ;
 wire \cs_registers_i/_0388_ ;
 wire \cs_registers_i/_0389_ ;
 wire \cs_registers_i/_0390_ ;
 wire \cs_registers_i/_0391_ ;
 wire \cs_registers_i/_0392_ ;
 wire \cs_registers_i/_0393_ ;
 wire \cs_registers_i/_0394_ ;
 wire \cs_registers_i/_0395_ ;
 wire \cs_registers_i/_0396_ ;
 wire \cs_registers_i/_0397_ ;
 wire \cs_registers_i/_0398_ ;
 wire \cs_registers_i/_0399_ ;
 wire \cs_registers_i/_0400_ ;
 wire \cs_registers_i/_0401_ ;
 wire \cs_registers_i/_0402_ ;
 wire \cs_registers_i/_0403_ ;
 wire \cs_registers_i/_0404_ ;
 wire \cs_registers_i/_0405_ ;
 wire \cs_registers_i/_0406_ ;
 wire \cs_registers_i/_0407_ ;
 wire \cs_registers_i/_0408_ ;
 wire \cs_registers_i/_0409_ ;
 wire \cs_registers_i/_0410_ ;
 wire \cs_registers_i/_0411_ ;
 wire \cs_registers_i/_0412_ ;
 wire \cs_registers_i/_0413_ ;
 wire \cs_registers_i/_0414_ ;
 wire \cs_registers_i/_0415_ ;
 wire \cs_registers_i/_0416_ ;
 wire \cs_registers_i/_0417_ ;
 wire \cs_registers_i/_0418_ ;
 wire \cs_registers_i/_0419_ ;
 wire \cs_registers_i/_0420_ ;
 wire \cs_registers_i/_0421_ ;
 wire \cs_registers_i/_0422_ ;
 wire \cs_registers_i/_0423_ ;
 wire \cs_registers_i/_0424_ ;
 wire \cs_registers_i/_0425_ ;
 wire \cs_registers_i/_0426_ ;
 wire \cs_registers_i/_0427_ ;
 wire \cs_registers_i/_0428_ ;
 wire \cs_registers_i/_0429_ ;
 wire \cs_registers_i/_0430_ ;
 wire \cs_registers_i/_0431_ ;
 wire \cs_registers_i/_0432_ ;
 wire \cs_registers_i/_0433_ ;
 wire \cs_registers_i/_0434_ ;
 wire \cs_registers_i/_0435_ ;
 wire \cs_registers_i/_0436_ ;
 wire \cs_registers_i/_0437_ ;
 wire \cs_registers_i/_0438_ ;
 wire \cs_registers_i/_0439_ ;
 wire \cs_registers_i/_0440_ ;
 wire \cs_registers_i/_0441_ ;
 wire \cs_registers_i/_0442_ ;
 wire \cs_registers_i/_0443_ ;
 wire \cs_registers_i/_0444_ ;
 wire \cs_registers_i/_0445_ ;
 wire \cs_registers_i/_0446_ ;
 wire \cs_registers_i/_0447_ ;
 wire \cs_registers_i/_0448_ ;
 wire \cs_registers_i/_0449_ ;
 wire \cs_registers_i/_0450_ ;
 wire \cs_registers_i/_0451_ ;
 wire \cs_registers_i/_0452_ ;
 wire \cs_registers_i/_0453_ ;
 wire \cs_registers_i/_0454_ ;
 wire \cs_registers_i/_0455_ ;
 wire \cs_registers_i/_0456_ ;
 wire \cs_registers_i/_0457_ ;
 wire \cs_registers_i/_0458_ ;
 wire \cs_registers_i/_0459_ ;
 wire \cs_registers_i/_0460_ ;
 wire \cs_registers_i/_0461_ ;
 wire \cs_registers_i/_0462_ ;
 wire \cs_registers_i/_0463_ ;
 wire \cs_registers_i/_0464_ ;
 wire \cs_registers_i/_0465_ ;
 wire \cs_registers_i/_0466_ ;
 wire \cs_registers_i/_0467_ ;
 wire \cs_registers_i/_0468_ ;
 wire \cs_registers_i/_0469_ ;
 wire \cs_registers_i/_0470_ ;
 wire \cs_registers_i/_0471_ ;
 wire \cs_registers_i/_0472_ ;
 wire net658;
 wire net657;
 wire net656;
 wire \cs_registers_i/_0476_ ;
 wire \cs_registers_i/_0477_ ;
 wire net655;
 wire net654;
 wire net653;
 wire \cs_registers_i/_0481_ ;
 wire net652;
 wire net651;
 wire \cs_registers_i/_0484_ ;
 wire \cs_registers_i/_0485_ ;
 wire \cs_registers_i/_0486_ ;
 wire net650;
 wire net649;
 wire net648;
 wire \cs_registers_i/_0490_ ;
 wire net647;
 wire \cs_registers_i/_0492_ ;
 wire \cs_registers_i/_0493_ ;
 wire net646;
 wire net645;
 wire net644;
 wire \cs_registers_i/_0497_ ;
 wire \cs_registers_i/_0498_ ;
 wire net643;
 wire \cs_registers_i/_0500_ ;
 wire \cs_registers_i/_0501_ ;
 wire \cs_registers_i/_0502_ ;
 wire \cs_registers_i/_0503_ ;
 wire \cs_registers_i/_0504_ ;
 wire \cs_registers_i/_0505_ ;
 wire \cs_registers_i/_0506_ ;
 wire \cs_registers_i/_0507_ ;
 wire \cs_registers_i/_0508_ ;
 wire \cs_registers_i/_0509_ ;
 wire \cs_registers_i/_0510_ ;
 wire \cs_registers_i/_0511_ ;
 wire \cs_registers_i/_0512_ ;
 wire \cs_registers_i/_0513_ ;
 wire net642;
 wire \cs_registers_i/_0515_ ;
 wire \cs_registers_i/_0516_ ;
 wire \cs_registers_i/_0517_ ;
 wire \cs_registers_i/_0518_ ;
 wire \cs_registers_i/_0519_ ;
 wire \cs_registers_i/_0520_ ;
 wire \cs_registers_i/_0521_ ;
 wire \cs_registers_i/_0522_ ;
 wire net641;
 wire \cs_registers_i/_0524_ ;
 wire \cs_registers_i/_0525_ ;
 wire \cs_registers_i/_0526_ ;
 wire \cs_registers_i/_0527_ ;
 wire \cs_registers_i/_0528_ ;
 wire \cs_registers_i/_0529_ ;
 wire \cs_registers_i/_0530_ ;
 wire \cs_registers_i/_0531_ ;
 wire \cs_registers_i/_0532_ ;
 wire \cs_registers_i/_0533_ ;
 wire \cs_registers_i/_0534_ ;
 wire \cs_registers_i/_0535_ ;
 wire \cs_registers_i/_0536_ ;
 wire \cs_registers_i/_0537_ ;
 wire \cs_registers_i/_0538_ ;
 wire \cs_registers_i/_0539_ ;
 wire \cs_registers_i/_0540_ ;
 wire \cs_registers_i/_0541_ ;
 wire \cs_registers_i/_0542_ ;
 wire \cs_registers_i/_0543_ ;
 wire \cs_registers_i/_0544_ ;
 wire \cs_registers_i/_0545_ ;
 wire \cs_registers_i/_0546_ ;
 wire net640;
 wire \cs_registers_i/_0548_ ;
 wire \cs_registers_i/_0549_ ;
 wire \cs_registers_i/_0550_ ;
 wire \cs_registers_i/_0551_ ;
 wire \cs_registers_i/_0552_ ;
 wire \cs_registers_i/_0553_ ;
 wire \cs_registers_i/_0554_ ;
 wire \cs_registers_i/_0555_ ;
 wire \cs_registers_i/_0556_ ;
 wire \cs_registers_i/_0557_ ;
 wire \cs_registers_i/_0558_ ;
 wire \cs_registers_i/_0559_ ;
 wire \cs_registers_i/_0560_ ;
 wire \cs_registers_i/_0561_ ;
 wire \cs_registers_i/_0562_ ;
 wire \cs_registers_i/_0563_ ;
 wire \cs_registers_i/_0564_ ;
 wire \cs_registers_i/_0565_ ;
 wire \cs_registers_i/_0566_ ;
 wire \cs_registers_i/_0567_ ;
 wire \cs_registers_i/_0568_ ;
 wire net639;
 wire \cs_registers_i/_0570_ ;
 wire \cs_registers_i/_0571_ ;
 wire \cs_registers_i/_0572_ ;
 wire \cs_registers_i/_0573_ ;
 wire \cs_registers_i/_0574_ ;
 wire \cs_registers_i/_0575_ ;
 wire \cs_registers_i/_0576_ ;
 wire \cs_registers_i/_0577_ ;
 wire \cs_registers_i/_0578_ ;
 wire \cs_registers_i/_0579_ ;
 wire \cs_registers_i/_0580_ ;
 wire \cs_registers_i/_0581_ ;
 wire net638;
 wire \cs_registers_i/_0583_ ;
 wire \cs_registers_i/_0584_ ;
 wire net637;
 wire net636;
 wire net635;
 wire \cs_registers_i/_0588_ ;
 wire net634;
 wire \cs_registers_i/_0590_ ;
 wire net633;
 wire \cs_registers_i/_0592_ ;
 wire \cs_registers_i/_0593_ ;
 wire \cs_registers_i/_0594_ ;
 wire net632;
 wire \cs_registers_i/_0596_ ;
 wire net631;
 wire \cs_registers_i/_0598_ ;
 wire \cs_registers_i/_0599_ ;
 wire \cs_registers_i/_0600_ ;
 wire \cs_registers_i/_0601_ ;
 wire net630;
 wire \cs_registers_i/_0603_ ;
 wire \cs_registers_i/_0604_ ;
 wire \cs_registers_i/_0605_ ;
 wire net629;
 wire net628;
 wire net627;
 wire net626;
 wire net625;
 wire net624;
 wire \cs_registers_i/_0612_ ;
 wire \cs_registers_i/_0613_ ;
 wire net623;
 wire net622;
 wire net621;
 wire net620;
 wire net619;
 wire \cs_registers_i/_0619_ ;
 wire \cs_registers_i/_0620_ ;
 wire \cs_registers_i/_0621_ ;
 wire net618;
 wire net617;
 wire \cs_registers_i/_0624_ ;
 wire \cs_registers_i/_0625_ ;
 wire \cs_registers_i/_0626_ ;
 wire \cs_registers_i/_0627_ ;
 wire \cs_registers_i/_0628_ ;
 wire \cs_registers_i/_0629_ ;
 wire \cs_registers_i/_0630_ ;
 wire \cs_registers_i/_0631_ ;
 wire net616;
 wire net615;
 wire \cs_registers_i/_0634_ ;
 wire \cs_registers_i/_0635_ ;
 wire \cs_registers_i/_0636_ ;
 wire net614;
 wire net613;
 wire \cs_registers_i/_0639_ ;
 wire \cs_registers_i/_0640_ ;
 wire net612;
 wire \cs_registers_i/_0642_ ;
 wire net611;
 wire \cs_registers_i/_0644_ ;
 wire \cs_registers_i/_0645_ ;
 wire net610;
 wire net609;
 wire \cs_registers_i/_0648_ ;
 wire \cs_registers_i/_0649_ ;
 wire \cs_registers_i/_0650_ ;
 wire \cs_registers_i/_0651_ ;
 wire \cs_registers_i/_0652_ ;
 wire \cs_registers_i/_0653_ ;
 wire net608;
 wire \cs_registers_i/_0655_ ;
 wire \cs_registers_i/_0656_ ;
 wire net607;
 wire net606;
 wire \cs_registers_i/_0659_ ;
 wire \cs_registers_i/_0660_ ;
 wire \cs_registers_i/_0661_ ;
 wire net605;
 wire net604;
 wire \cs_registers_i/_0664_ ;
 wire \cs_registers_i/_0665_ ;
 wire net603;
 wire \cs_registers_i/_0667_ ;
 wire \cs_registers_i/_0668_ ;
 wire \cs_registers_i/_0669_ ;
 wire \cs_registers_i/_0670_ ;
 wire \cs_registers_i/_0671_ ;
 wire \cs_registers_i/_0672_ ;
 wire \cs_registers_i/_0673_ ;
 wire \cs_registers_i/_0674_ ;
 wire \cs_registers_i/_0675_ ;
 wire \cs_registers_i/_0676_ ;
 wire \cs_registers_i/_0677_ ;
 wire \cs_registers_i/_0678_ ;
 wire \cs_registers_i/_0679_ ;
 wire \cs_registers_i/_0680_ ;
 wire net602;
 wire net601;
 wire \cs_registers_i/_0683_ ;
 wire net600;
 wire \cs_registers_i/_0685_ ;
 wire \cs_registers_i/_0686_ ;
 wire net599;
 wire \cs_registers_i/_0688_ ;
 wire \cs_registers_i/_0689_ ;
 wire net598;
 wire \cs_registers_i/_0691_ ;
 wire net597;
 wire \cs_registers_i/_0693_ ;
 wire \cs_registers_i/_0694_ ;
 wire \cs_registers_i/_0695_ ;
 wire \cs_registers_i/_0696_ ;
 wire \cs_registers_i/_0697_ ;
 wire \cs_registers_i/_0698_ ;
 wire net596;
 wire \cs_registers_i/_0700_ ;
 wire \cs_registers_i/_0701_ ;
 wire \cs_registers_i/_0702_ ;
 wire net595;
 wire net594;
 wire net593;
 wire net592;
 wire \cs_registers_i/_0707_ ;
 wire \cs_registers_i/_0708_ ;
 wire \cs_registers_i/_0709_ ;
 wire \cs_registers_i/_0710_ ;
 wire \cs_registers_i/_0711_ ;
 wire \cs_registers_i/_0712_ ;
 wire \cs_registers_i/_0713_ ;
 wire \cs_registers_i/_0714_ ;
 wire \cs_registers_i/_0715_ ;
 wire net591;
 wire \cs_registers_i/_0717_ ;
 wire \cs_registers_i/_0718_ ;
 wire \cs_registers_i/_0719_ ;
 wire \cs_registers_i/_0720_ ;
 wire \cs_registers_i/_0721_ ;
 wire \cs_registers_i/_0722_ ;
 wire \cs_registers_i/_0723_ ;
 wire \cs_registers_i/_0724_ ;
 wire \cs_registers_i/_0725_ ;
 wire \cs_registers_i/_0726_ ;
 wire net590;
 wire \cs_registers_i/_0728_ ;
 wire net589;
 wire \cs_registers_i/_0730_ ;
 wire \cs_registers_i/_0731_ ;
 wire \cs_registers_i/_0732_ ;
 wire \cs_registers_i/_0733_ ;
 wire \cs_registers_i/_0734_ ;
 wire \cs_registers_i/_0735_ ;
 wire \cs_registers_i/_0736_ ;
 wire \cs_registers_i/_0737_ ;
 wire \cs_registers_i/_0738_ ;
 wire net588;
 wire \cs_registers_i/_0740_ ;
 wire \cs_registers_i/_0741_ ;
 wire \cs_registers_i/_0742_ ;
 wire net587;
 wire net586;
 wire net585;
 wire net584;
 wire \cs_registers_i/_0747_ ;
 wire \cs_registers_i/_0748_ ;
 wire \cs_registers_i/_0749_ ;
 wire \cs_registers_i/_0750_ ;
 wire \cs_registers_i/_0751_ ;
 wire \cs_registers_i/_0752_ ;
 wire net583;
 wire \cs_registers_i/_0754_ ;
 wire \cs_registers_i/_0755_ ;
 wire net582;
 wire \cs_registers_i/_0757_ ;
 wire \cs_registers_i/_0758_ ;
 wire \cs_registers_i/_0759_ ;
 wire \cs_registers_i/_0760_ ;
 wire \cs_registers_i/_0761_ ;
 wire \cs_registers_i/_0762_ ;
 wire \cs_registers_i/_0763_ ;
 wire \cs_registers_i/_0764_ ;
 wire net581;
 wire \cs_registers_i/_0766_ ;
 wire \cs_registers_i/_0767_ ;
 wire \cs_registers_i/_0768_ ;
 wire net580;
 wire \cs_registers_i/_0770_ ;
 wire net579;
 wire \cs_registers_i/_0772_ ;
 wire \cs_registers_i/_0773_ ;
 wire net578;
 wire \cs_registers_i/_0775_ ;
 wire \cs_registers_i/_0776_ ;
 wire \cs_registers_i/_0777_ ;
 wire net577;
 wire \cs_registers_i/_0779_ ;
 wire \cs_registers_i/_0780_ ;
 wire \cs_registers_i/_0781_ ;
 wire \cs_registers_i/_0782_ ;
 wire \cs_registers_i/_0783_ ;
 wire net576;
 wire \cs_registers_i/_0785_ ;
 wire \cs_registers_i/_0786_ ;
 wire \cs_registers_i/_0787_ ;
 wire \cs_registers_i/_0788_ ;
 wire \cs_registers_i/_0789_ ;
 wire \cs_registers_i/_0790_ ;
 wire net575;
 wire \cs_registers_i/_0792_ ;
 wire \cs_registers_i/_0793_ ;
 wire \cs_registers_i/_0794_ ;
 wire \cs_registers_i/_0795_ ;
 wire \cs_registers_i/_0796_ ;
 wire \cs_registers_i/_0797_ ;
 wire \cs_registers_i/_0798_ ;
 wire \cs_registers_i/_0799_ ;
 wire \cs_registers_i/_0800_ ;
 wire \cs_registers_i/_0801_ ;
 wire \cs_registers_i/_0802_ ;
 wire \cs_registers_i/_0803_ ;
 wire \cs_registers_i/_0804_ ;
 wire \cs_registers_i/_0805_ ;
 wire \cs_registers_i/_0806_ ;
 wire \cs_registers_i/_0807_ ;
 wire \cs_registers_i/_0808_ ;
 wire net574;
 wire \cs_registers_i/_0810_ ;
 wire \cs_registers_i/_0811_ ;
 wire net573;
 wire \cs_registers_i/_0813_ ;
 wire \cs_registers_i/_0814_ ;
 wire \cs_registers_i/_0815_ ;
 wire \cs_registers_i/_0816_ ;
 wire \cs_registers_i/_0817_ ;
 wire \cs_registers_i/_0818_ ;
 wire \cs_registers_i/_0819_ ;
 wire \cs_registers_i/_0820_ ;
 wire \cs_registers_i/_0821_ ;
 wire \cs_registers_i/_0822_ ;
 wire \cs_registers_i/_0823_ ;
 wire \cs_registers_i/_0824_ ;
 wire \cs_registers_i/_0825_ ;
 wire \cs_registers_i/_0826_ ;
 wire \cs_registers_i/_0827_ ;
 wire \cs_registers_i/_0828_ ;
 wire \cs_registers_i/_0829_ ;
 wire \cs_registers_i/_0830_ ;
 wire \cs_registers_i/_0831_ ;
 wire \cs_registers_i/_0832_ ;
 wire \cs_registers_i/_0833_ ;
 wire \cs_registers_i/_0834_ ;
 wire net572;
 wire \cs_registers_i/_0836_ ;
 wire \cs_registers_i/_0837_ ;
 wire net571;
 wire net570;
 wire \cs_registers_i/_0840_ ;
 wire net569;
 wire \cs_registers_i/_0842_ ;
 wire \cs_registers_i/_0843_ ;
 wire \cs_registers_i/_0844_ ;
 wire \cs_registers_i/_0845_ ;
 wire \cs_registers_i/_0846_ ;
 wire \cs_registers_i/_0847_ ;
 wire \cs_registers_i/_0848_ ;
 wire \cs_registers_i/_0849_ ;
 wire \cs_registers_i/_0850_ ;
 wire \cs_registers_i/_0851_ ;
 wire \cs_registers_i/_0852_ ;
 wire \cs_registers_i/_0853_ ;
 wire \cs_registers_i/_0854_ ;
 wire \cs_registers_i/_0855_ ;
 wire \cs_registers_i/_0856_ ;
 wire \cs_registers_i/_0857_ ;
 wire \cs_registers_i/_0858_ ;
 wire \cs_registers_i/_0859_ ;
 wire \cs_registers_i/_0860_ ;
 wire net568;
 wire \cs_registers_i/_0862_ ;
 wire \cs_registers_i/_0863_ ;
 wire \cs_registers_i/_0864_ ;
 wire \cs_registers_i/_0865_ ;
 wire \cs_registers_i/_0866_ ;
 wire net567;
 wire net566;
 wire \cs_registers_i/_0869_ ;
 wire \cs_registers_i/_0870_ ;
 wire \cs_registers_i/_0871_ ;
 wire \cs_registers_i/_0872_ ;
 wire net565;
 wire \cs_registers_i/_0874_ ;
 wire \cs_registers_i/_0875_ ;
 wire \cs_registers_i/_0876_ ;
 wire \cs_registers_i/_0877_ ;
 wire \cs_registers_i/_0878_ ;
 wire \cs_registers_i/_0879_ ;
 wire \cs_registers_i/_0880_ ;
 wire \cs_registers_i/_0881_ ;
 wire \cs_registers_i/_0882_ ;
 wire \cs_registers_i/_0883_ ;
 wire net564;
 wire \cs_registers_i/_0885_ ;
 wire \cs_registers_i/_0886_ ;
 wire \cs_registers_i/_0887_ ;
 wire \cs_registers_i/_0888_ ;
 wire \cs_registers_i/_0889_ ;
 wire \cs_registers_i/_0890_ ;
 wire \cs_registers_i/_0891_ ;
 wire \cs_registers_i/_0892_ ;
 wire \cs_registers_i/_0893_ ;
 wire \cs_registers_i/_0894_ ;
 wire \cs_registers_i/_0895_ ;
 wire \cs_registers_i/_0896_ ;
 wire \cs_registers_i/_0897_ ;
 wire \cs_registers_i/_0898_ ;
 wire \cs_registers_i/_0899_ ;
 wire \cs_registers_i/_0900_ ;
 wire \cs_registers_i/_0901_ ;
 wire \cs_registers_i/_0902_ ;
 wire \cs_registers_i/_0903_ ;
 wire net563;
 wire \cs_registers_i/_0905_ ;
 wire net562;
 wire \cs_registers_i/_0907_ ;
 wire \cs_registers_i/_0908_ ;
 wire \cs_registers_i/_0909_ ;
 wire \cs_registers_i/_0910_ ;
 wire \cs_registers_i/_0911_ ;
 wire \cs_registers_i/_0912_ ;
 wire \cs_registers_i/_0913_ ;
 wire \cs_registers_i/_0914_ ;
 wire \cs_registers_i/_0915_ ;
 wire \cs_registers_i/_0916_ ;
 wire \cs_registers_i/_0917_ ;
 wire \cs_registers_i/_0918_ ;
 wire \cs_registers_i/_0919_ ;
 wire \cs_registers_i/_0920_ ;
 wire \cs_registers_i/_0921_ ;
 wire \cs_registers_i/_0922_ ;
 wire \cs_registers_i/_0923_ ;
 wire \cs_registers_i/_0924_ ;
 wire \cs_registers_i/_0925_ ;
 wire \cs_registers_i/_0926_ ;
 wire \cs_registers_i/_0927_ ;
 wire \cs_registers_i/_0928_ ;
 wire \cs_registers_i/_0929_ ;
 wire \cs_registers_i/_0930_ ;
 wire \cs_registers_i/_0931_ ;
 wire \cs_registers_i/_0932_ ;
 wire net561;
 wire net560;
 wire \cs_registers_i/_0935_ ;
 wire \cs_registers_i/_0936_ ;
 wire \cs_registers_i/_0937_ ;
 wire \cs_registers_i/_0938_ ;
 wire \cs_registers_i/_0939_ ;
 wire \cs_registers_i/_0940_ ;
 wire \cs_registers_i/_0941_ ;
 wire \cs_registers_i/_0942_ ;
 wire \cs_registers_i/_0943_ ;
 wire \cs_registers_i/_0944_ ;
 wire \cs_registers_i/_0945_ ;
 wire \cs_registers_i/_0946_ ;
 wire \cs_registers_i/_0947_ ;
 wire \cs_registers_i/_0948_ ;
 wire \cs_registers_i/_0949_ ;
 wire \cs_registers_i/_0950_ ;
 wire \cs_registers_i/_0951_ ;
 wire \cs_registers_i/_0952_ ;
 wire \cs_registers_i/_0953_ ;
 wire \cs_registers_i/_0954_ ;
 wire \cs_registers_i/_0955_ ;
 wire \cs_registers_i/_0956_ ;
 wire \cs_registers_i/_0957_ ;
 wire \cs_registers_i/_0958_ ;
 wire \cs_registers_i/_0959_ ;
 wire \cs_registers_i/_0960_ ;
 wire \cs_registers_i/_0961_ ;
 wire net559;
 wire \cs_registers_i/_0963_ ;
 wire \cs_registers_i/_0964_ ;
 wire \cs_registers_i/_0965_ ;
 wire \cs_registers_i/_0966_ ;
 wire \cs_registers_i/_0967_ ;
 wire \cs_registers_i/_0968_ ;
 wire \cs_registers_i/_0969_ ;
 wire \cs_registers_i/_0970_ ;
 wire \cs_registers_i/_0971_ ;
 wire \cs_registers_i/_0972_ ;
 wire \cs_registers_i/_0973_ ;
 wire \cs_registers_i/_0974_ ;
 wire \cs_registers_i/_0975_ ;
 wire \cs_registers_i/_0976_ ;
 wire \cs_registers_i/_0977_ ;
 wire \cs_registers_i/_0978_ ;
 wire \cs_registers_i/_0979_ ;
 wire \cs_registers_i/_0980_ ;
 wire \cs_registers_i/_0981_ ;
 wire \cs_registers_i/_0982_ ;
 wire \cs_registers_i/_0983_ ;
 wire net558;
 wire \cs_registers_i/_0985_ ;
 wire \cs_registers_i/_0986_ ;
 wire \cs_registers_i/_0987_ ;
 wire \cs_registers_i/_0988_ ;
 wire \cs_registers_i/_0989_ ;
 wire \cs_registers_i/_0990_ ;
 wire \cs_registers_i/_0991_ ;
 wire \cs_registers_i/_0992_ ;
 wire \cs_registers_i/_0993_ ;
 wire \cs_registers_i/_0994_ ;
 wire \cs_registers_i/_0995_ ;
 wire \cs_registers_i/_0996_ ;
 wire \cs_registers_i/_0997_ ;
 wire \cs_registers_i/_0998_ ;
 wire \cs_registers_i/_0999_ ;
 wire \cs_registers_i/_1000_ ;
 wire \cs_registers_i/_1001_ ;
 wire \cs_registers_i/_1002_ ;
 wire \cs_registers_i/_1003_ ;
 wire \cs_registers_i/_1004_ ;
 wire \cs_registers_i/_1005_ ;
 wire \cs_registers_i/_1006_ ;
 wire \cs_registers_i/_1007_ ;
 wire \cs_registers_i/_1008_ ;
 wire \cs_registers_i/_1009_ ;
 wire net557;
 wire \cs_registers_i/_1011_ ;
 wire \cs_registers_i/_1012_ ;
 wire \cs_registers_i/_1013_ ;
 wire \cs_registers_i/_1014_ ;
 wire \cs_registers_i/_1015_ ;
 wire \cs_registers_i/_1016_ ;
 wire \cs_registers_i/_1017_ ;
 wire \cs_registers_i/_1018_ ;
 wire \cs_registers_i/_1019_ ;
 wire \cs_registers_i/_1020_ ;
 wire \cs_registers_i/_1021_ ;
 wire \cs_registers_i/_1022_ ;
 wire \cs_registers_i/_1023_ ;
 wire \cs_registers_i/_1024_ ;
 wire \cs_registers_i/_1025_ ;
 wire \cs_registers_i/_1026_ ;
 wire \cs_registers_i/_1027_ ;
 wire \cs_registers_i/_1028_ ;
 wire \cs_registers_i/_1029_ ;
 wire \cs_registers_i/_1030_ ;
 wire \cs_registers_i/_1031_ ;
 wire \cs_registers_i/_1032_ ;
 wire \cs_registers_i/_1033_ ;
 wire \cs_registers_i/_1034_ ;
 wire \cs_registers_i/_1035_ ;
 wire \cs_registers_i/_1036_ ;
 wire \cs_registers_i/_1037_ ;
 wire \cs_registers_i/_1038_ ;
 wire \cs_registers_i/_1039_ ;
 wire \cs_registers_i/_1040_ ;
 wire \cs_registers_i/_1041_ ;
 wire \cs_registers_i/_1042_ ;
 wire \cs_registers_i/_1043_ ;
 wire \cs_registers_i/_1044_ ;
 wire \cs_registers_i/_1045_ ;
 wire \cs_registers_i/_1046_ ;
 wire \cs_registers_i/_1047_ ;
 wire \cs_registers_i/_1048_ ;
 wire \cs_registers_i/_1049_ ;
 wire \cs_registers_i/_1050_ ;
 wire \cs_registers_i/_1051_ ;
 wire \cs_registers_i/_1052_ ;
 wire net556;
 wire \cs_registers_i/_1054_ ;
 wire \cs_registers_i/_1055_ ;
 wire \cs_registers_i/_1056_ ;
 wire \cs_registers_i/_1057_ ;
 wire \cs_registers_i/_1058_ ;
 wire \cs_registers_i/_1059_ ;
 wire \cs_registers_i/_1060_ ;
 wire \cs_registers_i/_1061_ ;
 wire \cs_registers_i/_1062_ ;
 wire \cs_registers_i/_1063_ ;
 wire \cs_registers_i/_1064_ ;
 wire \cs_registers_i/_1065_ ;
 wire \cs_registers_i/_1066_ ;
 wire \cs_registers_i/_1067_ ;
 wire \cs_registers_i/_1068_ ;
 wire \cs_registers_i/_1069_ ;
 wire \cs_registers_i/_1070_ ;
 wire \cs_registers_i/_1071_ ;
 wire \cs_registers_i/_1072_ ;
 wire \cs_registers_i/_1073_ ;
 wire \cs_registers_i/_1074_ ;
 wire \cs_registers_i/_1075_ ;
 wire \cs_registers_i/_1076_ ;
 wire \cs_registers_i/_1077_ ;
 wire \cs_registers_i/_1078_ ;
 wire \cs_registers_i/_1079_ ;
 wire net555;
 wire \cs_registers_i/_1081_ ;
 wire \cs_registers_i/_1082_ ;
 wire net554;
 wire \cs_registers_i/_1084_ ;
 wire \cs_registers_i/_1085_ ;
 wire \cs_registers_i/_1086_ ;
 wire \cs_registers_i/_1087_ ;
 wire \cs_registers_i/_1088_ ;
 wire \cs_registers_i/_1089_ ;
 wire \cs_registers_i/_1090_ ;
 wire \cs_registers_i/_1091_ ;
 wire \cs_registers_i/_1092_ ;
 wire \cs_registers_i/_1093_ ;
 wire \cs_registers_i/_1094_ ;
 wire \cs_registers_i/_1095_ ;
 wire \cs_registers_i/_1096_ ;
 wire \cs_registers_i/_1097_ ;
 wire \cs_registers_i/_1098_ ;
 wire \cs_registers_i/_1099_ ;
 wire \cs_registers_i/_1100_ ;
 wire net553;
 wire \cs_registers_i/_1102_ ;
 wire \cs_registers_i/_1103_ ;
 wire \cs_registers_i/_1104_ ;
 wire \cs_registers_i/_1105_ ;
 wire \cs_registers_i/_1106_ ;
 wire \cs_registers_i/_1107_ ;
 wire \cs_registers_i/_1108_ ;
 wire \cs_registers_i/_1109_ ;
 wire \cs_registers_i/_1110_ ;
 wire \cs_registers_i/_1111_ ;
 wire \cs_registers_i/_1112_ ;
 wire \cs_registers_i/_1113_ ;
 wire \cs_registers_i/_1114_ ;
 wire \cs_registers_i/_1115_ ;
 wire \cs_registers_i/_1116_ ;
 wire \cs_registers_i/_1117_ ;
 wire \cs_registers_i/_1118_ ;
 wire \cs_registers_i/_1119_ ;
 wire \cs_registers_i/_1120_ ;
 wire \cs_registers_i/_1121_ ;
 wire \cs_registers_i/_1122_ ;
 wire \cs_registers_i/_1123_ ;
 wire \cs_registers_i/_1124_ ;
 wire \cs_registers_i/_1125_ ;
 wire \cs_registers_i/_1126_ ;
 wire \cs_registers_i/_1127_ ;
 wire \cs_registers_i/_1128_ ;
 wire net552;
 wire \cs_registers_i/_1130_ ;
 wire \cs_registers_i/_1131_ ;
 wire \cs_registers_i/_1132_ ;
 wire \cs_registers_i/_1133_ ;
 wire \cs_registers_i/_1134_ ;
 wire \cs_registers_i/_1135_ ;
 wire \cs_registers_i/_1136_ ;
 wire \cs_registers_i/_1137_ ;
 wire \cs_registers_i/_1138_ ;
 wire \cs_registers_i/_1139_ ;
 wire \cs_registers_i/_1140_ ;
 wire \cs_registers_i/_1141_ ;
 wire \cs_registers_i/_1142_ ;
 wire \cs_registers_i/_1143_ ;
 wire \cs_registers_i/_1144_ ;
 wire \cs_registers_i/_1145_ ;
 wire \cs_registers_i/_1146_ ;
 wire \cs_registers_i/_1147_ ;
 wire \cs_registers_i/_1148_ ;
 wire \cs_registers_i/_1149_ ;
 wire \cs_registers_i/_1150_ ;
 wire \cs_registers_i/_1151_ ;
 wire \cs_registers_i/_1152_ ;
 wire net551;
 wire \cs_registers_i/_1154_ ;
 wire net550;
 wire \cs_registers_i/_1156_ ;
 wire \cs_registers_i/_1157_ ;
 wire \cs_registers_i/_1158_ ;
 wire \cs_registers_i/_1159_ ;
 wire \cs_registers_i/_1160_ ;
 wire \cs_registers_i/_1161_ ;
 wire \cs_registers_i/_1162_ ;
 wire \cs_registers_i/_1163_ ;
 wire \cs_registers_i/_1164_ ;
 wire \cs_registers_i/_1165_ ;
 wire \cs_registers_i/_1166_ ;
 wire \cs_registers_i/_1167_ ;
 wire \cs_registers_i/_1168_ ;
 wire \cs_registers_i/_1169_ ;
 wire \cs_registers_i/_1170_ ;
 wire \cs_registers_i/_1171_ ;
 wire \cs_registers_i/_1172_ ;
 wire \cs_registers_i/_1173_ ;
 wire \cs_registers_i/_1174_ ;
 wire \cs_registers_i/_1175_ ;
 wire \cs_registers_i/_1176_ ;
 wire \cs_registers_i/_1177_ ;
 wire \cs_registers_i/_1178_ ;
 wire \cs_registers_i/_1179_ ;
 wire \cs_registers_i/_1180_ ;
 wire \cs_registers_i/_1181_ ;
 wire net549;
 wire net548;
 wire \cs_registers_i/_1184_ ;
 wire \cs_registers_i/_1185_ ;
 wire \cs_registers_i/_1186_ ;
 wire \cs_registers_i/_1187_ ;
 wire \cs_registers_i/_1188_ ;
 wire \cs_registers_i/_1189_ ;
 wire \cs_registers_i/_1190_ ;
 wire \cs_registers_i/_1191_ ;
 wire \cs_registers_i/_1192_ ;
 wire \cs_registers_i/_1193_ ;
 wire \cs_registers_i/_1194_ ;
 wire \cs_registers_i/_1195_ ;
 wire \cs_registers_i/_1196_ ;
 wire \cs_registers_i/_1197_ ;
 wire \cs_registers_i/_1198_ ;
 wire \cs_registers_i/_1199_ ;
 wire \cs_registers_i/_1200_ ;
 wire \cs_registers_i/_1201_ ;
 wire \cs_registers_i/_1202_ ;
 wire \cs_registers_i/_1203_ ;
 wire net547;
 wire \cs_registers_i/_1205_ ;
 wire \cs_registers_i/_1206_ ;
 wire \cs_registers_i/_1207_ ;
 wire \cs_registers_i/_1208_ ;
 wire \cs_registers_i/_1209_ ;
 wire \cs_registers_i/_1210_ ;
 wire \cs_registers_i/_1211_ ;
 wire \cs_registers_i/_1212_ ;
 wire \cs_registers_i/_1213_ ;
 wire \cs_registers_i/_1214_ ;
 wire \cs_registers_i/_1215_ ;
 wire \cs_registers_i/_1216_ ;
 wire \cs_registers_i/_1217_ ;
 wire \cs_registers_i/_1218_ ;
 wire \cs_registers_i/_1219_ ;
 wire \cs_registers_i/_1220_ ;
 wire \cs_registers_i/_1221_ ;
 wire \cs_registers_i/_1222_ ;
 wire \cs_registers_i/_1223_ ;
 wire \cs_registers_i/_1224_ ;
 wire net546;
 wire \cs_registers_i/_1226_ ;
 wire \cs_registers_i/_1227_ ;
 wire \cs_registers_i/_1228_ ;
 wire \cs_registers_i/_1229_ ;
 wire \cs_registers_i/_1230_ ;
 wire \cs_registers_i/_1231_ ;
 wire \cs_registers_i/_1232_ ;
 wire \cs_registers_i/_1233_ ;
 wire \cs_registers_i/_1234_ ;
 wire \cs_registers_i/_1235_ ;
 wire \cs_registers_i/_1236_ ;
 wire \cs_registers_i/_1237_ ;
 wire \cs_registers_i/_1238_ ;
 wire \cs_registers_i/_1239_ ;
 wire \cs_registers_i/_1240_ ;
 wire \cs_registers_i/_1241_ ;
 wire \cs_registers_i/_1242_ ;
 wire \cs_registers_i/_1243_ ;
 wire \cs_registers_i/_1244_ ;
 wire net545;
 wire \cs_registers_i/_1246_ ;
 wire \cs_registers_i/_1247_ ;
 wire \cs_registers_i/_1248_ ;
 wire \cs_registers_i/_1249_ ;
 wire \cs_registers_i/_1250_ ;
 wire \cs_registers_i/_1251_ ;
 wire \cs_registers_i/_1252_ ;
 wire \cs_registers_i/_1253_ ;
 wire \cs_registers_i/_1254_ ;
 wire \cs_registers_i/_1255_ ;
 wire \cs_registers_i/_1256_ ;
 wire \cs_registers_i/_1257_ ;
 wire \cs_registers_i/_1258_ ;
 wire \cs_registers_i/_1259_ ;
 wire \cs_registers_i/_1260_ ;
 wire \cs_registers_i/_1261_ ;
 wire \cs_registers_i/_1262_ ;
 wire \cs_registers_i/_1263_ ;
 wire \cs_registers_i/_1264_ ;
 wire \cs_registers_i/_1265_ ;
 wire \cs_registers_i/_1266_ ;
 wire \cs_registers_i/_1267_ ;
 wire \cs_registers_i/_1268_ ;
 wire \cs_registers_i/_1269_ ;
 wire \cs_registers_i/_1270_ ;
 wire \cs_registers_i/_1271_ ;
 wire \cs_registers_i/_1272_ ;
 wire net544;
 wire \cs_registers_i/_1274_ ;
 wire \cs_registers_i/_1275_ ;
 wire \cs_registers_i/_1276_ ;
 wire \cs_registers_i/_1277_ ;
 wire \cs_registers_i/_1278_ ;
 wire \cs_registers_i/_1279_ ;
 wire \cs_registers_i/_1280_ ;
 wire \cs_registers_i/_1281_ ;
 wire \cs_registers_i/_1282_ ;
 wire \cs_registers_i/_1283_ ;
 wire \cs_registers_i/_1284_ ;
 wire \cs_registers_i/_1285_ ;
 wire \cs_registers_i/_1286_ ;
 wire \cs_registers_i/_1287_ ;
 wire \cs_registers_i/_1288_ ;
 wire \cs_registers_i/_1289_ ;
 wire \cs_registers_i/_1290_ ;
 wire \cs_registers_i/_1291_ ;
 wire \cs_registers_i/_1292_ ;
 wire \cs_registers_i/_1293_ ;
 wire \cs_registers_i/_1294_ ;
 wire \cs_registers_i/_1295_ ;
 wire \cs_registers_i/_1296_ ;
 wire \cs_registers_i/_1297_ ;
 wire \cs_registers_i/_1298_ ;
 wire \cs_registers_i/_1299_ ;
 wire \cs_registers_i/_1300_ ;
 wire \cs_registers_i/_1301_ ;
 wire \cs_registers_i/_1302_ ;
 wire \cs_registers_i/_1303_ ;
 wire \cs_registers_i/_1304_ ;
 wire net543;
 wire \cs_registers_i/_1306_ ;
 wire \cs_registers_i/_1307_ ;
 wire \cs_registers_i/_1308_ ;
 wire \cs_registers_i/_1309_ ;
 wire \cs_registers_i/_1310_ ;
 wire \cs_registers_i/_1311_ ;
 wire \cs_registers_i/_1312_ ;
 wire \cs_registers_i/_1313_ ;
 wire \cs_registers_i/_1314_ ;
 wire \cs_registers_i/_1315_ ;
 wire \cs_registers_i/_1316_ ;
 wire \cs_registers_i/_1317_ ;
 wire \cs_registers_i/_1318_ ;
 wire \cs_registers_i/_1319_ ;
 wire \cs_registers_i/_1320_ ;
 wire \cs_registers_i/_1321_ ;
 wire \cs_registers_i/_1322_ ;
 wire net542;
 wire \cs_registers_i/_1324_ ;
 wire \cs_registers_i/_1325_ ;
 wire \cs_registers_i/_1326_ ;
 wire \cs_registers_i/_1327_ ;
 wire \cs_registers_i/_1328_ ;
 wire \cs_registers_i/_1329_ ;
 wire \cs_registers_i/_1330_ ;
 wire \cs_registers_i/_1331_ ;
 wire \cs_registers_i/_1332_ ;
 wire \cs_registers_i/_1333_ ;
 wire \cs_registers_i/_1334_ ;
 wire \cs_registers_i/_1335_ ;
 wire \cs_registers_i/_1336_ ;
 wire \cs_registers_i/_1337_ ;
 wire \cs_registers_i/_1338_ ;
 wire \cs_registers_i/_1339_ ;
 wire \cs_registers_i/_1340_ ;
 wire \cs_registers_i/_1341_ ;
 wire \cs_registers_i/_1342_ ;
 wire \cs_registers_i/_1343_ ;
 wire \cs_registers_i/_1344_ ;
 wire \cs_registers_i/_1345_ ;
 wire \cs_registers_i/_1346_ ;
 wire \cs_registers_i/_1347_ ;
 wire \cs_registers_i/_1348_ ;
 wire net541;
 wire \cs_registers_i/_1350_ ;
 wire \cs_registers_i/_1351_ ;
 wire \cs_registers_i/_1352_ ;
 wire \cs_registers_i/_1353_ ;
 wire \cs_registers_i/_1354_ ;
 wire \cs_registers_i/_1355_ ;
 wire \cs_registers_i/_1356_ ;
 wire \cs_registers_i/_1357_ ;
 wire \cs_registers_i/_1358_ ;
 wire \cs_registers_i/_1359_ ;
 wire \cs_registers_i/_1360_ ;
 wire \cs_registers_i/_1361_ ;
 wire \cs_registers_i/_1362_ ;
 wire \cs_registers_i/_1363_ ;
 wire \cs_registers_i/_1364_ ;
 wire \cs_registers_i/_1365_ ;
 wire \cs_registers_i/_1366_ ;
 wire \cs_registers_i/_1367_ ;
 wire \cs_registers_i/_1368_ ;
 wire \cs_registers_i/_1369_ ;
 wire net540;
 wire \cs_registers_i/_1371_ ;
 wire \cs_registers_i/_1372_ ;
 wire \cs_registers_i/_1373_ ;
 wire \cs_registers_i/_1374_ ;
 wire \cs_registers_i/_1375_ ;
 wire \cs_registers_i/_1376_ ;
 wire \cs_registers_i/_1377_ ;
 wire \cs_registers_i/_1378_ ;
 wire \cs_registers_i/_1379_ ;
 wire \cs_registers_i/_1380_ ;
 wire \cs_registers_i/_1381_ ;
 wire \cs_registers_i/_1382_ ;
 wire \cs_registers_i/_1383_ ;
 wire \cs_registers_i/_1384_ ;
 wire \cs_registers_i/_1385_ ;
 wire \cs_registers_i/_1386_ ;
 wire \cs_registers_i/_1387_ ;
 wire \cs_registers_i/_1388_ ;
 wire \cs_registers_i/_1389_ ;
 wire \cs_registers_i/_1390_ ;
 wire \cs_registers_i/_1391_ ;
 wire \cs_registers_i/_1392_ ;
 wire \cs_registers_i/_1393_ ;
 wire \cs_registers_i/_1394_ ;
 wire \cs_registers_i/_1395_ ;
 wire \cs_registers_i/_1396_ ;
 wire net539;
 wire \cs_registers_i/_1398_ ;
 wire \cs_registers_i/_1399_ ;
 wire \cs_registers_i/_1400_ ;
 wire net538;
 wire net537;
 wire net536;
 wire \cs_registers_i/_1404_ ;
 wire net535;
 wire net534;
 wire \cs_registers_i/_1407_ ;
 wire \cs_registers_i/_1408_ ;
 wire net533;
 wire \cs_registers_i/_1410_ ;
 wire \cs_registers_i/_1411_ ;
 wire \cs_registers_i/_1412_ ;
 wire net532;
 wire net531;
 wire \cs_registers_i/_1415_ ;
 wire net530;
 wire \cs_registers_i/_1417_ ;
 wire net529;
 wire \cs_registers_i/_1419_ ;
 wire \cs_registers_i/_1420_ ;
 wire \cs_registers_i/_1421_ ;
 wire net528;
 wire net527;
 wire net526;
 wire \cs_registers_i/_1425_ ;
 wire \cs_registers_i/_1426_ ;
 wire \cs_registers_i/_1427_ ;
 wire \cs_registers_i/_1428_ ;
 wire net525;
 wire \cs_registers_i/_1430_ ;
 wire \cs_registers_i/_1431_ ;
 wire \cs_registers_i/_1432_ ;
 wire \cs_registers_i/_1433_ ;
 wire \cs_registers_i/_1434_ ;
 wire \cs_registers_i/_1435_ ;
 wire \cs_registers_i/_1436_ ;
 wire \cs_registers_i/_1437_ ;
 wire \cs_registers_i/_1438_ ;
 wire \cs_registers_i/_1439_ ;
 wire \cs_registers_i/_1440_ ;
 wire \cs_registers_i/_1441_ ;
 wire \cs_registers_i/_1442_ ;
 wire \cs_registers_i/_1443_ ;
 wire \cs_registers_i/_1444_ ;
 wire \cs_registers_i/_1445_ ;
 wire \cs_registers_i/_1446_ ;
 wire \cs_registers_i/_1447_ ;
 wire \cs_registers_i/_1448_ ;
 wire \cs_registers_i/_1449_ ;
 wire \cs_registers_i/_1450_ ;
 wire \cs_registers_i/_1451_ ;
 wire \cs_registers_i/_1452_ ;
 wire net524;
 wire net523;
 wire \cs_registers_i/_1455_ ;
 wire net522;
 wire \cs_registers_i/_1457_ ;
 wire net521;
 wire net520;
 wire \cs_registers_i/_1460_ ;
 wire \cs_registers_i/_1461_ ;
 wire \cs_registers_i/_1462_ ;
 wire \cs_registers_i/_1463_ ;
 wire \cs_registers_i/_1464_ ;
 wire \cs_registers_i/_1465_ ;
 wire \cs_registers_i/_1466_ ;
 wire \cs_registers_i/_1467_ ;
 wire \cs_registers_i/_1468_ ;
 wire net519;
 wire \cs_registers_i/_1470_ ;
 wire \cs_registers_i/_1471_ ;
 wire net518;
 wire \cs_registers_i/_1473_ ;
 wire \cs_registers_i/_1474_ ;
 wire \cs_registers_i/_1475_ ;
 wire \cs_registers_i/_1476_ ;
 wire \cs_registers_i/_1477_ ;
 wire \cs_registers_i/_1478_ ;
 wire net517;
 wire \cs_registers_i/_1480_ ;
 wire \cs_registers_i/_1481_ ;
 wire \cs_registers_i/_1482_ ;
 wire \cs_registers_i/_1483_ ;
 wire \cs_registers_i/_1484_ ;
 wire \cs_registers_i/_1485_ ;
 wire \cs_registers_i/_1486_ ;
 wire \cs_registers_i/_1487_ ;
 wire \cs_registers_i/_1488_ ;
 wire \cs_registers_i/_1489_ ;
 wire \cs_registers_i/_1490_ ;
 wire \cs_registers_i/_1491_ ;
 wire \cs_registers_i/_1492_ ;
 wire \cs_registers_i/_1493_ ;
 wire \cs_registers_i/_1494_ ;
 wire \cs_registers_i/_1495_ ;
 wire \cs_registers_i/_1496_ ;
 wire \cs_registers_i/_1497_ ;
 wire \cs_registers_i/_1498_ ;
 wire \cs_registers_i/_1499_ ;
 wire \cs_registers_i/_1500_ ;
 wire \cs_registers_i/_1501_ ;
 wire \cs_registers_i/_1502_ ;
 wire \cs_registers_i/_1503_ ;
 wire \cs_registers_i/_1504_ ;
 wire \cs_registers_i/_1505_ ;
 wire \cs_registers_i/_1506_ ;
 wire net516;
 wire \cs_registers_i/_1508_ ;
 wire \cs_registers_i/_1509_ ;
 wire \cs_registers_i/_1510_ ;
 wire \cs_registers_i/_1511_ ;
 wire \cs_registers_i/_1512_ ;
 wire \cs_registers_i/_1513_ ;
 wire \cs_registers_i/_1514_ ;
 wire \cs_registers_i/_1515_ ;
 wire \cs_registers_i/_1516_ ;
 wire \cs_registers_i/_1517_ ;
 wire \cs_registers_i/_1518_ ;
 wire \cs_registers_i/_1519_ ;
 wire \cs_registers_i/_1520_ ;
 wire net515;
 wire \cs_registers_i/_1522_ ;
 wire \cs_registers_i/_1523_ ;
 wire \cs_registers_i/_1524_ ;
 wire \cs_registers_i/_1525_ ;
 wire \cs_registers_i/_1526_ ;
 wire \cs_registers_i/_1527_ ;
 wire net514;
 wire \cs_registers_i/_1529_ ;
 wire \cs_registers_i/_1530_ ;
 wire \cs_registers_i/_1531_ ;
 wire \cs_registers_i/_1532_ ;
 wire \cs_registers_i/_1533_ ;
 wire \cs_registers_i/_1534_ ;
 wire \cs_registers_i/_1535_ ;
 wire \cs_registers_i/_1536_ ;
 wire \cs_registers_i/_1537_ ;
 wire \cs_registers_i/_1538_ ;
 wire \cs_registers_i/_1539_ ;
 wire net513;
 wire \cs_registers_i/_1541_ ;
 wire \cs_registers_i/_1542_ ;
 wire \cs_registers_i/_1543_ ;
 wire \cs_registers_i/_1544_ ;
 wire \cs_registers_i/_1545_ ;
 wire \cs_registers_i/_1546_ ;
 wire \cs_registers_i/_1547_ ;
 wire \cs_registers_i/_1548_ ;
 wire \cs_registers_i/_1549_ ;
 wire \cs_registers_i/_1550_ ;
 wire \cs_registers_i/_1551_ ;
 wire \cs_registers_i/_1552_ ;
 wire \cs_registers_i/_1553_ ;
 wire \cs_registers_i/_1554_ ;
 wire \cs_registers_i/_1555_ ;
 wire \cs_registers_i/_1556_ ;
 wire \cs_registers_i/_1557_ ;
 wire \cs_registers_i/_1558_ ;
 wire \cs_registers_i/_1559_ ;
 wire \cs_registers_i/_1560_ ;
 wire \cs_registers_i/_1561_ ;
 wire \cs_registers_i/_1562_ ;
 wire \cs_registers_i/_1563_ ;
 wire \cs_registers_i/_1564_ ;
 wire \cs_registers_i/_1565_ ;
 wire \cs_registers_i/_1566_ ;
 wire \cs_registers_i/_1567_ ;
 wire \cs_registers_i/_1568_ ;
 wire \cs_registers_i/_1569_ ;
 wire \cs_registers_i/_1570_ ;
 wire \cs_registers_i/_1571_ ;
 wire \cs_registers_i/_1572_ ;
 wire \cs_registers_i/_1573_ ;
 wire \cs_registers_i/_1574_ ;
 wire \cs_registers_i/_1575_ ;
 wire \cs_registers_i/_1576_ ;
 wire \cs_registers_i/_1577_ ;
 wire \cs_registers_i/_1578_ ;
 wire net512;
 wire net511;
 wire \cs_registers_i/_1581_ ;
 wire \cs_registers_i/_1582_ ;
 wire \cs_registers_i/_1583_ ;
 wire net510;
 wire \cs_registers_i/_1585_ ;
 wire \cs_registers_i/_1586_ ;
 wire \cs_registers_i/_1587_ ;
 wire \cs_registers_i/_1588_ ;
 wire net509;
 wire net508;
 wire \cs_registers_i/_1591_ ;
 wire net507;
 wire net506;
 wire net505;
 wire \cs_registers_i/_1595_ ;
 wire \cs_registers_i/_1596_ ;
 wire \cs_registers_i/_1597_ ;
 wire \cs_registers_i/_1598_ ;
 wire \cs_registers_i/_1599_ ;
 wire net504;
 wire \cs_registers_i/_1601_ ;
 wire \cs_registers_i/_1602_ ;
 wire \cs_registers_i/_1603_ ;
 wire \cs_registers_i/_1604_ ;
 wire \cs_registers_i/_1605_ ;
 wire \cs_registers_i/_1606_ ;
 wire \cs_registers_i/_1607_ ;
 wire \cs_registers_i/_1608_ ;
 wire \cs_registers_i/_1609_ ;
 wire \cs_registers_i/_1610_ ;
 wire \cs_registers_i/_1611_ ;
 wire \cs_registers_i/_1612_ ;
 wire \cs_registers_i/_1613_ ;
 wire net503;
 wire \cs_registers_i/_1615_ ;
 wire \cs_registers_i/_1616_ ;
 wire \cs_registers_i/_1617_ ;
 wire \cs_registers_i/_1618_ ;
 wire \cs_registers_i/_1619_ ;
 wire net502;
 wire \cs_registers_i/_1621_ ;
 wire \cs_registers_i/_1622_ ;
 wire \cs_registers_i/_1623_ ;
 wire \cs_registers_i/_1624_ ;
 wire \cs_registers_i/_1625_ ;
 wire \cs_registers_i/_1626_ ;
 wire \cs_registers_i/_1627_ ;
 wire net501;
 wire net500;
 wire \cs_registers_i/_1630_ ;
 wire \cs_registers_i/_1631_ ;
 wire \cs_registers_i/_1632_ ;
 wire \cs_registers_i/_1633_ ;
 wire \cs_registers_i/_1634_ ;
 wire \cs_registers_i/_1635_ ;
 wire \cs_registers_i/_1636_ ;
 wire \cs_registers_i/_1637_ ;
 wire \cs_registers_i/_1638_ ;
 wire \cs_registers_i/_1639_ ;
 wire \cs_registers_i/_1640_ ;
 wire \cs_registers_i/_1641_ ;
 wire \cs_registers_i/_1642_ ;
 wire \cs_registers_i/_1643_ ;
 wire \cs_registers_i/_1644_ ;
 wire \cs_registers_i/_1645_ ;
 wire \cs_registers_i/_1646_ ;
 wire \cs_registers_i/_1647_ ;
 wire \cs_registers_i/_1648_ ;
 wire \cs_registers_i/_1649_ ;
 wire \cs_registers_i/_1650_ ;
 wire \cs_registers_i/_1651_ ;
 wire \cs_registers_i/_1652_ ;
 wire \cs_registers_i/_1653_ ;
 wire \cs_registers_i/_1654_ ;
 wire \cs_registers_i/_1655_ ;
 wire \cs_registers_i/_1656_ ;
 wire \cs_registers_i/_1657_ ;
 wire \cs_registers_i/_1658_ ;
 wire \cs_registers_i/_1659_ ;
 wire \cs_registers_i/_1660_ ;
 wire \cs_registers_i/_1661_ ;
 wire \cs_registers_i/_1662_ ;
 wire \cs_registers_i/_1663_ ;
 wire \cs_registers_i/_1664_ ;
 wire \cs_registers_i/_1665_ ;
 wire \cs_registers_i/_1666_ ;
 wire \cs_registers_i/_1667_ ;
 wire \cs_registers_i/_1668_ ;
 wire \cs_registers_i/_1669_ ;
 wire \cs_registers_i/_1670_ ;
 wire \cs_registers_i/_1671_ ;
 wire net499;
 wire net498;
 wire net497;
 wire \cs_registers_i/_1675_ ;
 wire \cs_registers_i/_1676_ ;
 wire \cs_registers_i/_1677_ ;
 wire \cs_registers_i/_1678_ ;
 wire \cs_registers_i/_1679_ ;
 wire \cs_registers_i/_1680_ ;
 wire \cs_registers_i/_1681_ ;
 wire \cs_registers_i/_1682_ ;
 wire \cs_registers_i/_1683_ ;
 wire \cs_registers_i/_1684_ ;
 wire \cs_registers_i/_1685_ ;
 wire \cs_registers_i/_1686_ ;
 wire \cs_registers_i/_1687_ ;
 wire \cs_registers_i/_1688_ ;
 wire \cs_registers_i/_1689_ ;
 wire \cs_registers_i/_1690_ ;
 wire net496;
 wire \cs_registers_i/_1692_ ;
 wire \cs_registers_i/_1693_ ;
 wire \cs_registers_i/_1694_ ;
 wire \cs_registers_i/_1695_ ;
 wire \cs_registers_i/_1696_ ;
 wire net495;
 wire \cs_registers_i/_1698_ ;
 wire \cs_registers_i/_1699_ ;
 wire \cs_registers_i/_1700_ ;
 wire net494;
 wire \cs_registers_i/_1702_ ;
 wire \cs_registers_i/_1703_ ;
 wire net493;
 wire net492;
 wire net491;
 wire \cs_registers_i/_1707_ ;
 wire net490;
 wire net489;
 wire net488;
 wire \cs_registers_i/_1711_ ;
 wire \cs_registers_i/_1712_ ;
 wire \cs_registers_i/_1713_ ;
 wire \cs_registers_i/_1714_ ;
 wire \cs_registers_i/_1715_ ;
 wire \cs_registers_i/_1716_ ;
 wire \cs_registers_i/_1717_ ;
 wire \cs_registers_i/_1718_ ;
 wire \cs_registers_i/_1719_ ;
 wire \cs_registers_i/_1720_ ;
 wire \cs_registers_i/_1721_ ;
 wire \cs_registers_i/_1722_ ;
 wire \cs_registers_i/_1723_ ;
 wire \cs_registers_i/_1724_ ;
 wire \cs_registers_i/_1725_ ;
 wire \cs_registers_i/_1726_ ;
 wire \cs_registers_i/_1727_ ;
 wire net487;
 wire \cs_registers_i/_1729_ ;
 wire \cs_registers_i/_1730_ ;
 wire \cs_registers_i/_1731_ ;
 wire \cs_registers_i/_1732_ ;
 wire \cs_registers_i/_1733_ ;
 wire \cs_registers_i/_1734_ ;
 wire \cs_registers_i/_1735_ ;
 wire \cs_registers_i/_1736_ ;
 wire \cs_registers_i/_1737_ ;
 wire \cs_registers_i/_1738_ ;
 wire \cs_registers_i/_1739_ ;
 wire \cs_registers_i/_1740_ ;
 wire \cs_registers_i/_1741_ ;
 wire \cs_registers_i/_1742_ ;
 wire \cs_registers_i/_1743_ ;
 wire \cs_registers_i/_1744_ ;
 wire \cs_registers_i/_1745_ ;
 wire \cs_registers_i/_1746_ ;
 wire \cs_registers_i/_1747_ ;
 wire \cs_registers_i/_1748_ ;
 wire \cs_registers_i/_1749_ ;
 wire \cs_registers_i/_1750_ ;
 wire \cs_registers_i/_1751_ ;
 wire \cs_registers_i/_1752_ ;
 wire \cs_registers_i/_1753_ ;
 wire \cs_registers_i/_1754_ ;
 wire \cs_registers_i/_1755_ ;
 wire \cs_registers_i/_1756_ ;
 wire \cs_registers_i/_1757_ ;
 wire \cs_registers_i/_1758_ ;
 wire \cs_registers_i/_1759_ ;
 wire \cs_registers_i/_1760_ ;
 wire \cs_registers_i/_1761_ ;
 wire net486;
 wire \cs_registers_i/_1763_ ;
 wire net485;
 wire net484;
 wire \cs_registers_i/_1766_ ;
 wire \cs_registers_i/_1767_ ;
 wire \cs_registers_i/_1768_ ;
 wire \cs_registers_i/_1769_ ;
 wire net483;
 wire \cs_registers_i/_1771_ ;
 wire net482;
 wire \cs_registers_i/_1773_ ;
 wire \cs_registers_i/_1774_ ;
 wire net481;
 wire \cs_registers_i/_1776_ ;
 wire \cs_registers_i/_1777_ ;
 wire \cs_registers_i/_1778_ ;
 wire net480;
 wire \cs_registers_i/_1780_ ;
 wire \cs_registers_i/_1781_ ;
 wire \cs_registers_i/_1782_ ;
 wire net479;
 wire \cs_registers_i/_1784_ ;
 wire \cs_registers_i/_1785_ ;
 wire \cs_registers_i/_1786_ ;
 wire \cs_registers_i/_1787_ ;
 wire \cs_registers_i/_1788_ ;
 wire \cs_registers_i/_1789_ ;
 wire \cs_registers_i/_1790_ ;
 wire \cs_registers_i/_1791_ ;
 wire net478;
 wire net477;
 wire \cs_registers_i/_1794_ ;
 wire \cs_registers_i/_1795_ ;
 wire \cs_registers_i/_1796_ ;
 wire \cs_registers_i/_1797_ ;
 wire \cs_registers_i/_1798_ ;
 wire \cs_registers_i/_1799_ ;
 wire \cs_registers_i/_1800_ ;
 wire net476;
 wire \cs_registers_i/_1802_ ;
 wire \cs_registers_i/_1803_ ;
 wire \cs_registers_i/_1804_ ;
 wire \cs_registers_i/_1805_ ;
 wire \cs_registers_i/_1806_ ;
 wire \cs_registers_i/_1807_ ;
 wire \cs_registers_i/_1808_ ;
 wire \cs_registers_i/_1809_ ;
 wire \cs_registers_i/_1810_ ;
 wire net475;
 wire \cs_registers_i/_1812_ ;
 wire \cs_registers_i/_1813_ ;
 wire \cs_registers_i/_1814_ ;
 wire \cs_registers_i/_1815_ ;
 wire \cs_registers_i/_1816_ ;
 wire \cs_registers_i/_1817_ ;
 wire \cs_registers_i/_1818_ ;
 wire \cs_registers_i/_1819_ ;
 wire \cs_registers_i/_1820_ ;
 wire \cs_registers_i/_1821_ ;
 wire \cs_registers_i/_1822_ ;
 wire \cs_registers_i/_1823_ ;
 wire \cs_registers_i/_1824_ ;
 wire \cs_registers_i/_1825_ ;
 wire net474;
 wire \cs_registers_i/_1827_ ;
 wire \cs_registers_i/_1828_ ;
 wire \cs_registers_i/_1829_ ;
 wire \cs_registers_i/_1830_ ;
 wire \cs_registers_i/_1831_ ;
 wire net473;
 wire \cs_registers_i/_1833_ ;
 wire \cs_registers_i/_1834_ ;
 wire \cs_registers_i/_1835_ ;
 wire \cs_registers_i/_1836_ ;
 wire \cs_registers_i/_1837_ ;
 wire \cs_registers_i/_1838_ ;
 wire \cs_registers_i/_1839_ ;
 wire \cs_registers_i/_1840_ ;
 wire \cs_registers_i/_1841_ ;
 wire \cs_registers_i/_1842_ ;
 wire \cs_registers_i/_1843_ ;
 wire \cs_registers_i/_1844_ ;
 wire \cs_registers_i/_1845_ ;
 wire \cs_registers_i/_1846_ ;
 wire \cs_registers_i/_1847_ ;
 wire \cs_registers_i/_1848_ ;
 wire \cs_registers_i/_1849_ ;
 wire \cs_registers_i/_1850_ ;
 wire \cs_registers_i/_1851_ ;
 wire \cs_registers_i/_1852_ ;
 wire \cs_registers_i/_1853_ ;
 wire \cs_registers_i/_1854_ ;
 wire \cs_registers_i/_1855_ ;
 wire \cs_registers_i/_1856_ ;
 wire \cs_registers_i/_1857_ ;
 wire \cs_registers_i/_1858_ ;
 wire \cs_registers_i/_1859_ ;
 wire \cs_registers_i/_1860_ ;
 wire \cs_registers_i/_1861_ ;
 wire \cs_registers_i/_1862_ ;
 wire \cs_registers_i/_1863_ ;
 wire \cs_registers_i/_1864_ ;
 wire \cs_registers_i/_1865_ ;
 wire \cs_registers_i/_1866_ ;
 wire \cs_registers_i/_1867_ ;
 wire \cs_registers_i/_1868_ ;
 wire \cs_registers_i/_1869_ ;
 wire \cs_registers_i/_1870_ ;
 wire \cs_registers_i/_1871_ ;
 wire \cs_registers_i/_1872_ ;
 wire \cs_registers_i/_1873_ ;
 wire \cs_registers_i/_1874_ ;
 wire \cs_registers_i/_1875_ ;
 wire \cs_registers_i/_1876_ ;
 wire \cs_registers_i/_1877_ ;
 wire \cs_registers_i/_1878_ ;
 wire \cs_registers_i/_1879_ ;
 wire \cs_registers_i/_1880_ ;
 wire \cs_registers_i/_1881_ ;
 wire \cs_registers_i/_1882_ ;
 wire \cs_registers_i/_1883_ ;
 wire \cs_registers_i/_1884_ ;
 wire \cs_registers_i/_1885_ ;
 wire \cs_registers_i/_1886_ ;
 wire \cs_registers_i/_1887_ ;
 wire \cs_registers_i/_1888_ ;
 wire \cs_registers_i/_1889_ ;
 wire \cs_registers_i/_1890_ ;
 wire \cs_registers_i/_1891_ ;
 wire \cs_registers_i/_1892_ ;
 wire \cs_registers_i/_1893_ ;
 wire \cs_registers_i/_1894_ ;
 wire \cs_registers_i/_1895_ ;
 wire \cs_registers_i/_1896_ ;
 wire \cs_registers_i/_1897_ ;
 wire \cs_registers_i/_1898_ ;
 wire net472;
 wire \cs_registers_i/_1900_ ;
 wire \cs_registers_i/_1901_ ;
 wire \cs_registers_i/_1902_ ;
 wire \cs_registers_i/_1903_ ;
 wire \cs_registers_i/_1904_ ;
 wire \cs_registers_i/_1905_ ;
 wire \cs_registers_i/_1906_ ;
 wire \cs_registers_i/_1907_ ;
 wire \cs_registers_i/_1908_ ;
 wire \cs_registers_i/_1909_ ;
 wire \cs_registers_i/_1910_ ;
 wire \cs_registers_i/_1911_ ;
 wire \cs_registers_i/_1912_ ;
 wire \cs_registers_i/_1913_ ;
 wire net471;
 wire \cs_registers_i/_1915_ ;
 wire \cs_registers_i/_1916_ ;
 wire \cs_registers_i/_1917_ ;
 wire \cs_registers_i/_1918_ ;
 wire \cs_registers_i/_1919_ ;
 wire \cs_registers_i/_1920_ ;
 wire \cs_registers_i/_1921_ ;
 wire \cs_registers_i/_1922_ ;
 wire \cs_registers_i/_1923_ ;
 wire \cs_registers_i/_1924_ ;
 wire \cs_registers_i/_1925_ ;
 wire \cs_registers_i/_1926_ ;
 wire net470;
 wire \cs_registers_i/_1928_ ;
 wire \cs_registers_i/_1929_ ;
 wire \cs_registers_i/_1930_ ;
 wire \cs_registers_i/_1931_ ;
 wire \cs_registers_i/_1932_ ;
 wire \cs_registers_i/_1933_ ;
 wire \cs_registers_i/_1934_ ;
 wire net469;
 wire \cs_registers_i/_1936_ ;
 wire \cs_registers_i/_1937_ ;
 wire \cs_registers_i/_1938_ ;
 wire \cs_registers_i/_1939_ ;
 wire \cs_registers_i/_1940_ ;
 wire \cs_registers_i/_1941_ ;
 wire \cs_registers_i/_1942_ ;
 wire \cs_registers_i/_1943_ ;
 wire \cs_registers_i/_1944_ ;
 wire \cs_registers_i/_1945_ ;
 wire \cs_registers_i/_1946_ ;
 wire \cs_registers_i/_1947_ ;
 wire \cs_registers_i/_1948_ ;
 wire \cs_registers_i/_1949_ ;
 wire \cs_registers_i/_1950_ ;
 wire \cs_registers_i/_1951_ ;
 wire \cs_registers_i/_1952_ ;
 wire \cs_registers_i/_1953_ ;
 wire \cs_registers_i/_1954_ ;
 wire \cs_registers_i/_1955_ ;
 wire \cs_registers_i/_1956_ ;
 wire \cs_registers_i/_1957_ ;
 wire \cs_registers_i/_1958_ ;
 wire \cs_registers_i/_1959_ ;
 wire \cs_registers_i/_1960_ ;
 wire \cs_registers_i/_1961_ ;
 wire net468;
 wire \cs_registers_i/_1963_ ;
 wire \cs_registers_i/_1964_ ;
 wire \cs_registers_i/_1965_ ;
 wire \cs_registers_i/_1966_ ;
 wire \cs_registers_i/_1967_ ;
 wire \cs_registers_i/_1968_ ;
 wire \cs_registers_i/_1969_ ;
 wire \cs_registers_i/_1970_ ;
 wire \cs_registers_i/_1971_ ;
 wire \cs_registers_i/_1972_ ;
 wire \cs_registers_i/_1973_ ;
 wire \cs_registers_i/_1974_ ;
 wire \cs_registers_i/_1975_ ;
 wire \cs_registers_i/_1976_ ;
 wire \cs_registers_i/_1977_ ;
 wire \cs_registers_i/_1978_ ;
 wire \cs_registers_i/_1979_ ;
 wire \cs_registers_i/_1980_ ;
 wire \cs_registers_i/_1981_ ;
 wire \cs_registers_i/_1982_ ;
 wire \cs_registers_i/_1983_ ;
 wire \cs_registers_i/_1984_ ;
 wire \cs_registers_i/_1985_ ;
 wire \cs_registers_i/_1986_ ;
 wire \cs_registers_i/_1987_ ;
 wire \cs_registers_i/_1988_ ;
 wire \cs_registers_i/_1989_ ;
 wire \cs_registers_i/_1990_ ;
 wire \cs_registers_i/_1991_ ;
 wire \cs_registers_i/_1992_ ;
 wire \cs_registers_i/_1993_ ;
 wire \cs_registers_i/_1994_ ;
 wire \cs_registers_i/_1995_ ;
 wire \cs_registers_i/_1996_ ;
 wire \cs_registers_i/_1997_ ;
 wire \cs_registers_i/_1998_ ;
 wire \cs_registers_i/_1999_ ;
 wire \cs_registers_i/_2000_ ;
 wire \cs_registers_i/_2001_ ;
 wire \cs_registers_i/_2002_ ;
 wire \cs_registers_i/_2003_ ;
 wire \cs_registers_i/_2004_ ;
 wire \cs_registers_i/_2005_ ;
 wire \cs_registers_i/_2006_ ;
 wire \cs_registers_i/_2007_ ;
 wire \cs_registers_i/_2008_ ;
 wire \cs_registers_i/_2009_ ;
 wire \cs_registers_i/_2010_ ;
 wire \cs_registers_i/_2011_ ;
 wire \cs_registers_i/_2012_ ;
 wire \cs_registers_i/_2013_ ;
 wire \cs_registers_i/_2014_ ;
 wire \cs_registers_i/_2015_ ;
 wire \cs_registers_i/_2016_ ;
 wire \cs_registers_i/_2017_ ;
 wire \cs_registers_i/_2018_ ;
 wire \cs_registers_i/_2019_ ;
 wire \cs_registers_i/_2020_ ;
 wire \cs_registers_i/_2021_ ;
 wire \cs_registers_i/_2022_ ;
 wire \cs_registers_i/_2023_ ;
 wire \cs_registers_i/_2024_ ;
 wire \cs_registers_i/_2025_ ;
 wire \cs_registers_i/_2026_ ;
 wire \cs_registers_i/_2027_ ;
 wire \cs_registers_i/_2028_ ;
 wire \cs_registers_i/_2029_ ;
 wire \cs_registers_i/_2030_ ;
 wire \cs_registers_i/_2031_ ;
 wire \cs_registers_i/_2032_ ;
 wire \cs_registers_i/_2033_ ;
 wire \cs_registers_i/_2034_ ;
 wire \cs_registers_i/_2035_ ;
 wire \cs_registers_i/_2036_ ;
 wire \cs_registers_i/_2037_ ;
 wire \cs_registers_i/_2038_ ;
 wire \cs_registers_i/_2039_ ;
 wire \cs_registers_i/_2040_ ;
 wire \cs_registers_i/_2041_ ;
 wire \cs_registers_i/_2042_ ;
 wire \cs_registers_i/_2043_ ;
 wire \cs_registers_i/_2044_ ;
 wire \cs_registers_i/_2045_ ;
 wire \cs_registers_i/_2046_ ;
 wire \cs_registers_i/_2047_ ;
 wire \cs_registers_i/_2048_ ;
 wire \cs_registers_i/_2049_ ;
 wire \cs_registers_i/_2050_ ;
 wire \cs_registers_i/_2051_ ;
 wire \cs_registers_i/_2052_ ;
 wire \cs_registers_i/_2053_ ;
 wire \cs_registers_i/_2054_ ;
 wire \cs_registers_i/_2055_ ;
 wire \cs_registers_i/_2056_ ;
 wire \cs_registers_i/_2057_ ;
 wire \cs_registers_i/_2058_ ;
 wire \cs_registers_i/_2059_ ;
 wire \cs_registers_i/_2060_ ;
 wire \cs_registers_i/_2061_ ;
 wire \cs_registers_i/_2062_ ;
 wire \cs_registers_i/_2063_ ;
 wire \cs_registers_i/_2064_ ;
 wire \cs_registers_i/_2065_ ;
 wire \cs_registers_i/_2066_ ;
 wire \cs_registers_i/_2067_ ;
 wire \cs_registers_i/_2068_ ;
 wire net467;
 wire net466;
 wire net465;
 wire \cs_registers_i/_2072_ ;
 wire \cs_registers_i/_2073_ ;
 wire \cs_registers_i/_2074_ ;
 wire \cs_registers_i/_2075_ ;
 wire \cs_registers_i/_2076_ ;
 wire net464;
 wire \cs_registers_i/_2078_ ;
 wire \cs_registers_i/_2079_ ;
 wire \cs_registers_i/_2080_ ;
 wire \cs_registers_i/_2081_ ;
 wire \cs_registers_i/_2082_ ;
 wire \cs_registers_i/_2083_ ;
 wire \cs_registers_i/_2084_ ;
 wire \cs_registers_i/_2085_ ;
 wire \cs_registers_i/_2086_ ;
 wire \cs_registers_i/_2087_ ;
 wire \cs_registers_i/_2088_ ;
 wire \cs_registers_i/_2089_ ;
 wire \cs_registers_i/_2090_ ;
 wire \cs_registers_i/_2091_ ;
 wire \cs_registers_i/_2092_ ;
 wire \cs_registers_i/_2093_ ;
 wire net463;
 wire \cs_registers_i/_2095_ ;
 wire \cs_registers_i/_2096_ ;
 wire \cs_registers_i/_2097_ ;
 wire \cs_registers_i/_2098_ ;
 wire \cs_registers_i/_2099_ ;
 wire \cs_registers_i/_2100_ ;
 wire \cs_registers_i/_2101_ ;
 wire \cs_registers_i/_2102_ ;
 wire \cs_registers_i/_2103_ ;
 wire \cs_registers_i/_2104_ ;
 wire \cs_registers_i/_2105_ ;
 wire \cs_registers_i/_2106_ ;
 wire \cs_registers_i/_2107_ ;
 wire \cs_registers_i/_2108_ ;
 wire \cs_registers_i/_2109_ ;
 wire \cs_registers_i/_2110_ ;
 wire net462;
 wire \cs_registers_i/_2112_ ;
 wire \cs_registers_i/_2113_ ;
 wire \cs_registers_i/_2114_ ;
 wire \cs_registers_i/_2115_ ;
 wire \cs_registers_i/_2116_ ;
 wire \cs_registers_i/_2117_ ;
 wire \cs_registers_i/_2118_ ;
 wire \cs_registers_i/_2119_ ;
 wire \cs_registers_i/_2120_ ;
 wire \cs_registers_i/_2121_ ;
 wire \cs_registers_i/_2122_ ;
 wire \cs_registers_i/_2123_ ;
 wire \cs_registers_i/_2124_ ;
 wire \cs_registers_i/_2125_ ;
 wire \cs_registers_i/_2126_ ;
 wire \cs_registers_i/_2127_ ;
 wire \cs_registers_i/_2128_ ;
 wire \cs_registers_i/_2129_ ;
 wire \cs_registers_i/_2130_ ;
 wire \cs_registers_i/_2131_ ;
 wire \cs_registers_i/_2132_ ;
 wire \cs_registers_i/_2133_ ;
 wire \cs_registers_i/_2134_ ;
 wire \cs_registers_i/_2135_ ;
 wire \cs_registers_i/_2136_ ;
 wire \cs_registers_i/_2137_ ;
 wire \cs_registers_i/_2138_ ;
 wire \cs_registers_i/_2139_ ;
 wire net461;
 wire \cs_registers_i/_2141_ ;
 wire \cs_registers_i/_2142_ ;
 wire \cs_registers_i/_2143_ ;
 wire \cs_registers_i/_2144_ ;
 wire \cs_registers_i/_2145_ ;
 wire \cs_registers_i/_2146_ ;
 wire \cs_registers_i/_2147_ ;
 wire \cs_registers_i/_2148_ ;
 wire \cs_registers_i/_2149_ ;
 wire \cs_registers_i/_2150_ ;
 wire \cs_registers_i/_2151_ ;
 wire \cs_registers_i/_2152_ ;
 wire \cs_registers_i/_2153_ ;
 wire \cs_registers_i/_2154_ ;
 wire \cs_registers_i/_2155_ ;
 wire \cs_registers_i/_2156_ ;
 wire \cs_registers_i/_2157_ ;
 wire \cs_registers_i/_2158_ ;
 wire \cs_registers_i/_2159_ ;
 wire \cs_registers_i/_2160_ ;
 wire \cs_registers_i/_2161_ ;
 wire \cs_registers_i/_2162_ ;
 wire \cs_registers_i/_2163_ ;
 wire \cs_registers_i/_2164_ ;
 wire \cs_registers_i/_2165_ ;
 wire \cs_registers_i/_2166_ ;
 wire net460;
 wire \cs_registers_i/_2168_ ;
 wire \cs_registers_i/_2169_ ;
 wire \cs_registers_i/_2170_ ;
 wire \cs_registers_i/_2171_ ;
 wire \cs_registers_i/_2172_ ;
 wire \cs_registers_i/_2173_ ;
 wire \cs_registers_i/_2174_ ;
 wire \cs_registers_i/_2175_ ;
 wire \cs_registers_i/_2176_ ;
 wire \cs_registers_i/_2177_ ;
 wire \cs_registers_i/_2178_ ;
 wire net459;
 wire \cs_registers_i/_2180_ ;
 wire \cs_registers_i/_2181_ ;
 wire \cs_registers_i/_2182_ ;
 wire \cs_registers_i/_2183_ ;
 wire \cs_registers_i/_2184_ ;
 wire net458;
 wire \cs_registers_i/_2186_ ;
 wire \cs_registers_i/_2187_ ;
 wire \cs_registers_i/_2188_ ;
 wire \cs_registers_i/_2189_ ;
 wire \cs_registers_i/_2190_ ;
 wire \cs_registers_i/_2191_ ;
 wire net457;
 wire \cs_registers_i/_2193_ ;
 wire \cs_registers_i/_2194_ ;
 wire \cs_registers_i/_2195_ ;
 wire net456;
 wire \cs_registers_i/_2197_ ;
 wire \cs_registers_i/_2198_ ;
 wire \cs_registers_i/_2199_ ;
 wire \cs_registers_i/_2200_ ;
 wire \cs_registers_i/_2201_ ;
 wire \cs_registers_i/_2202_ ;
 wire \cs_registers_i/_2203_ ;
 wire \cs_registers_i/_2204_ ;
 wire \cs_registers_i/_2205_ ;
 wire \cs_registers_i/_2206_ ;
 wire \cs_registers_i/_2207_ ;
 wire \cs_registers_i/_2208_ ;
 wire \cs_registers_i/_2209_ ;
 wire \cs_registers_i/_2210_ ;
 wire \cs_registers_i/_2211_ ;
 wire \cs_registers_i/_2212_ ;
 wire \cs_registers_i/_2213_ ;
 wire \cs_registers_i/_2214_ ;
 wire \cs_registers_i/_2215_ ;
 wire \cs_registers_i/_2216_ ;
 wire \cs_registers_i/_2217_ ;
 wire \cs_registers_i/_2218_ ;
 wire \cs_registers_i/_2219_ ;
 wire \cs_registers_i/_2220_ ;
 wire \cs_registers_i/_2221_ ;
 wire \cs_registers_i/_2222_ ;
 wire \cs_registers_i/_2223_ ;
 wire \cs_registers_i/_2224_ ;
 wire \cs_registers_i/_2225_ ;
 wire \cs_registers_i/_2226_ ;
 wire \cs_registers_i/_2227_ ;
 wire \cs_registers_i/_2228_ ;
 wire \cs_registers_i/_2229_ ;
 wire \cs_registers_i/_2230_ ;
 wire \cs_registers_i/_2231_ ;
 wire \cs_registers_i/_2232_ ;
 wire \cs_registers_i/_2233_ ;
 wire \cs_registers_i/_2234_ ;
 wire \cs_registers_i/_2235_ ;
 wire \cs_registers_i/_2236_ ;
 wire \cs_registers_i/_2237_ ;
 wire \cs_registers_i/_2238_ ;
 wire \cs_registers_i/_2239_ ;
 wire \cs_registers_i/_2240_ ;
 wire \cs_registers_i/_2241_ ;
 wire \cs_registers_i/_2242_ ;
 wire \cs_registers_i/_2243_ ;
 wire \cs_registers_i/_2244_ ;
 wire \cs_registers_i/_2245_ ;
 wire \cs_registers_i/_2246_ ;
 wire \cs_registers_i/_2247_ ;
 wire \cs_registers_i/_2248_ ;
 wire \cs_registers_i/_2249_ ;
 wire \cs_registers_i/_2250_ ;
 wire \cs_registers_i/_2251_ ;
 wire \cs_registers_i/_2252_ ;
 wire \cs_registers_i/_2253_ ;
 wire \cs_registers_i/_2254_ ;
 wire \cs_registers_i/_2255_ ;
 wire \cs_registers_i/_2256_ ;
 wire \cs_registers_i/_2257_ ;
 wire \cs_registers_i/_2258_ ;
 wire \cs_registers_i/_2259_ ;
 wire \cs_registers_i/_2260_ ;
 wire \cs_registers_i/_2261_ ;
 wire \cs_registers_i/_2262_ ;
 wire \cs_registers_i/_2263_ ;
 wire \cs_registers_i/_2264_ ;
 wire \cs_registers_i/_2265_ ;
 wire \cs_registers_i/_2266_ ;
 wire \cs_registers_i/_2267_ ;
 wire \cs_registers_i/_2268_ ;
 wire \cs_registers_i/_2269_ ;
 wire \cs_registers_i/_2270_ ;
 wire \cs_registers_i/_2271_ ;
 wire \cs_registers_i/_2272_ ;
 wire \cs_registers_i/_2273_ ;
 wire \cs_registers_i/_2274_ ;
 wire \cs_registers_i/_2275_ ;
 wire \cs_registers_i/_2276_ ;
 wire \cs_registers_i/_2277_ ;
 wire \cs_registers_i/_2278_ ;
 wire \cs_registers_i/_2279_ ;
 wire \cs_registers_i/_2280_ ;
 wire \cs_registers_i/_2281_ ;
 wire \cs_registers_i/_2282_ ;
 wire \cs_registers_i/_2283_ ;
 wire \cs_registers_i/_2284_ ;
 wire \cs_registers_i/_2285_ ;
 wire \cs_registers_i/_2286_ ;
 wire \cs_registers_i/_2287_ ;
 wire \cs_registers_i/_2288_ ;
 wire \cs_registers_i/_2289_ ;
 wire \cs_registers_i/_2290_ ;
 wire \cs_registers_i/_2291_ ;
 wire \cs_registers_i/_2292_ ;
 wire \cs_registers_i/_2293_ ;
 wire \cs_registers_i/_2294_ ;
 wire \cs_registers_i/_2295_ ;
 wire \cs_registers_i/_2296_ ;
 wire \cs_registers_i/_2297_ ;
 wire \cs_registers_i/_2298_ ;
 wire \cs_registers_i/_2299_ ;
 wire \cs_registers_i/_2300_ ;
 wire \cs_registers_i/_2301_ ;
 wire \cs_registers_i/_2302_ ;
 wire \cs_registers_i/_2303_ ;
 wire \cs_registers_i/_2304_ ;
 wire \cs_registers_i/_2305_ ;
 wire \cs_registers_i/_2306_ ;
 wire \cs_registers_i/_2307_ ;
 wire \cs_registers_i/_2308_ ;
 wire \cs_registers_i/_2309_ ;
 wire \cs_registers_i/_2310_ ;
 wire \cs_registers_i/_2311_ ;
 wire \cs_registers_i/_2312_ ;
 wire \cs_registers_i/_2313_ ;
 wire \cs_registers_i/_2314_ ;
 wire \cs_registers_i/_2315_ ;
 wire \cs_registers_i/_2316_ ;
 wire \cs_registers_i/_2317_ ;
 wire \cs_registers_i/_2318_ ;
 wire \cs_registers_i/_2319_ ;
 wire \cs_registers_i/_2320_ ;
 wire \cs_registers_i/_2321_ ;
 wire \cs_registers_i/_2322_ ;
 wire \cs_registers_i/_2323_ ;
 wire \cs_registers_i/_2324_ ;
 wire \cs_registers_i/_2325_ ;
 wire \cs_registers_i/_2326_ ;
 wire \cs_registers_i/_2327_ ;
 wire \cs_registers_i/_2328_ ;
 wire \cs_registers_i/_2329_ ;
 wire \cs_registers_i/_2330_ ;
 wire net455;
 wire net454;
 wire \cs_registers_i/_2333_ ;
 wire net453;
 wire net452;
 wire net451;
 wire net450;
 wire net449;
 wire net448;
 wire net447;
 wire \cs_registers_i/_2341_ ;
 wire \cs_registers_i/_2342_ ;
 wire \cs_registers_i/_2343_ ;
 wire \cs_registers_i/_2344_ ;
 wire \cs_registers_i/_2345_ ;
 wire \cs_registers_i/_2346_ ;
 wire \cs_registers_i/_2347_ ;
 wire \cs_registers_i/_2348_ ;
 wire \cs_registers_i/_2349_ ;
 wire \cs_registers_i/_2350_ ;
 wire \cs_registers_i/_2351_ ;
 wire \cs_registers_i/_2352_ ;
 wire \cs_registers_i/_2353_ ;
 wire \cs_registers_i/_2354_ ;
 wire \cs_registers_i/_2355_ ;
 wire \cs_registers_i/_2356_ ;
 wire \cs_registers_i/_2357_ ;
 wire \cs_registers_i/_2358_ ;
 wire \cs_registers_i/_2359_ ;
 wire net446;
 wire \cs_registers_i/_2361_ ;
 wire net445;
 wire net444;
 wire net443;
 wire \cs_registers_i/_2365_ ;
 wire \cs_registers_i/_2366_ ;
 wire net442;
 wire \cs_registers_i/_2368_ ;
 wire \cs_registers_i/_2369_ ;
 wire \cs_registers_i/_2370_ ;
 wire \cs_registers_i/_2371_ ;
 wire \cs_registers_i/_2372_ ;
 wire \cs_registers_i/_2373_ ;
 wire \cs_registers_i/_2374_ ;
 wire \cs_registers_i/_2375_ ;
 wire \cs_registers_i/_2376_ ;
 wire \cs_registers_i/_2377_ ;
 wire \cs_registers_i/_2378_ ;
 wire \cs_registers_i/_2379_ ;
 wire \cs_registers_i/_2380_ ;
 wire \cs_registers_i/_2381_ ;
 wire \cs_registers_i/_2382_ ;
 wire \cs_registers_i/_2383_ ;
 wire \cs_registers_i/_2384_ ;
 wire \cs_registers_i/_2385_ ;
 wire \cs_registers_i/_2386_ ;
 wire \cs_registers_i/_2387_ ;
 wire \cs_registers_i/_2388_ ;
 wire \cs_registers_i/_2389_ ;
 wire net441;
 wire \cs_registers_i/_2391_ ;
 wire \cs_registers_i/_2392_ ;
 wire net440;
 wire \cs_registers_i/_2394_ ;
 wire \cs_registers_i/_2395_ ;
 wire \cs_registers_i/_2396_ ;
 wire \cs_registers_i/_2397_ ;
 wire net439;
 wire net438;
 wire \cs_registers_i/_2400_ ;
 wire \cs_registers_i/_2401_ ;
 wire \cs_registers_i/_2402_ ;
 wire \cs_registers_i/_2403_ ;
 wire \cs_registers_i/_2404_ ;
 wire \cs_registers_i/_2405_ ;
 wire \cs_registers_i/_2406_ ;
 wire \cs_registers_i/_2407_ ;
 wire \cs_registers_i/_2408_ ;
 wire \cs_registers_i/_2409_ ;
 wire \cs_registers_i/_2410_ ;
 wire \cs_registers_i/_2411_ ;
 wire \cs_registers_i/_2412_ ;
 wire \cs_registers_i/_2413_ ;
 wire \cs_registers_i/_2414_ ;
 wire \cs_registers_i/_2415_ ;
 wire \cs_registers_i/_2416_ ;
 wire \cs_registers_i/_2417_ ;
 wire \cs_registers_i/_2418_ ;
 wire \cs_registers_i/_2419_ ;
 wire \cs_registers_i/_2420_ ;
 wire \cs_registers_i/_2421_ ;
 wire \cs_registers_i/_2422_ ;
 wire \cs_registers_i/_2423_ ;
 wire net437;
 wire \cs_registers_i/_2425_ ;
 wire \cs_registers_i/_2426_ ;
 wire net436;
 wire \cs_registers_i/_2428_ ;
 wire \cs_registers_i/_2429_ ;
 wire \cs_registers_i/_2430_ ;
 wire \cs_registers_i/_2431_ ;
 wire net435;
 wire net434;
 wire \cs_registers_i/_2434_ ;
 wire \cs_registers_i/_2435_ ;
 wire \cs_registers_i/_2436_ ;
 wire \cs_registers_i/_2437_ ;
 wire \cs_registers_i/_2438_ ;
 wire \cs_registers_i/_2439_ ;
 wire \cs_registers_i/_2440_ ;
 wire \cs_registers_i/_2441_ ;
 wire \cs_registers_i/_2442_ ;
 wire \cs_registers_i/_2443_ ;
 wire \cs_registers_i/_2444_ ;
 wire \cs_registers_i/_2445_ ;
 wire \cs_registers_i/_2446_ ;
 wire \cs_registers_i/_2447_ ;
 wire \cs_registers_i/_2448_ ;
 wire \cs_registers_i/_2449_ ;
 wire \cs_registers_i/_2450_ ;
 wire \cs_registers_i/_2451_ ;
 wire \cs_registers_i/_2452_ ;
 wire \cs_registers_i/_2453_ ;
 wire \cs_registers_i/_2454_ ;
 wire \cs_registers_i/_2455_ ;
 wire \cs_registers_i/_2456_ ;
 wire \cs_registers_i/_2457_ ;
 wire \cs_registers_i/_2458_ ;
 wire \cs_registers_i/_2459_ ;
 wire \cs_registers_i/_2460_ ;
 wire \cs_registers_i/_2461_ ;
 wire \cs_registers_i/_2462_ ;
 wire \cs_registers_i/_2463_ ;
 wire \cs_registers_i/_2464_ ;
 wire \cs_registers_i/_2465_ ;
 wire \cs_registers_i/_2466_ ;
 wire \cs_registers_i/_2467_ ;
 wire \cs_registers_i/_2468_ ;
 wire \cs_registers_i/_2469_ ;
 wire \cs_registers_i/_2470_ ;
 wire \cs_registers_i/_2471_ ;
 wire \cs_registers_i/_2472_ ;
 wire \cs_registers_i/_2473_ ;
 wire \cs_registers_i/_2474_ ;
 wire \cs_registers_i/_2475_ ;
 wire \cs_registers_i/_2476_ ;
 wire \cs_registers_i/_2477_ ;
 wire \cs_registers_i/_2478_ ;
 wire \cs_registers_i/_2479_ ;
 wire \cs_registers_i/_2480_ ;
 wire \cs_registers_i/_2481_ ;
 wire \cs_registers_i/_2482_ ;
 wire \cs_registers_i/_2483_ ;
 wire \cs_registers_i/_2484_ ;
 wire \cs_registers_i/_2485_ ;
 wire \cs_registers_i/_2486_ ;
 wire \cs_registers_i/_2487_ ;
 wire \cs_registers_i/_2488_ ;
 wire \cs_registers_i/_2489_ ;
 wire \cs_registers_i/_2490_ ;
 wire \cs_registers_i/_2491_ ;
 wire \cs_registers_i/_2492_ ;
 wire \cs_registers_i/_2493_ ;
 wire \cs_registers_i/_2494_ ;
 wire \cs_registers_i/_2495_ ;
 wire \cs_registers_i/_2496_ ;
 wire \cs_registers_i/_2497_ ;
 wire \cs_registers_i/_2498_ ;
 wire \cs_registers_i/_2499_ ;
 wire \cs_registers_i/_2500_ ;
 wire \cs_registers_i/_2501_ ;
 wire \cs_registers_i/_2502_ ;
 wire \cs_registers_i/_2503_ ;
 wire \cs_registers_i/_2504_ ;
 wire \cs_registers_i/_2505_ ;
 wire \cs_registers_i/_2506_ ;
 wire \cs_registers_i/_2507_ ;
 wire \cs_registers_i/_2508_ ;
 wire \cs_registers_i/_2509_ ;
 wire \cs_registers_i/_2510_ ;
 wire \cs_registers_i/_2511_ ;
 wire \cs_registers_i/_2512_ ;
 wire \cs_registers_i/_2513_ ;
 wire \cs_registers_i/_2514_ ;
 wire \cs_registers_i/_2515_ ;
 wire \cs_registers_i/_2516_ ;
 wire \cs_registers_i/_2517_ ;
 wire \cs_registers_i/_2518_ ;
 wire \cs_registers_i/_2519_ ;
 wire \cs_registers_i/_2520_ ;
 wire \cs_registers_i/_2521_ ;
 wire \cs_registers_i/_2522_ ;
 wire \cs_registers_i/_2523_ ;
 wire \cs_registers_i/_2524_ ;
 wire \cs_registers_i/_2525_ ;
 wire \cs_registers_i/_2526_ ;
 wire \cs_registers_i/_2527_ ;
 wire \cs_registers_i/_2528_ ;
 wire \cs_registers_i/_2529_ ;
 wire \cs_registers_i/_2530_ ;
 wire \cs_registers_i/_2531_ ;
 wire \cs_registers_i/_2532_ ;
 wire \cs_registers_i/_2533_ ;
 wire \cs_registers_i/_2534_ ;
 wire \cs_registers_i/_2535_ ;
 wire \cs_registers_i/_2536_ ;
 wire \cs_registers_i/_2537_ ;
 wire \cs_registers_i/_2538_ ;
 wire \cs_registers_i/_2539_ ;
 wire \cs_registers_i/_2540_ ;
 wire \cs_registers_i/_2541_ ;
 wire \cs_registers_i/_2542_ ;
 wire \cs_registers_i/_2543_ ;
 wire \cs_registers_i/_2544_ ;
 wire \cs_registers_i/_2545_ ;
 wire \cs_registers_i/_2546_ ;
 wire \cs_registers_i/_2547_ ;
 wire \cs_registers_i/_2548_ ;
 wire \cs_registers_i/_2549_ ;
 wire \cs_registers_i/_2550_ ;
 wire \cs_registers_i/_2551_ ;
 wire \cs_registers_i/_2552_ ;
 wire \cs_registers_i/_2553_ ;
 wire \cs_registers_i/_2554_ ;
 wire \cs_registers_i/_2555_ ;
 wire \cs_registers_i/_2556_ ;
 wire \cs_registers_i/_2557_ ;
 wire \cs_registers_i/_2558_ ;
 wire \cs_registers_i/_2559_ ;
 wire \cs_registers_i/_2560_ ;
 wire \cs_registers_i/_2561_ ;
 wire \cs_registers_i/_2562_ ;
 wire \cs_registers_i/_2563_ ;
 wire \cs_registers_i/_2564_ ;
 wire \cs_registers_i/_2565_ ;
 wire \cs_registers_i/_2566_ ;
 wire \cs_registers_i/_2567_ ;
 wire \cs_registers_i/_2568_ ;
 wire \cs_registers_i/_2569_ ;
 wire \cs_registers_i/_2570_ ;
 wire \cs_registers_i/_2571_ ;
 wire \cs_registers_i/_2572_ ;
 wire \cs_registers_i/_2573_ ;
 wire \cs_registers_i/_2574_ ;
 wire \cs_registers_i/_2575_ ;
 wire \cs_registers_i/_2576_ ;
 wire \cs_registers_i/_2577_ ;
 wire \cs_registers_i/_2578_ ;
 wire \cs_registers_i/_2579_ ;
 wire \cs_registers_i/_2580_ ;
 wire \cs_registers_i/_2581_ ;
 wire \cs_registers_i/_2582_ ;
 wire \cs_registers_i/_2583_ ;
 wire \cs_registers_i/_2584_ ;
 wire \cs_registers_i/_2585_ ;
 wire \cs_registers_i/_2586_ ;
 wire \cs_registers_i/_2587_ ;
 wire \cs_registers_i/_2588_ ;
 wire \cs_registers_i/_2589_ ;
 wire \cs_registers_i/_2590_ ;
 wire \cs_registers_i/_2591_ ;
 wire \cs_registers_i/_2592_ ;
 wire \cs_registers_i/_2593_ ;
 wire \cs_registers_i/_2594_ ;
 wire \cs_registers_i/_2595_ ;
 wire \cs_registers_i/_2596_ ;
 wire \cs_registers_i/_2597_ ;
 wire \cs_registers_i/_2598_ ;
 wire \cs_registers_i/_2599_ ;
 wire \cs_registers_i/_2600_ ;
 wire \cs_registers_i/_2601_ ;
 wire \cs_registers_i/_2602_ ;
 wire \cs_registers_i/_2603_ ;
 wire \cs_registers_i/_2604_ ;
 wire \cs_registers_i/_2605_ ;
 wire \cs_registers_i/_2606_ ;
 wire \cs_registers_i/_2607_ ;
 wire \cs_registers_i/_2608_ ;
 wire \cs_registers_i/_2609_ ;
 wire \cs_registers_i/_2610_ ;
 wire \cs_registers_i/_2611_ ;
 wire \cs_registers_i/_2612_ ;
 wire \cs_registers_i/_2613_ ;
 wire \cs_registers_i/_2614_ ;
 wire \cs_registers_i/_2615_ ;
 wire \cs_registers_i/_2616_ ;
 wire \cs_registers_i/_2617_ ;
 wire \cs_registers_i/_2618_ ;
 wire \cs_registers_i/_2619_ ;
 wire \cs_registers_i/_2620_ ;
 wire \cs_registers_i/_2621_ ;
 wire \cs_registers_i/_2622_ ;
 wire \cs_registers_i/_2623_ ;
 wire \cs_registers_i/_2624_ ;
 wire \cs_registers_i/_2625_ ;
 wire \cs_registers_i/_2626_ ;
 wire \cs_registers_i/_2627_ ;
 wire \cs_registers_i/_2628_ ;
 wire \cs_registers_i/_2629_ ;
 wire \cs_registers_i/_2630_ ;
 wire \cs_registers_i/_2631_ ;
 wire \cs_registers_i/_2632_ ;
 wire \cs_registers_i/_2633_ ;
 wire \cs_registers_i/_2634_ ;
 wire \cs_registers_i/_2635_ ;
 wire \cs_registers_i/_2636_ ;
 wire \cs_registers_i/_2637_ ;
 wire \cs_registers_i/_2638_ ;
 wire \cs_registers_i/_2639_ ;
 wire \cs_registers_i/_2640_ ;
 wire \cs_registers_i/_2641_ ;
 wire \cs_registers_i/_2642_ ;
 wire \cs_registers_i/_2643_ ;
 wire \cs_registers_i/_2644_ ;
 wire \cs_registers_i/_2645_ ;
 wire \cs_registers_i/_2646_ ;
 wire \cs_registers_i/_2647_ ;
 wire \cs_registers_i/_2648_ ;
 wire \cs_registers_i/_2649_ ;
 wire \cs_registers_i/_2650_ ;
 wire \cs_registers_i/_2651_ ;
 wire \cs_registers_i/_2652_ ;
 wire \cs_registers_i/_2653_ ;
 wire \cs_registers_i/_2654_ ;
 wire \cs_registers_i/_2655_ ;
 wire \cs_registers_i/_2656_ ;
 wire \cs_registers_i/_2657_ ;
 wire \cs_registers_i/_2658_ ;
 wire \cs_registers_i/_2659_ ;
 wire \cs_registers_i/_2660_ ;
 wire \cs_registers_i/_2661_ ;
 wire \cs_registers_i/_2662_ ;
 wire \cs_registers_i/_2663_ ;
 wire \cs_registers_i/_2664_ ;
 wire \cs_registers_i/_2665_ ;
 wire \cs_registers_i/_2666_ ;
 wire \cs_registers_i/_2667_ ;
 wire \cs_registers_i/_2668_ ;
 wire \cs_registers_i/_2669_ ;
 wire \cs_registers_i/_2670_ ;
 wire \cs_registers_i/_2671_ ;
 wire \cs_registers_i/_2672_ ;
 wire \cs_registers_i/_2673_ ;
 wire \cs_registers_i/_2674_ ;
 wire \cs_registers_i/_2675_ ;
 wire \cs_registers_i/_2676_ ;
 wire \cs_registers_i/_2677_ ;
 wire \cs_registers_i/_2678_ ;
 wire \cs_registers_i/_2679_ ;
 wire \cs_registers_i/_2680_ ;
 wire \cs_registers_i/_2681_ ;
 wire \cs_registers_i/_2682_ ;
 wire \cs_registers_i/_2683_ ;
 wire \cs_registers_i/_2684_ ;
 wire \cs_registers_i/_2685_ ;
 wire \cs_registers_i/_2686_ ;
 wire \cs_registers_i/_2687_ ;
 wire \cs_registers_i/_2688_ ;
 wire \cs_registers_i/_2689_ ;
 wire \cs_registers_i/_2690_ ;
 wire \cs_registers_i/_2691_ ;
 wire \cs_registers_i/_2692_ ;
 wire \cs_registers_i/_2693_ ;
 wire \cs_registers_i/_2694_ ;
 wire \cs_registers_i/_2695_ ;
 wire \cs_registers_i/_2696_ ;
 wire \cs_registers_i/_2697_ ;
 wire \cs_registers_i/_2698_ ;
 wire \cs_registers_i/_2699_ ;
 wire \cs_registers_i/_2700_ ;
 wire \cs_registers_i/_2701_ ;
 wire \cs_registers_i/_2702_ ;
 wire \cs_registers_i/_2703_ ;
 wire \cs_registers_i/_2704_ ;
 wire \cs_registers_i/_2705_ ;
 wire \cs_registers_i/_2706_ ;
 wire \cs_registers_i/_2707_ ;
 wire \cs_registers_i/_2708_ ;
 wire \cs_registers_i/_2709_ ;
 wire \cs_registers_i/_2710_ ;
 wire \cs_registers_i/_2711_ ;
 wire \cs_registers_i/_2712_ ;
 wire \cs_registers_i/_2713_ ;
 wire \cs_registers_i/_2714_ ;
 wire \cs_registers_i/_2715_ ;
 wire \cs_registers_i/_2716_ ;
 wire \cs_registers_i/_2717_ ;
 wire \cs_registers_i/_2718_ ;
 wire \cs_registers_i/_2719_ ;
 wire \cs_registers_i/_2720_ ;
 wire \cs_registers_i/_2721_ ;
 wire \cs_registers_i/_2722_ ;
 wire \cs_registers_i/_2723_ ;
 wire \cs_registers_i/_2724_ ;
 wire \cs_registers_i/_2725_ ;
 wire \cs_registers_i/_2726_ ;
 wire \cs_registers_i/_2727_ ;
 wire \cs_registers_i/_2728_ ;
 wire \cs_registers_i/_2729_ ;
 wire \cs_registers_i/_2730_ ;
 wire \cs_registers_i/_2731_ ;
 wire \cs_registers_i/_2732_ ;
 wire \cs_registers_i/_2733_ ;
 wire \cs_registers_i/_2734_ ;
 wire \cs_registers_i/_2735_ ;
 wire \cs_registers_i/_2736_ ;
 wire \cs_registers_i/_2737_ ;
 wire \cs_registers_i/_2738_ ;
 wire \cs_registers_i/_2739_ ;
 wire \cs_registers_i/_2740_ ;
 wire \cs_registers_i/_2741_ ;
 wire \cs_registers_i/_2742_ ;
 wire \cs_registers_i/_2743_ ;
 wire \cs_registers_i/_2744_ ;
 wire \cs_registers_i/_2745_ ;
 wire \cs_registers_i/_2746_ ;
 wire \cs_registers_i/_2747_ ;
 wire \cs_registers_i/_2748_ ;
 wire \cs_registers_i/_2749_ ;
 wire \cs_registers_i/_2750_ ;
 wire \cs_registers_i/_2751_ ;
 wire \cs_registers_i/_2752_ ;
 wire \cs_registers_i/_2753_ ;
 wire \cs_registers_i/_2754_ ;
 wire \cs_registers_i/_2755_ ;
 wire \cs_registers_i/_2756_ ;
 wire \cs_registers_i/_2757_ ;
 wire \cs_registers_i/_2758_ ;
 wire \cs_registers_i/_2759_ ;
 wire \cs_registers_i/_2760_ ;
 wire \cs_registers_i/_2761_ ;
 wire \cs_registers_i/_2762_ ;
 wire \cs_registers_i/_2763_ ;
 wire \cs_registers_i/_2764_ ;
 wire \cs_registers_i/_2765_ ;
 wire \cs_registers_i/_2766_ ;
 wire \cs_registers_i/_2767_ ;
 wire \cs_registers_i/_2768_ ;
 wire \cs_registers_i/_2769_ ;
 wire \cs_registers_i/_2770_ ;
 wire \cs_registers_i/_2771_ ;
 wire \cs_registers_i/_2772_ ;
 wire \cs_registers_i/_2773_ ;
 wire \cs_registers_i/_2774_ ;
 wire \cs_registers_i/_2775_ ;
 wire \cs_registers_i/_2776_ ;
 wire \cs_registers_i/_2777_ ;
 wire \cs_registers_i/_2778_ ;
 wire \cs_registers_i/_2779_ ;
 wire \cs_registers_i/_2780_ ;
 wire \cs_registers_i/_2781_ ;
 wire \cs_registers_i/_2782_ ;
 wire \cs_registers_i/_2783_ ;
 wire \cs_registers_i/_2784_ ;
 wire \cs_registers_i/_2785_ ;
 wire \cs_registers_i/_2786_ ;
 wire \cs_registers_i/_2787_ ;
 wire \cs_registers_i/_2788_ ;
 wire \cs_registers_i/_2789_ ;
 wire \cs_registers_i/_2790_ ;
 wire \cs_registers_i/_2791_ ;
 wire \cs_registers_i/_2792_ ;
 wire \cs_registers_i/_2793_ ;
 wire \cs_registers_i/_2794_ ;
 wire \cs_registers_i/_2795_ ;
 wire \cs_registers_i/_2796_ ;
 wire \cs_registers_i/_2797_ ;
 wire \cs_registers_i/_2798_ ;
 wire \cs_registers_i/_2799_ ;
 wire \cs_registers_i/_2800_ ;
 wire \cs_registers_i/_2801_ ;
 wire \cs_registers_i/_2802_ ;
 wire \cs_registers_i/_2803_ ;
 wire \cs_registers_i/_2804_ ;
 wire \cs_registers_i/_2805_ ;
 wire \cs_registers_i/_2806_ ;
 wire \cs_registers_i/_2807_ ;
 wire \cs_registers_i/_2808_ ;
 wire \cs_registers_i/_2809_ ;
 wire \cs_registers_i/_2810_ ;
 wire \cs_registers_i/_2811_ ;
 wire \cs_registers_i/_2812_ ;
 wire \cs_registers_i/_2813_ ;
 wire \cs_registers_i/_2814_ ;
 wire \cs_registers_i/_2815_ ;
 wire \cs_registers_i/_2816_ ;
 wire \cs_registers_i/_2817_ ;
 wire \cs_registers_i/_2818_ ;
 wire \cs_registers_i/_2819_ ;
 wire \cs_registers_i/_2820_ ;
 wire \cs_registers_i/_2821_ ;
 wire \cs_registers_i/_2822_ ;
 wire \cs_registers_i/_2823_ ;
 wire \cs_registers_i/_2824_ ;
 wire \cs_registers_i/_2825_ ;
 wire \cs_registers_i/_2826_ ;
 wire \cs_registers_i/_2827_ ;
 wire \cs_registers_i/_2828_ ;
 wire \cs_registers_i/_2829_ ;
 wire \cs_registers_i/_2830_ ;
 wire \cs_registers_i/_2831_ ;
 wire \cs_registers_i/_2832_ ;
 wire \cs_registers_i/_2833_ ;
 wire \cs_registers_i/_2834_ ;
 wire \cs_registers_i/_2835_ ;
 wire \cs_registers_i/_2836_ ;
 wire \cs_registers_i/_2837_ ;
 wire \cs_registers_i/_2838_ ;
 wire \cs_registers_i/_2839_ ;
 wire \cs_registers_i/_2840_ ;
 wire \cs_registers_i/_2841_ ;
 wire \cs_registers_i/_2842_ ;
 wire \cs_registers_i/_2843_ ;
 wire \cs_registers_i/_2844_ ;
 wire \cs_registers_i/_2845_ ;
 wire \cs_registers_i/_2846_ ;
 wire \cs_registers_i/_2847_ ;
 wire \cs_registers_i/_2848_ ;
 wire \cs_registers_i/_2849_ ;
 wire \cs_registers_i/_2850_ ;
 wire \cs_registers_i/_2851_ ;
 wire \cs_registers_i/_2852_ ;
 wire \cs_registers_i/_2853_ ;
 wire \cs_registers_i/_2854_ ;
 wire \cs_registers_i/_2855_ ;
 wire \cs_registers_i/_2856_ ;
 wire \cs_registers_i/_2857_ ;
 wire \cs_registers_i/_2858_ ;
 wire \cs_registers_i/_2859_ ;
 wire \cs_registers_i/_2860_ ;
 wire \cs_registers_i/_2861_ ;
 wire \cs_registers_i/_2862_ ;
 wire \cs_registers_i/_2863_ ;
 wire \cs_registers_i/_2864_ ;
 wire \cs_registers_i/_2865_ ;
 wire \cs_registers_i/_2866_ ;
 wire \cs_registers_i/_2867_ ;
 wire \cs_registers_i/_2868_ ;
 wire \cs_registers_i/_2869_ ;
 wire \cs_registers_i/_2870_ ;
 wire \cs_registers_i/_2871_ ;
 wire \cs_registers_i/_2872_ ;
 wire \cs_registers_i/_2873_ ;
 wire \cs_registers_i/_2874_ ;
 wire \cs_registers_i/_2875_ ;
 wire \cs_registers_i/_2876_ ;
 wire \cs_registers_i/_2877_ ;
 wire \cs_registers_i/_2878_ ;
 wire \cs_registers_i/_2879_ ;
 wire \cs_registers_i/_2880_ ;
 wire \cs_registers_i/_2881_ ;
 wire \cs_registers_i/_2882_ ;
 wire \cs_registers_i/_2883_ ;
 wire \cs_registers_i/_2884_ ;
 wire \cs_registers_i/_2885_ ;
 wire \cs_registers_i/_2886_ ;
 wire \cs_registers_i/_2887_ ;
 wire \cs_registers_i/_2888_ ;
 wire \cs_registers_i/_2889_ ;
 wire \cs_registers_i/_2890_ ;
 wire \cs_registers_i/_2891_ ;
 wire \cs_registers_i/_2892_ ;
 wire \cs_registers_i/_2893_ ;
 wire \cs_registers_i/_2894_ ;
 wire \cs_registers_i/_2895_ ;
 wire \cs_registers_i/_2896_ ;
 wire \cs_registers_i/_2897_ ;
 wire \cs_registers_i/_2898_ ;
 wire \cs_registers_i/_2899_ ;
 wire \cs_registers_i/_2900_ ;
 wire \cs_registers_i/_2901_ ;
 wire \cs_registers_i/_2902_ ;
 wire \cs_registers_i/_2903_ ;
 wire \cs_registers_i/_2904_ ;
 wire \cs_registers_i/_2905_ ;
 wire \cs_registers_i/_2906_ ;
 wire \cs_registers_i/_2907_ ;
 wire \cs_registers_i/_2908_ ;
 wire \cs_registers_i/_2909_ ;
 wire \cs_registers_i/_2910_ ;
 wire \cs_registers_i/_2911_ ;
 wire \cs_registers_i/_2912_ ;
 wire \cs_registers_i/_2913_ ;
 wire \cs_registers_i/_2914_ ;
 wire \cs_registers_i/_2915_ ;
 wire \cs_registers_i/_2916_ ;
 wire \cs_registers_i/_2917_ ;
 wire \cs_registers_i/_2918_ ;
 wire \cs_registers_i/_2919_ ;
 wire \cs_registers_i/_2920_ ;
 wire \cs_registers_i/_2921_ ;
 wire \cs_registers_i/dcsr_q_0_ ;
 wire \cs_registers_i/dcsr_q_10_ ;
 wire \cs_registers_i/dcsr_q_11_ ;
 wire \cs_registers_i/dcsr_q_13_ ;
 wire \cs_registers_i/dcsr_q_14_ ;
 wire \cs_registers_i/dcsr_q_16_ ;
 wire \cs_registers_i/dcsr_q_17_ ;
 wire \cs_registers_i/dcsr_q_18_ ;
 wire \cs_registers_i/dcsr_q_19_ ;
 wire \cs_registers_i/dcsr_q_1_ ;
 wire \cs_registers_i/dcsr_q_20_ ;
 wire \cs_registers_i/dcsr_q_21_ ;
 wire \cs_registers_i/dcsr_q_22_ ;
 wire \cs_registers_i/dcsr_q_23_ ;
 wire \cs_registers_i/dcsr_q_24_ ;
 wire \cs_registers_i/dcsr_q_25_ ;
 wire \cs_registers_i/dcsr_q_26_ ;
 wire \cs_registers_i/dcsr_q_27_ ;
 wire \cs_registers_i/dcsr_q_28_ ;
 wire \cs_registers_i/dcsr_q_29_ ;
 wire \cs_registers_i/dcsr_q_30_ ;
 wire \cs_registers_i/dcsr_q_31_ ;
 wire \cs_registers_i/dcsr_q_3_ ;
 wire \cs_registers_i/dcsr_q_4_ ;
 wire \cs_registers_i/dcsr_q_5_ ;
 wire \cs_registers_i/dcsr_q_6_ ;
 wire \cs_registers_i/dcsr_q_7_ ;
 wire \cs_registers_i/dcsr_q_8_ ;
 wire \cs_registers_i/dcsr_q_9_ ;
 wire \cs_registers_i/dscratch0_q_0_ ;
 wire \cs_registers_i/dscratch0_q_10_ ;
 wire \cs_registers_i/dscratch0_q_11_ ;
 wire \cs_registers_i/dscratch0_q_12_ ;
 wire \cs_registers_i/dscratch0_q_13_ ;
 wire \cs_registers_i/dscratch0_q_14_ ;
 wire \cs_registers_i/dscratch0_q_15_ ;
 wire \cs_registers_i/dscratch0_q_16_ ;
 wire \cs_registers_i/dscratch0_q_17_ ;
 wire \cs_registers_i/dscratch0_q_18_ ;
 wire \cs_registers_i/dscratch0_q_19_ ;
 wire \cs_registers_i/dscratch0_q_1_ ;
 wire \cs_registers_i/dscratch0_q_20_ ;
 wire \cs_registers_i/dscratch0_q_21_ ;
 wire \cs_registers_i/dscratch0_q_22_ ;
 wire \cs_registers_i/dscratch0_q_23_ ;
 wire \cs_registers_i/dscratch0_q_24_ ;
 wire \cs_registers_i/dscratch0_q_25_ ;
 wire \cs_registers_i/dscratch0_q_26_ ;
 wire \cs_registers_i/dscratch0_q_27_ ;
 wire \cs_registers_i/dscratch0_q_28_ ;
 wire \cs_registers_i/dscratch0_q_29_ ;
 wire \cs_registers_i/dscratch0_q_2_ ;
 wire \cs_registers_i/dscratch0_q_30_ ;
 wire \cs_registers_i/dscratch0_q_31_ ;
 wire \cs_registers_i/dscratch0_q_3_ ;
 wire \cs_registers_i/dscratch0_q_4_ ;
 wire \cs_registers_i/dscratch0_q_5_ ;
 wire \cs_registers_i/dscratch0_q_6_ ;
 wire \cs_registers_i/dscratch0_q_7_ ;
 wire \cs_registers_i/dscratch0_q_8_ ;
 wire \cs_registers_i/dscratch0_q_9_ ;
 wire \cs_registers_i/dscratch1_q_0_ ;
 wire \cs_registers_i/dscratch1_q_10_ ;
 wire \cs_registers_i/dscratch1_q_11_ ;
 wire \cs_registers_i/dscratch1_q_12_ ;
 wire \cs_registers_i/dscratch1_q_13_ ;
 wire \cs_registers_i/dscratch1_q_14_ ;
 wire \cs_registers_i/dscratch1_q_15_ ;
 wire \cs_registers_i/dscratch1_q_16_ ;
 wire \cs_registers_i/dscratch1_q_17_ ;
 wire \cs_registers_i/dscratch1_q_18_ ;
 wire \cs_registers_i/dscratch1_q_19_ ;
 wire \cs_registers_i/dscratch1_q_1_ ;
 wire \cs_registers_i/dscratch1_q_20_ ;
 wire \cs_registers_i/dscratch1_q_21_ ;
 wire \cs_registers_i/dscratch1_q_22_ ;
 wire \cs_registers_i/dscratch1_q_23_ ;
 wire \cs_registers_i/dscratch1_q_24_ ;
 wire \cs_registers_i/dscratch1_q_25_ ;
 wire \cs_registers_i/dscratch1_q_26_ ;
 wire \cs_registers_i/dscratch1_q_27_ ;
 wire \cs_registers_i/dscratch1_q_28_ ;
 wire \cs_registers_i/dscratch1_q_29_ ;
 wire \cs_registers_i/dscratch1_q_2_ ;
 wire \cs_registers_i/dscratch1_q_30_ ;
 wire \cs_registers_i/dscratch1_q_31_ ;
 wire \cs_registers_i/dscratch1_q_3_ ;
 wire \cs_registers_i/dscratch1_q_4_ ;
 wire \cs_registers_i/dscratch1_q_5_ ;
 wire \cs_registers_i/dscratch1_q_6_ ;
 wire \cs_registers_i/dscratch1_q_7_ ;
 wire \cs_registers_i/dscratch1_q_8_ ;
 wire \cs_registers_i/dscratch1_q_9_ ;
 wire \cs_registers_i/mcause_q_0_ ;
 wire \cs_registers_i/mcause_q_1_ ;
 wire \cs_registers_i/mcause_q_2_ ;
 wire \cs_registers_i/mcause_q_3_ ;
 wire \cs_registers_i/mcause_q_4_ ;
 wire \cs_registers_i/mcause_q_5_ ;
 wire \cs_registers_i/mcause_q_6_ ;
 wire \cs_registers_i/mcountinhibit_0_ ;
 wire \cs_registers_i/mcountinhibit_2_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_inc_i ;
 wire \cs_registers_i/mcycle_counter_i.counter_upd_0_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_0_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_10_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_11_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_12_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_13_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_14_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_15_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_16_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_17_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_18_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_19_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_1_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_20_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_21_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_22_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_23_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_24_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_25_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_26_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_27_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_28_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_29_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_2_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_30_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_31_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_32_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_33_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_34_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_35_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_36_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_37_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_38_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_39_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_3_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_40_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_41_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_42_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_43_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_44_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_45_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_46_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_47_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_48_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_49_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_4_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_50_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_51_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_52_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_53_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_54_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_55_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_56_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_57_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_58_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_59_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_5_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_60_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_61_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_62_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_63_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_6_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_7_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_8_ ;
 wire \cs_registers_i/mcycle_counter_i.counter_val_o_9_ ;
 wire \cs_registers_i/mhpmcounter_1856_ ;
 wire \cs_registers_i/mhpmcounter_1857_ ;
 wire \cs_registers_i/mhpmcounter_1858_ ;
 wire \cs_registers_i/mhpmcounter_1859_ ;
 wire \cs_registers_i/mhpmcounter_1860_ ;
 wire \cs_registers_i/mhpmcounter_1861_ ;
 wire \cs_registers_i/mhpmcounter_1862_ ;
 wire \cs_registers_i/mhpmcounter_1863_ ;
 wire \cs_registers_i/mhpmcounter_1864_ ;
 wire \cs_registers_i/mhpmcounter_1865_ ;
 wire \cs_registers_i/mhpmcounter_1866_ ;
 wire \cs_registers_i/mhpmcounter_1867_ ;
 wire \cs_registers_i/mhpmcounter_1868_ ;
 wire \cs_registers_i/mhpmcounter_1869_ ;
 wire \cs_registers_i/mhpmcounter_1870_ ;
 wire \cs_registers_i/mhpmcounter_1871_ ;
 wire \cs_registers_i/mhpmcounter_1872_ ;
 wire \cs_registers_i/mhpmcounter_1873_ ;
 wire \cs_registers_i/mhpmcounter_1874_ ;
 wire \cs_registers_i/mhpmcounter_1875_ ;
 wire \cs_registers_i/mhpmcounter_1876_ ;
 wire \cs_registers_i/mhpmcounter_1877_ ;
 wire \cs_registers_i/mhpmcounter_1878_ ;
 wire \cs_registers_i/mhpmcounter_1879_ ;
 wire \cs_registers_i/mhpmcounter_1880_ ;
 wire \cs_registers_i/mhpmcounter_1881_ ;
 wire \cs_registers_i/mhpmcounter_1882_ ;
 wire \cs_registers_i/mhpmcounter_1883_ ;
 wire \cs_registers_i/mhpmcounter_1884_ ;
 wire \cs_registers_i/mhpmcounter_1885_ ;
 wire \cs_registers_i/mhpmcounter_1886_ ;
 wire \cs_registers_i/mhpmcounter_1887_ ;
 wire \cs_registers_i/mhpmcounter_1888_ ;
 wire \cs_registers_i/mhpmcounter_1889_ ;
 wire \cs_registers_i/mhpmcounter_1890_ ;
 wire \cs_registers_i/mhpmcounter_1891_ ;
 wire \cs_registers_i/mhpmcounter_1892_ ;
 wire \cs_registers_i/mhpmcounter_1893_ ;
 wire \cs_registers_i/mhpmcounter_1894_ ;
 wire \cs_registers_i/mhpmcounter_1895_ ;
 wire \cs_registers_i/mhpmcounter_1896_ ;
 wire \cs_registers_i/mhpmcounter_1897_ ;
 wire \cs_registers_i/mhpmcounter_1898_ ;
 wire \cs_registers_i/mhpmcounter_1899_ ;
 wire \cs_registers_i/mhpmcounter_1900_ ;
 wire \cs_registers_i/mhpmcounter_1901_ ;
 wire \cs_registers_i/mhpmcounter_1902_ ;
 wire \cs_registers_i/mhpmcounter_1903_ ;
 wire \cs_registers_i/mhpmcounter_1904_ ;
 wire \cs_registers_i/mhpmcounter_1905_ ;
 wire \cs_registers_i/mhpmcounter_1906_ ;
 wire \cs_registers_i/mhpmcounter_1907_ ;
 wire \cs_registers_i/mhpmcounter_1908_ ;
 wire \cs_registers_i/mhpmcounter_1909_ ;
 wire \cs_registers_i/mhpmcounter_1910_ ;
 wire \cs_registers_i/mhpmcounter_1911_ ;
 wire \cs_registers_i/mhpmcounter_1912_ ;
 wire \cs_registers_i/mhpmcounter_1913_ ;
 wire \cs_registers_i/mhpmcounter_1914_ ;
 wire \cs_registers_i/mhpmcounter_1915_ ;
 wire \cs_registers_i/mhpmcounter_1916_ ;
 wire \cs_registers_i/mhpmcounter_1917_ ;
 wire \cs_registers_i/mhpmcounter_1918_ ;
 wire \cs_registers_i/mhpmcounter_1919_ ;
 wire \cs_registers_i/mie_q_0_ ;
 wire \cs_registers_i/mie_q_10_ ;
 wire \cs_registers_i/mie_q_11_ ;
 wire \cs_registers_i/mie_q_12_ ;
 wire \cs_registers_i/mie_q_13_ ;
 wire \cs_registers_i/mie_q_14_ ;
 wire \cs_registers_i/mie_q_15_ ;
 wire \cs_registers_i/mie_q_16_ ;
 wire \cs_registers_i/mie_q_17_ ;
 wire \cs_registers_i/mie_q_18_ ;
 wire \cs_registers_i/mie_q_1_ ;
 wire \cs_registers_i/mie_q_2_ ;
 wire \cs_registers_i/mie_q_3_ ;
 wire \cs_registers_i/mie_q_4_ ;
 wire \cs_registers_i/mie_q_5_ ;
 wire \cs_registers_i/mie_q_6_ ;
 wire \cs_registers_i/mie_q_7_ ;
 wire \cs_registers_i/mie_q_8_ ;
 wire \cs_registers_i/mie_q_9_ ;
 wire \cs_registers_i/minstret_counter_i.counter_inc_i_$_AND__Y_B ;
 wire \cs_registers_i/minstret_counter_i.counter_val_upd_o_0_ ;
 wire \cs_registers_i/mscratch_q_0_ ;
 wire \cs_registers_i/mscratch_q_10_ ;
 wire \cs_registers_i/mscratch_q_11_ ;
 wire \cs_registers_i/mscratch_q_12_ ;
 wire \cs_registers_i/mscratch_q_13_ ;
 wire \cs_registers_i/mscratch_q_14_ ;
 wire \cs_registers_i/mscratch_q_15_ ;
 wire \cs_registers_i/mscratch_q_16_ ;
 wire \cs_registers_i/mscratch_q_17_ ;
 wire \cs_registers_i/mscratch_q_18_ ;
 wire \cs_registers_i/mscratch_q_19_ ;
 wire \cs_registers_i/mscratch_q_1_ ;
 wire \cs_registers_i/mscratch_q_20_ ;
 wire \cs_registers_i/mscratch_q_21_ ;
 wire \cs_registers_i/mscratch_q_22_ ;
 wire \cs_registers_i/mscratch_q_23_ ;
 wire \cs_registers_i/mscratch_q_24_ ;
 wire \cs_registers_i/mscratch_q_25_ ;
 wire \cs_registers_i/mscratch_q_26_ ;
 wire \cs_registers_i/mscratch_q_27_ ;
 wire \cs_registers_i/mscratch_q_28_ ;
 wire \cs_registers_i/mscratch_q_29_ ;
 wire \cs_registers_i/mscratch_q_2_ ;
 wire \cs_registers_i/mscratch_q_30_ ;
 wire \cs_registers_i/mscratch_q_31_ ;
 wire \cs_registers_i/mscratch_q_3_ ;
 wire \cs_registers_i/mscratch_q_4_ ;
 wire \cs_registers_i/mscratch_q_5_ ;
 wire \cs_registers_i/mscratch_q_6_ ;
 wire \cs_registers_i/mscratch_q_7_ ;
 wire \cs_registers_i/mscratch_q_8_ ;
 wire \cs_registers_i/mscratch_q_9_ ;
 wire \cs_registers_i/mstack_cause_q_0_ ;
 wire \cs_registers_i/mstack_cause_q_1_ ;
 wire \cs_registers_i/mstack_cause_q_2_ ;
 wire \cs_registers_i/mstack_cause_q_3_ ;
 wire \cs_registers_i/mstack_cause_q_4_ ;
 wire \cs_registers_i/mstack_cause_q_5_ ;
 wire \cs_registers_i/mstack_cause_q_6_ ;
 wire \cs_registers_i/mstack_epc_q_0_ ;
 wire \cs_registers_i/mstack_epc_q_10_ ;
 wire \cs_registers_i/mstack_epc_q_11_ ;
 wire \cs_registers_i/mstack_epc_q_12_ ;
 wire \cs_registers_i/mstack_epc_q_13_ ;
 wire \cs_registers_i/mstack_epc_q_14_ ;
 wire \cs_registers_i/mstack_epc_q_15_ ;
 wire \cs_registers_i/mstack_epc_q_16_ ;
 wire \cs_registers_i/mstack_epc_q_17_ ;
 wire \cs_registers_i/mstack_epc_q_18_ ;
 wire \cs_registers_i/mstack_epc_q_19_ ;
 wire \cs_registers_i/mstack_epc_q_1_ ;
 wire \cs_registers_i/mstack_epc_q_20_ ;
 wire \cs_registers_i/mstack_epc_q_21_ ;
 wire \cs_registers_i/mstack_epc_q_22_ ;
 wire \cs_registers_i/mstack_epc_q_23_ ;
 wire \cs_registers_i/mstack_epc_q_24_ ;
 wire \cs_registers_i/mstack_epc_q_25_ ;
 wire \cs_registers_i/mstack_epc_q_26_ ;
 wire \cs_registers_i/mstack_epc_q_27_ ;
 wire \cs_registers_i/mstack_epc_q_28_ ;
 wire \cs_registers_i/mstack_epc_q_29_ ;
 wire \cs_registers_i/mstack_epc_q_2_ ;
 wire \cs_registers_i/mstack_epc_q_30_ ;
 wire \cs_registers_i/mstack_epc_q_31_ ;
 wire \cs_registers_i/mstack_epc_q_3_ ;
 wire \cs_registers_i/mstack_epc_q_4_ ;
 wire \cs_registers_i/mstack_epc_q_5_ ;
 wire \cs_registers_i/mstack_epc_q_6_ ;
 wire \cs_registers_i/mstack_epc_q_7_ ;
 wire \cs_registers_i/mstack_epc_q_8_ ;
 wire \cs_registers_i/mstack_epc_q_9_ ;
 wire \cs_registers_i/mstack_q_0_ ;
 wire \cs_registers_i/mstack_q_1_ ;
 wire \cs_registers_i/mstack_q_2_ ;
 wire \cs_registers_i/mstatus_q_1_ ;
 wire \cs_registers_i/mstatus_q_2_ ;
 wire \cs_registers_i/mstatus_q_3_ ;
 wire \cs_registers_i/mstatus_q_4_ ;
 wire \cs_registers_i/mtval_q_0_ ;
 wire \cs_registers_i/mtval_q_10_ ;
 wire \cs_registers_i/mtval_q_11_ ;
 wire \cs_registers_i/mtval_q_12_ ;
 wire \cs_registers_i/mtval_q_13_ ;
 wire \cs_registers_i/mtval_q_14_ ;
 wire \cs_registers_i/mtval_q_15_ ;
 wire \cs_registers_i/mtval_q_16_ ;
 wire \cs_registers_i/mtval_q_17_ ;
 wire \cs_registers_i/mtval_q_18_ ;
 wire \cs_registers_i/mtval_q_19_ ;
 wire \cs_registers_i/mtval_q_1_ ;
 wire \cs_registers_i/mtval_q_20_ ;
 wire \cs_registers_i/mtval_q_21_ ;
 wire \cs_registers_i/mtval_q_22_ ;
 wire \cs_registers_i/mtval_q_23_ ;
 wire \cs_registers_i/mtval_q_24_ ;
 wire \cs_registers_i/mtval_q_25_ ;
 wire \cs_registers_i/mtval_q_26_ ;
 wire \cs_registers_i/mtval_q_27_ ;
 wire \cs_registers_i/mtval_q_28_ ;
 wire \cs_registers_i/mtval_q_29_ ;
 wire \cs_registers_i/mtval_q_2_ ;
 wire \cs_registers_i/mtval_q_30_ ;
 wire \cs_registers_i/mtval_q_31_ ;
 wire \cs_registers_i/mtval_q_3_ ;
 wire \cs_registers_i/mtval_q_4_ ;
 wire \cs_registers_i/mtval_q_5_ ;
 wire \cs_registers_i/mtval_q_6_ ;
 wire \cs_registers_i/mtval_q_7_ ;
 wire \cs_registers_i/mtval_q_8_ ;
 wire \cs_registers_i/mtval_q_9_ ;
 wire \register_file_i/_0000_ ;
 wire \register_file_i/_0001_ ;
 wire \register_file_i/_0002_ ;
 wire \register_file_i/_0003_ ;
 wire \register_file_i/_0004_ ;
 wire \register_file_i/_0005_ ;
 wire \register_file_i/_0006_ ;
 wire \register_file_i/_0007_ ;
 wire \register_file_i/_0008_ ;
 wire \register_file_i/_0009_ ;
 wire \register_file_i/_0010_ ;
 wire \register_file_i/_0011_ ;
 wire \register_file_i/_0012_ ;
 wire \register_file_i/_0013_ ;
 wire \register_file_i/_0014_ ;
 wire \register_file_i/_0015_ ;
 wire \register_file_i/_0016_ ;
 wire \register_file_i/_0017_ ;
 wire \register_file_i/_0018_ ;
 wire \register_file_i/_0019_ ;
 wire \register_file_i/_0020_ ;
 wire \register_file_i/_0021_ ;
 wire \register_file_i/_0022_ ;
 wire \register_file_i/_0023_ ;
 wire \register_file_i/_0024_ ;
 wire \register_file_i/_0025_ ;
 wire \register_file_i/_0026_ ;
 wire \register_file_i/_0027_ ;
 wire \register_file_i/_0028_ ;
 wire \register_file_i/_0029_ ;
 wire \register_file_i/_0030_ ;
 wire \register_file_i/_0031_ ;
 wire \register_file_i/_0032_ ;
 wire \register_file_i/_0033_ ;
 wire \register_file_i/_0034_ ;
 wire \register_file_i/_0035_ ;
 wire \register_file_i/_0036_ ;
 wire \register_file_i/_0037_ ;
 wire \register_file_i/_0038_ ;
 wire \register_file_i/_0039_ ;
 wire \register_file_i/_0040_ ;
 wire \register_file_i/_0041_ ;
 wire \register_file_i/_0042_ ;
 wire \register_file_i/_0043_ ;
 wire \register_file_i/_0044_ ;
 wire \register_file_i/_0045_ ;
 wire \register_file_i/_0046_ ;
 wire \register_file_i/_0047_ ;
 wire \register_file_i/_0048_ ;
 wire \register_file_i/_0049_ ;
 wire \register_file_i/_0050_ ;
 wire \register_file_i/_0051_ ;
 wire \register_file_i/_0052_ ;
 wire \register_file_i/_0053_ ;
 wire \register_file_i/_0054_ ;
 wire \register_file_i/_0055_ ;
 wire \register_file_i/_0056_ ;
 wire \register_file_i/_0057_ ;
 wire \register_file_i/_0058_ ;
 wire \register_file_i/_0059_ ;
 wire \register_file_i/_0060_ ;
 wire \register_file_i/_0061_ ;
 wire \register_file_i/_0062_ ;
 wire \register_file_i/_0063_ ;
 wire \register_file_i/_0064_ ;
 wire \register_file_i/_0065_ ;
 wire \register_file_i/_0066_ ;
 wire \register_file_i/_0067_ ;
 wire \register_file_i/_0068_ ;
 wire \register_file_i/_0069_ ;
 wire \register_file_i/_0070_ ;
 wire \register_file_i/_0071_ ;
 wire \register_file_i/_0072_ ;
 wire \register_file_i/_0073_ ;
 wire \register_file_i/_0074_ ;
 wire \register_file_i/_0075_ ;
 wire \register_file_i/_0076_ ;
 wire \register_file_i/_0077_ ;
 wire \register_file_i/_0078_ ;
 wire \register_file_i/_0079_ ;
 wire \register_file_i/_0080_ ;
 wire \register_file_i/_0081_ ;
 wire \register_file_i/_0082_ ;
 wire \register_file_i/_0083_ ;
 wire \register_file_i/_0084_ ;
 wire \register_file_i/_0085_ ;
 wire \register_file_i/_0086_ ;
 wire \register_file_i/_0087_ ;
 wire \register_file_i/_0088_ ;
 wire \register_file_i/_0089_ ;
 wire \register_file_i/_0090_ ;
 wire \register_file_i/_0091_ ;
 wire \register_file_i/_0092_ ;
 wire \register_file_i/_0093_ ;
 wire \register_file_i/_0094_ ;
 wire \register_file_i/_0095_ ;
 wire \register_file_i/_0096_ ;
 wire \register_file_i/_0097_ ;
 wire \register_file_i/_0098_ ;
 wire \register_file_i/_0099_ ;
 wire \register_file_i/_0100_ ;
 wire \register_file_i/_0101_ ;
 wire \register_file_i/_0102_ ;
 wire \register_file_i/_0103_ ;
 wire \register_file_i/_0104_ ;
 wire \register_file_i/_0105_ ;
 wire \register_file_i/_0106_ ;
 wire \register_file_i/_0107_ ;
 wire \register_file_i/_0108_ ;
 wire \register_file_i/_0109_ ;
 wire \register_file_i/_0110_ ;
 wire \register_file_i/_0111_ ;
 wire \register_file_i/_0112_ ;
 wire \register_file_i/_0113_ ;
 wire \register_file_i/_0114_ ;
 wire \register_file_i/_0115_ ;
 wire \register_file_i/_0116_ ;
 wire \register_file_i/_0117_ ;
 wire \register_file_i/_0118_ ;
 wire \register_file_i/_0119_ ;
 wire \register_file_i/_0120_ ;
 wire \register_file_i/_0121_ ;
 wire \register_file_i/_0122_ ;
 wire \register_file_i/_0123_ ;
 wire \register_file_i/_0124_ ;
 wire \register_file_i/_0125_ ;
 wire \register_file_i/_0126_ ;
 wire \register_file_i/_0127_ ;
 wire \register_file_i/_0128_ ;
 wire \register_file_i/_0129_ ;
 wire \register_file_i/_0130_ ;
 wire \register_file_i/_0131_ ;
 wire \register_file_i/_0132_ ;
 wire \register_file_i/_0133_ ;
 wire \register_file_i/_0134_ ;
 wire \register_file_i/_0135_ ;
 wire \register_file_i/_0136_ ;
 wire \register_file_i/_0137_ ;
 wire \register_file_i/_0138_ ;
 wire \register_file_i/_0139_ ;
 wire \register_file_i/_0140_ ;
 wire \register_file_i/_0141_ ;
 wire \register_file_i/_0142_ ;
 wire \register_file_i/_0143_ ;
 wire \register_file_i/_0144_ ;
 wire \register_file_i/_0145_ ;
 wire \register_file_i/_0146_ ;
 wire \register_file_i/_0147_ ;
 wire \register_file_i/_0148_ ;
 wire \register_file_i/_0149_ ;
 wire \register_file_i/_0150_ ;
 wire \register_file_i/_0151_ ;
 wire \register_file_i/_0152_ ;
 wire \register_file_i/_0153_ ;
 wire \register_file_i/_0154_ ;
 wire \register_file_i/_0155_ ;
 wire \register_file_i/_0156_ ;
 wire \register_file_i/_0157_ ;
 wire \register_file_i/_0158_ ;
 wire \register_file_i/_0159_ ;
 wire \register_file_i/_0160_ ;
 wire \register_file_i/_0161_ ;
 wire \register_file_i/_0162_ ;
 wire \register_file_i/_0163_ ;
 wire \register_file_i/_0164_ ;
 wire \register_file_i/_0165_ ;
 wire \register_file_i/_0166_ ;
 wire \register_file_i/_0167_ ;
 wire \register_file_i/_0168_ ;
 wire \register_file_i/_0169_ ;
 wire \register_file_i/_0170_ ;
 wire \register_file_i/_0171_ ;
 wire \register_file_i/_0172_ ;
 wire \register_file_i/_0173_ ;
 wire \register_file_i/_0174_ ;
 wire \register_file_i/_0175_ ;
 wire \register_file_i/_0176_ ;
 wire \register_file_i/_0177_ ;
 wire \register_file_i/_0178_ ;
 wire \register_file_i/_0179_ ;
 wire \register_file_i/_0180_ ;
 wire \register_file_i/_0181_ ;
 wire \register_file_i/_0182_ ;
 wire \register_file_i/_0183_ ;
 wire \register_file_i/_0184_ ;
 wire \register_file_i/_0185_ ;
 wire \register_file_i/_0186_ ;
 wire \register_file_i/_0187_ ;
 wire \register_file_i/_0188_ ;
 wire \register_file_i/_0189_ ;
 wire \register_file_i/_0190_ ;
 wire \register_file_i/_0191_ ;
 wire \register_file_i/_0192_ ;
 wire \register_file_i/_0193_ ;
 wire \register_file_i/_0194_ ;
 wire \register_file_i/_0195_ ;
 wire \register_file_i/_0196_ ;
 wire \register_file_i/_0197_ ;
 wire \register_file_i/_0198_ ;
 wire \register_file_i/_0199_ ;
 wire \register_file_i/_0200_ ;
 wire \register_file_i/_0201_ ;
 wire \register_file_i/_0202_ ;
 wire \register_file_i/_0203_ ;
 wire \register_file_i/_0204_ ;
 wire \register_file_i/_0205_ ;
 wire \register_file_i/_0206_ ;
 wire \register_file_i/_0207_ ;
 wire \register_file_i/_0208_ ;
 wire \register_file_i/_0209_ ;
 wire \register_file_i/_0210_ ;
 wire \register_file_i/_0211_ ;
 wire \register_file_i/_0212_ ;
 wire \register_file_i/_0213_ ;
 wire \register_file_i/_0214_ ;
 wire \register_file_i/_0215_ ;
 wire \register_file_i/_0216_ ;
 wire \register_file_i/_0217_ ;
 wire \register_file_i/_0218_ ;
 wire \register_file_i/_0219_ ;
 wire \register_file_i/_0220_ ;
 wire \register_file_i/_0221_ ;
 wire \register_file_i/_0222_ ;
 wire \register_file_i/_0223_ ;
 wire \register_file_i/_0224_ ;
 wire \register_file_i/_0225_ ;
 wire \register_file_i/_0226_ ;
 wire \register_file_i/_0227_ ;
 wire \register_file_i/_0228_ ;
 wire \register_file_i/_0229_ ;
 wire \register_file_i/_0230_ ;
 wire \register_file_i/_0231_ ;
 wire \register_file_i/_0232_ ;
 wire \register_file_i/_0233_ ;
 wire \register_file_i/_0234_ ;
 wire \register_file_i/_0235_ ;
 wire \register_file_i/_0236_ ;
 wire \register_file_i/_0237_ ;
 wire \register_file_i/_0238_ ;
 wire \register_file_i/_0239_ ;
 wire \register_file_i/_0240_ ;
 wire \register_file_i/_0241_ ;
 wire \register_file_i/_0242_ ;
 wire \register_file_i/_0243_ ;
 wire \register_file_i/_0244_ ;
 wire \register_file_i/_0245_ ;
 wire \register_file_i/_0246_ ;
 wire \register_file_i/_0247_ ;
 wire \register_file_i/_0248_ ;
 wire \register_file_i/_0249_ ;
 wire \register_file_i/_0250_ ;
 wire \register_file_i/_0251_ ;
 wire \register_file_i/_0252_ ;
 wire \register_file_i/_0253_ ;
 wire \register_file_i/_0254_ ;
 wire \register_file_i/_0255_ ;
 wire \register_file_i/_0256_ ;
 wire \register_file_i/_0257_ ;
 wire \register_file_i/_0258_ ;
 wire \register_file_i/_0259_ ;
 wire \register_file_i/_0260_ ;
 wire \register_file_i/_0261_ ;
 wire \register_file_i/_0262_ ;
 wire \register_file_i/_0263_ ;
 wire \register_file_i/_0264_ ;
 wire \register_file_i/_0265_ ;
 wire \register_file_i/_0266_ ;
 wire \register_file_i/_0267_ ;
 wire \register_file_i/_0268_ ;
 wire \register_file_i/_0269_ ;
 wire \register_file_i/_0270_ ;
 wire \register_file_i/_0271_ ;
 wire \register_file_i/_0272_ ;
 wire \register_file_i/_0273_ ;
 wire \register_file_i/_0274_ ;
 wire \register_file_i/_0275_ ;
 wire \register_file_i/_0276_ ;
 wire \register_file_i/_0277_ ;
 wire \register_file_i/_0278_ ;
 wire \register_file_i/_0279_ ;
 wire \register_file_i/_0280_ ;
 wire \register_file_i/_0281_ ;
 wire \register_file_i/_0282_ ;
 wire \register_file_i/_0283_ ;
 wire \register_file_i/_0284_ ;
 wire \register_file_i/_0285_ ;
 wire \register_file_i/_0286_ ;
 wire \register_file_i/_0287_ ;
 wire \register_file_i/_0288_ ;
 wire \register_file_i/_0289_ ;
 wire \register_file_i/_0290_ ;
 wire \register_file_i/_0291_ ;
 wire \register_file_i/_0292_ ;
 wire \register_file_i/_0293_ ;
 wire \register_file_i/_0294_ ;
 wire \register_file_i/_0295_ ;
 wire \register_file_i/_0296_ ;
 wire \register_file_i/_0297_ ;
 wire \register_file_i/_0298_ ;
 wire \register_file_i/_0299_ ;
 wire \register_file_i/_0300_ ;
 wire \register_file_i/_0301_ ;
 wire \register_file_i/_0302_ ;
 wire \register_file_i/_0303_ ;
 wire \register_file_i/_0304_ ;
 wire \register_file_i/_0305_ ;
 wire \register_file_i/_0306_ ;
 wire \register_file_i/_0307_ ;
 wire \register_file_i/_0308_ ;
 wire \register_file_i/_0309_ ;
 wire \register_file_i/_0310_ ;
 wire \register_file_i/_0311_ ;
 wire \register_file_i/_0312_ ;
 wire \register_file_i/_0313_ ;
 wire \register_file_i/_0314_ ;
 wire \register_file_i/_0315_ ;
 wire \register_file_i/_0316_ ;
 wire \register_file_i/_0317_ ;
 wire \register_file_i/_0318_ ;
 wire \register_file_i/_0319_ ;
 wire \register_file_i/_0320_ ;
 wire \register_file_i/_0321_ ;
 wire \register_file_i/_0322_ ;
 wire \register_file_i/_0323_ ;
 wire \register_file_i/_0324_ ;
 wire \register_file_i/_0325_ ;
 wire \register_file_i/_0326_ ;
 wire \register_file_i/_0327_ ;
 wire \register_file_i/_0328_ ;
 wire \register_file_i/_0329_ ;
 wire \register_file_i/_0330_ ;
 wire \register_file_i/_0331_ ;
 wire \register_file_i/_0332_ ;
 wire \register_file_i/_0333_ ;
 wire \register_file_i/_0334_ ;
 wire \register_file_i/_0335_ ;
 wire \register_file_i/_0336_ ;
 wire \register_file_i/_0337_ ;
 wire \register_file_i/_0338_ ;
 wire \register_file_i/_0339_ ;
 wire \register_file_i/_0340_ ;
 wire \register_file_i/_0341_ ;
 wire \register_file_i/_0342_ ;
 wire \register_file_i/_0343_ ;
 wire \register_file_i/_0344_ ;
 wire \register_file_i/_0345_ ;
 wire \register_file_i/_0346_ ;
 wire \register_file_i/_0347_ ;
 wire \register_file_i/_0348_ ;
 wire \register_file_i/_0349_ ;
 wire \register_file_i/_0350_ ;
 wire \register_file_i/_0351_ ;
 wire \register_file_i/_0352_ ;
 wire \register_file_i/_0353_ ;
 wire \register_file_i/_0354_ ;
 wire \register_file_i/_0355_ ;
 wire \register_file_i/_0356_ ;
 wire \register_file_i/_0357_ ;
 wire \register_file_i/_0358_ ;
 wire \register_file_i/_0359_ ;
 wire \register_file_i/_0360_ ;
 wire \register_file_i/_0361_ ;
 wire \register_file_i/_0362_ ;
 wire \register_file_i/_0363_ ;
 wire \register_file_i/_0364_ ;
 wire \register_file_i/_0365_ ;
 wire \register_file_i/_0366_ ;
 wire \register_file_i/_0367_ ;
 wire \register_file_i/_0368_ ;
 wire \register_file_i/_0369_ ;
 wire \register_file_i/_0370_ ;
 wire \register_file_i/_0371_ ;
 wire \register_file_i/_0372_ ;
 wire \register_file_i/_0373_ ;
 wire \register_file_i/_0374_ ;
 wire \register_file_i/_0375_ ;
 wire \register_file_i/_0376_ ;
 wire \register_file_i/_0377_ ;
 wire \register_file_i/_0378_ ;
 wire \register_file_i/_0379_ ;
 wire \register_file_i/_0380_ ;
 wire \register_file_i/_0381_ ;
 wire \register_file_i/_0382_ ;
 wire \register_file_i/_0383_ ;
 wire \register_file_i/_0384_ ;
 wire \register_file_i/_0385_ ;
 wire \register_file_i/_0386_ ;
 wire \register_file_i/_0387_ ;
 wire \register_file_i/_0388_ ;
 wire \register_file_i/_0389_ ;
 wire \register_file_i/_0390_ ;
 wire \register_file_i/_0391_ ;
 wire \register_file_i/_0392_ ;
 wire \register_file_i/_0393_ ;
 wire \register_file_i/_0394_ ;
 wire \register_file_i/_0395_ ;
 wire \register_file_i/_0396_ ;
 wire \register_file_i/_0397_ ;
 wire \register_file_i/_0398_ ;
 wire \register_file_i/_0399_ ;
 wire \register_file_i/_0400_ ;
 wire \register_file_i/_0401_ ;
 wire \register_file_i/_0402_ ;
 wire \register_file_i/_0403_ ;
 wire \register_file_i/_0404_ ;
 wire \register_file_i/_0405_ ;
 wire \register_file_i/_0406_ ;
 wire \register_file_i/_0407_ ;
 wire \register_file_i/_0408_ ;
 wire \register_file_i/_0409_ ;
 wire \register_file_i/_0410_ ;
 wire \register_file_i/_0411_ ;
 wire \register_file_i/_0412_ ;
 wire \register_file_i/_0413_ ;
 wire \register_file_i/_0414_ ;
 wire \register_file_i/_0415_ ;
 wire \register_file_i/_0416_ ;
 wire \register_file_i/_0417_ ;
 wire \register_file_i/_0418_ ;
 wire \register_file_i/_0419_ ;
 wire \register_file_i/_0420_ ;
 wire \register_file_i/_0421_ ;
 wire \register_file_i/_0422_ ;
 wire \register_file_i/_0423_ ;
 wire \register_file_i/_0424_ ;
 wire \register_file_i/_0425_ ;
 wire \register_file_i/_0426_ ;
 wire \register_file_i/_0427_ ;
 wire \register_file_i/_0428_ ;
 wire \register_file_i/_0429_ ;
 wire \register_file_i/_0430_ ;
 wire \register_file_i/_0431_ ;
 wire \register_file_i/_0432_ ;
 wire \register_file_i/_0433_ ;
 wire \register_file_i/_0434_ ;
 wire \register_file_i/_0435_ ;
 wire \register_file_i/_0436_ ;
 wire \register_file_i/_0437_ ;
 wire \register_file_i/_0438_ ;
 wire \register_file_i/_0439_ ;
 wire \register_file_i/_0440_ ;
 wire \register_file_i/_0441_ ;
 wire \register_file_i/_0442_ ;
 wire \register_file_i/_0443_ ;
 wire \register_file_i/_0444_ ;
 wire \register_file_i/_0445_ ;
 wire \register_file_i/_0446_ ;
 wire \register_file_i/_0447_ ;
 wire \register_file_i/_0448_ ;
 wire \register_file_i/_0449_ ;
 wire \register_file_i/_0450_ ;
 wire \register_file_i/_0451_ ;
 wire \register_file_i/_0452_ ;
 wire \register_file_i/_0453_ ;
 wire \register_file_i/_0454_ ;
 wire \register_file_i/_0455_ ;
 wire \register_file_i/_0456_ ;
 wire \register_file_i/_0457_ ;
 wire \register_file_i/_0458_ ;
 wire \register_file_i/_0459_ ;
 wire \register_file_i/_0460_ ;
 wire \register_file_i/_0461_ ;
 wire \register_file_i/_0462_ ;
 wire \register_file_i/_0463_ ;
 wire \register_file_i/_0464_ ;
 wire \register_file_i/_0465_ ;
 wire \register_file_i/_0466_ ;
 wire \register_file_i/_0467_ ;
 wire \register_file_i/_0468_ ;
 wire \register_file_i/_0469_ ;
 wire \register_file_i/_0470_ ;
 wire \register_file_i/_0471_ ;
 wire \register_file_i/_0472_ ;
 wire \register_file_i/_0473_ ;
 wire \register_file_i/_0474_ ;
 wire \register_file_i/_0475_ ;
 wire \register_file_i/_0476_ ;
 wire \register_file_i/_0477_ ;
 wire \register_file_i/_0478_ ;
 wire \register_file_i/_0479_ ;
 wire \register_file_i/_0480_ ;
 wire \register_file_i/_0481_ ;
 wire \register_file_i/_0482_ ;
 wire \register_file_i/_0483_ ;
 wire \register_file_i/_0484_ ;
 wire \register_file_i/_0485_ ;
 wire \register_file_i/_0486_ ;
 wire \register_file_i/_0487_ ;
 wire \register_file_i/_0488_ ;
 wire \register_file_i/_0489_ ;
 wire \register_file_i/_0490_ ;
 wire \register_file_i/_0491_ ;
 wire \register_file_i/_0492_ ;
 wire \register_file_i/_0493_ ;
 wire \register_file_i/_0494_ ;
 wire \register_file_i/_0495_ ;
 wire \register_file_i/_0496_ ;
 wire \register_file_i/_0497_ ;
 wire \register_file_i/_0498_ ;
 wire \register_file_i/_0499_ ;
 wire \register_file_i/_0500_ ;
 wire \register_file_i/_0501_ ;
 wire \register_file_i/_0502_ ;
 wire \register_file_i/_0503_ ;
 wire \register_file_i/_0504_ ;
 wire \register_file_i/_0505_ ;
 wire \register_file_i/_0506_ ;
 wire \register_file_i/_0507_ ;
 wire \register_file_i/_0508_ ;
 wire \register_file_i/_0509_ ;
 wire \register_file_i/_0510_ ;
 wire \register_file_i/_0511_ ;
 wire \register_file_i/_0512_ ;
 wire \register_file_i/_0513_ ;
 wire \register_file_i/_0514_ ;
 wire \register_file_i/_0515_ ;
 wire \register_file_i/_0516_ ;
 wire \register_file_i/_0517_ ;
 wire \register_file_i/_0518_ ;
 wire \register_file_i/_0519_ ;
 wire \register_file_i/_0520_ ;
 wire \register_file_i/_0521_ ;
 wire \register_file_i/_0522_ ;
 wire \register_file_i/_0523_ ;
 wire \register_file_i/_0524_ ;
 wire \register_file_i/_0525_ ;
 wire \register_file_i/_0526_ ;
 wire \register_file_i/_0527_ ;
 wire \register_file_i/_0528_ ;
 wire \register_file_i/_0529_ ;
 wire \register_file_i/_0530_ ;
 wire \register_file_i/_0531_ ;
 wire \register_file_i/_0532_ ;
 wire \register_file_i/_0533_ ;
 wire \register_file_i/_0534_ ;
 wire \register_file_i/_0535_ ;
 wire \register_file_i/_0536_ ;
 wire \register_file_i/_0537_ ;
 wire \register_file_i/_0538_ ;
 wire \register_file_i/_0539_ ;
 wire \register_file_i/_0540_ ;
 wire \register_file_i/_0541_ ;
 wire \register_file_i/_0542_ ;
 wire \register_file_i/_0543_ ;
 wire \register_file_i/_0544_ ;
 wire \register_file_i/_0545_ ;
 wire \register_file_i/_0546_ ;
 wire \register_file_i/_0547_ ;
 wire \register_file_i/_0548_ ;
 wire \register_file_i/_0549_ ;
 wire \register_file_i/_0550_ ;
 wire \register_file_i/_0551_ ;
 wire \register_file_i/_0552_ ;
 wire \register_file_i/_0553_ ;
 wire \register_file_i/_0554_ ;
 wire \register_file_i/_0555_ ;
 wire \register_file_i/_0556_ ;
 wire \register_file_i/_0557_ ;
 wire \register_file_i/_0558_ ;
 wire \register_file_i/_0559_ ;
 wire \register_file_i/_0560_ ;
 wire \register_file_i/_0561_ ;
 wire \register_file_i/_0562_ ;
 wire \register_file_i/_0563_ ;
 wire \register_file_i/_0564_ ;
 wire \register_file_i/_0565_ ;
 wire \register_file_i/_0566_ ;
 wire \register_file_i/_0567_ ;
 wire \register_file_i/_0568_ ;
 wire \register_file_i/_0569_ ;
 wire \register_file_i/_0570_ ;
 wire \register_file_i/_0571_ ;
 wire \register_file_i/_0572_ ;
 wire \register_file_i/_0573_ ;
 wire \register_file_i/_0574_ ;
 wire \register_file_i/_0575_ ;
 wire \register_file_i/_0576_ ;
 wire \register_file_i/_0577_ ;
 wire \register_file_i/_0578_ ;
 wire \register_file_i/_0579_ ;
 wire \register_file_i/_0580_ ;
 wire \register_file_i/_0581_ ;
 wire \register_file_i/_0582_ ;
 wire \register_file_i/_0583_ ;
 wire \register_file_i/_0584_ ;
 wire \register_file_i/_0585_ ;
 wire \register_file_i/_0586_ ;
 wire \register_file_i/_0587_ ;
 wire \register_file_i/_0588_ ;
 wire \register_file_i/_0589_ ;
 wire \register_file_i/_0590_ ;
 wire \register_file_i/_0591_ ;
 wire \register_file_i/_0592_ ;
 wire \register_file_i/_0593_ ;
 wire \register_file_i/_0594_ ;
 wire \register_file_i/_0595_ ;
 wire \register_file_i/_0596_ ;
 wire \register_file_i/_0597_ ;
 wire \register_file_i/_0598_ ;
 wire \register_file_i/_0599_ ;
 wire \register_file_i/_0600_ ;
 wire \register_file_i/_0601_ ;
 wire \register_file_i/_0602_ ;
 wire \register_file_i/_0603_ ;
 wire \register_file_i/_0604_ ;
 wire \register_file_i/_0605_ ;
 wire \register_file_i/_0606_ ;
 wire \register_file_i/_0607_ ;
 wire \register_file_i/_0608_ ;
 wire \register_file_i/_0609_ ;
 wire \register_file_i/_0610_ ;
 wire \register_file_i/_0611_ ;
 wire \register_file_i/_0612_ ;
 wire \register_file_i/_0613_ ;
 wire \register_file_i/_0614_ ;
 wire \register_file_i/_0615_ ;
 wire \register_file_i/_0616_ ;
 wire \register_file_i/_0617_ ;
 wire \register_file_i/_0618_ ;
 wire \register_file_i/_0619_ ;
 wire \register_file_i/_0620_ ;
 wire \register_file_i/_0621_ ;
 wire \register_file_i/_0622_ ;
 wire \register_file_i/_0623_ ;
 wire \register_file_i/_0624_ ;
 wire \register_file_i/_0625_ ;
 wire \register_file_i/_0626_ ;
 wire \register_file_i/_0627_ ;
 wire \register_file_i/_0628_ ;
 wire \register_file_i/_0629_ ;
 wire \register_file_i/_0630_ ;
 wire \register_file_i/_0631_ ;
 wire \register_file_i/_0632_ ;
 wire \register_file_i/_0633_ ;
 wire \register_file_i/_0634_ ;
 wire \register_file_i/_0635_ ;
 wire \register_file_i/_0636_ ;
 wire \register_file_i/_0637_ ;
 wire \register_file_i/_0638_ ;
 wire \register_file_i/_0639_ ;
 wire \register_file_i/_0640_ ;
 wire \register_file_i/_0641_ ;
 wire \register_file_i/_0642_ ;
 wire \register_file_i/_0643_ ;
 wire \register_file_i/_0644_ ;
 wire \register_file_i/_0645_ ;
 wire \register_file_i/_0646_ ;
 wire \register_file_i/_0647_ ;
 wire \register_file_i/_0648_ ;
 wire \register_file_i/_0649_ ;
 wire \register_file_i/_0650_ ;
 wire \register_file_i/_0651_ ;
 wire \register_file_i/_0652_ ;
 wire \register_file_i/_0653_ ;
 wire \register_file_i/_0654_ ;
 wire \register_file_i/_0655_ ;
 wire \register_file_i/_0656_ ;
 wire \register_file_i/_0657_ ;
 wire \register_file_i/_0658_ ;
 wire \register_file_i/_0659_ ;
 wire \register_file_i/_0660_ ;
 wire \register_file_i/_0661_ ;
 wire \register_file_i/_0662_ ;
 wire \register_file_i/_0663_ ;
 wire \register_file_i/_0664_ ;
 wire \register_file_i/_0665_ ;
 wire \register_file_i/_0666_ ;
 wire \register_file_i/_0667_ ;
 wire \register_file_i/_0668_ ;
 wire \register_file_i/_0669_ ;
 wire \register_file_i/_0670_ ;
 wire \register_file_i/_0671_ ;
 wire \register_file_i/_0672_ ;
 wire \register_file_i/_0673_ ;
 wire \register_file_i/_0674_ ;
 wire \register_file_i/_0675_ ;
 wire \register_file_i/_0676_ ;
 wire \register_file_i/_0677_ ;
 wire \register_file_i/_0678_ ;
 wire \register_file_i/_0679_ ;
 wire \register_file_i/_0680_ ;
 wire \register_file_i/_0681_ ;
 wire \register_file_i/_0682_ ;
 wire \register_file_i/_0683_ ;
 wire \register_file_i/_0684_ ;
 wire \register_file_i/_0685_ ;
 wire \register_file_i/_0686_ ;
 wire \register_file_i/_0687_ ;
 wire \register_file_i/_0688_ ;
 wire \register_file_i/_0689_ ;
 wire \register_file_i/_0690_ ;
 wire \register_file_i/_0691_ ;
 wire \register_file_i/_0692_ ;
 wire \register_file_i/_0693_ ;
 wire \register_file_i/_0694_ ;
 wire \register_file_i/_0695_ ;
 wire \register_file_i/_0696_ ;
 wire \register_file_i/_0697_ ;
 wire \register_file_i/_0698_ ;
 wire \register_file_i/_0699_ ;
 wire \register_file_i/_0700_ ;
 wire \register_file_i/_0701_ ;
 wire \register_file_i/_0702_ ;
 wire \register_file_i/_0703_ ;
 wire \register_file_i/_0704_ ;
 wire \register_file_i/_0705_ ;
 wire \register_file_i/_0706_ ;
 wire \register_file_i/_0707_ ;
 wire \register_file_i/_0708_ ;
 wire \register_file_i/_0709_ ;
 wire \register_file_i/_0710_ ;
 wire \register_file_i/_0711_ ;
 wire \register_file_i/_0712_ ;
 wire \register_file_i/_0713_ ;
 wire \register_file_i/_0714_ ;
 wire \register_file_i/_0715_ ;
 wire \register_file_i/_0716_ ;
 wire \register_file_i/_0717_ ;
 wire \register_file_i/_0718_ ;
 wire \register_file_i/_0719_ ;
 wire \register_file_i/_0720_ ;
 wire \register_file_i/_0721_ ;
 wire \register_file_i/_0722_ ;
 wire \register_file_i/_0723_ ;
 wire \register_file_i/_0724_ ;
 wire \register_file_i/_0725_ ;
 wire \register_file_i/_0726_ ;
 wire \register_file_i/_0727_ ;
 wire \register_file_i/_0728_ ;
 wire \register_file_i/_0729_ ;
 wire \register_file_i/_0730_ ;
 wire \register_file_i/_0731_ ;
 wire \register_file_i/_0732_ ;
 wire \register_file_i/_0733_ ;
 wire \register_file_i/_0734_ ;
 wire \register_file_i/_0735_ ;
 wire \register_file_i/_0736_ ;
 wire \register_file_i/_0737_ ;
 wire \register_file_i/_0738_ ;
 wire \register_file_i/_0739_ ;
 wire \register_file_i/_0740_ ;
 wire \register_file_i/_0741_ ;
 wire \register_file_i/_0742_ ;
 wire \register_file_i/_0743_ ;
 wire \register_file_i/_0744_ ;
 wire \register_file_i/_0745_ ;
 wire \register_file_i/_0746_ ;
 wire \register_file_i/_0747_ ;
 wire \register_file_i/_0748_ ;
 wire \register_file_i/_0749_ ;
 wire \register_file_i/_0750_ ;
 wire \register_file_i/_0751_ ;
 wire \register_file_i/_0752_ ;
 wire \register_file_i/_0753_ ;
 wire \register_file_i/_0754_ ;
 wire \register_file_i/_0755_ ;
 wire \register_file_i/_0756_ ;
 wire \register_file_i/_0757_ ;
 wire \register_file_i/_0758_ ;
 wire \register_file_i/_0759_ ;
 wire \register_file_i/_0760_ ;
 wire \register_file_i/_0761_ ;
 wire \register_file_i/_0762_ ;
 wire \register_file_i/_0763_ ;
 wire \register_file_i/_0764_ ;
 wire \register_file_i/_0765_ ;
 wire \register_file_i/_0766_ ;
 wire \register_file_i/_0767_ ;
 wire \register_file_i/_0768_ ;
 wire \register_file_i/_0769_ ;
 wire \register_file_i/_0770_ ;
 wire \register_file_i/_0771_ ;
 wire \register_file_i/_0772_ ;
 wire \register_file_i/_0773_ ;
 wire \register_file_i/_0774_ ;
 wire \register_file_i/_0775_ ;
 wire \register_file_i/_0776_ ;
 wire \register_file_i/_0777_ ;
 wire \register_file_i/_0778_ ;
 wire \register_file_i/_0779_ ;
 wire \register_file_i/_0780_ ;
 wire \register_file_i/_0781_ ;
 wire \register_file_i/_0782_ ;
 wire \register_file_i/_0783_ ;
 wire \register_file_i/_0784_ ;
 wire \register_file_i/_0785_ ;
 wire \register_file_i/_0786_ ;
 wire \register_file_i/_0787_ ;
 wire \register_file_i/_0788_ ;
 wire \register_file_i/_0789_ ;
 wire \register_file_i/_0790_ ;
 wire \register_file_i/_0791_ ;
 wire \register_file_i/_0792_ ;
 wire \register_file_i/_0793_ ;
 wire \register_file_i/_0794_ ;
 wire \register_file_i/_0795_ ;
 wire \register_file_i/_0796_ ;
 wire \register_file_i/_0797_ ;
 wire \register_file_i/_0798_ ;
 wire \register_file_i/_0799_ ;
 wire \register_file_i/_0800_ ;
 wire \register_file_i/_0801_ ;
 wire \register_file_i/_0802_ ;
 wire \register_file_i/_0803_ ;
 wire \register_file_i/_0804_ ;
 wire \register_file_i/_0805_ ;
 wire \register_file_i/_0806_ ;
 wire \register_file_i/_0807_ ;
 wire \register_file_i/_0808_ ;
 wire \register_file_i/_0809_ ;
 wire \register_file_i/_0810_ ;
 wire \register_file_i/_0811_ ;
 wire \register_file_i/_0812_ ;
 wire \register_file_i/_0813_ ;
 wire \register_file_i/_0814_ ;
 wire \register_file_i/_0815_ ;
 wire \register_file_i/_0816_ ;
 wire \register_file_i/_0817_ ;
 wire \register_file_i/_0818_ ;
 wire \register_file_i/_0819_ ;
 wire \register_file_i/_0820_ ;
 wire \register_file_i/_0821_ ;
 wire \register_file_i/_0822_ ;
 wire \register_file_i/_0823_ ;
 wire \register_file_i/_0824_ ;
 wire \register_file_i/_0825_ ;
 wire \register_file_i/_0826_ ;
 wire \register_file_i/_0827_ ;
 wire \register_file_i/_0828_ ;
 wire \register_file_i/_0829_ ;
 wire \register_file_i/_0830_ ;
 wire \register_file_i/_0831_ ;
 wire \register_file_i/_0832_ ;
 wire \register_file_i/_0833_ ;
 wire \register_file_i/_0834_ ;
 wire \register_file_i/_0835_ ;
 wire \register_file_i/_0836_ ;
 wire \register_file_i/_0837_ ;
 wire \register_file_i/_0838_ ;
 wire \register_file_i/_0839_ ;
 wire \register_file_i/_0840_ ;
 wire \register_file_i/_0841_ ;
 wire \register_file_i/_0842_ ;
 wire \register_file_i/_0843_ ;
 wire \register_file_i/_0844_ ;
 wire \register_file_i/_0845_ ;
 wire \register_file_i/_0846_ ;
 wire \register_file_i/_0847_ ;
 wire \register_file_i/_0848_ ;
 wire \register_file_i/_0849_ ;
 wire \register_file_i/_0850_ ;
 wire \register_file_i/_0851_ ;
 wire \register_file_i/_0852_ ;
 wire \register_file_i/_0853_ ;
 wire \register_file_i/_0854_ ;
 wire \register_file_i/_0855_ ;
 wire \register_file_i/_0856_ ;
 wire \register_file_i/_0857_ ;
 wire \register_file_i/_0858_ ;
 wire \register_file_i/_0859_ ;
 wire \register_file_i/_0860_ ;
 wire \register_file_i/_0861_ ;
 wire \register_file_i/_0862_ ;
 wire \register_file_i/_0863_ ;
 wire \register_file_i/_0864_ ;
 wire \register_file_i/_0865_ ;
 wire \register_file_i/_0866_ ;
 wire \register_file_i/_0867_ ;
 wire \register_file_i/_0868_ ;
 wire \register_file_i/_0869_ ;
 wire \register_file_i/_0870_ ;
 wire \register_file_i/_0871_ ;
 wire \register_file_i/_0872_ ;
 wire \register_file_i/_0873_ ;
 wire \register_file_i/_0874_ ;
 wire \register_file_i/_0875_ ;
 wire \register_file_i/_0876_ ;
 wire \register_file_i/_0877_ ;
 wire \register_file_i/_0878_ ;
 wire \register_file_i/_0879_ ;
 wire \register_file_i/_0880_ ;
 wire \register_file_i/_0881_ ;
 wire \register_file_i/_0882_ ;
 wire \register_file_i/_0883_ ;
 wire \register_file_i/_0884_ ;
 wire \register_file_i/_0885_ ;
 wire \register_file_i/_0886_ ;
 wire \register_file_i/_0887_ ;
 wire \register_file_i/_0888_ ;
 wire \register_file_i/_0889_ ;
 wire \register_file_i/_0890_ ;
 wire \register_file_i/_0891_ ;
 wire \register_file_i/_0892_ ;
 wire \register_file_i/_0893_ ;
 wire \register_file_i/_0894_ ;
 wire \register_file_i/_0895_ ;
 wire \register_file_i/_0896_ ;
 wire \register_file_i/_0897_ ;
 wire \register_file_i/_0898_ ;
 wire \register_file_i/_0899_ ;
 wire \register_file_i/_0900_ ;
 wire \register_file_i/_0901_ ;
 wire \register_file_i/_0902_ ;
 wire \register_file_i/_0903_ ;
 wire \register_file_i/_0904_ ;
 wire \register_file_i/_0905_ ;
 wire \register_file_i/_0906_ ;
 wire \register_file_i/_0907_ ;
 wire \register_file_i/_0908_ ;
 wire \register_file_i/_0909_ ;
 wire \register_file_i/_0910_ ;
 wire \register_file_i/_0911_ ;
 wire \register_file_i/_0912_ ;
 wire \register_file_i/_0913_ ;
 wire \register_file_i/_0914_ ;
 wire \register_file_i/_0915_ ;
 wire \register_file_i/_0916_ ;
 wire \register_file_i/_0917_ ;
 wire \register_file_i/_0918_ ;
 wire \register_file_i/_0919_ ;
 wire \register_file_i/_0920_ ;
 wire \register_file_i/_0921_ ;
 wire \register_file_i/_0922_ ;
 wire \register_file_i/_0923_ ;
 wire \register_file_i/_0924_ ;
 wire \register_file_i/_0925_ ;
 wire \register_file_i/_0926_ ;
 wire \register_file_i/_0927_ ;
 wire \register_file_i/_0928_ ;
 wire \register_file_i/_0929_ ;
 wire \register_file_i/_0930_ ;
 wire \register_file_i/_0931_ ;
 wire \register_file_i/_0932_ ;
 wire \register_file_i/_0933_ ;
 wire \register_file_i/_0934_ ;
 wire \register_file_i/_0935_ ;
 wire \register_file_i/_0936_ ;
 wire \register_file_i/_0937_ ;
 wire \register_file_i/_0938_ ;
 wire \register_file_i/_0939_ ;
 wire \register_file_i/_0940_ ;
 wire \register_file_i/_0941_ ;
 wire \register_file_i/_0942_ ;
 wire \register_file_i/_0943_ ;
 wire \register_file_i/_0944_ ;
 wire \register_file_i/_0945_ ;
 wire \register_file_i/_0946_ ;
 wire \register_file_i/_0947_ ;
 wire \register_file_i/_0948_ ;
 wire \register_file_i/_0949_ ;
 wire \register_file_i/_0950_ ;
 wire \register_file_i/_0951_ ;
 wire \register_file_i/_0952_ ;
 wire \register_file_i/_0953_ ;
 wire \register_file_i/_0954_ ;
 wire \register_file_i/_0955_ ;
 wire \register_file_i/_0956_ ;
 wire \register_file_i/_0957_ ;
 wire \register_file_i/_0958_ ;
 wire \register_file_i/_0959_ ;
 wire \register_file_i/_0960_ ;
 wire \register_file_i/_0961_ ;
 wire \register_file_i/_0962_ ;
 wire \register_file_i/_0963_ ;
 wire \register_file_i/_0964_ ;
 wire \register_file_i/_0965_ ;
 wire \register_file_i/_0966_ ;
 wire \register_file_i/_0967_ ;
 wire \register_file_i/_0968_ ;
 wire \register_file_i/_0969_ ;
 wire \register_file_i/_0970_ ;
 wire \register_file_i/_0971_ ;
 wire \register_file_i/_0972_ ;
 wire \register_file_i/_0973_ ;
 wire \register_file_i/_0974_ ;
 wire \register_file_i/_0975_ ;
 wire \register_file_i/_0976_ ;
 wire \register_file_i/_0977_ ;
 wire \register_file_i/_0978_ ;
 wire \register_file_i/_0979_ ;
 wire \register_file_i/_0980_ ;
 wire \register_file_i/_0981_ ;
 wire \register_file_i/_0982_ ;
 wire \register_file_i/_0983_ ;
 wire \register_file_i/_0984_ ;
 wire \register_file_i/_0985_ ;
 wire \register_file_i/_0986_ ;
 wire \register_file_i/_0987_ ;
 wire \register_file_i/_0988_ ;
 wire \register_file_i/_0989_ ;
 wire \register_file_i/_0990_ ;
 wire \register_file_i/_0991_ ;
 wire net433;
 wire net432;
 wire \register_file_i/_0994_ ;
 wire net431;
 wire net430;
 wire net429;
 wire net428;
 wire net427;
 wire \register_file_i/_1000_ ;
 wire net426;
 wire \register_file_i/_1002_ ;
 wire \register_file_i/_1003_ ;
 wire net425;
 wire net424;
 wire net423;
 wire \register_file_i/_1007_ ;
 wire \register_file_i/_1008_ ;
 wire net422;
 wire net421;
 wire \register_file_i/_1011_ ;
 wire net420;
 wire \register_file_i/_1013_ ;
 wire \register_file_i/_1014_ ;
 wire net419;
 wire net418;
 wire \register_file_i/_1017_ ;
 wire \register_file_i/_1018_ ;
 wire net417;
 wire \register_file_i/_1020_ ;
 wire \register_file_i/_1021_ ;
 wire net416;
 wire net415;
 wire net414;
 wire net413;
 wire net412;
 wire \register_file_i/_1027_ ;
 wire net411;
 wire \register_file_i/_1029_ ;
 wire net410;
 wire \register_file_i/_1031_ ;
 wire net409;
 wire net408;
 wire \register_file_i/_1034_ ;
 wire net407;
 wire \register_file_i/_1036_ ;
 wire net406;
 wire \register_file_i/_1038_ ;
 wire \register_file_i/_1039_ ;
 wire \register_file_i/_1040_ ;
 wire \register_file_i/_1041_ ;
 wire \register_file_i/_1042_ ;
 wire net405;
 wire net404;
 wire net403;
 wire net402;
 wire \register_file_i/_1047_ ;
 wire \register_file_i/_1048_ ;
 wire \register_file_i/_1049_ ;
 wire net401;
 wire net400;
 wire \register_file_i/_1052_ ;
 wire net399;
 wire net398;
 wire \register_file_i/_1055_ ;
 wire net397;
 wire net396;
 wire \register_file_i/_1058_ ;
 wire \register_file_i/_1059_ ;
 wire net395;
 wire \register_file_i/_1061_ ;
 wire net394;
 wire \register_file_i/_1063_ ;
 wire net393;
 wire \register_file_i/_1065_ ;
 wire \register_file_i/_1066_ ;
 wire net392;
 wire \register_file_i/_1068_ ;
 wire \register_file_i/_1069_ ;
 wire \register_file_i/_1070_ ;
 wire \register_file_i/_1071_ ;
 wire \register_file_i/_1072_ ;
 wire net391;
 wire \register_file_i/_1074_ ;
 wire \register_file_i/_1075_ ;
 wire \register_file_i/_1076_ ;
 wire \register_file_i/_1077_ ;
 wire \register_file_i/_1078_ ;
 wire net390;
 wire \register_file_i/_1080_ ;
 wire \register_file_i/_1081_ ;
 wire \register_file_i/_1082_ ;
 wire \register_file_i/_1083_ ;
 wire \register_file_i/_1084_ ;
 wire \register_file_i/_1085_ ;
 wire \register_file_i/_1086_ ;
 wire net389;
 wire net388;
 wire \register_file_i/_1089_ ;
 wire net387;
 wire \register_file_i/_1091_ ;
 wire \register_file_i/_1092_ ;
 wire net386;
 wire \register_file_i/_1094_ ;
 wire net385;
 wire \register_file_i/_1096_ ;
 wire \register_file_i/_1097_ ;
 wire \register_file_i/_1098_ ;
 wire \register_file_i/_1099_ ;
 wire \register_file_i/_1100_ ;
 wire \register_file_i/_1101_ ;
 wire \register_file_i/_1102_ ;
 wire \register_file_i/_1103_ ;
 wire \register_file_i/_1104_ ;
 wire \register_file_i/_1105_ ;
 wire \register_file_i/_1106_ ;
 wire \register_file_i/_1107_ ;
 wire \register_file_i/_1108_ ;
 wire \register_file_i/_1109_ ;
 wire \register_file_i/_1110_ ;
 wire \register_file_i/_1111_ ;
 wire \register_file_i/_1112_ ;
 wire \register_file_i/_1113_ ;
 wire \register_file_i/_1114_ ;
 wire \register_file_i/_1115_ ;
 wire \register_file_i/_1116_ ;
 wire net384;
 wire \register_file_i/_1118_ ;
 wire \register_file_i/_1119_ ;
 wire \register_file_i/_1120_ ;
 wire \register_file_i/_1121_ ;
 wire \register_file_i/_1122_ ;
 wire \register_file_i/_1123_ ;
 wire \register_file_i/_1124_ ;
 wire \register_file_i/_1125_ ;
 wire net383;
 wire \register_file_i/_1127_ ;
 wire \register_file_i/_1128_ ;
 wire \register_file_i/_1129_ ;
 wire \register_file_i/_1130_ ;
 wire \register_file_i/_1131_ ;
 wire \register_file_i/_1132_ ;
 wire \register_file_i/_1133_ ;
 wire \register_file_i/_1134_ ;
 wire \register_file_i/_1135_ ;
 wire \register_file_i/_1136_ ;
 wire \register_file_i/_1137_ ;
 wire \register_file_i/_1138_ ;
 wire \register_file_i/_1139_ ;
 wire \register_file_i/_1140_ ;
 wire \register_file_i/_1141_ ;
 wire \register_file_i/_1142_ ;
 wire \register_file_i/_1143_ ;
 wire \register_file_i/_1144_ ;
 wire \register_file_i/_1145_ ;
 wire \register_file_i/_1146_ ;
 wire net382;
 wire \register_file_i/_1148_ ;
 wire \register_file_i/_1149_ ;
 wire \register_file_i/_1150_ ;
 wire \register_file_i/_1151_ ;
 wire \register_file_i/_1152_ ;
 wire \register_file_i/_1153_ ;
 wire \register_file_i/_1154_ ;
 wire \register_file_i/_1155_ ;
 wire \register_file_i/_1156_ ;
 wire \register_file_i/_1157_ ;
 wire \register_file_i/_1158_ ;
 wire \register_file_i/_1159_ ;
 wire \register_file_i/_1160_ ;
 wire net381;
 wire \register_file_i/_1162_ ;
 wire \register_file_i/_1163_ ;
 wire \register_file_i/_1164_ ;
 wire \register_file_i/_1165_ ;
 wire \register_file_i/_1166_ ;
 wire net380;
 wire \register_file_i/_1168_ ;
 wire \register_file_i/_1169_ ;
 wire \register_file_i/_1170_ ;
 wire \register_file_i/_1171_ ;
 wire \register_file_i/_1172_ ;
 wire \register_file_i/_1173_ ;
 wire \register_file_i/_1174_ ;
 wire \register_file_i/_1175_ ;
 wire \register_file_i/_1176_ ;
 wire \register_file_i/_1177_ ;
 wire \register_file_i/_1178_ ;
 wire \register_file_i/_1179_ ;
 wire \register_file_i/_1180_ ;
 wire \register_file_i/_1181_ ;
 wire net379;
 wire \register_file_i/_1183_ ;
 wire \register_file_i/_1184_ ;
 wire \register_file_i/_1185_ ;
 wire \register_file_i/_1186_ ;
 wire \register_file_i/_1187_ ;
 wire \register_file_i/_1188_ ;
 wire \register_file_i/_1189_ ;
 wire \register_file_i/_1190_ ;
 wire \register_file_i/_1191_ ;
 wire \register_file_i/_1192_ ;
 wire \register_file_i/_1193_ ;
 wire net378;
 wire \register_file_i/_1195_ ;
 wire \register_file_i/_1196_ ;
 wire net377;
 wire \register_file_i/_1198_ ;
 wire \register_file_i/_1199_ ;
 wire \register_file_i/_1200_ ;
 wire \register_file_i/_1201_ ;
 wire \register_file_i/_1202_ ;
 wire \register_file_i/_1203_ ;
 wire \register_file_i/_1204_ ;
 wire \register_file_i/_1205_ ;
 wire \register_file_i/_1206_ ;
 wire \register_file_i/_1207_ ;
 wire \register_file_i/_1208_ ;
 wire \register_file_i/_1209_ ;
 wire \register_file_i/_1210_ ;
 wire \register_file_i/_1211_ ;
 wire \register_file_i/_1212_ ;
 wire \register_file_i/_1213_ ;
 wire \register_file_i/_1214_ ;
 wire \register_file_i/_1215_ ;
 wire \register_file_i/_1216_ ;
 wire \register_file_i/_1217_ ;
 wire \register_file_i/_1218_ ;
 wire net376;
 wire \register_file_i/_1220_ ;
 wire \register_file_i/_1221_ ;
 wire \register_file_i/_1222_ ;
 wire \register_file_i/_1223_ ;
 wire \register_file_i/_1224_ ;
 wire \register_file_i/_1225_ ;
 wire \register_file_i/_1226_ ;
 wire \register_file_i/_1227_ ;
 wire net375;
 wire \register_file_i/_1229_ ;
 wire \register_file_i/_1230_ ;
 wire \register_file_i/_1231_ ;
 wire \register_file_i/_1232_ ;
 wire \register_file_i/_1233_ ;
 wire \register_file_i/_1234_ ;
 wire \register_file_i/_1235_ ;
 wire \register_file_i/_1236_ ;
 wire \register_file_i/_1237_ ;
 wire net374;
 wire \register_file_i/_1239_ ;
 wire \register_file_i/_1240_ ;
 wire net373;
 wire \register_file_i/_1242_ ;
 wire \register_file_i/_1243_ ;
 wire \register_file_i/_1244_ ;
 wire \register_file_i/_1245_ ;
 wire \register_file_i/_1246_ ;
 wire \register_file_i/_1247_ ;
 wire \register_file_i/_1248_ ;
 wire \register_file_i/_1249_ ;
 wire \register_file_i/_1250_ ;
 wire net372;
 wire \register_file_i/_1252_ ;
 wire \register_file_i/_1253_ ;
 wire \register_file_i/_1254_ ;
 wire \register_file_i/_1255_ ;
 wire \register_file_i/_1256_ ;
 wire \register_file_i/_1257_ ;
 wire \register_file_i/_1258_ ;
 wire net371;
 wire \register_file_i/_1260_ ;
 wire \register_file_i/_1261_ ;
 wire \register_file_i/_1262_ ;
 wire \register_file_i/_1263_ ;
 wire \register_file_i/_1264_ ;
 wire \register_file_i/_1265_ ;
 wire \register_file_i/_1266_ ;
 wire \register_file_i/_1267_ ;
 wire \register_file_i/_1268_ ;
 wire \register_file_i/_1269_ ;
 wire net370;
 wire \register_file_i/_1271_ ;
 wire \register_file_i/_1272_ ;
 wire \register_file_i/_1273_ ;
 wire \register_file_i/_1274_ ;
 wire \register_file_i/_1275_ ;
 wire \register_file_i/_1276_ ;
 wire \register_file_i/_1277_ ;
 wire \register_file_i/_1278_ ;
 wire \register_file_i/_1279_ ;
 wire \register_file_i/_1280_ ;
 wire net369;
 wire \register_file_i/_1282_ ;
 wire \register_file_i/_1283_ ;
 wire \register_file_i/_1284_ ;
 wire \register_file_i/_1285_ ;
 wire \register_file_i/_1286_ ;
 wire \register_file_i/_1287_ ;
 wire \register_file_i/_1288_ ;
 wire \register_file_i/_1289_ ;
 wire \register_file_i/_1290_ ;
 wire \register_file_i/_1291_ ;
 wire \register_file_i/_1292_ ;
 wire \register_file_i/_1293_ ;
 wire \register_file_i/_1294_ ;
 wire net368;
 wire \register_file_i/_1296_ ;
 wire \register_file_i/_1297_ ;
 wire \register_file_i/_1298_ ;
 wire \register_file_i/_1299_ ;
 wire \register_file_i/_1300_ ;
 wire \register_file_i/_1301_ ;
 wire \register_file_i/_1302_ ;
 wire \register_file_i/_1303_ ;
 wire \register_file_i/_1304_ ;
 wire net367;
 wire net366;
 wire \register_file_i/_1307_ ;
 wire \register_file_i/_1308_ ;
 wire \register_file_i/_1309_ ;
 wire \register_file_i/_1310_ ;
 wire \register_file_i/_1311_ ;
 wire net365;
 wire \register_file_i/_1313_ ;
 wire \register_file_i/_1314_ ;
 wire net364;
 wire \register_file_i/_1316_ ;
 wire net363;
 wire \register_file_i/_1318_ ;
 wire \register_file_i/_1319_ ;
 wire net362;
 wire \register_file_i/_1321_ ;
 wire net361;
 wire \register_file_i/_1323_ ;
 wire net360;
 wire net359;
 wire net358;
 wire \register_file_i/_1327_ ;
 wire \register_file_i/_1328_ ;
 wire \register_file_i/_1329_ ;
 wire \register_file_i/_1330_ ;
 wire \register_file_i/_1331_ ;
 wire \register_file_i/_1332_ ;
 wire \register_file_i/_1333_ ;
 wire net357;
 wire \register_file_i/_1335_ ;
 wire \register_file_i/_1336_ ;
 wire net356;
 wire \register_file_i/_1338_ ;
 wire \register_file_i/_1339_ ;
 wire \register_file_i/_1340_ ;
 wire \register_file_i/_1341_ ;
 wire \register_file_i/_1342_ ;
 wire \register_file_i/_1343_ ;
 wire \register_file_i/_1344_ ;
 wire \register_file_i/_1345_ ;
 wire \register_file_i/_1346_ ;
 wire \register_file_i/_1347_ ;
 wire \register_file_i/_1348_ ;
 wire net355;
 wire \register_file_i/_1350_ ;
 wire \register_file_i/_1351_ ;
 wire \register_file_i/_1352_ ;
 wire \register_file_i/_1353_ ;
 wire \register_file_i/_1354_ ;
 wire net354;
 wire \register_file_i/_1356_ ;
 wire \register_file_i/_1357_ ;
 wire \register_file_i/_1358_ ;
 wire \register_file_i/_1359_ ;
 wire \register_file_i/_1360_ ;
 wire \register_file_i/_1361_ ;
 wire \register_file_i/_1362_ ;
 wire net353;
 wire \register_file_i/_1364_ ;
 wire net352;
 wire \register_file_i/_1366_ ;
 wire \register_file_i/_1367_ ;
 wire \register_file_i/_1368_ ;
 wire \register_file_i/_1369_ ;
 wire \register_file_i/_1370_ ;
 wire \register_file_i/_1371_ ;
 wire \register_file_i/_1372_ ;
 wire \register_file_i/_1373_ ;
 wire \register_file_i/_1374_ ;
 wire \register_file_i/_1375_ ;
 wire \register_file_i/_1376_ ;
 wire \register_file_i/_1377_ ;
 wire \register_file_i/_1378_ ;
 wire \register_file_i/_1379_ ;
 wire \register_file_i/_1380_ ;
 wire \register_file_i/_1381_ ;
 wire \register_file_i/_1382_ ;
 wire \register_file_i/_1383_ ;
 wire \register_file_i/_1384_ ;
 wire \register_file_i/_1385_ ;
 wire \register_file_i/_1386_ ;
 wire \register_file_i/_1387_ ;
 wire \register_file_i/_1388_ ;
 wire \register_file_i/_1389_ ;
 wire net351;
 wire \register_file_i/_1391_ ;
 wire \register_file_i/_1392_ ;
 wire \register_file_i/_1393_ ;
 wire \register_file_i/_1394_ ;
 wire \register_file_i/_1395_ ;
 wire \register_file_i/_1396_ ;
 wire \register_file_i/_1397_ ;
 wire \register_file_i/_1398_ ;
 wire net350;
 wire \register_file_i/_1400_ ;
 wire \register_file_i/_1401_ ;
 wire \register_file_i/_1402_ ;
 wire \register_file_i/_1403_ ;
 wire \register_file_i/_1404_ ;
 wire \register_file_i/_1405_ ;
 wire \register_file_i/_1406_ ;
 wire \register_file_i/_1407_ ;
 wire \register_file_i/_1408_ ;
 wire \register_file_i/_1409_ ;
 wire \register_file_i/_1410_ ;
 wire \register_file_i/_1411_ ;
 wire \register_file_i/_1412_ ;
 wire \register_file_i/_1413_ ;
 wire \register_file_i/_1414_ ;
 wire \register_file_i/_1415_ ;
 wire \register_file_i/_1416_ ;
 wire \register_file_i/_1417_ ;
 wire \register_file_i/_1418_ ;
 wire \register_file_i/_1419_ ;
 wire net349;
 wire \register_file_i/_1421_ ;
 wire \register_file_i/_1422_ ;
 wire \register_file_i/_1423_ ;
 wire \register_file_i/_1424_ ;
 wire \register_file_i/_1425_ ;
 wire \register_file_i/_1426_ ;
 wire \register_file_i/_1427_ ;
 wire \register_file_i/_1428_ ;
 wire \register_file_i/_1429_ ;
 wire \register_file_i/_1430_ ;
 wire \register_file_i/_1431_ ;
 wire \register_file_i/_1432_ ;
 wire \register_file_i/_1433_ ;
 wire net348;
 wire \register_file_i/_1435_ ;
 wire \register_file_i/_1436_ ;
 wire \register_file_i/_1437_ ;
 wire \register_file_i/_1438_ ;
 wire \register_file_i/_1439_ ;
 wire net347;
 wire \register_file_i/_1441_ ;
 wire \register_file_i/_1442_ ;
 wire \register_file_i/_1443_ ;
 wire \register_file_i/_1444_ ;
 wire \register_file_i/_1445_ ;
 wire \register_file_i/_1446_ ;
 wire \register_file_i/_1447_ ;
 wire \register_file_i/_1448_ ;
 wire \register_file_i/_1449_ ;
 wire \register_file_i/_1450_ ;
 wire \register_file_i/_1451_ ;
 wire \register_file_i/_1452_ ;
 wire \register_file_i/_1453_ ;
 wire \register_file_i/_1454_ ;
 wire net346;
 wire \register_file_i/_1456_ ;
 wire \register_file_i/_1457_ ;
 wire \register_file_i/_1458_ ;
 wire \register_file_i/_1459_ ;
 wire \register_file_i/_1460_ ;
 wire \register_file_i/_1461_ ;
 wire \register_file_i/_1462_ ;
 wire \register_file_i/_1463_ ;
 wire \register_file_i/_1464_ ;
 wire \register_file_i/_1465_ ;
 wire \register_file_i/_1466_ ;
 wire net345;
 wire \register_file_i/_1468_ ;
 wire \register_file_i/_1469_ ;
 wire net344;
 wire \register_file_i/_1471_ ;
 wire \register_file_i/_1472_ ;
 wire \register_file_i/_1473_ ;
 wire \register_file_i/_1474_ ;
 wire \register_file_i/_1475_ ;
 wire \register_file_i/_1476_ ;
 wire \register_file_i/_1477_ ;
 wire \register_file_i/_1478_ ;
 wire \register_file_i/_1479_ ;
 wire \register_file_i/_1480_ ;
 wire \register_file_i/_1481_ ;
 wire \register_file_i/_1482_ ;
 wire \register_file_i/_1483_ ;
 wire \register_file_i/_1484_ ;
 wire \register_file_i/_1485_ ;
 wire \register_file_i/_1486_ ;
 wire \register_file_i/_1487_ ;
 wire \register_file_i/_1488_ ;
 wire \register_file_i/_1489_ ;
 wire \register_file_i/_1490_ ;
 wire \register_file_i/_1491_ ;
 wire net343;
 wire \register_file_i/_1493_ ;
 wire \register_file_i/_1494_ ;
 wire \register_file_i/_1495_ ;
 wire \register_file_i/_1496_ ;
 wire \register_file_i/_1497_ ;
 wire \register_file_i/_1498_ ;
 wire \register_file_i/_1499_ ;
 wire \register_file_i/_1500_ ;
 wire net342;
 wire \register_file_i/_1502_ ;
 wire \register_file_i/_1503_ ;
 wire \register_file_i/_1504_ ;
 wire \register_file_i/_1505_ ;
 wire \register_file_i/_1506_ ;
 wire \register_file_i/_1507_ ;
 wire \register_file_i/_1508_ ;
 wire \register_file_i/_1509_ ;
 wire \register_file_i/_1510_ ;
 wire net341;
 wire \register_file_i/_1512_ ;
 wire \register_file_i/_1513_ ;
 wire net340;
 wire \register_file_i/_1515_ ;
 wire \register_file_i/_1516_ ;
 wire \register_file_i/_1517_ ;
 wire \register_file_i/_1518_ ;
 wire \register_file_i/_1519_ ;
 wire \register_file_i/_1520_ ;
 wire \register_file_i/_1521_ ;
 wire \register_file_i/_1522_ ;
 wire \register_file_i/_1523_ ;
 wire net339;
 wire \register_file_i/_1525_ ;
 wire \register_file_i/_1526_ ;
 wire \register_file_i/_1527_ ;
 wire \register_file_i/_1528_ ;
 wire \register_file_i/_1529_ ;
 wire \register_file_i/_1530_ ;
 wire \register_file_i/_1531_ ;
 wire net338;
 wire \register_file_i/_1533_ ;
 wire \register_file_i/_1534_ ;
 wire \register_file_i/_1535_ ;
 wire \register_file_i/_1536_ ;
 wire \register_file_i/_1537_ ;
 wire \register_file_i/_1538_ ;
 wire \register_file_i/_1539_ ;
 wire \register_file_i/_1540_ ;
 wire \register_file_i/_1541_ ;
 wire \register_file_i/_1542_ ;
 wire net337;
 wire \register_file_i/_1544_ ;
 wire \register_file_i/_1545_ ;
 wire \register_file_i/_1546_ ;
 wire \register_file_i/_1547_ ;
 wire \register_file_i/_1548_ ;
 wire \register_file_i/_1549_ ;
 wire \register_file_i/_1550_ ;
 wire \register_file_i/_1551_ ;
 wire \register_file_i/_1552_ ;
 wire \register_file_i/_1553_ ;
 wire net336;
 wire \register_file_i/_1555_ ;
 wire \register_file_i/_1556_ ;
 wire \register_file_i/_1557_ ;
 wire \register_file_i/_1558_ ;
 wire \register_file_i/_1559_ ;
 wire \register_file_i/_1560_ ;
 wire \register_file_i/_1561_ ;
 wire \register_file_i/_1562_ ;
 wire \register_file_i/_1563_ ;
 wire \register_file_i/_1564_ ;
 wire \register_file_i/_1565_ ;
 wire \register_file_i/_1566_ ;
 wire \register_file_i/_1567_ ;
 wire net335;
 wire \register_file_i/_1569_ ;
 wire \register_file_i/_1570_ ;
 wire \register_file_i/_1571_ ;
 wire \register_file_i/_1572_ ;
 wire \register_file_i/_1573_ ;
 wire \register_file_i/_1574_ ;
 wire \register_file_i/_1575_ ;
 wire \register_file_i/_1576_ ;
 wire \register_file_i/_1577_ ;
 wire net334;
 wire net333;
 wire \register_file_i/_1580_ ;
 wire \register_file_i/_1581_ ;
 wire \register_file_i/_1582_ ;
 wire \register_file_i/_1583_ ;
 wire \register_file_i/_1584_ ;
 wire net332;
 wire \register_file_i/_1586_ ;
 wire \register_file_i/_1587_ ;
 wire net331;
 wire \register_file_i/_1589_ ;
 wire net330;
 wire \register_file_i/_1591_ ;
 wire \register_file_i/_1592_ ;
 wire net329;
 wire \register_file_i/_1594_ ;
 wire net328;
 wire \register_file_i/_1596_ ;
 wire net327;
 wire net326;
 wire \register_file_i/_1599_ ;
 wire \register_file_i/_1600_ ;
 wire \register_file_i/_1601_ ;
 wire \register_file_i/_1602_ ;
 wire \register_file_i/_1603_ ;
 wire \register_file_i/_1604_ ;
 wire \register_file_i/_1605_ ;
 wire net325;
 wire \register_file_i/_1607_ ;
 wire \register_file_i/_1608_ ;
 wire net324;
 wire \register_file_i/_1610_ ;
 wire \register_file_i/_1611_ ;
 wire \register_file_i/_1612_ ;
 wire \register_file_i/_1613_ ;
 wire \register_file_i/_1614_ ;
 wire \register_file_i/_1615_ ;
 wire \register_file_i/_1616_ ;
 wire \register_file_i/_1617_ ;
 wire \register_file_i/_1618_ ;
 wire \register_file_i/_1619_ ;
 wire \register_file_i/_1620_ ;
 wire net323;
 wire \register_file_i/_1622_ ;
 wire \register_file_i/_1623_ ;
 wire \register_file_i/_1624_ ;
 wire \register_file_i/_1625_ ;
 wire net322;
 wire \register_file_i/_1627_ ;
 wire \register_file_i/_1628_ ;
 wire \register_file_i/_1629_ ;
 wire \register_file_i/_1630_ ;
 wire \register_file_i/_1631_ ;
 wire \register_file_i/_1632_ ;
 wire \register_file_i/_1633_ ;
 wire \register_file_i/_1634_ ;
 wire \register_file_i/_1635_ ;
 wire \register_file_i/_1636_ ;
 wire net321;
 wire \register_file_i/_1638_ ;
 wire net320;
 wire \register_file_i/_1640_ ;
 wire \register_file_i/_1641_ ;
 wire \register_file_i/_1642_ ;
 wire \register_file_i/_1643_ ;
 wire \register_file_i/_1644_ ;
 wire \register_file_i/_1645_ ;
 wire \register_file_i/_1646_ ;
 wire \register_file_i/_1647_ ;
 wire \register_file_i/_1648_ ;
 wire \register_file_i/_1649_ ;
 wire \register_file_i/_1650_ ;
 wire \register_file_i/_1651_ ;
 wire \register_file_i/_1652_ ;
 wire \register_file_i/_1653_ ;
 wire \register_file_i/_1654_ ;
 wire \register_file_i/_1655_ ;
 wire \register_file_i/_1656_ ;
 wire \register_file_i/_1657_ ;
 wire \register_file_i/_1658_ ;
 wire \register_file_i/_1659_ ;
 wire \register_file_i/_1660_ ;
 wire \register_file_i/_1661_ ;
 wire \register_file_i/_1662_ ;
 wire \register_file_i/_1663_ ;
 wire \register_file_i/_1664_ ;
 wire \register_file_i/_1665_ ;
 wire \register_file_i/_1666_ ;
 wire \register_file_i/_1667_ ;
 wire \register_file_i/_1668_ ;
 wire \register_file_i/_1669_ ;
 wire \register_file_i/_1670_ ;
 wire \register_file_i/_1671_ ;
 wire \register_file_i/_1672_ ;
 wire \register_file_i/_1673_ ;
 wire \register_file_i/_1674_ ;
 wire \register_file_i/_1675_ ;
 wire \register_file_i/_1676_ ;
 wire \register_file_i/_1677_ ;
 wire \register_file_i/_1678_ ;
 wire \register_file_i/_1679_ ;
 wire \register_file_i/_1680_ ;
 wire \register_file_i/_1681_ ;
 wire \register_file_i/_1682_ ;
 wire \register_file_i/_1683_ ;
 wire \register_file_i/_1684_ ;
 wire \register_file_i/_1685_ ;
 wire \register_file_i/_1686_ ;
 wire \register_file_i/_1687_ ;
 wire \register_file_i/_1688_ ;
 wire \register_file_i/_1689_ ;
 wire \register_file_i/_1690_ ;
 wire \register_file_i/_1691_ ;
 wire \register_file_i/_1692_ ;
 wire \register_file_i/_1693_ ;
 wire \register_file_i/_1694_ ;
 wire \register_file_i/_1695_ ;
 wire \register_file_i/_1696_ ;
 wire \register_file_i/_1697_ ;
 wire \register_file_i/_1698_ ;
 wire \register_file_i/_1699_ ;
 wire \register_file_i/_1700_ ;
 wire \register_file_i/_1701_ ;
 wire \register_file_i/_1702_ ;
 wire \register_file_i/_1703_ ;
 wire \register_file_i/_1704_ ;
 wire \register_file_i/_1705_ ;
 wire \register_file_i/_1706_ ;
 wire \register_file_i/_1707_ ;
 wire \register_file_i/_1708_ ;
 wire \register_file_i/_1709_ ;
 wire \register_file_i/_1710_ ;
 wire \register_file_i/_1711_ ;
 wire \register_file_i/_1712_ ;
 wire \register_file_i/_1713_ ;
 wire \register_file_i/_1714_ ;
 wire \register_file_i/_1715_ ;
 wire \register_file_i/_1716_ ;
 wire \register_file_i/_1717_ ;
 wire \register_file_i/_1718_ ;
 wire \register_file_i/_1719_ ;
 wire \register_file_i/_1720_ ;
 wire \register_file_i/_1721_ ;
 wire \register_file_i/_1722_ ;
 wire \register_file_i/_1723_ ;
 wire \register_file_i/_1724_ ;
 wire \register_file_i/_1725_ ;
 wire \register_file_i/_1726_ ;
 wire \register_file_i/_1727_ ;
 wire \register_file_i/_1728_ ;
 wire \register_file_i/_1729_ ;
 wire \register_file_i/_1730_ ;
 wire \register_file_i/_1731_ ;
 wire \register_file_i/_1732_ ;
 wire \register_file_i/_1733_ ;
 wire \register_file_i/_1734_ ;
 wire \register_file_i/_1735_ ;
 wire \register_file_i/_1736_ ;
 wire \register_file_i/_1737_ ;
 wire \register_file_i/_1738_ ;
 wire \register_file_i/_1739_ ;
 wire \register_file_i/_1740_ ;
 wire \register_file_i/_1741_ ;
 wire \register_file_i/_1742_ ;
 wire \register_file_i/_1743_ ;
 wire \register_file_i/_1744_ ;
 wire \register_file_i/_1745_ ;
 wire \register_file_i/_1746_ ;
 wire \register_file_i/_1747_ ;
 wire \register_file_i/_1748_ ;
 wire \register_file_i/_1749_ ;
 wire \register_file_i/_1750_ ;
 wire \register_file_i/_1751_ ;
 wire \register_file_i/_1752_ ;
 wire \register_file_i/_1753_ ;
 wire \register_file_i/_1754_ ;
 wire \register_file_i/_1755_ ;
 wire \register_file_i/_1756_ ;
 wire \register_file_i/_1757_ ;
 wire \register_file_i/_1758_ ;
 wire \register_file_i/_1759_ ;
 wire \register_file_i/_1760_ ;
 wire \register_file_i/_1761_ ;
 wire \register_file_i/_1762_ ;
 wire \register_file_i/_1763_ ;
 wire \register_file_i/_1764_ ;
 wire \register_file_i/_1765_ ;
 wire \register_file_i/_1766_ ;
 wire \register_file_i/_1767_ ;
 wire \register_file_i/_1768_ ;
 wire \register_file_i/_1769_ ;
 wire \register_file_i/_1770_ ;
 wire \register_file_i/_1771_ ;
 wire \register_file_i/_1772_ ;
 wire \register_file_i/_1773_ ;
 wire \register_file_i/_1774_ ;
 wire \register_file_i/_1775_ ;
 wire \register_file_i/_1776_ ;
 wire \register_file_i/_1777_ ;
 wire \register_file_i/_1778_ ;
 wire \register_file_i/_1779_ ;
 wire \register_file_i/_1780_ ;
 wire \register_file_i/_1781_ ;
 wire \register_file_i/_1782_ ;
 wire \register_file_i/_1783_ ;
 wire \register_file_i/_1784_ ;
 wire \register_file_i/_1785_ ;
 wire \register_file_i/_1786_ ;
 wire \register_file_i/_1787_ ;
 wire \register_file_i/_1788_ ;
 wire \register_file_i/_1789_ ;
 wire \register_file_i/_1790_ ;
 wire \register_file_i/_1791_ ;
 wire \register_file_i/_1792_ ;
 wire \register_file_i/_1793_ ;
 wire \register_file_i/_1794_ ;
 wire \register_file_i/_1795_ ;
 wire \register_file_i/_1796_ ;
 wire \register_file_i/_1797_ ;
 wire \register_file_i/_1798_ ;
 wire \register_file_i/_1799_ ;
 wire \register_file_i/_1800_ ;
 wire \register_file_i/_1801_ ;
 wire \register_file_i/_1802_ ;
 wire \register_file_i/_1803_ ;
 wire \register_file_i/_1804_ ;
 wire \register_file_i/_1805_ ;
 wire \register_file_i/_1806_ ;
 wire \register_file_i/_1807_ ;
 wire \register_file_i/_1808_ ;
 wire \register_file_i/_1809_ ;
 wire \register_file_i/_1810_ ;
 wire \register_file_i/_1811_ ;
 wire \register_file_i/_1812_ ;
 wire \register_file_i/_1813_ ;
 wire \register_file_i/_1814_ ;
 wire \register_file_i/_1815_ ;
 wire \register_file_i/_1816_ ;
 wire \register_file_i/_1817_ ;
 wire \register_file_i/_1818_ ;
 wire \register_file_i/_1819_ ;
 wire \register_file_i/_1820_ ;
 wire \register_file_i/_1821_ ;
 wire \register_file_i/_1822_ ;
 wire \register_file_i/_1823_ ;
 wire \register_file_i/_1824_ ;
 wire \register_file_i/_1825_ ;
 wire \register_file_i/_1826_ ;
 wire \register_file_i/_1827_ ;
 wire \register_file_i/_1828_ ;
 wire \register_file_i/_1829_ ;
 wire \register_file_i/_1830_ ;
 wire \register_file_i/_1831_ ;
 wire \register_file_i/_1832_ ;
 wire \register_file_i/_1833_ ;
 wire \register_file_i/_1834_ ;
 wire \register_file_i/_1835_ ;
 wire \register_file_i/_1836_ ;
 wire \register_file_i/_1837_ ;
 wire \register_file_i/_1838_ ;
 wire \register_file_i/_1839_ ;
 wire \register_file_i/_1840_ ;
 wire \register_file_i/_1841_ ;
 wire \register_file_i/_1842_ ;
 wire \register_file_i/_1843_ ;
 wire \register_file_i/_1844_ ;
 wire \register_file_i/_1845_ ;
 wire \register_file_i/_1846_ ;
 wire \register_file_i/_1847_ ;
 wire \register_file_i/_1848_ ;
 wire \register_file_i/_1849_ ;
 wire \register_file_i/_1850_ ;
 wire \register_file_i/_1851_ ;
 wire \register_file_i/_1852_ ;
 wire \register_file_i/_1853_ ;
 wire \register_file_i/_1854_ ;
 wire \register_file_i/_1855_ ;
 wire \register_file_i/_1856_ ;
 wire \register_file_i/_1857_ ;
 wire \register_file_i/_1858_ ;
 wire \register_file_i/_1859_ ;
 wire \register_file_i/_1860_ ;
 wire \register_file_i/_1861_ ;
 wire \register_file_i/_1862_ ;
 wire \register_file_i/_1863_ ;
 wire \register_file_i/_1864_ ;
 wire \register_file_i/_1865_ ;
 wire \register_file_i/_1866_ ;
 wire \register_file_i/_1867_ ;
 wire \register_file_i/_1868_ ;
 wire \register_file_i/_1869_ ;
 wire \register_file_i/_1870_ ;
 wire \register_file_i/_1871_ ;
 wire \register_file_i/_1872_ ;
 wire \register_file_i/_1873_ ;
 wire \register_file_i/_1874_ ;
 wire \register_file_i/_1875_ ;
 wire \register_file_i/_1876_ ;
 wire \register_file_i/_1877_ ;
 wire \register_file_i/_1878_ ;
 wire \register_file_i/_1879_ ;
 wire \register_file_i/_1880_ ;
 wire \register_file_i/_1881_ ;
 wire \register_file_i/_1882_ ;
 wire \register_file_i/_1883_ ;
 wire \register_file_i/_1884_ ;
 wire \register_file_i/_1885_ ;
 wire \register_file_i/_1886_ ;
 wire \register_file_i/_1887_ ;
 wire \register_file_i/_1888_ ;
 wire \register_file_i/_1889_ ;
 wire \register_file_i/_1890_ ;
 wire \register_file_i/_1891_ ;
 wire \register_file_i/_1892_ ;
 wire \register_file_i/_1893_ ;
 wire net319;
 wire net318;
 wire \register_file_i/_1896_ ;
 wire net317;
 wire net316;
 wire net315;
 wire net314;
 wire net313;
 wire \register_file_i/_1902_ ;
 wire net312;
 wire \register_file_i/_1904_ ;
 wire \register_file_i/_1905_ ;
 wire net311;
 wire net310;
 wire net309;
 wire \register_file_i/_1909_ ;
 wire \register_file_i/_1910_ ;
 wire net308;
 wire net307;
 wire \register_file_i/_1913_ ;
 wire net306;
 wire \register_file_i/_1915_ ;
 wire \register_file_i/_1916_ ;
 wire net305;
 wire net304;
 wire \register_file_i/_1919_ ;
 wire \register_file_i/_1920_ ;
 wire net303;
 wire \register_file_i/_1922_ ;
 wire \register_file_i/_1923_ ;
 wire net302;
 wire net301;
 wire net300;
 wire net299;
 wire net298;
 wire \register_file_i/_1929_ ;
 wire net297;
 wire \register_file_i/_1931_ ;
 wire net296;
 wire \register_file_i/_1933_ ;
 wire net295;
 wire net294;
 wire \register_file_i/_1936_ ;
 wire net293;
 wire \register_file_i/_1938_ ;
 wire net292;
 wire \register_file_i/_1940_ ;
 wire \register_file_i/_1941_ ;
 wire \register_file_i/_1942_ ;
 wire \register_file_i/_1943_ ;
 wire \register_file_i/_1944_ ;
 wire net291;
 wire net290;
 wire net289;
 wire net288;
 wire \register_file_i/_1949_ ;
 wire \register_file_i/_1950_ ;
 wire \register_file_i/_1951_ ;
 wire net287;
 wire net286;
 wire \register_file_i/_1954_ ;
 wire net285;
 wire net284;
 wire \register_file_i/_1957_ ;
 wire net283;
 wire net282;
 wire \register_file_i/_1960_ ;
 wire \register_file_i/_1961_ ;
 wire net281;
 wire \register_file_i/_1963_ ;
 wire net280;
 wire \register_file_i/_1965_ ;
 wire net279;
 wire \register_file_i/_1967_ ;
 wire \register_file_i/_1968_ ;
 wire net278;
 wire \register_file_i/_1970_ ;
 wire \register_file_i/_1971_ ;
 wire \register_file_i/_1972_ ;
 wire \register_file_i/_1973_ ;
 wire \register_file_i/_1974_ ;
 wire net277;
 wire \register_file_i/_1976_ ;
 wire \register_file_i/_1977_ ;
 wire \register_file_i/_1978_ ;
 wire \register_file_i/_1979_ ;
 wire \register_file_i/_1980_ ;
 wire net276;
 wire \register_file_i/_1982_ ;
 wire \register_file_i/_1983_ ;
 wire \register_file_i/_1984_ ;
 wire \register_file_i/_1985_ ;
 wire \register_file_i/_1986_ ;
 wire \register_file_i/_1987_ ;
 wire \register_file_i/_1988_ ;
 wire net275;
 wire net274;
 wire \register_file_i/_1991_ ;
 wire net273;
 wire \register_file_i/_1993_ ;
 wire \register_file_i/_1994_ ;
 wire net272;
 wire \register_file_i/_1996_ ;
 wire net271;
 wire \register_file_i/_1998_ ;
 wire \register_file_i/_1999_ ;
 wire \register_file_i/_2000_ ;
 wire \register_file_i/_2001_ ;
 wire \register_file_i/_2002_ ;
 wire \register_file_i/_2003_ ;
 wire \register_file_i/_2004_ ;
 wire \register_file_i/_2005_ ;
 wire \register_file_i/_2006_ ;
 wire \register_file_i/_2007_ ;
 wire \register_file_i/_2008_ ;
 wire \register_file_i/_2009_ ;
 wire \register_file_i/_2010_ ;
 wire \register_file_i/_2011_ ;
 wire \register_file_i/_2012_ ;
 wire \register_file_i/_2013_ ;
 wire \register_file_i/_2014_ ;
 wire \register_file_i/_2015_ ;
 wire \register_file_i/_2016_ ;
 wire \register_file_i/_2017_ ;
 wire \register_file_i/_2018_ ;
 wire net270;
 wire \register_file_i/_2020_ ;
 wire \register_file_i/_2021_ ;
 wire \register_file_i/_2022_ ;
 wire \register_file_i/_2023_ ;
 wire \register_file_i/_2024_ ;
 wire \register_file_i/_2025_ ;
 wire \register_file_i/_2026_ ;
 wire \register_file_i/_2027_ ;
 wire net269;
 wire \register_file_i/_2029_ ;
 wire \register_file_i/_2030_ ;
 wire \register_file_i/_2031_ ;
 wire \register_file_i/_2032_ ;
 wire \register_file_i/_2033_ ;
 wire \register_file_i/_2034_ ;
 wire \register_file_i/_2035_ ;
 wire \register_file_i/_2036_ ;
 wire \register_file_i/_2037_ ;
 wire \register_file_i/_2038_ ;
 wire \register_file_i/_2039_ ;
 wire \register_file_i/_2040_ ;
 wire \register_file_i/_2041_ ;
 wire \register_file_i/_2042_ ;
 wire \register_file_i/_2043_ ;
 wire \register_file_i/_2044_ ;
 wire \register_file_i/_2045_ ;
 wire \register_file_i/_2046_ ;
 wire \register_file_i/_2047_ ;
 wire \register_file_i/_2048_ ;
 wire net268;
 wire \register_file_i/_2050_ ;
 wire \register_file_i/_2051_ ;
 wire \register_file_i/_2052_ ;
 wire \register_file_i/_2053_ ;
 wire \register_file_i/_2054_ ;
 wire \register_file_i/_2055_ ;
 wire \register_file_i/_2056_ ;
 wire \register_file_i/_2057_ ;
 wire \register_file_i/_2058_ ;
 wire \register_file_i/_2059_ ;
 wire \register_file_i/_2060_ ;
 wire \register_file_i/_2061_ ;
 wire \register_file_i/_2062_ ;
 wire net267;
 wire \register_file_i/_2064_ ;
 wire \register_file_i/_2065_ ;
 wire \register_file_i/_2066_ ;
 wire \register_file_i/_2067_ ;
 wire \register_file_i/_2068_ ;
 wire net266;
 wire \register_file_i/_2070_ ;
 wire \register_file_i/_2071_ ;
 wire \register_file_i/_2072_ ;
 wire \register_file_i/_2073_ ;
 wire \register_file_i/_2074_ ;
 wire \register_file_i/_2075_ ;
 wire \register_file_i/_2076_ ;
 wire \register_file_i/_2077_ ;
 wire \register_file_i/_2078_ ;
 wire \register_file_i/_2079_ ;
 wire \register_file_i/_2080_ ;
 wire \register_file_i/_2081_ ;
 wire \register_file_i/_2082_ ;
 wire \register_file_i/_2083_ ;
 wire net265;
 wire \register_file_i/_2085_ ;
 wire \register_file_i/_2086_ ;
 wire \register_file_i/_2087_ ;
 wire \register_file_i/_2088_ ;
 wire \register_file_i/_2089_ ;
 wire \register_file_i/_2090_ ;
 wire \register_file_i/_2091_ ;
 wire \register_file_i/_2092_ ;
 wire \register_file_i/_2093_ ;
 wire \register_file_i/_2094_ ;
 wire \register_file_i/_2095_ ;
 wire net264;
 wire \register_file_i/_2097_ ;
 wire \register_file_i/_2098_ ;
 wire net263;
 wire \register_file_i/_2100_ ;
 wire \register_file_i/_2101_ ;
 wire \register_file_i/_2102_ ;
 wire \register_file_i/_2103_ ;
 wire \register_file_i/_2104_ ;
 wire \register_file_i/_2105_ ;
 wire \register_file_i/_2106_ ;
 wire \register_file_i/_2107_ ;
 wire \register_file_i/_2108_ ;
 wire \register_file_i/_2109_ ;
 wire \register_file_i/_2110_ ;
 wire \register_file_i/_2111_ ;
 wire \register_file_i/_2112_ ;
 wire \register_file_i/_2113_ ;
 wire \register_file_i/_2114_ ;
 wire \register_file_i/_2115_ ;
 wire \register_file_i/_2116_ ;
 wire \register_file_i/_2117_ ;
 wire \register_file_i/_2118_ ;
 wire \register_file_i/_2119_ ;
 wire \register_file_i/_2120_ ;
 wire net262;
 wire \register_file_i/_2122_ ;
 wire \register_file_i/_2123_ ;
 wire \register_file_i/_2124_ ;
 wire \register_file_i/_2125_ ;
 wire \register_file_i/_2126_ ;
 wire \register_file_i/_2127_ ;
 wire \register_file_i/_2128_ ;
 wire \register_file_i/_2129_ ;
 wire net261;
 wire \register_file_i/_2131_ ;
 wire \register_file_i/_2132_ ;
 wire \register_file_i/_2133_ ;
 wire \register_file_i/_2134_ ;
 wire \register_file_i/_2135_ ;
 wire \register_file_i/_2136_ ;
 wire \register_file_i/_2137_ ;
 wire \register_file_i/_2138_ ;
 wire \register_file_i/_2139_ ;
 wire net260;
 wire \register_file_i/_2141_ ;
 wire \register_file_i/_2142_ ;
 wire net259;
 wire \register_file_i/_2144_ ;
 wire \register_file_i/_2145_ ;
 wire \register_file_i/_2146_ ;
 wire \register_file_i/_2147_ ;
 wire \register_file_i/_2148_ ;
 wire \register_file_i/_2149_ ;
 wire \register_file_i/_2150_ ;
 wire \register_file_i/_2151_ ;
 wire \register_file_i/_2152_ ;
 wire net258;
 wire \register_file_i/_2154_ ;
 wire \register_file_i/_2155_ ;
 wire \register_file_i/_2156_ ;
 wire \register_file_i/_2157_ ;
 wire \register_file_i/_2158_ ;
 wire \register_file_i/_2159_ ;
 wire \register_file_i/_2160_ ;
 wire net257;
 wire \register_file_i/_2162_ ;
 wire \register_file_i/_2163_ ;
 wire \register_file_i/_2164_ ;
 wire \register_file_i/_2165_ ;
 wire \register_file_i/_2166_ ;
 wire \register_file_i/_2167_ ;
 wire \register_file_i/_2168_ ;
 wire \register_file_i/_2169_ ;
 wire \register_file_i/_2170_ ;
 wire \register_file_i/_2171_ ;
 wire net256;
 wire \register_file_i/_2173_ ;
 wire \register_file_i/_2174_ ;
 wire \register_file_i/_2175_ ;
 wire \register_file_i/_2176_ ;
 wire \register_file_i/_2177_ ;
 wire \register_file_i/_2178_ ;
 wire \register_file_i/_2179_ ;
 wire \register_file_i/_2180_ ;
 wire \register_file_i/_2181_ ;
 wire \register_file_i/_2182_ ;
 wire net255;
 wire \register_file_i/_2184_ ;
 wire \register_file_i/_2185_ ;
 wire \register_file_i/_2186_ ;
 wire \register_file_i/_2187_ ;
 wire \register_file_i/_2188_ ;
 wire \register_file_i/_2189_ ;
 wire \register_file_i/_2190_ ;
 wire \register_file_i/_2191_ ;
 wire \register_file_i/_2192_ ;
 wire \register_file_i/_2193_ ;
 wire \register_file_i/_2194_ ;
 wire \register_file_i/_2195_ ;
 wire \register_file_i/_2196_ ;
 wire net254;
 wire \register_file_i/_2198_ ;
 wire \register_file_i/_2199_ ;
 wire \register_file_i/_2200_ ;
 wire \register_file_i/_2201_ ;
 wire \register_file_i/_2202_ ;
 wire \register_file_i/_2203_ ;
 wire \register_file_i/_2204_ ;
 wire \register_file_i/_2205_ ;
 wire \register_file_i/_2206_ ;
 wire net253;
 wire net252;
 wire \register_file_i/_2209_ ;
 wire \register_file_i/_2210_ ;
 wire \register_file_i/_2211_ ;
 wire \register_file_i/_2212_ ;
 wire \register_file_i/_2213_ ;
 wire net251;
 wire \register_file_i/_2215_ ;
 wire \register_file_i/_2216_ ;
 wire net250;
 wire \register_file_i/_2218_ ;
 wire net249;
 wire \register_file_i/_2220_ ;
 wire \register_file_i/_2221_ ;
 wire net248;
 wire \register_file_i/_2223_ ;
 wire net247;
 wire \register_file_i/_2225_ ;
 wire net246;
 wire net245;
 wire net244;
 wire \register_file_i/_2229_ ;
 wire \register_file_i/_2230_ ;
 wire \register_file_i/_2231_ ;
 wire \register_file_i/_2232_ ;
 wire \register_file_i/_2233_ ;
 wire \register_file_i/_2234_ ;
 wire \register_file_i/_2235_ ;
 wire net243;
 wire \register_file_i/_2237_ ;
 wire \register_file_i/_2238_ ;
 wire net242;
 wire \register_file_i/_2240_ ;
 wire \register_file_i/_2241_ ;
 wire \register_file_i/_2242_ ;
 wire \register_file_i/_2243_ ;
 wire \register_file_i/_2244_ ;
 wire \register_file_i/_2245_ ;
 wire \register_file_i/_2246_ ;
 wire \register_file_i/_2247_ ;
 wire \register_file_i/_2248_ ;
 wire \register_file_i/_2249_ ;
 wire \register_file_i/_2250_ ;
 wire net241;
 wire \register_file_i/_2252_ ;
 wire \register_file_i/_2253_ ;
 wire \register_file_i/_2254_ ;
 wire \register_file_i/_2255_ ;
 wire \register_file_i/_2256_ ;
 wire net240;
 wire \register_file_i/_2258_ ;
 wire \register_file_i/_2259_ ;
 wire \register_file_i/_2260_ ;
 wire \register_file_i/_2261_ ;
 wire \register_file_i/_2262_ ;
 wire \register_file_i/_2263_ ;
 wire \register_file_i/_2264_ ;
 wire net239;
 wire \register_file_i/_2266_ ;
 wire net238;
 wire \register_file_i/_2268_ ;
 wire \register_file_i/_2269_ ;
 wire \register_file_i/_2270_ ;
 wire \register_file_i/_2271_ ;
 wire \register_file_i/_2272_ ;
 wire \register_file_i/_2273_ ;
 wire \register_file_i/_2274_ ;
 wire \register_file_i/_2275_ ;
 wire \register_file_i/_2276_ ;
 wire \register_file_i/_2277_ ;
 wire \register_file_i/_2278_ ;
 wire \register_file_i/_2279_ ;
 wire \register_file_i/_2280_ ;
 wire \register_file_i/_2281_ ;
 wire \register_file_i/_2282_ ;
 wire \register_file_i/_2283_ ;
 wire \register_file_i/_2284_ ;
 wire \register_file_i/_2285_ ;
 wire \register_file_i/_2286_ ;
 wire \register_file_i/_2287_ ;
 wire \register_file_i/_2288_ ;
 wire \register_file_i/_2289_ ;
 wire \register_file_i/_2290_ ;
 wire \register_file_i/_2291_ ;
 wire net237;
 wire \register_file_i/_2293_ ;
 wire \register_file_i/_2294_ ;
 wire \register_file_i/_2295_ ;
 wire \register_file_i/_2296_ ;
 wire \register_file_i/_2297_ ;
 wire \register_file_i/_2298_ ;
 wire \register_file_i/_2299_ ;
 wire \register_file_i/_2300_ ;
 wire net236;
 wire \register_file_i/_2302_ ;
 wire \register_file_i/_2303_ ;
 wire \register_file_i/_2304_ ;
 wire \register_file_i/_2305_ ;
 wire \register_file_i/_2306_ ;
 wire \register_file_i/_2307_ ;
 wire \register_file_i/_2308_ ;
 wire \register_file_i/_2309_ ;
 wire \register_file_i/_2310_ ;
 wire \register_file_i/_2311_ ;
 wire \register_file_i/_2312_ ;
 wire \register_file_i/_2313_ ;
 wire \register_file_i/_2314_ ;
 wire \register_file_i/_2315_ ;
 wire \register_file_i/_2316_ ;
 wire \register_file_i/_2317_ ;
 wire \register_file_i/_2318_ ;
 wire \register_file_i/_2319_ ;
 wire \register_file_i/_2320_ ;
 wire \register_file_i/_2321_ ;
 wire net235;
 wire \register_file_i/_2323_ ;
 wire \register_file_i/_2324_ ;
 wire \register_file_i/_2325_ ;
 wire \register_file_i/_2326_ ;
 wire \register_file_i/_2327_ ;
 wire \register_file_i/_2328_ ;
 wire \register_file_i/_2329_ ;
 wire \register_file_i/_2330_ ;
 wire \register_file_i/_2331_ ;
 wire \register_file_i/_2332_ ;
 wire \register_file_i/_2333_ ;
 wire \register_file_i/_2334_ ;
 wire \register_file_i/_2335_ ;
 wire net234;
 wire \register_file_i/_2337_ ;
 wire \register_file_i/_2338_ ;
 wire \register_file_i/_2339_ ;
 wire \register_file_i/_2340_ ;
 wire \register_file_i/_2341_ ;
 wire net233;
 wire \register_file_i/_2343_ ;
 wire \register_file_i/_2344_ ;
 wire \register_file_i/_2345_ ;
 wire \register_file_i/_2346_ ;
 wire \register_file_i/_2347_ ;
 wire \register_file_i/_2348_ ;
 wire \register_file_i/_2349_ ;
 wire \register_file_i/_2350_ ;
 wire \register_file_i/_2351_ ;
 wire \register_file_i/_2352_ ;
 wire \register_file_i/_2353_ ;
 wire \register_file_i/_2354_ ;
 wire \register_file_i/_2355_ ;
 wire \register_file_i/_2356_ ;
 wire net232;
 wire \register_file_i/_2358_ ;
 wire \register_file_i/_2359_ ;
 wire \register_file_i/_2360_ ;
 wire \register_file_i/_2361_ ;
 wire \register_file_i/_2362_ ;
 wire \register_file_i/_2363_ ;
 wire \register_file_i/_2364_ ;
 wire \register_file_i/_2365_ ;
 wire \register_file_i/_2366_ ;
 wire \register_file_i/_2367_ ;
 wire \register_file_i/_2368_ ;
 wire net231;
 wire \register_file_i/_2370_ ;
 wire \register_file_i/_2371_ ;
 wire net230;
 wire \register_file_i/_2373_ ;
 wire \register_file_i/_2374_ ;
 wire \register_file_i/_2375_ ;
 wire \register_file_i/_2376_ ;
 wire \register_file_i/_2377_ ;
 wire \register_file_i/_2378_ ;
 wire \register_file_i/_2379_ ;
 wire \register_file_i/_2380_ ;
 wire \register_file_i/_2381_ ;
 wire \register_file_i/_2382_ ;
 wire \register_file_i/_2383_ ;
 wire \register_file_i/_2384_ ;
 wire \register_file_i/_2385_ ;
 wire \register_file_i/_2386_ ;
 wire \register_file_i/_2387_ ;
 wire \register_file_i/_2388_ ;
 wire \register_file_i/_2389_ ;
 wire \register_file_i/_2390_ ;
 wire \register_file_i/_2391_ ;
 wire \register_file_i/_2392_ ;
 wire \register_file_i/_2393_ ;
 wire net229;
 wire \register_file_i/_2395_ ;
 wire \register_file_i/_2396_ ;
 wire \register_file_i/_2397_ ;
 wire \register_file_i/_2398_ ;
 wire \register_file_i/_2399_ ;
 wire \register_file_i/_2400_ ;
 wire \register_file_i/_2401_ ;
 wire \register_file_i/_2402_ ;
 wire net228;
 wire \register_file_i/_2404_ ;
 wire \register_file_i/_2405_ ;
 wire \register_file_i/_2406_ ;
 wire \register_file_i/_2407_ ;
 wire \register_file_i/_2408_ ;
 wire \register_file_i/_2409_ ;
 wire \register_file_i/_2410_ ;
 wire \register_file_i/_2411_ ;
 wire \register_file_i/_2412_ ;
 wire net227;
 wire \register_file_i/_2414_ ;
 wire \register_file_i/_2415_ ;
 wire net226;
 wire \register_file_i/_2417_ ;
 wire \register_file_i/_2418_ ;
 wire \register_file_i/_2419_ ;
 wire \register_file_i/_2420_ ;
 wire \register_file_i/_2421_ ;
 wire \register_file_i/_2422_ ;
 wire \register_file_i/_2423_ ;
 wire \register_file_i/_2424_ ;
 wire \register_file_i/_2425_ ;
 wire net225;
 wire \register_file_i/_2427_ ;
 wire \register_file_i/_2428_ ;
 wire \register_file_i/_2429_ ;
 wire \register_file_i/_2430_ ;
 wire \register_file_i/_2431_ ;
 wire \register_file_i/_2432_ ;
 wire \register_file_i/_2433_ ;
 wire net224;
 wire \register_file_i/_2435_ ;
 wire \register_file_i/_2436_ ;
 wire \register_file_i/_2437_ ;
 wire \register_file_i/_2438_ ;
 wire \register_file_i/_2439_ ;
 wire \register_file_i/_2440_ ;
 wire \register_file_i/_2441_ ;
 wire \register_file_i/_2442_ ;
 wire \register_file_i/_2443_ ;
 wire \register_file_i/_2444_ ;
 wire net223;
 wire \register_file_i/_2446_ ;
 wire \register_file_i/_2447_ ;
 wire \register_file_i/_2448_ ;
 wire \register_file_i/_2449_ ;
 wire \register_file_i/_2450_ ;
 wire \register_file_i/_2451_ ;
 wire \register_file_i/_2452_ ;
 wire \register_file_i/_2453_ ;
 wire \register_file_i/_2454_ ;
 wire \register_file_i/_2455_ ;
 wire net222;
 wire \register_file_i/_2457_ ;
 wire \register_file_i/_2458_ ;
 wire \register_file_i/_2459_ ;
 wire \register_file_i/_2460_ ;
 wire \register_file_i/_2461_ ;
 wire \register_file_i/_2462_ ;
 wire \register_file_i/_2463_ ;
 wire \register_file_i/_2464_ ;
 wire \register_file_i/_2465_ ;
 wire \register_file_i/_2466_ ;
 wire \register_file_i/_2467_ ;
 wire \register_file_i/_2468_ ;
 wire \register_file_i/_2469_ ;
 wire net221;
 wire \register_file_i/_2471_ ;
 wire \register_file_i/_2472_ ;
 wire \register_file_i/_2473_ ;
 wire \register_file_i/_2474_ ;
 wire \register_file_i/_2475_ ;
 wire \register_file_i/_2476_ ;
 wire \register_file_i/_2477_ ;
 wire \register_file_i/_2478_ ;
 wire \register_file_i/_2479_ ;
 wire net220;
 wire net219;
 wire \register_file_i/_2482_ ;
 wire \register_file_i/_2483_ ;
 wire \register_file_i/_2484_ ;
 wire \register_file_i/_2485_ ;
 wire \register_file_i/_2486_ ;
 wire net218;
 wire \register_file_i/_2488_ ;
 wire \register_file_i/_2489_ ;
 wire net217;
 wire \register_file_i/_2491_ ;
 wire net216;
 wire \register_file_i/_2493_ ;
 wire \register_file_i/_2494_ ;
 wire net215;
 wire \register_file_i/_2496_ ;
 wire net214;
 wire \register_file_i/_2498_ ;
 wire net213;
 wire net212;
 wire \register_file_i/_2501_ ;
 wire \register_file_i/_2502_ ;
 wire \register_file_i/_2503_ ;
 wire \register_file_i/_2504_ ;
 wire \register_file_i/_2505_ ;
 wire \register_file_i/_2506_ ;
 wire \register_file_i/_2507_ ;
 wire net211;
 wire \register_file_i/_2509_ ;
 wire \register_file_i/_2510_ ;
 wire net210;
 wire \register_file_i/_2512_ ;
 wire \register_file_i/_2513_ ;
 wire \register_file_i/_2514_ ;
 wire \register_file_i/_2515_ ;
 wire \register_file_i/_2516_ ;
 wire \register_file_i/_2517_ ;
 wire \register_file_i/_2518_ ;
 wire \register_file_i/_2519_ ;
 wire \register_file_i/_2520_ ;
 wire \register_file_i/_2521_ ;
 wire \register_file_i/_2522_ ;
 wire net209;
 wire \register_file_i/_2524_ ;
 wire \register_file_i/_2525_ ;
 wire \register_file_i/_2526_ ;
 wire \register_file_i/_2527_ ;
 wire net208;
 wire \register_file_i/_2529_ ;
 wire \register_file_i/_2530_ ;
 wire \register_file_i/_2531_ ;
 wire \register_file_i/_2532_ ;
 wire \register_file_i/_2533_ ;
 wire \register_file_i/_2534_ ;
 wire \register_file_i/_2535_ ;
 wire \register_file_i/_2536_ ;
 wire \register_file_i/_2537_ ;
 wire \register_file_i/_2538_ ;
 wire net207;
 wire \register_file_i/_2540_ ;
 wire net206;
 wire \register_file_i/_2542_ ;
 wire \register_file_i/_2543_ ;
 wire \register_file_i/_2544_ ;
 wire \register_file_i/_2545_ ;
 wire \register_file_i/_2546_ ;
 wire \register_file_i/_2547_ ;
 wire \register_file_i/_2548_ ;
 wire \register_file_i/_2549_ ;
 wire \register_file_i/_2550_ ;
 wire \register_file_i/_2551_ ;
 wire \register_file_i/_2552_ ;
 wire \register_file_i/_2553_ ;
 wire \register_file_i/_2554_ ;
 wire \register_file_i/_2555_ ;
 wire \register_file_i/_2556_ ;
 wire \register_file_i/_2557_ ;
 wire \register_file_i/_2558_ ;
 wire \register_file_i/_2559_ ;
 wire \register_file_i/_2560_ ;
 wire \register_file_i/_2561_ ;
 wire \register_file_i/_2562_ ;
 wire \register_file_i/_2563_ ;
 wire \register_file_i/_2564_ ;
 wire \register_file_i/_2565_ ;
 wire \register_file_i/_2566_ ;
 wire \register_file_i/_2567_ ;
 wire \register_file_i/_2568_ ;
 wire \register_file_i/_2569_ ;
 wire \register_file_i/_2570_ ;
 wire \register_file_i/_2571_ ;
 wire \register_file_i/_2572_ ;
 wire \register_file_i/_2573_ ;
 wire \register_file_i/_2574_ ;
 wire \register_file_i/_2575_ ;
 wire \register_file_i/_2576_ ;
 wire \register_file_i/_2577_ ;
 wire \register_file_i/_2578_ ;
 wire \register_file_i/_2579_ ;
 wire \register_file_i/_2580_ ;
 wire \register_file_i/_2581_ ;
 wire \register_file_i/_2582_ ;
 wire \register_file_i/_2583_ ;
 wire \register_file_i/_2584_ ;
 wire \register_file_i/_2585_ ;
 wire \register_file_i/_2586_ ;
 wire \register_file_i/_2587_ ;
 wire \register_file_i/_2588_ ;
 wire \register_file_i/_2589_ ;
 wire \register_file_i/_2590_ ;
 wire \register_file_i/_2591_ ;
 wire \register_file_i/_2592_ ;
 wire \register_file_i/_2593_ ;
 wire \register_file_i/_2594_ ;
 wire \register_file_i/_2595_ ;
 wire \register_file_i/_2596_ ;
 wire \register_file_i/_2597_ ;
 wire \register_file_i/_2598_ ;
 wire \register_file_i/_2599_ ;
 wire \register_file_i/_2600_ ;
 wire \register_file_i/_2601_ ;
 wire \register_file_i/_2602_ ;
 wire \register_file_i/_2603_ ;
 wire \register_file_i/_2604_ ;
 wire \register_file_i/_2605_ ;
 wire \register_file_i/_2606_ ;
 wire \register_file_i/_2607_ ;
 wire \register_file_i/_2608_ ;
 wire \register_file_i/_2609_ ;
 wire \register_file_i/_2610_ ;
 wire \register_file_i/_2611_ ;
 wire \register_file_i/_2612_ ;
 wire \register_file_i/_2613_ ;
 wire \register_file_i/_2614_ ;
 wire \register_file_i/_2615_ ;
 wire \register_file_i/_2616_ ;
 wire \register_file_i/_2617_ ;
 wire \register_file_i/_2618_ ;
 wire \register_file_i/_2619_ ;
 wire \register_file_i/_2620_ ;
 wire \register_file_i/_2621_ ;
 wire \register_file_i/_2622_ ;
 wire \register_file_i/_2623_ ;
 wire \register_file_i/_2624_ ;
 wire \register_file_i/_2625_ ;
 wire \register_file_i/_2626_ ;
 wire \register_file_i/_2627_ ;
 wire \register_file_i/_2628_ ;
 wire \register_file_i/_2629_ ;
 wire \register_file_i/_2630_ ;
 wire \register_file_i/_2631_ ;
 wire \register_file_i/_2632_ ;
 wire \register_file_i/_2633_ ;
 wire \register_file_i/_2634_ ;
 wire \register_file_i/_2635_ ;
 wire \register_file_i/_2636_ ;
 wire \register_file_i/_2637_ ;
 wire \register_file_i/_2638_ ;
 wire \register_file_i/_2639_ ;
 wire \register_file_i/_2640_ ;
 wire \register_file_i/_2641_ ;
 wire \register_file_i/_2642_ ;
 wire \register_file_i/_2643_ ;
 wire \register_file_i/_2644_ ;
 wire \register_file_i/_2645_ ;
 wire \register_file_i/_2646_ ;
 wire \register_file_i/_2647_ ;
 wire \register_file_i/_2648_ ;
 wire \register_file_i/_2649_ ;
 wire \register_file_i/_2650_ ;
 wire \register_file_i/_2651_ ;
 wire \register_file_i/_2652_ ;
 wire \register_file_i/_2653_ ;
 wire \register_file_i/_2654_ ;
 wire \register_file_i/_2655_ ;
 wire \register_file_i/_2656_ ;
 wire \register_file_i/_2657_ ;
 wire \register_file_i/_2658_ ;
 wire \register_file_i/_2659_ ;
 wire \register_file_i/_2660_ ;
 wire \register_file_i/_2661_ ;
 wire \register_file_i/_2662_ ;
 wire \register_file_i/_2663_ ;
 wire \register_file_i/_2664_ ;
 wire \register_file_i/_2665_ ;
 wire \register_file_i/_2666_ ;
 wire \register_file_i/_2667_ ;
 wire \register_file_i/_2668_ ;
 wire \register_file_i/_2669_ ;
 wire \register_file_i/_2670_ ;
 wire \register_file_i/_2671_ ;
 wire \register_file_i/_2672_ ;
 wire \register_file_i/_2673_ ;
 wire \register_file_i/_2674_ ;
 wire \register_file_i/_2675_ ;
 wire \register_file_i/_2676_ ;
 wire \register_file_i/_2677_ ;
 wire \register_file_i/_2678_ ;
 wire \register_file_i/_2679_ ;
 wire \register_file_i/_2680_ ;
 wire \register_file_i/_2681_ ;
 wire \register_file_i/_2682_ ;
 wire \register_file_i/_2683_ ;
 wire \register_file_i/_2684_ ;
 wire \register_file_i/_2685_ ;
 wire \register_file_i/_2686_ ;
 wire \register_file_i/_2687_ ;
 wire \register_file_i/_2688_ ;
 wire \register_file_i/_2689_ ;
 wire \register_file_i/_2690_ ;
 wire \register_file_i/_2691_ ;
 wire \register_file_i/_2692_ ;
 wire \register_file_i/_2693_ ;
 wire \register_file_i/_2694_ ;
 wire \register_file_i/_2695_ ;
 wire \register_file_i/_2696_ ;
 wire \register_file_i/_2697_ ;
 wire \register_file_i/_2698_ ;
 wire \register_file_i/_2699_ ;
 wire \register_file_i/_2700_ ;
 wire \register_file_i/_2701_ ;
 wire \register_file_i/_2702_ ;
 wire \register_file_i/_2703_ ;
 wire \register_file_i/_2704_ ;
 wire \register_file_i/_2705_ ;
 wire \register_file_i/_2706_ ;
 wire \register_file_i/_2707_ ;
 wire \register_file_i/_2708_ ;
 wire \register_file_i/_2709_ ;
 wire \register_file_i/_2710_ ;
 wire \register_file_i/_2711_ ;
 wire \register_file_i/_2712_ ;
 wire \register_file_i/_2713_ ;
 wire \register_file_i/_2714_ ;
 wire \register_file_i/_2715_ ;
 wire \register_file_i/_2716_ ;
 wire \register_file_i/_2717_ ;
 wire \register_file_i/_2718_ ;
 wire \register_file_i/_2719_ ;
 wire \register_file_i/_2720_ ;
 wire \register_file_i/_2721_ ;
 wire \register_file_i/_2722_ ;
 wire \register_file_i/_2723_ ;
 wire \register_file_i/_2724_ ;
 wire \register_file_i/_2725_ ;
 wire \register_file_i/_2726_ ;
 wire \register_file_i/_2727_ ;
 wire \register_file_i/_2728_ ;
 wire \register_file_i/_2729_ ;
 wire \register_file_i/_2730_ ;
 wire \register_file_i/_2731_ ;
 wire \register_file_i/_2732_ ;
 wire \register_file_i/_2733_ ;
 wire \register_file_i/_2734_ ;
 wire \register_file_i/_2735_ ;
 wire \register_file_i/_2736_ ;
 wire \register_file_i/_2737_ ;
 wire \register_file_i/_2738_ ;
 wire \register_file_i/_2739_ ;
 wire \register_file_i/_2740_ ;
 wire \register_file_i/_2741_ ;
 wire \register_file_i/_2742_ ;
 wire \register_file_i/_2743_ ;
 wire \register_file_i/_2744_ ;
 wire \register_file_i/_2745_ ;
 wire \register_file_i/_2746_ ;
 wire \register_file_i/_2747_ ;
 wire \register_file_i/_2748_ ;
 wire \register_file_i/_2749_ ;
 wire \register_file_i/_2750_ ;
 wire \register_file_i/_2751_ ;
 wire \register_file_i/_2752_ ;
 wire \register_file_i/_2753_ ;
 wire \register_file_i/_2754_ ;
 wire \register_file_i/_2755_ ;
 wire \register_file_i/_2756_ ;
 wire \register_file_i/_2757_ ;
 wire \register_file_i/_2758_ ;
 wire \register_file_i/_2759_ ;
 wire \register_file_i/_2760_ ;
 wire \register_file_i/_2761_ ;
 wire \register_file_i/_2762_ ;
 wire \register_file_i/_2763_ ;
 wire \register_file_i/_2764_ ;
 wire \register_file_i/_2765_ ;
 wire \register_file_i/_2766_ ;
 wire \register_file_i/_2767_ ;
 wire \register_file_i/_2768_ ;
 wire \register_file_i/_2769_ ;
 wire \register_file_i/_2770_ ;
 wire \register_file_i/_2771_ ;
 wire \register_file_i/_2772_ ;
 wire \register_file_i/_2773_ ;
 wire \register_file_i/_2774_ ;
 wire \register_file_i/_2775_ ;
 wire \register_file_i/_2776_ ;
 wire \register_file_i/_2777_ ;
 wire \register_file_i/_2778_ ;
 wire \register_file_i/_2779_ ;
 wire \register_file_i/_2780_ ;
 wire \register_file_i/_2781_ ;
 wire \register_file_i/_2782_ ;
 wire \register_file_i/_2783_ ;
 wire \register_file_i/_2784_ ;
 wire \register_file_i/_2785_ ;
 wire \register_file_i/_2786_ ;
 wire \register_file_i/_2787_ ;
 wire \register_file_i/_2788_ ;
 wire \register_file_i/_2789_ ;
 wire \register_file_i/_2790_ ;
 wire \register_file_i/_2791_ ;
 wire \register_file_i/_2792_ ;
 wire \register_file_i/_2793_ ;
 wire \register_file_i/_2794_ ;
 wire \register_file_i/_2795_ ;
 wire net205;
 wire net204;
 wire net203;
 wire \register_file_i/_2799_ ;
 wire \register_file_i/_2800_ ;
 wire \register_file_i/_2801_ ;
 wire net202;
 wire net201;
 wire net200;
 wire net199;
 wire net198;
 wire net197;
 wire net196;
 wire net195;
 wire net194;
 wire net193;
 wire net192;
 wire \register_file_i/_2813_ ;
 wire \register_file_i/_2814_ ;
 wire \register_file_i/_2815_ ;
 wire \register_file_i/_2816_ ;
 wire \register_file_i/_2817_ ;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire net173;
 wire net172;
 wire net171;
 wire net170;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire net162;
 wire net161;
 wire net160;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net155;
 wire net154;
 wire net153;
 wire net152;
 wire net151;
 wire net150;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire net144;
 wire \register_file_i/_2866_ ;
 wire \register_file_i/_2867_ ;
 wire \register_file_i/_2868_ ;
 wire \register_file_i/_2869_ ;
 wire \register_file_i/_2870_ ;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire \register_file_i/_2877_ ;
 wire \register_file_i/_2878_ ;
 wire \register_file_i/_2879_ ;
 wire net137;
 wire net136;
 wire net135;
 wire \register_file_i/_2883_ ;
 wire \register_file_i/_2884_ ;
 wire \register_file_i/_2885_ ;
 wire net134;
 wire net133;
 wire net132;
 wire net131;
 wire \register_file_i/_2890_ ;
 wire net130;
 wire net129;
 wire net128;
 wire net127;
 wire net126;
 wire net125;
 wire net124;
 wire net123;
 wire net122;
 wire net121;
 wire \register_file_i/_2901_ ;
 wire \register_file_i/_2902_ ;
 wire \register_file_i/_2903_ ;
 wire net120;
 wire net119;
 wire net118;
 wire \register_file_i/_2907_ ;
 wire net117;
 wire net116;
 wire net115;
 wire \register_file_i/_2911_ ;
 wire net114;
 wire \register_file_i/_2913_ ;
 wire net113;
 wire net112;
 wire net111;
 wire \register_file_i/_2917_ ;
 wire net110;
 wire net109;
 wire net108;
 wire \register_file_i/_2921_ ;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire \register_file_i/_2926_ ;
 wire \register_file_i/_2927_ ;
 wire net103;
 wire net102;
 wire net101;
 wire net100;
 wire \register_file_i/_2932_ ;
 wire net99;
 wire net98;
 wire net97;
 wire \register_file_i/_2936_ ;
 wire net96;
 wire net95;
 wire net94;
 wire \register_file_i/_2940_ ;
 wire \register_file_i/_2941_ ;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire \register_file_i/_2946_ ;
 wire \register_file_i/_2947_ ;
 wire net89;
 wire net88;
 wire net87;
 wire \register_file_i/_2951_ ;
 wire \register_file_i/_2952_ ;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire \register_file_i/_2981_ ;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire \register_file_i/_2992_ ;
 wire net48;
 wire net47;
 wire \register_file_i/_2995_ ;
 wire net46;
 wire net45;
 wire net44;
 wire \register_file_i/_2999_ ;
 wire net43;
 wire net42;
 wire net41;
 wire \register_file_i/_3003_ ;
 wire net40;
 wire net39;
 wire net38;
 wire \register_file_i/_3007_ ;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire \register_file_i/_3012_ ;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire \register_file_i/_3017_ ;
 wire net29;
 wire net28;
 wire net27;
 wire \register_file_i/_3021_ ;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire \register_file_i/_3026_ ;
 wire net22;
 wire net21;
 wire net20;
 wire \register_file_i/_3030_ ;
 wire net19;
 wire net18;
 wire net17;
 wire \register_file_i/_3034_ ;
 wire net16;
 wire net15;
 wire net14;
 wire \register_file_i/_3038_ ;
 wire net13;
 wire net12;
 wire net11;
 wire \register_file_i/_3042_ ;
 wire \register_file_i/_3043_ ;
 wire \register_file_i/_3044_ ;
 wire \register_file_i/_3045_ ;
 wire \register_file_i/_3046_ ;
 wire \register_file_i/_3047_ ;
 wire \register_file_i/_3048_ ;
 wire \register_file_i/_3049_ ;
 wire \register_file_i/_3050_ ;
 wire \register_file_i/_3051_ ;
 wire \register_file_i/_3052_ ;
 wire \register_file_i/_3053_ ;
 wire \register_file_i/_3054_ ;
 wire \register_file_i/_3055_ ;
 wire \register_file_i/_3056_ ;
 wire \register_file_i/_3057_ ;
 wire \register_file_i/_3058_ ;
 wire \register_file_i/_3059_ ;
 wire \register_file_i/_3060_ ;
 wire \register_file_i/_3061_ ;
 wire \register_file_i/_3062_ ;
 wire \register_file_i/_3063_ ;
 wire \register_file_i/_3064_ ;
 wire \register_file_i/_3065_ ;
 wire \register_file_i/_3066_ ;
 wire \register_file_i/_3067_ ;
 wire \register_file_i/_3068_ ;
 wire \register_file_i/_3069_ ;
 wire \register_file_i/_3070_ ;
 wire \register_file_i/_3071_ ;
 wire \register_file_i/_3072_ ;
 wire \register_file_i/_3073_ ;
 wire \register_file_i/_3074_ ;
 wire \register_file_i/_3075_ ;
 wire \register_file_i/_3076_ ;
 wire \register_file_i/_3077_ ;
 wire \register_file_i/_3078_ ;
 wire \register_file_i/_3079_ ;
 wire \register_file_i/_3080_ ;
 wire \register_file_i/_3081_ ;
 wire \register_file_i/_3082_ ;
 wire \register_file_i/_3083_ ;
 wire \register_file_i/_3084_ ;
 wire \register_file_i/_3085_ ;
 wire \register_file_i/_3086_ ;
 wire \register_file_i/_3087_ ;
 wire \register_file_i/_3088_ ;
 wire \register_file_i/_3089_ ;
 wire \register_file_i/_3090_ ;
 wire \register_file_i/_3091_ ;
 wire \register_file_i/_3092_ ;
 wire \register_file_i/_3093_ ;
 wire \register_file_i/_3094_ ;
 wire \register_file_i/_3095_ ;
 wire \register_file_i/_3096_ ;
 wire \register_file_i/_3097_ ;
 wire \register_file_i/_3098_ ;
 wire \register_file_i/_3099_ ;
 wire \register_file_i/_3100_ ;
 wire \register_file_i/_3101_ ;
 wire \register_file_i/_3102_ ;
 wire \register_file_i/_3103_ ;
 wire \register_file_i/_3104_ ;
 wire \register_file_i/_3105_ ;
 wire \register_file_i/_3106_ ;
 wire \register_file_i/_3107_ ;
 wire \register_file_i/_3108_ ;
 wire \register_file_i/_3109_ ;
 wire \register_file_i/_3110_ ;
 wire \register_file_i/_3111_ ;
 wire \register_file_i/_3112_ ;
 wire \register_file_i/_3113_ ;
 wire \register_file_i/_3114_ ;
 wire \register_file_i/_3115_ ;
 wire \register_file_i/_3116_ ;
 wire \register_file_i/_3117_ ;
 wire \register_file_i/_3118_ ;
 wire \register_file_i/_3119_ ;
 wire \register_file_i/_3120_ ;
 wire \register_file_i/_3121_ ;
 wire \register_file_i/_3122_ ;
 wire \register_file_i/_3123_ ;
 wire \register_file_i/_3124_ ;
 wire \register_file_i/_3125_ ;
 wire \register_file_i/_3126_ ;
 wire \register_file_i/_3127_ ;
 wire \register_file_i/_3128_ ;
 wire \register_file_i/_3129_ ;
 wire \register_file_i/_3130_ ;
 wire \register_file_i/_3131_ ;
 wire \register_file_i/_3132_ ;
 wire \register_file_i/_3133_ ;
 wire \register_file_i/_3134_ ;
 wire \register_file_i/_3135_ ;
 wire \register_file_i/_3136_ ;
 wire \register_file_i/_3137_ ;
 wire \register_file_i/_3138_ ;
 wire \register_file_i/_3139_ ;
 wire \register_file_i/_3140_ ;
 wire \register_file_i/_3141_ ;
 wire \register_file_i/_3142_ ;
 wire \register_file_i/_3143_ ;
 wire \register_file_i/_3144_ ;
 wire \register_file_i/_3145_ ;
 wire \register_file_i/_3146_ ;
 wire \register_file_i/_3147_ ;
 wire \register_file_i/_3148_ ;
 wire \register_file_i/_3149_ ;
 wire \register_file_i/_3150_ ;
 wire \register_file_i/_3151_ ;
 wire \register_file_i/_3152_ ;
 wire \register_file_i/_3153_ ;
 wire \register_file_i/_3154_ ;
 wire \register_file_i/_3155_ ;
 wire \register_file_i/_3156_ ;
 wire \register_file_i/_3157_ ;
 wire \register_file_i/_3158_ ;
 wire \register_file_i/_3159_ ;
 wire \register_file_i/_3160_ ;
 wire \register_file_i/_3161_ ;
 wire \register_file_i/_3162_ ;
 wire \register_file_i/_3163_ ;
 wire \register_file_i/_3164_ ;
 wire \register_file_i/_3165_ ;
 wire \register_file_i/_3166_ ;
 wire \register_file_i/_3167_ ;
 wire \register_file_i/_3168_ ;
 wire \register_file_i/_3169_ ;
 wire \register_file_i/_3170_ ;
 wire \register_file_i/_3171_ ;
 wire \register_file_i/_3172_ ;
 wire \register_file_i/_3173_ ;
 wire \register_file_i/_3174_ ;
 wire \register_file_i/_3175_ ;
 wire \register_file_i/_3176_ ;
 wire \register_file_i/_3177_ ;
 wire \register_file_i/_3178_ ;
 wire \register_file_i/_3179_ ;
 wire \register_file_i/_3180_ ;
 wire \register_file_i/_3181_ ;
 wire \register_file_i/_3182_ ;
 wire \register_file_i/_3183_ ;
 wire \register_file_i/_3184_ ;
 wire \register_file_i/_3185_ ;
 wire \register_file_i/_3186_ ;
 wire \register_file_i/_3187_ ;
 wire \register_file_i/_3188_ ;
 wire \register_file_i/_3189_ ;
 wire \register_file_i/_3190_ ;
 wire \register_file_i/_3191_ ;
 wire \register_file_i/_3192_ ;
 wire \register_file_i/_3193_ ;
 wire \register_file_i/_3194_ ;
 wire \register_file_i/_3195_ ;
 wire \register_file_i/_3196_ ;
 wire \register_file_i/_3197_ ;
 wire \register_file_i/_3198_ ;
 wire \register_file_i/_3199_ ;
 wire \register_file_i/_3200_ ;
 wire \register_file_i/_3201_ ;
 wire \register_file_i/_3202_ ;
 wire \register_file_i/_3203_ ;
 wire \register_file_i/_3204_ ;
 wire \register_file_i/_3205_ ;
 wire \register_file_i/_3206_ ;
 wire \register_file_i/_3207_ ;
 wire \register_file_i/_3208_ ;
 wire \register_file_i/_3209_ ;
 wire \register_file_i/_3210_ ;
 wire \register_file_i/_3211_ ;
 wire \register_file_i/_3212_ ;
 wire \register_file_i/_3213_ ;
 wire \register_file_i/_3214_ ;
 wire \register_file_i/_3215_ ;
 wire \register_file_i/_3216_ ;
 wire \register_file_i/_3217_ ;
 wire \register_file_i/_3218_ ;
 wire \register_file_i/_3219_ ;
 wire \register_file_i/_3220_ ;
 wire \register_file_i/_3221_ ;
 wire \register_file_i/_3222_ ;
 wire \register_file_i/_3223_ ;
 wire \register_file_i/_3224_ ;
 wire \register_file_i/_3225_ ;
 wire \register_file_i/_3226_ ;
 wire \register_file_i/_3227_ ;
 wire \register_file_i/_3228_ ;
 wire \register_file_i/_3229_ ;
 wire \register_file_i/_3230_ ;
 wire \register_file_i/_3231_ ;
 wire \register_file_i/_3232_ ;
 wire \register_file_i/_3233_ ;
 wire \register_file_i/_3234_ ;
 wire \register_file_i/_3235_ ;
 wire \register_file_i/_3236_ ;
 wire \register_file_i/_3237_ ;
 wire \register_file_i/_3238_ ;
 wire \register_file_i/_3239_ ;
 wire \register_file_i/_3240_ ;
 wire \register_file_i/_3241_ ;
 wire \register_file_i/_3242_ ;
 wire \register_file_i/_3243_ ;
 wire \register_file_i/_3244_ ;
 wire \register_file_i/_3245_ ;
 wire \register_file_i/_3246_ ;
 wire \register_file_i/_3247_ ;
 wire \register_file_i/_3248_ ;
 wire \register_file_i/_3249_ ;
 wire \register_file_i/_3250_ ;
 wire \register_file_i/_3251_ ;
 wire \register_file_i/_3252_ ;
 wire \register_file_i/_3253_ ;
 wire \register_file_i/_3254_ ;
 wire \register_file_i/_3255_ ;
 wire \register_file_i/_3256_ ;
 wire \register_file_i/_3257_ ;
 wire \register_file_i/_3258_ ;
 wire \register_file_i/_3259_ ;
 wire \register_file_i/_3260_ ;
 wire \register_file_i/_3261_ ;
 wire \register_file_i/_3262_ ;
 wire \register_file_i/_3263_ ;
 wire \register_file_i/_3264_ ;
 wire \register_file_i/_3265_ ;
 wire \register_file_i/_3266_ ;
 wire \register_file_i/_3267_ ;
 wire \register_file_i/_3268_ ;
 wire \register_file_i/_3269_ ;
 wire \register_file_i/_3270_ ;
 wire \register_file_i/_3271_ ;
 wire \register_file_i/_3272_ ;
 wire \register_file_i/_3273_ ;
 wire \register_file_i/_3274_ ;
 wire \register_file_i/_3275_ ;
 wire \register_file_i/_3276_ ;
 wire \register_file_i/_3277_ ;
 wire \register_file_i/_3278_ ;
 wire \register_file_i/_3279_ ;
 wire \register_file_i/_3280_ ;
 wire \register_file_i/_3281_ ;
 wire \register_file_i/_3282_ ;
 wire \register_file_i/_3283_ ;
 wire \register_file_i/_3284_ ;
 wire \register_file_i/_3285_ ;
 wire \register_file_i/_3286_ ;
 wire \register_file_i/_3287_ ;
 wire \register_file_i/_3288_ ;
 wire \register_file_i/_3289_ ;
 wire \register_file_i/_3290_ ;
 wire \register_file_i/_3291_ ;
 wire \register_file_i/_3292_ ;
 wire \register_file_i/_3293_ ;
 wire \register_file_i/_3294_ ;
 wire \register_file_i/_3295_ ;
 wire \register_file_i/_3296_ ;
 wire \register_file_i/_3297_ ;
 wire \register_file_i/_3298_ ;
 wire \register_file_i/_3299_ ;
 wire \register_file_i/_3300_ ;
 wire \register_file_i/_3301_ ;
 wire \register_file_i/_3302_ ;
 wire \register_file_i/_3303_ ;
 wire \register_file_i/_3304_ ;
 wire \register_file_i/_3305_ ;
 wire \register_file_i/_3306_ ;
 wire \register_file_i/_3307_ ;
 wire \register_file_i/_3308_ ;
 wire \register_file_i/_3309_ ;
 wire \register_file_i/_3310_ ;
 wire \register_file_i/_3311_ ;
 wire \register_file_i/_3312_ ;
 wire \register_file_i/_3313_ ;
 wire \register_file_i/_3314_ ;
 wire \register_file_i/_3315_ ;
 wire \register_file_i/_3316_ ;
 wire \register_file_i/_3317_ ;
 wire \register_file_i/_3318_ ;
 wire \register_file_i/_3319_ ;
 wire \register_file_i/_3320_ ;
 wire \register_file_i/_3321_ ;
 wire \register_file_i/_3322_ ;
 wire \register_file_i/_3323_ ;
 wire \register_file_i/_3324_ ;
 wire \register_file_i/_3325_ ;
 wire \register_file_i/_3326_ ;
 wire \register_file_i/_3327_ ;
 wire \register_file_i/_3328_ ;
 wire \register_file_i/_3329_ ;
 wire \register_file_i/_3330_ ;
 wire \register_file_i/_3331_ ;
 wire \register_file_i/_3332_ ;
 wire \register_file_i/_3333_ ;
 wire \register_file_i/_3334_ ;
 wire \register_file_i/_3335_ ;
 wire \register_file_i/_3336_ ;
 wire \register_file_i/_3337_ ;
 wire \register_file_i/_3338_ ;
 wire \register_file_i/_3339_ ;
 wire \register_file_i/_3340_ ;
 wire \register_file_i/_3341_ ;
 wire \register_file_i/_3342_ ;
 wire \register_file_i/_3343_ ;
 wire \register_file_i/_3344_ ;
 wire \register_file_i/_3345_ ;
 wire \register_file_i/_3346_ ;
 wire \register_file_i/_3347_ ;
 wire \register_file_i/_3348_ ;
 wire \register_file_i/_3349_ ;
 wire \register_file_i/_3350_ ;
 wire \register_file_i/_3351_ ;
 wire \register_file_i/_3352_ ;
 wire \register_file_i/_3353_ ;
 wire \register_file_i/_3354_ ;
 wire \register_file_i/_3355_ ;
 wire \register_file_i/_3356_ ;
 wire \register_file_i/_3357_ ;
 wire \register_file_i/_3358_ ;
 wire \register_file_i/_3359_ ;
 wire \register_file_i/_3360_ ;
 wire \register_file_i/_3361_ ;
 wire \register_file_i/_3362_ ;
 wire \register_file_i/_3363_ ;
 wire \register_file_i/_3364_ ;
 wire \register_file_i/_3365_ ;
 wire \register_file_i/_3366_ ;
 wire \register_file_i/_3367_ ;
 wire \register_file_i/_3368_ ;
 wire \register_file_i/_3369_ ;
 wire \register_file_i/_3370_ ;
 wire \register_file_i/_3371_ ;
 wire \register_file_i/_3372_ ;
 wire \register_file_i/_3373_ ;
 wire \register_file_i/_3374_ ;
 wire \register_file_i/_3375_ ;
 wire \register_file_i/_3376_ ;
 wire \register_file_i/_3377_ ;
 wire \register_file_i/_3378_ ;
 wire \register_file_i/_3379_ ;
 wire \register_file_i/_3380_ ;
 wire \register_file_i/_3381_ ;
 wire \register_file_i/_3382_ ;
 wire \register_file_i/_3383_ ;
 wire \register_file_i/_3384_ ;
 wire \register_file_i/_3385_ ;
 wire \register_file_i/_3386_ ;
 wire \register_file_i/_3387_ ;
 wire \register_file_i/_3388_ ;
 wire \register_file_i/_3389_ ;
 wire \register_file_i/_3390_ ;
 wire \register_file_i/_3391_ ;
 wire \register_file_i/_3392_ ;
 wire \register_file_i/_3393_ ;
 wire \register_file_i/_3394_ ;
 wire \register_file_i/_3395_ ;
 wire \register_file_i/_3396_ ;
 wire \register_file_i/_3397_ ;
 wire \register_file_i/_3398_ ;
 wire \register_file_i/_3399_ ;
 wire \register_file_i/_3400_ ;
 wire \register_file_i/_3401_ ;
 wire \register_file_i/_3402_ ;
 wire \register_file_i/_3403_ ;
 wire \register_file_i/_3404_ ;
 wire \register_file_i/_3405_ ;
 wire \register_file_i/_3406_ ;
 wire \register_file_i/_3407_ ;
 wire \register_file_i/_3408_ ;
 wire \register_file_i/_3409_ ;
 wire \register_file_i/_3410_ ;
 wire \register_file_i/_3411_ ;
 wire \register_file_i/_3412_ ;
 wire \register_file_i/_3413_ ;
 wire \register_file_i/_3414_ ;
 wire \register_file_i/_3415_ ;
 wire \register_file_i/_3416_ ;
 wire \register_file_i/_3417_ ;
 wire \register_file_i/_3418_ ;
 wire \register_file_i/_3419_ ;
 wire \register_file_i/_3420_ ;
 wire \register_file_i/_3421_ ;
 wire \register_file_i/_3422_ ;
 wire \register_file_i/_3423_ ;
 wire \register_file_i/_3424_ ;
 wire \register_file_i/_3425_ ;
 wire \register_file_i/_3426_ ;
 wire \register_file_i/_3427_ ;
 wire \register_file_i/_3428_ ;
 wire \register_file_i/_3429_ ;
 wire \register_file_i/_3430_ ;
 wire \register_file_i/_3431_ ;
 wire \register_file_i/_3432_ ;
 wire \register_file_i/_3433_ ;
 wire \register_file_i/_3434_ ;
 wire \register_file_i/_3435_ ;
 wire \register_file_i/_3436_ ;
 wire \register_file_i/_3437_ ;
 wire \register_file_i/_3438_ ;
 wire \register_file_i/_3439_ ;
 wire \register_file_i/_3440_ ;
 wire \register_file_i/_3441_ ;
 wire \register_file_i/_3442_ ;
 wire \register_file_i/_3443_ ;
 wire \register_file_i/_3444_ ;
 wire \register_file_i/_3445_ ;
 wire \register_file_i/_3446_ ;
 wire \register_file_i/_3447_ ;
 wire \register_file_i/_3448_ ;
 wire \register_file_i/_3449_ ;
 wire \register_file_i/_3450_ ;
 wire \register_file_i/_3451_ ;
 wire \register_file_i/_3452_ ;
 wire \register_file_i/_3453_ ;
 wire \register_file_i/_3454_ ;
 wire \register_file_i/_3455_ ;
 wire \register_file_i/_3456_ ;
 wire \register_file_i/_3457_ ;
 wire \register_file_i/_3458_ ;
 wire \register_file_i/_3459_ ;
 wire \register_file_i/_3460_ ;
 wire \register_file_i/_3461_ ;
 wire \register_file_i/_3462_ ;
 wire \register_file_i/_3463_ ;
 wire \register_file_i/_3464_ ;
 wire \register_file_i/_3465_ ;
 wire \register_file_i/_3466_ ;
 wire \register_file_i/_3467_ ;
 wire \register_file_i/_3468_ ;
 wire \register_file_i/_3469_ ;
 wire \register_file_i/_3470_ ;
 wire \register_file_i/_3471_ ;
 wire \register_file_i/_3472_ ;
 wire \register_file_i/_3473_ ;
 wire \register_file_i/_3474_ ;
 wire \register_file_i/_3475_ ;
 wire \register_file_i/_3476_ ;
 wire \register_file_i/_3477_ ;
 wire \register_file_i/_3478_ ;
 wire \register_file_i/_3479_ ;
 wire \register_file_i/_3480_ ;
 wire \register_file_i/_3481_ ;
 wire \register_file_i/_3482_ ;
 wire \register_file_i/_3483_ ;
 wire \register_file_i/_3484_ ;
 wire \register_file_i/_3485_ ;
 wire \register_file_i/_3486_ ;
 wire \register_file_i/_3487_ ;
 wire \register_file_i/_3488_ ;
 wire \register_file_i/_3489_ ;
 wire \register_file_i/_3490_ ;
 wire \register_file_i/_3491_ ;
 wire \register_file_i/_3492_ ;
 wire \register_file_i/_3493_ ;
 wire \register_file_i/_3494_ ;
 wire \register_file_i/_3495_ ;
 wire \register_file_i/_3496_ ;
 wire \register_file_i/_3497_ ;
 wire \register_file_i/_3498_ ;
 wire \register_file_i/_3499_ ;
 wire \register_file_i/_3500_ ;
 wire \register_file_i/_3501_ ;
 wire \register_file_i/_3502_ ;
 wire \register_file_i/_3503_ ;
 wire \register_file_i/_3504_ ;
 wire \register_file_i/_3505_ ;
 wire \register_file_i/_3506_ ;
 wire \register_file_i/_3507_ ;
 wire \register_file_i/_3508_ ;
 wire \register_file_i/_3509_ ;
 wire \register_file_i/_3510_ ;
 wire \register_file_i/_3511_ ;
 wire \register_file_i/_3512_ ;
 wire \register_file_i/_3513_ ;
 wire \register_file_i/_3514_ ;
 wire \register_file_i/_3515_ ;
 wire \register_file_i/_3516_ ;
 wire \register_file_i/_3517_ ;
 wire \register_file_i/_3518_ ;
 wire \register_file_i/_3519_ ;
 wire \register_file_i/_3520_ ;
 wire \register_file_i/_3521_ ;
 wire \register_file_i/_3522_ ;
 wire \register_file_i/_3523_ ;
 wire \register_file_i/_3524_ ;
 wire \register_file_i/_3525_ ;
 wire \register_file_i/_3526_ ;
 wire \register_file_i/_3527_ ;
 wire \register_file_i/_3528_ ;
 wire \register_file_i/_3529_ ;
 wire \register_file_i/_3530_ ;
 wire \register_file_i/_3531_ ;
 wire \register_file_i/_3532_ ;
 wire \register_file_i/_3533_ ;
 wire \register_file_i/_3534_ ;
 wire \register_file_i/_3535_ ;
 wire \register_file_i/_3536_ ;
 wire \register_file_i/_3537_ ;
 wire \register_file_i/_3538_ ;
 wire \register_file_i/_3539_ ;
 wire \register_file_i/_3540_ ;
 wire \register_file_i/_3541_ ;
 wire \register_file_i/_3542_ ;
 wire \register_file_i/_3543_ ;
 wire \register_file_i/_3544_ ;
 wire \register_file_i/_3545_ ;
 wire \register_file_i/_3546_ ;
 wire \register_file_i/_3547_ ;
 wire \register_file_i/_3548_ ;
 wire \register_file_i/_3549_ ;
 wire \register_file_i/_3550_ ;
 wire \register_file_i/_3551_ ;
 wire \register_file_i/_3552_ ;
 wire \register_file_i/_3553_ ;
 wire \register_file_i/_3554_ ;
 wire \register_file_i/_3555_ ;
 wire \register_file_i/_3556_ ;
 wire \register_file_i/_3557_ ;
 wire \register_file_i/_3558_ ;
 wire \register_file_i/_3559_ ;
 wire \register_file_i/_3560_ ;
 wire \register_file_i/_3561_ ;
 wire \register_file_i/_3562_ ;
 wire \register_file_i/_3563_ ;
 wire \register_file_i/_3564_ ;
 wire \register_file_i/_3565_ ;
 wire \register_file_i/_3566_ ;
 wire \register_file_i/_3567_ ;
 wire \register_file_i/_3568_ ;
 wire \register_file_i/_3569_ ;
 wire \register_file_i/_3570_ ;
 wire \register_file_i/_3571_ ;
 wire \register_file_i/_3572_ ;
 wire \register_file_i/_3573_ ;
 wire \register_file_i/_3574_ ;
 wire \register_file_i/_3575_ ;
 wire \register_file_i/_3576_ ;
 wire \register_file_i/_3577_ ;
 wire \register_file_i/_3578_ ;
 wire \register_file_i/_3579_ ;
 wire \register_file_i/_3580_ ;
 wire \register_file_i/_3581_ ;
 wire \register_file_i/_3582_ ;
 wire \register_file_i/_3583_ ;
 wire \register_file_i/_3584_ ;
 wire \register_file_i/_3585_ ;
 wire \register_file_i/_3586_ ;
 wire \register_file_i/_3587_ ;
 wire \register_file_i/_3588_ ;
 wire \register_file_i/_3589_ ;
 wire \register_file_i/_3590_ ;
 wire \register_file_i/_3591_ ;
 wire \register_file_i/_3592_ ;
 wire \register_file_i/_3593_ ;
 wire \register_file_i/_3594_ ;
 wire \register_file_i/_3595_ ;
 wire \register_file_i/_3596_ ;
 wire \register_file_i/_3597_ ;
 wire \register_file_i/_3598_ ;
 wire \register_file_i/_3599_ ;
 wire \register_file_i/_3600_ ;
 wire \register_file_i/_3601_ ;
 wire \register_file_i/_3602_ ;
 wire \register_file_i/_3603_ ;
 wire \register_file_i/_3604_ ;
 wire \register_file_i/_3605_ ;
 wire \register_file_i/_3606_ ;
 wire \register_file_i/_3607_ ;
 wire \register_file_i/_3608_ ;
 wire \register_file_i/_3609_ ;
 wire \register_file_i/_3610_ ;
 wire \register_file_i/_3611_ ;
 wire \register_file_i/_3612_ ;
 wire \register_file_i/_3613_ ;
 wire \register_file_i/_3614_ ;
 wire \register_file_i/_3615_ ;
 wire \register_file_i/_3616_ ;
 wire \register_file_i/_3617_ ;
 wire \register_file_i/_3618_ ;
 wire \register_file_i/_3619_ ;
 wire \register_file_i/_3620_ ;
 wire \register_file_i/_3621_ ;
 wire \register_file_i/_3622_ ;
 wire \register_file_i/_3623_ ;
 wire \register_file_i/_3624_ ;
 wire \register_file_i/_3625_ ;
 wire \register_file_i/_3626_ ;
 wire \register_file_i/_3627_ ;
 wire \register_file_i/_3628_ ;
 wire \register_file_i/_3629_ ;
 wire \register_file_i/_3630_ ;
 wire \register_file_i/_3631_ ;
 wire \register_file_i/_3632_ ;
 wire \register_file_i/_3633_ ;
 wire \register_file_i/_3634_ ;
 wire \register_file_i/_3635_ ;
 wire \register_file_i/_3636_ ;
 wire \register_file_i/_3637_ ;
 wire \register_file_i/_3638_ ;
 wire \register_file_i/_3639_ ;
 wire \register_file_i/_3640_ ;
 wire \register_file_i/_3641_ ;
 wire \register_file_i/_3642_ ;
 wire \register_file_i/_3643_ ;
 wire \register_file_i/_3644_ ;
 wire \register_file_i/_3645_ ;
 wire \register_file_i/_3646_ ;
 wire \register_file_i/_3647_ ;
 wire \register_file_i/_3648_ ;
 wire \register_file_i/_3649_ ;
 wire \register_file_i/_3650_ ;
 wire \register_file_i/_3651_ ;
 wire \register_file_i/_3652_ ;
 wire \register_file_i/_3653_ ;
 wire \register_file_i/_3654_ ;
 wire \register_file_i/_3655_ ;
 wire \register_file_i/_3656_ ;
 wire \register_file_i/_3657_ ;
 wire \register_file_i/_3658_ ;
 wire \register_file_i/_3659_ ;
 wire \register_file_i/_3660_ ;
 wire \register_file_i/_3661_ ;
 wire \register_file_i/_3662_ ;
 wire \register_file_i/_3663_ ;
 wire \register_file_i/_3664_ ;
 wire \register_file_i/_3665_ ;
 wire \register_file_i/_3666_ ;
 wire \register_file_i/_3667_ ;
 wire \register_file_i/_3668_ ;
 wire \register_file_i/_3669_ ;
 wire \register_file_i/_3670_ ;
 wire \register_file_i/_3671_ ;
 wire \register_file_i/_3672_ ;
 wire \register_file_i/_3673_ ;
 wire \register_file_i/_3674_ ;
 wire \register_file_i/_3675_ ;
 wire \register_file_i/_3676_ ;
 wire \register_file_i/_3677_ ;
 wire \register_file_i/_3678_ ;
 wire \register_file_i/_3679_ ;
 wire \register_file_i/_3680_ ;
 wire \register_file_i/_3681_ ;
 wire \register_file_i/_3682_ ;
 wire \register_file_i/_3683_ ;
 wire \register_file_i/_3684_ ;
 wire \register_file_i/_3685_ ;
 wire \register_file_i/_3686_ ;
 wire \register_file_i/_3687_ ;
 wire \register_file_i/_3688_ ;
 wire \register_file_i/_3689_ ;
 wire \register_file_i/_3690_ ;
 wire \register_file_i/_3691_ ;
 wire \register_file_i/_3692_ ;
 wire \register_file_i/_3693_ ;
 wire \register_file_i/_3694_ ;
 wire \register_file_i/_3695_ ;
 wire \register_file_i/_3696_ ;
 wire \register_file_i/_3697_ ;
 wire \register_file_i/_3698_ ;
 wire \register_file_i/_3699_ ;
 wire \register_file_i/_3700_ ;
 wire \register_file_i/_3701_ ;
 wire \register_file_i/_3702_ ;
 wire \register_file_i/_3703_ ;
 wire \register_file_i/_3704_ ;
 wire \register_file_i/_3705_ ;
 wire \register_file_i/_3706_ ;
 wire \register_file_i/_3707_ ;
 wire \register_file_i/_3708_ ;
 wire \register_file_i/_3709_ ;
 wire \register_file_i/_3710_ ;
 wire \register_file_i/_3711_ ;
 wire \register_file_i/_3712_ ;
 wire \register_file_i/_3713_ ;
 wire \register_file_i/_3714_ ;
 wire \register_file_i/_3715_ ;
 wire \register_file_i/_3716_ ;
 wire \register_file_i/_3717_ ;
 wire \register_file_i/_3718_ ;
 wire \register_file_i/_3719_ ;
 wire \register_file_i/_3720_ ;
 wire \register_file_i/_3721_ ;
 wire \register_file_i/_3722_ ;
 wire \register_file_i/_3723_ ;
 wire \register_file_i/_3724_ ;
 wire \register_file_i/_3725_ ;
 wire \register_file_i/_3726_ ;
 wire \register_file_i/_3727_ ;
 wire \register_file_i/_3728_ ;
 wire \register_file_i/_3729_ ;
 wire \register_file_i/_3730_ ;
 wire \register_file_i/_3731_ ;
 wire \register_file_i/_3732_ ;
 wire \register_file_i/_3733_ ;
 wire \register_file_i/_3734_ ;
 wire \register_file_i/_3735_ ;
 wire \register_file_i/_3736_ ;
 wire \register_file_i/_3737_ ;
 wire \register_file_i/_3738_ ;
 wire \register_file_i/_3739_ ;
 wire \register_file_i/_3740_ ;
 wire \register_file_i/_3741_ ;
 wire \register_file_i/_3742_ ;
 wire \register_file_i/_3743_ ;
 wire \register_file_i/_3744_ ;
 wire \register_file_i/_3745_ ;
 wire \register_file_i/_3746_ ;
 wire \register_file_i/_3747_ ;
 wire \register_file_i/_3748_ ;
 wire \register_file_i/_3749_ ;
 wire \register_file_i/_3750_ ;
 wire \register_file_i/_3751_ ;
 wire \register_file_i/_3752_ ;
 wire \register_file_i/_3753_ ;
 wire \register_file_i/_3754_ ;
 wire \register_file_i/_3755_ ;
 wire \register_file_i/_3756_ ;
 wire \register_file_i/_3757_ ;
 wire \register_file_i/_3758_ ;
 wire \register_file_i/_3759_ ;
 wire \register_file_i/_3760_ ;
 wire \register_file_i/_3761_ ;
 wire \register_file_i/_3762_ ;
 wire \register_file_i/_3763_ ;
 wire \register_file_i/_3764_ ;
 wire \register_file_i/_3765_ ;
 wire \register_file_i/_3766_ ;
 wire \register_file_i/_3767_ ;
 wire \register_file_i/_3768_ ;
 wire \register_file_i/_3769_ ;
 wire \register_file_i/_3770_ ;
 wire \register_file_i/_3771_ ;
 wire \register_file_i/_3772_ ;
 wire \register_file_i/_3773_ ;
 wire \register_file_i/_3774_ ;
 wire \register_file_i/_3775_ ;
 wire \register_file_i/_3776_ ;
 wire \register_file_i/_3777_ ;
 wire \register_file_i/_3778_ ;
 wire \register_file_i/_3779_ ;
 wire \register_file_i/_3780_ ;
 wire \register_file_i/_3781_ ;
 wire \register_file_i/_3782_ ;
 wire \register_file_i/_3783_ ;
 wire \register_file_i/_3784_ ;
 wire \register_file_i/_3785_ ;
 wire \register_file_i/_3786_ ;
 wire \register_file_i/_3787_ ;
 wire \register_file_i/_3788_ ;
 wire \register_file_i/_3789_ ;
 wire \register_file_i/_3790_ ;
 wire \register_file_i/_3791_ ;
 wire \register_file_i/_3792_ ;
 wire \register_file_i/_3793_ ;
 wire \register_file_i/_3794_ ;
 wire \register_file_i/_3795_ ;
 wire \register_file_i/_3796_ ;
 wire \register_file_i/_3797_ ;
 wire \register_file_i/_3798_ ;
 wire \register_file_i/_3799_ ;
 wire \register_file_i/_3800_ ;
 wire \register_file_i/_3801_ ;
 wire \register_file_i/_3802_ ;
 wire \register_file_i/_3803_ ;
 wire \register_file_i/_3804_ ;
 wire \register_file_i/_3805_ ;
 wire \register_file_i/_3806_ ;
 wire \register_file_i/_3807_ ;
 wire \register_file_i/_3808_ ;
 wire \register_file_i/_3809_ ;
 wire \register_file_i/_3810_ ;
 wire \register_file_i/_3811_ ;
 wire \register_file_i/_3812_ ;
 wire \register_file_i/_3813_ ;
 wire \register_file_i/_3814_ ;
 wire \register_file_i/_3815_ ;
 wire \register_file_i/_3816_ ;
 wire \register_file_i/_3817_ ;
 wire \register_file_i/_3818_ ;
 wire \register_file_i/_3819_ ;
 wire \register_file_i/_3820_ ;
 wire \register_file_i/_3821_ ;
 wire \register_file_i/_3822_ ;
 wire \register_file_i/_3823_ ;
 wire \register_file_i/_3824_ ;
 wire \register_file_i/_3825_ ;
 wire \register_file_i/_3826_ ;
 wire \register_file_i/_3827_ ;
 wire \register_file_i/_3828_ ;
 wire \register_file_i/_3829_ ;
 wire \register_file_i/_3830_ ;
 wire \register_file_i/_3831_ ;
 wire \register_file_i/_3832_ ;
 wire \register_file_i/_3833_ ;
 wire \register_file_i/_3834_ ;
 wire \register_file_i/_3835_ ;
 wire \register_file_i/_3836_ ;
 wire \register_file_i/_3837_ ;
 wire \register_file_i/_3838_ ;
 wire \register_file_i/_3839_ ;
 wire \register_file_i/_3840_ ;
 wire \register_file_i/_3841_ ;
 wire \register_file_i/_3842_ ;
 wire \register_file_i/_3843_ ;
 wire \register_file_i/_3844_ ;
 wire \register_file_i/_3845_ ;
 wire \register_file_i/_3846_ ;
 wire \register_file_i/_3847_ ;
 wire \register_file_i/_3848_ ;
 wire \register_file_i/_3849_ ;
 wire \register_file_i/_3850_ ;
 wire \register_file_i/_3851_ ;
 wire \register_file_i/_3852_ ;
 wire \register_file_i/_3853_ ;
 wire \register_file_i/_3854_ ;
 wire \register_file_i/_3855_ ;
 wire \register_file_i/_3856_ ;
 wire \register_file_i/_3857_ ;
 wire \register_file_i/_3858_ ;
 wire \register_file_i/_3859_ ;
 wire \register_file_i/_3860_ ;
 wire \register_file_i/_3861_ ;
 wire \register_file_i/_3862_ ;
 wire \register_file_i/_3863_ ;
 wire \register_file_i/_3864_ ;
 wire \register_file_i/_3865_ ;
 wire \register_file_i/_3866_ ;
 wire \register_file_i/_3867_ ;
 wire \register_file_i/_3868_ ;
 wire \register_file_i/_3869_ ;
 wire \register_file_i/_3870_ ;
 wire \register_file_i/_3871_ ;
 wire \register_file_i/_3872_ ;
 wire \register_file_i/_3873_ ;
 wire \register_file_i/_3874_ ;
 wire \register_file_i/_3875_ ;
 wire \register_file_i/_3876_ ;
 wire \register_file_i/_3877_ ;
 wire \register_file_i/_3878_ ;
 wire \register_file_i/_3879_ ;
 wire \register_file_i/_3880_ ;
 wire \register_file_i/_3881_ ;
 wire \register_file_i/_3882_ ;
 wire \register_file_i/_3883_ ;
 wire \register_file_i/_3884_ ;
 wire \register_file_i/_3885_ ;
 wire \register_file_i/_3886_ ;
 wire \register_file_i/_3887_ ;
 wire \register_file_i/_3888_ ;
 wire \register_file_i/_3889_ ;
 wire \register_file_i/_3890_ ;
 wire \register_file_i/_3891_ ;
 wire \register_file_i/_3892_ ;
 wire \register_file_i/_3893_ ;
 wire \register_file_i/_3894_ ;
 wire \register_file_i/_3895_ ;
 wire \register_file_i/_3896_ ;
 wire \register_file_i/_3897_ ;
 wire \register_file_i/_3898_ ;
 wire \register_file_i/_3899_ ;
 wire \register_file_i/_3900_ ;
 wire \register_file_i/_3901_ ;
 wire \register_file_i/_3902_ ;
 wire \register_file_i/_3903_ ;
 wire \register_file_i/_3904_ ;
 wire \register_file_i/_3905_ ;
 wire \register_file_i/_3906_ ;
 wire \register_file_i/_3907_ ;
 wire \register_file_i/_3908_ ;
 wire \register_file_i/_3909_ ;
 wire \register_file_i/_3910_ ;
 wire \register_file_i/_3911_ ;
 wire \register_file_i/_3912_ ;
 wire \register_file_i/_3913_ ;
 wire \register_file_i/_3914_ ;
 wire \register_file_i/_3915_ ;
 wire \register_file_i/_3916_ ;
 wire \register_file_i/_3917_ ;
 wire \register_file_i/_3918_ ;
 wire \register_file_i/_3919_ ;
 wire \register_file_i/_3920_ ;
 wire \register_file_i/_3921_ ;
 wire \register_file_i/_3922_ ;
 wire \register_file_i/_3923_ ;
 wire \register_file_i/_3924_ ;
 wire \register_file_i/_3925_ ;
 wire \register_file_i/_3926_ ;
 wire \register_file_i/_3927_ ;
 wire \register_file_i/_3928_ ;
 wire \register_file_i/_3929_ ;
 wire \register_file_i/_3930_ ;
 wire \register_file_i/_3931_ ;
 wire \register_file_i/_3932_ ;
 wire \register_file_i/_3933_ ;
 wire \register_file_i/_3934_ ;
 wire \register_file_i/_3935_ ;
 wire \register_file_i/_3936_ ;
 wire \register_file_i/_3937_ ;
 wire \register_file_i/_3938_ ;
 wire \register_file_i/_3939_ ;
 wire \register_file_i/_3940_ ;
 wire \register_file_i/_3941_ ;
 wire \register_file_i/_3942_ ;
 wire \register_file_i/_3943_ ;
 wire \register_file_i/_3944_ ;
 wire \register_file_i/_3945_ ;
 wire \register_file_i/_3946_ ;
 wire \register_file_i/_3947_ ;
 wire \register_file_i/_3948_ ;
 wire \register_file_i/_3949_ ;
 wire \register_file_i/_3950_ ;
 wire \register_file_i/_3951_ ;
 wire \register_file_i/_3952_ ;
 wire \register_file_i/_3953_ ;
 wire \register_file_i/_3954_ ;
 wire \register_file_i/_3955_ ;
 wire \register_file_i/_3956_ ;
 wire \register_file_i/_3957_ ;
 wire \register_file_i/_3958_ ;
 wire \register_file_i/_3959_ ;
 wire \register_file_i/_3960_ ;
 wire \register_file_i/_3961_ ;
 wire \register_file_i/_3962_ ;
 wire \register_file_i/_3963_ ;
 wire \register_file_i/_3964_ ;
 wire \register_file_i/_3965_ ;
 wire \register_file_i/_3966_ ;
 wire \register_file_i/_3967_ ;
 wire \register_file_i/_3968_ ;
 wire \register_file_i/_3969_ ;
 wire \register_file_i/_3970_ ;
 wire \register_file_i/_3971_ ;
 wire \register_file_i/_3972_ ;
 wire \register_file_i/_3973_ ;
 wire \register_file_i/_3974_ ;
 wire \register_file_i/_3975_ ;
 wire \register_file_i/_3976_ ;
 wire \register_file_i/_3977_ ;
 wire \register_file_i/_3978_ ;
 wire \register_file_i/_3979_ ;
 wire \register_file_i/_3980_ ;
 wire \register_file_i/_3981_ ;
 wire \register_file_i/_3982_ ;
 wire \register_file_i/_3983_ ;
 wire \register_file_i/_3984_ ;
 wire \register_file_i/_3985_ ;
 wire \register_file_i/_3986_ ;
 wire \register_file_i/_3987_ ;
 wire \register_file_i/_3988_ ;
 wire \register_file_i/_3989_ ;
 wire \register_file_i/_3990_ ;
 wire \register_file_i/_3991_ ;
 wire \register_file_i/_3992_ ;
 wire \register_file_i/_3993_ ;
 wire \register_file_i/_3994_ ;
 wire \register_file_i/_3995_ ;
 wire \register_file_i/_3996_ ;
 wire \register_file_i/_3997_ ;
 wire \register_file_i/_3998_ ;
 wire \register_file_i/_3999_ ;
 wire \register_file_i/_4000_ ;
 wire \register_file_i/_4001_ ;
 wire \register_file_i/_4002_ ;
 wire \register_file_i/_4003_ ;
 wire \register_file_i/_4004_ ;
 wire \register_file_i/_4005_ ;
 wire \register_file_i/_4006_ ;
 wire \register_file_i/_4007_ ;
 wire \register_file_i/_4008_ ;
 wire \register_file_i/_4009_ ;
 wire \register_file_i/_4010_ ;
 wire \register_file_i/_4011_ ;
 wire \register_file_i/_4012_ ;
 wire \register_file_i/_4013_ ;
 wire \register_file_i/_4014_ ;
 wire \register_file_i/_4015_ ;
 wire \register_file_i/_4016_ ;
 wire \register_file_i/_4017_ ;
 wire \register_file_i/_4018_ ;
 wire \register_file_i/_4019_ ;
 wire \register_file_i/_4020_ ;
 wire \register_file_i/_4021_ ;
 wire \register_file_i/_4022_ ;
 wire \register_file_i/_4023_ ;
 wire \register_file_i/_4024_ ;
 wire \register_file_i/_4025_ ;
 wire \register_file_i/_4026_ ;
 wire \register_file_i/_4027_ ;
 wire \register_file_i/_4028_ ;
 wire \register_file_i/_4029_ ;
 wire \register_file_i/_4030_ ;
 wire \register_file_i/_4031_ ;
 wire \register_file_i/_4032_ ;
 wire \register_file_i/_4033_ ;
 wire \register_file_i/rf_reg_1000_ ;
 wire \register_file_i/rf_reg_1001_ ;
 wire \register_file_i/rf_reg_1002_ ;
 wire \register_file_i/rf_reg_1003_ ;
 wire \register_file_i/rf_reg_1004_ ;
 wire \register_file_i/rf_reg_1005_ ;
 wire \register_file_i/rf_reg_1006_ ;
 wire \register_file_i/rf_reg_1007_ ;
 wire \register_file_i/rf_reg_1008_ ;
 wire \register_file_i/rf_reg_1009_ ;
 wire \register_file_i/rf_reg_100_ ;
 wire \register_file_i/rf_reg_1010_ ;
 wire \register_file_i/rf_reg_1011_ ;
 wire \register_file_i/rf_reg_1012_ ;
 wire \register_file_i/rf_reg_1013_ ;
 wire \register_file_i/rf_reg_1014_ ;
 wire \register_file_i/rf_reg_1015_ ;
 wire \register_file_i/rf_reg_1016_ ;
 wire \register_file_i/rf_reg_1017_ ;
 wire \register_file_i/rf_reg_1018_ ;
 wire \register_file_i/rf_reg_1019_ ;
 wire \register_file_i/rf_reg_101_ ;
 wire \register_file_i/rf_reg_1020_ ;
 wire \register_file_i/rf_reg_1021_ ;
 wire \register_file_i/rf_reg_1022_ ;
 wire \register_file_i/rf_reg_1023_ ;
 wire \register_file_i/rf_reg_102_ ;
 wire \register_file_i/rf_reg_103_ ;
 wire \register_file_i/rf_reg_104_ ;
 wire \register_file_i/rf_reg_105_ ;
 wire \register_file_i/rf_reg_106_ ;
 wire \register_file_i/rf_reg_107_ ;
 wire \register_file_i/rf_reg_108_ ;
 wire \register_file_i/rf_reg_109_ ;
 wire \register_file_i/rf_reg_110_ ;
 wire \register_file_i/rf_reg_111_ ;
 wire \register_file_i/rf_reg_112_ ;
 wire \register_file_i/rf_reg_113_ ;
 wire \register_file_i/rf_reg_114_ ;
 wire \register_file_i/rf_reg_115_ ;
 wire \register_file_i/rf_reg_116_ ;
 wire \register_file_i/rf_reg_117_ ;
 wire \register_file_i/rf_reg_118_ ;
 wire \register_file_i/rf_reg_119_ ;
 wire \register_file_i/rf_reg_120_ ;
 wire \register_file_i/rf_reg_121_ ;
 wire \register_file_i/rf_reg_122_ ;
 wire \register_file_i/rf_reg_123_ ;
 wire \register_file_i/rf_reg_124_ ;
 wire \register_file_i/rf_reg_125_ ;
 wire \register_file_i/rf_reg_126_ ;
 wire \register_file_i/rf_reg_127_ ;
 wire \register_file_i/rf_reg_128_ ;
 wire \register_file_i/rf_reg_129_ ;
 wire \register_file_i/rf_reg_130_ ;
 wire \register_file_i/rf_reg_131_ ;
 wire \register_file_i/rf_reg_132_ ;
 wire \register_file_i/rf_reg_133_ ;
 wire \register_file_i/rf_reg_134_ ;
 wire \register_file_i/rf_reg_135_ ;
 wire \register_file_i/rf_reg_136_ ;
 wire \register_file_i/rf_reg_137_ ;
 wire \register_file_i/rf_reg_138_ ;
 wire \register_file_i/rf_reg_139_ ;
 wire \register_file_i/rf_reg_140_ ;
 wire \register_file_i/rf_reg_141_ ;
 wire \register_file_i/rf_reg_142_ ;
 wire \register_file_i/rf_reg_143_ ;
 wire \register_file_i/rf_reg_144_ ;
 wire \register_file_i/rf_reg_145_ ;
 wire \register_file_i/rf_reg_146_ ;
 wire \register_file_i/rf_reg_147_ ;
 wire \register_file_i/rf_reg_148_ ;
 wire \register_file_i/rf_reg_149_ ;
 wire \register_file_i/rf_reg_150_ ;
 wire \register_file_i/rf_reg_151_ ;
 wire \register_file_i/rf_reg_152_ ;
 wire \register_file_i/rf_reg_153_ ;
 wire \register_file_i/rf_reg_154_ ;
 wire \register_file_i/rf_reg_155_ ;
 wire \register_file_i/rf_reg_156_ ;
 wire \register_file_i/rf_reg_157_ ;
 wire \register_file_i/rf_reg_158_ ;
 wire \register_file_i/rf_reg_159_ ;
 wire \register_file_i/rf_reg_160_ ;
 wire \register_file_i/rf_reg_161_ ;
 wire \register_file_i/rf_reg_162_ ;
 wire \register_file_i/rf_reg_163_ ;
 wire \register_file_i/rf_reg_164_ ;
 wire \register_file_i/rf_reg_165_ ;
 wire \register_file_i/rf_reg_166_ ;
 wire \register_file_i/rf_reg_167_ ;
 wire \register_file_i/rf_reg_168_ ;
 wire \register_file_i/rf_reg_169_ ;
 wire \register_file_i/rf_reg_170_ ;
 wire \register_file_i/rf_reg_171_ ;
 wire \register_file_i/rf_reg_172_ ;
 wire \register_file_i/rf_reg_173_ ;
 wire \register_file_i/rf_reg_174_ ;
 wire \register_file_i/rf_reg_175_ ;
 wire \register_file_i/rf_reg_176_ ;
 wire \register_file_i/rf_reg_177_ ;
 wire \register_file_i/rf_reg_178_ ;
 wire \register_file_i/rf_reg_179_ ;
 wire \register_file_i/rf_reg_180_ ;
 wire \register_file_i/rf_reg_181_ ;
 wire \register_file_i/rf_reg_182_ ;
 wire \register_file_i/rf_reg_183_ ;
 wire \register_file_i/rf_reg_184_ ;
 wire \register_file_i/rf_reg_185_ ;
 wire \register_file_i/rf_reg_186_ ;
 wire \register_file_i/rf_reg_187_ ;
 wire \register_file_i/rf_reg_188_ ;
 wire \register_file_i/rf_reg_189_ ;
 wire \register_file_i/rf_reg_190_ ;
 wire \register_file_i/rf_reg_191_ ;
 wire \register_file_i/rf_reg_192_ ;
 wire \register_file_i/rf_reg_193_ ;
 wire \register_file_i/rf_reg_194_ ;
 wire \register_file_i/rf_reg_195_ ;
 wire \register_file_i/rf_reg_196_ ;
 wire \register_file_i/rf_reg_197_ ;
 wire \register_file_i/rf_reg_198_ ;
 wire \register_file_i/rf_reg_199_ ;
 wire \register_file_i/rf_reg_200_ ;
 wire \register_file_i/rf_reg_201_ ;
 wire \register_file_i/rf_reg_202_ ;
 wire \register_file_i/rf_reg_203_ ;
 wire \register_file_i/rf_reg_204_ ;
 wire \register_file_i/rf_reg_205_ ;
 wire \register_file_i/rf_reg_206_ ;
 wire \register_file_i/rf_reg_207_ ;
 wire \register_file_i/rf_reg_208_ ;
 wire \register_file_i/rf_reg_209_ ;
 wire \register_file_i/rf_reg_210_ ;
 wire \register_file_i/rf_reg_211_ ;
 wire \register_file_i/rf_reg_212_ ;
 wire \register_file_i/rf_reg_213_ ;
 wire \register_file_i/rf_reg_214_ ;
 wire \register_file_i/rf_reg_215_ ;
 wire \register_file_i/rf_reg_216_ ;
 wire \register_file_i/rf_reg_217_ ;
 wire \register_file_i/rf_reg_218_ ;
 wire \register_file_i/rf_reg_219_ ;
 wire \register_file_i/rf_reg_220_ ;
 wire \register_file_i/rf_reg_221_ ;
 wire \register_file_i/rf_reg_222_ ;
 wire \register_file_i/rf_reg_223_ ;
 wire \register_file_i/rf_reg_224_ ;
 wire \register_file_i/rf_reg_225_ ;
 wire \register_file_i/rf_reg_226_ ;
 wire \register_file_i/rf_reg_227_ ;
 wire \register_file_i/rf_reg_228_ ;
 wire \register_file_i/rf_reg_229_ ;
 wire \register_file_i/rf_reg_230_ ;
 wire \register_file_i/rf_reg_231_ ;
 wire \register_file_i/rf_reg_232_ ;
 wire \register_file_i/rf_reg_233_ ;
 wire \register_file_i/rf_reg_234_ ;
 wire \register_file_i/rf_reg_235_ ;
 wire \register_file_i/rf_reg_236_ ;
 wire \register_file_i/rf_reg_237_ ;
 wire \register_file_i/rf_reg_238_ ;
 wire \register_file_i/rf_reg_239_ ;
 wire \register_file_i/rf_reg_240_ ;
 wire \register_file_i/rf_reg_241_ ;
 wire \register_file_i/rf_reg_242_ ;
 wire \register_file_i/rf_reg_243_ ;
 wire \register_file_i/rf_reg_244_ ;
 wire \register_file_i/rf_reg_245_ ;
 wire \register_file_i/rf_reg_246_ ;
 wire \register_file_i/rf_reg_247_ ;
 wire \register_file_i/rf_reg_248_ ;
 wire \register_file_i/rf_reg_249_ ;
 wire \register_file_i/rf_reg_250_ ;
 wire \register_file_i/rf_reg_251_ ;
 wire \register_file_i/rf_reg_252_ ;
 wire \register_file_i/rf_reg_253_ ;
 wire \register_file_i/rf_reg_254_ ;
 wire \register_file_i/rf_reg_255_ ;
 wire \register_file_i/rf_reg_256_ ;
 wire \register_file_i/rf_reg_257_ ;
 wire \register_file_i/rf_reg_258_ ;
 wire \register_file_i/rf_reg_259_ ;
 wire \register_file_i/rf_reg_260_ ;
 wire \register_file_i/rf_reg_261_ ;
 wire \register_file_i/rf_reg_262_ ;
 wire \register_file_i/rf_reg_263_ ;
 wire \register_file_i/rf_reg_264_ ;
 wire \register_file_i/rf_reg_265_ ;
 wire \register_file_i/rf_reg_266_ ;
 wire \register_file_i/rf_reg_267_ ;
 wire \register_file_i/rf_reg_268_ ;
 wire \register_file_i/rf_reg_269_ ;
 wire \register_file_i/rf_reg_270_ ;
 wire \register_file_i/rf_reg_271_ ;
 wire \register_file_i/rf_reg_272_ ;
 wire \register_file_i/rf_reg_273_ ;
 wire \register_file_i/rf_reg_274_ ;
 wire \register_file_i/rf_reg_275_ ;
 wire \register_file_i/rf_reg_276_ ;
 wire \register_file_i/rf_reg_277_ ;
 wire \register_file_i/rf_reg_278_ ;
 wire \register_file_i/rf_reg_279_ ;
 wire \register_file_i/rf_reg_280_ ;
 wire \register_file_i/rf_reg_281_ ;
 wire \register_file_i/rf_reg_282_ ;
 wire \register_file_i/rf_reg_283_ ;
 wire \register_file_i/rf_reg_284_ ;
 wire \register_file_i/rf_reg_285_ ;
 wire \register_file_i/rf_reg_286_ ;
 wire \register_file_i/rf_reg_287_ ;
 wire \register_file_i/rf_reg_288_ ;
 wire \register_file_i/rf_reg_289_ ;
 wire \register_file_i/rf_reg_290_ ;
 wire \register_file_i/rf_reg_291_ ;
 wire \register_file_i/rf_reg_292_ ;
 wire \register_file_i/rf_reg_293_ ;
 wire \register_file_i/rf_reg_294_ ;
 wire \register_file_i/rf_reg_295_ ;
 wire \register_file_i/rf_reg_296_ ;
 wire \register_file_i/rf_reg_297_ ;
 wire \register_file_i/rf_reg_298_ ;
 wire \register_file_i/rf_reg_299_ ;
 wire \register_file_i/rf_reg_300_ ;
 wire \register_file_i/rf_reg_301_ ;
 wire \register_file_i/rf_reg_302_ ;
 wire \register_file_i/rf_reg_303_ ;
 wire \register_file_i/rf_reg_304_ ;
 wire \register_file_i/rf_reg_305_ ;
 wire \register_file_i/rf_reg_306_ ;
 wire \register_file_i/rf_reg_307_ ;
 wire \register_file_i/rf_reg_308_ ;
 wire \register_file_i/rf_reg_309_ ;
 wire \register_file_i/rf_reg_310_ ;
 wire \register_file_i/rf_reg_311_ ;
 wire \register_file_i/rf_reg_312_ ;
 wire \register_file_i/rf_reg_313_ ;
 wire \register_file_i/rf_reg_314_ ;
 wire \register_file_i/rf_reg_315_ ;
 wire \register_file_i/rf_reg_316_ ;
 wire \register_file_i/rf_reg_317_ ;
 wire \register_file_i/rf_reg_318_ ;
 wire \register_file_i/rf_reg_319_ ;
 wire \register_file_i/rf_reg_320_ ;
 wire \register_file_i/rf_reg_321_ ;
 wire \register_file_i/rf_reg_322_ ;
 wire \register_file_i/rf_reg_323_ ;
 wire \register_file_i/rf_reg_324_ ;
 wire \register_file_i/rf_reg_325_ ;
 wire \register_file_i/rf_reg_326_ ;
 wire \register_file_i/rf_reg_327_ ;
 wire \register_file_i/rf_reg_328_ ;
 wire \register_file_i/rf_reg_329_ ;
 wire \register_file_i/rf_reg_32_ ;
 wire \register_file_i/rf_reg_330_ ;
 wire \register_file_i/rf_reg_331_ ;
 wire \register_file_i/rf_reg_332_ ;
 wire \register_file_i/rf_reg_333_ ;
 wire \register_file_i/rf_reg_334_ ;
 wire \register_file_i/rf_reg_335_ ;
 wire \register_file_i/rf_reg_336_ ;
 wire \register_file_i/rf_reg_337_ ;
 wire \register_file_i/rf_reg_338_ ;
 wire \register_file_i/rf_reg_339_ ;
 wire \register_file_i/rf_reg_33_ ;
 wire \register_file_i/rf_reg_340_ ;
 wire \register_file_i/rf_reg_341_ ;
 wire \register_file_i/rf_reg_342_ ;
 wire \register_file_i/rf_reg_343_ ;
 wire \register_file_i/rf_reg_344_ ;
 wire \register_file_i/rf_reg_345_ ;
 wire \register_file_i/rf_reg_346_ ;
 wire \register_file_i/rf_reg_347_ ;
 wire \register_file_i/rf_reg_348_ ;
 wire \register_file_i/rf_reg_349_ ;
 wire \register_file_i/rf_reg_34_ ;
 wire \register_file_i/rf_reg_350_ ;
 wire \register_file_i/rf_reg_351_ ;
 wire \register_file_i/rf_reg_352_ ;
 wire \register_file_i/rf_reg_353_ ;
 wire \register_file_i/rf_reg_354_ ;
 wire \register_file_i/rf_reg_355_ ;
 wire \register_file_i/rf_reg_356_ ;
 wire \register_file_i/rf_reg_357_ ;
 wire \register_file_i/rf_reg_358_ ;
 wire \register_file_i/rf_reg_359_ ;
 wire \register_file_i/rf_reg_35_ ;
 wire \register_file_i/rf_reg_360_ ;
 wire \register_file_i/rf_reg_361_ ;
 wire \register_file_i/rf_reg_362_ ;
 wire \register_file_i/rf_reg_363_ ;
 wire \register_file_i/rf_reg_364_ ;
 wire \register_file_i/rf_reg_365_ ;
 wire \register_file_i/rf_reg_366_ ;
 wire \register_file_i/rf_reg_367_ ;
 wire \register_file_i/rf_reg_368_ ;
 wire \register_file_i/rf_reg_369_ ;
 wire \register_file_i/rf_reg_36_ ;
 wire \register_file_i/rf_reg_370_ ;
 wire \register_file_i/rf_reg_371_ ;
 wire \register_file_i/rf_reg_372_ ;
 wire \register_file_i/rf_reg_373_ ;
 wire \register_file_i/rf_reg_374_ ;
 wire \register_file_i/rf_reg_375_ ;
 wire \register_file_i/rf_reg_376_ ;
 wire \register_file_i/rf_reg_377_ ;
 wire \register_file_i/rf_reg_378_ ;
 wire \register_file_i/rf_reg_379_ ;
 wire \register_file_i/rf_reg_37_ ;
 wire \register_file_i/rf_reg_380_ ;
 wire \register_file_i/rf_reg_381_ ;
 wire \register_file_i/rf_reg_382_ ;
 wire \register_file_i/rf_reg_383_ ;
 wire \register_file_i/rf_reg_384_ ;
 wire \register_file_i/rf_reg_385_ ;
 wire \register_file_i/rf_reg_386_ ;
 wire \register_file_i/rf_reg_387_ ;
 wire \register_file_i/rf_reg_388_ ;
 wire \register_file_i/rf_reg_389_ ;
 wire \register_file_i/rf_reg_38_ ;
 wire \register_file_i/rf_reg_390_ ;
 wire \register_file_i/rf_reg_391_ ;
 wire \register_file_i/rf_reg_392_ ;
 wire \register_file_i/rf_reg_393_ ;
 wire \register_file_i/rf_reg_394_ ;
 wire \register_file_i/rf_reg_395_ ;
 wire \register_file_i/rf_reg_396_ ;
 wire \register_file_i/rf_reg_397_ ;
 wire \register_file_i/rf_reg_398_ ;
 wire \register_file_i/rf_reg_399_ ;
 wire \register_file_i/rf_reg_39_ ;
 wire \register_file_i/rf_reg_400_ ;
 wire \register_file_i/rf_reg_401_ ;
 wire \register_file_i/rf_reg_402_ ;
 wire \register_file_i/rf_reg_403_ ;
 wire \register_file_i/rf_reg_404_ ;
 wire \register_file_i/rf_reg_405_ ;
 wire \register_file_i/rf_reg_406_ ;
 wire \register_file_i/rf_reg_407_ ;
 wire \register_file_i/rf_reg_408_ ;
 wire \register_file_i/rf_reg_409_ ;
 wire \register_file_i/rf_reg_40_ ;
 wire \register_file_i/rf_reg_410_ ;
 wire \register_file_i/rf_reg_411_ ;
 wire \register_file_i/rf_reg_412_ ;
 wire \register_file_i/rf_reg_413_ ;
 wire \register_file_i/rf_reg_414_ ;
 wire \register_file_i/rf_reg_415_ ;
 wire \register_file_i/rf_reg_416_ ;
 wire \register_file_i/rf_reg_417_ ;
 wire \register_file_i/rf_reg_418_ ;
 wire \register_file_i/rf_reg_419_ ;
 wire \register_file_i/rf_reg_41_ ;
 wire \register_file_i/rf_reg_420_ ;
 wire \register_file_i/rf_reg_421_ ;
 wire \register_file_i/rf_reg_422_ ;
 wire \register_file_i/rf_reg_423_ ;
 wire \register_file_i/rf_reg_424_ ;
 wire \register_file_i/rf_reg_425_ ;
 wire \register_file_i/rf_reg_426_ ;
 wire \register_file_i/rf_reg_427_ ;
 wire \register_file_i/rf_reg_428_ ;
 wire \register_file_i/rf_reg_429_ ;
 wire \register_file_i/rf_reg_42_ ;
 wire \register_file_i/rf_reg_430_ ;
 wire \register_file_i/rf_reg_431_ ;
 wire \register_file_i/rf_reg_432_ ;
 wire \register_file_i/rf_reg_433_ ;
 wire \register_file_i/rf_reg_434_ ;
 wire \register_file_i/rf_reg_435_ ;
 wire \register_file_i/rf_reg_436_ ;
 wire \register_file_i/rf_reg_437_ ;
 wire \register_file_i/rf_reg_438_ ;
 wire \register_file_i/rf_reg_439_ ;
 wire \register_file_i/rf_reg_43_ ;
 wire \register_file_i/rf_reg_440_ ;
 wire \register_file_i/rf_reg_441_ ;
 wire \register_file_i/rf_reg_442_ ;
 wire \register_file_i/rf_reg_443_ ;
 wire \register_file_i/rf_reg_444_ ;
 wire \register_file_i/rf_reg_445_ ;
 wire \register_file_i/rf_reg_446_ ;
 wire \register_file_i/rf_reg_447_ ;
 wire \register_file_i/rf_reg_448_ ;
 wire \register_file_i/rf_reg_449_ ;
 wire \register_file_i/rf_reg_44_ ;
 wire \register_file_i/rf_reg_450_ ;
 wire \register_file_i/rf_reg_451_ ;
 wire \register_file_i/rf_reg_452_ ;
 wire \register_file_i/rf_reg_453_ ;
 wire \register_file_i/rf_reg_454_ ;
 wire \register_file_i/rf_reg_455_ ;
 wire \register_file_i/rf_reg_456_ ;
 wire \register_file_i/rf_reg_457_ ;
 wire \register_file_i/rf_reg_458_ ;
 wire \register_file_i/rf_reg_459_ ;
 wire \register_file_i/rf_reg_45_ ;
 wire \register_file_i/rf_reg_460_ ;
 wire \register_file_i/rf_reg_461_ ;
 wire \register_file_i/rf_reg_462_ ;
 wire \register_file_i/rf_reg_463_ ;
 wire \register_file_i/rf_reg_464_ ;
 wire \register_file_i/rf_reg_465_ ;
 wire \register_file_i/rf_reg_466_ ;
 wire \register_file_i/rf_reg_467_ ;
 wire \register_file_i/rf_reg_468_ ;
 wire \register_file_i/rf_reg_469_ ;
 wire \register_file_i/rf_reg_46_ ;
 wire \register_file_i/rf_reg_470_ ;
 wire \register_file_i/rf_reg_471_ ;
 wire \register_file_i/rf_reg_472_ ;
 wire \register_file_i/rf_reg_473_ ;
 wire \register_file_i/rf_reg_474_ ;
 wire \register_file_i/rf_reg_475_ ;
 wire \register_file_i/rf_reg_476_ ;
 wire \register_file_i/rf_reg_477_ ;
 wire \register_file_i/rf_reg_478_ ;
 wire \register_file_i/rf_reg_479_ ;
 wire \register_file_i/rf_reg_47_ ;
 wire \register_file_i/rf_reg_480_ ;
 wire \register_file_i/rf_reg_481_ ;
 wire \register_file_i/rf_reg_482_ ;
 wire \register_file_i/rf_reg_483_ ;
 wire \register_file_i/rf_reg_484_ ;
 wire \register_file_i/rf_reg_485_ ;
 wire \register_file_i/rf_reg_486_ ;
 wire \register_file_i/rf_reg_487_ ;
 wire \register_file_i/rf_reg_488_ ;
 wire \register_file_i/rf_reg_489_ ;
 wire \register_file_i/rf_reg_48_ ;
 wire \register_file_i/rf_reg_490_ ;
 wire \register_file_i/rf_reg_491_ ;
 wire \register_file_i/rf_reg_492_ ;
 wire \register_file_i/rf_reg_493_ ;
 wire \register_file_i/rf_reg_494_ ;
 wire \register_file_i/rf_reg_495_ ;
 wire \register_file_i/rf_reg_496_ ;
 wire \register_file_i/rf_reg_497_ ;
 wire \register_file_i/rf_reg_498_ ;
 wire \register_file_i/rf_reg_499_ ;
 wire \register_file_i/rf_reg_49_ ;
 wire \register_file_i/rf_reg_500_ ;
 wire \register_file_i/rf_reg_501_ ;
 wire \register_file_i/rf_reg_502_ ;
 wire \register_file_i/rf_reg_503_ ;
 wire \register_file_i/rf_reg_504_ ;
 wire \register_file_i/rf_reg_505_ ;
 wire \register_file_i/rf_reg_506_ ;
 wire \register_file_i/rf_reg_507_ ;
 wire \register_file_i/rf_reg_508_ ;
 wire \register_file_i/rf_reg_509_ ;
 wire \register_file_i/rf_reg_50_ ;
 wire \register_file_i/rf_reg_510_ ;
 wire \register_file_i/rf_reg_511_ ;
 wire \register_file_i/rf_reg_512_ ;
 wire \register_file_i/rf_reg_513_ ;
 wire \register_file_i/rf_reg_514_ ;
 wire \register_file_i/rf_reg_515_ ;
 wire \register_file_i/rf_reg_516_ ;
 wire \register_file_i/rf_reg_517_ ;
 wire \register_file_i/rf_reg_518_ ;
 wire \register_file_i/rf_reg_519_ ;
 wire \register_file_i/rf_reg_51_ ;
 wire \register_file_i/rf_reg_520_ ;
 wire \register_file_i/rf_reg_521_ ;
 wire \register_file_i/rf_reg_522_ ;
 wire \register_file_i/rf_reg_523_ ;
 wire \register_file_i/rf_reg_524_ ;
 wire \register_file_i/rf_reg_525_ ;
 wire \register_file_i/rf_reg_526_ ;
 wire \register_file_i/rf_reg_527_ ;
 wire \register_file_i/rf_reg_528_ ;
 wire \register_file_i/rf_reg_529_ ;
 wire \register_file_i/rf_reg_52_ ;
 wire \register_file_i/rf_reg_530_ ;
 wire \register_file_i/rf_reg_531_ ;
 wire \register_file_i/rf_reg_532_ ;
 wire \register_file_i/rf_reg_533_ ;
 wire \register_file_i/rf_reg_534_ ;
 wire \register_file_i/rf_reg_535_ ;
 wire \register_file_i/rf_reg_536_ ;
 wire \register_file_i/rf_reg_537_ ;
 wire \register_file_i/rf_reg_538_ ;
 wire \register_file_i/rf_reg_539_ ;
 wire \register_file_i/rf_reg_53_ ;
 wire \register_file_i/rf_reg_540_ ;
 wire \register_file_i/rf_reg_541_ ;
 wire \register_file_i/rf_reg_542_ ;
 wire \register_file_i/rf_reg_543_ ;
 wire \register_file_i/rf_reg_544_ ;
 wire \register_file_i/rf_reg_545_ ;
 wire \register_file_i/rf_reg_546_ ;
 wire \register_file_i/rf_reg_547_ ;
 wire \register_file_i/rf_reg_548_ ;
 wire \register_file_i/rf_reg_549_ ;
 wire \register_file_i/rf_reg_54_ ;
 wire \register_file_i/rf_reg_550_ ;
 wire \register_file_i/rf_reg_551_ ;
 wire \register_file_i/rf_reg_552_ ;
 wire \register_file_i/rf_reg_553_ ;
 wire \register_file_i/rf_reg_554_ ;
 wire \register_file_i/rf_reg_555_ ;
 wire \register_file_i/rf_reg_556_ ;
 wire \register_file_i/rf_reg_557_ ;
 wire \register_file_i/rf_reg_558_ ;
 wire \register_file_i/rf_reg_559_ ;
 wire \register_file_i/rf_reg_55_ ;
 wire \register_file_i/rf_reg_560_ ;
 wire \register_file_i/rf_reg_561_ ;
 wire \register_file_i/rf_reg_562_ ;
 wire \register_file_i/rf_reg_563_ ;
 wire \register_file_i/rf_reg_564_ ;
 wire \register_file_i/rf_reg_565_ ;
 wire \register_file_i/rf_reg_566_ ;
 wire \register_file_i/rf_reg_567_ ;
 wire \register_file_i/rf_reg_568_ ;
 wire \register_file_i/rf_reg_569_ ;
 wire \register_file_i/rf_reg_56_ ;
 wire \register_file_i/rf_reg_570_ ;
 wire \register_file_i/rf_reg_571_ ;
 wire \register_file_i/rf_reg_572_ ;
 wire \register_file_i/rf_reg_573_ ;
 wire \register_file_i/rf_reg_574_ ;
 wire \register_file_i/rf_reg_575_ ;
 wire \register_file_i/rf_reg_576_ ;
 wire \register_file_i/rf_reg_577_ ;
 wire \register_file_i/rf_reg_578_ ;
 wire \register_file_i/rf_reg_579_ ;
 wire \register_file_i/rf_reg_57_ ;
 wire \register_file_i/rf_reg_580_ ;
 wire \register_file_i/rf_reg_581_ ;
 wire \register_file_i/rf_reg_582_ ;
 wire \register_file_i/rf_reg_583_ ;
 wire \register_file_i/rf_reg_584_ ;
 wire \register_file_i/rf_reg_585_ ;
 wire \register_file_i/rf_reg_586_ ;
 wire \register_file_i/rf_reg_587_ ;
 wire \register_file_i/rf_reg_588_ ;
 wire \register_file_i/rf_reg_589_ ;
 wire \register_file_i/rf_reg_58_ ;
 wire \register_file_i/rf_reg_590_ ;
 wire \register_file_i/rf_reg_591_ ;
 wire \register_file_i/rf_reg_592_ ;
 wire \register_file_i/rf_reg_593_ ;
 wire \register_file_i/rf_reg_594_ ;
 wire \register_file_i/rf_reg_595_ ;
 wire \register_file_i/rf_reg_596_ ;
 wire \register_file_i/rf_reg_597_ ;
 wire \register_file_i/rf_reg_598_ ;
 wire \register_file_i/rf_reg_599_ ;
 wire \register_file_i/rf_reg_59_ ;
 wire \register_file_i/rf_reg_600_ ;
 wire \register_file_i/rf_reg_601_ ;
 wire \register_file_i/rf_reg_602_ ;
 wire \register_file_i/rf_reg_603_ ;
 wire \register_file_i/rf_reg_604_ ;
 wire \register_file_i/rf_reg_605_ ;
 wire \register_file_i/rf_reg_606_ ;
 wire \register_file_i/rf_reg_607_ ;
 wire \register_file_i/rf_reg_608_ ;
 wire \register_file_i/rf_reg_609_ ;
 wire \register_file_i/rf_reg_60_ ;
 wire \register_file_i/rf_reg_610_ ;
 wire \register_file_i/rf_reg_611_ ;
 wire \register_file_i/rf_reg_612_ ;
 wire \register_file_i/rf_reg_613_ ;
 wire \register_file_i/rf_reg_614_ ;
 wire \register_file_i/rf_reg_615_ ;
 wire \register_file_i/rf_reg_616_ ;
 wire \register_file_i/rf_reg_617_ ;
 wire \register_file_i/rf_reg_618_ ;
 wire \register_file_i/rf_reg_619_ ;
 wire \register_file_i/rf_reg_61_ ;
 wire \register_file_i/rf_reg_620_ ;
 wire \register_file_i/rf_reg_621_ ;
 wire \register_file_i/rf_reg_622_ ;
 wire \register_file_i/rf_reg_623_ ;
 wire \register_file_i/rf_reg_624_ ;
 wire \register_file_i/rf_reg_625_ ;
 wire \register_file_i/rf_reg_626_ ;
 wire \register_file_i/rf_reg_627_ ;
 wire \register_file_i/rf_reg_628_ ;
 wire \register_file_i/rf_reg_629_ ;
 wire \register_file_i/rf_reg_62_ ;
 wire \register_file_i/rf_reg_630_ ;
 wire \register_file_i/rf_reg_631_ ;
 wire \register_file_i/rf_reg_632_ ;
 wire \register_file_i/rf_reg_633_ ;
 wire \register_file_i/rf_reg_634_ ;
 wire \register_file_i/rf_reg_635_ ;
 wire \register_file_i/rf_reg_636_ ;
 wire \register_file_i/rf_reg_637_ ;
 wire \register_file_i/rf_reg_638_ ;
 wire \register_file_i/rf_reg_639_ ;
 wire \register_file_i/rf_reg_63_ ;
 wire \register_file_i/rf_reg_640_ ;
 wire \register_file_i/rf_reg_641_ ;
 wire \register_file_i/rf_reg_642_ ;
 wire \register_file_i/rf_reg_643_ ;
 wire \register_file_i/rf_reg_644_ ;
 wire \register_file_i/rf_reg_645_ ;
 wire \register_file_i/rf_reg_646_ ;
 wire \register_file_i/rf_reg_647_ ;
 wire \register_file_i/rf_reg_648_ ;
 wire \register_file_i/rf_reg_649_ ;
 wire \register_file_i/rf_reg_64_ ;
 wire \register_file_i/rf_reg_650_ ;
 wire \register_file_i/rf_reg_651_ ;
 wire \register_file_i/rf_reg_652_ ;
 wire \register_file_i/rf_reg_653_ ;
 wire \register_file_i/rf_reg_654_ ;
 wire \register_file_i/rf_reg_655_ ;
 wire \register_file_i/rf_reg_656_ ;
 wire \register_file_i/rf_reg_657_ ;
 wire \register_file_i/rf_reg_658_ ;
 wire \register_file_i/rf_reg_659_ ;
 wire \register_file_i/rf_reg_65_ ;
 wire \register_file_i/rf_reg_660_ ;
 wire \register_file_i/rf_reg_661_ ;
 wire \register_file_i/rf_reg_662_ ;
 wire \register_file_i/rf_reg_663_ ;
 wire \register_file_i/rf_reg_664_ ;
 wire \register_file_i/rf_reg_665_ ;
 wire \register_file_i/rf_reg_666_ ;
 wire \register_file_i/rf_reg_667_ ;
 wire \register_file_i/rf_reg_668_ ;
 wire \register_file_i/rf_reg_669_ ;
 wire \register_file_i/rf_reg_66_ ;
 wire \register_file_i/rf_reg_670_ ;
 wire \register_file_i/rf_reg_671_ ;
 wire \register_file_i/rf_reg_672_ ;
 wire \register_file_i/rf_reg_673_ ;
 wire \register_file_i/rf_reg_674_ ;
 wire \register_file_i/rf_reg_675_ ;
 wire \register_file_i/rf_reg_676_ ;
 wire \register_file_i/rf_reg_677_ ;
 wire \register_file_i/rf_reg_678_ ;
 wire \register_file_i/rf_reg_679_ ;
 wire \register_file_i/rf_reg_67_ ;
 wire \register_file_i/rf_reg_680_ ;
 wire \register_file_i/rf_reg_681_ ;
 wire \register_file_i/rf_reg_682_ ;
 wire \register_file_i/rf_reg_683_ ;
 wire \register_file_i/rf_reg_684_ ;
 wire \register_file_i/rf_reg_685_ ;
 wire \register_file_i/rf_reg_686_ ;
 wire \register_file_i/rf_reg_687_ ;
 wire \register_file_i/rf_reg_688_ ;
 wire \register_file_i/rf_reg_689_ ;
 wire \register_file_i/rf_reg_68_ ;
 wire \register_file_i/rf_reg_690_ ;
 wire \register_file_i/rf_reg_691_ ;
 wire \register_file_i/rf_reg_692_ ;
 wire \register_file_i/rf_reg_693_ ;
 wire \register_file_i/rf_reg_694_ ;
 wire \register_file_i/rf_reg_695_ ;
 wire \register_file_i/rf_reg_696_ ;
 wire \register_file_i/rf_reg_697_ ;
 wire \register_file_i/rf_reg_698_ ;
 wire \register_file_i/rf_reg_699_ ;
 wire \register_file_i/rf_reg_69_ ;
 wire \register_file_i/rf_reg_700_ ;
 wire \register_file_i/rf_reg_701_ ;
 wire \register_file_i/rf_reg_702_ ;
 wire \register_file_i/rf_reg_703_ ;
 wire \register_file_i/rf_reg_704_ ;
 wire \register_file_i/rf_reg_705_ ;
 wire \register_file_i/rf_reg_706_ ;
 wire \register_file_i/rf_reg_707_ ;
 wire \register_file_i/rf_reg_708_ ;
 wire \register_file_i/rf_reg_709_ ;
 wire \register_file_i/rf_reg_70_ ;
 wire \register_file_i/rf_reg_710_ ;
 wire \register_file_i/rf_reg_711_ ;
 wire \register_file_i/rf_reg_712_ ;
 wire \register_file_i/rf_reg_713_ ;
 wire \register_file_i/rf_reg_714_ ;
 wire \register_file_i/rf_reg_715_ ;
 wire \register_file_i/rf_reg_716_ ;
 wire \register_file_i/rf_reg_717_ ;
 wire \register_file_i/rf_reg_718_ ;
 wire \register_file_i/rf_reg_719_ ;
 wire \register_file_i/rf_reg_71_ ;
 wire \register_file_i/rf_reg_720_ ;
 wire \register_file_i/rf_reg_721_ ;
 wire \register_file_i/rf_reg_722_ ;
 wire \register_file_i/rf_reg_723_ ;
 wire \register_file_i/rf_reg_724_ ;
 wire \register_file_i/rf_reg_725_ ;
 wire \register_file_i/rf_reg_726_ ;
 wire \register_file_i/rf_reg_727_ ;
 wire \register_file_i/rf_reg_728_ ;
 wire \register_file_i/rf_reg_729_ ;
 wire \register_file_i/rf_reg_72_ ;
 wire \register_file_i/rf_reg_730_ ;
 wire \register_file_i/rf_reg_731_ ;
 wire \register_file_i/rf_reg_732_ ;
 wire \register_file_i/rf_reg_733_ ;
 wire \register_file_i/rf_reg_734_ ;
 wire \register_file_i/rf_reg_735_ ;
 wire \register_file_i/rf_reg_736_ ;
 wire \register_file_i/rf_reg_737_ ;
 wire \register_file_i/rf_reg_738_ ;
 wire \register_file_i/rf_reg_739_ ;
 wire \register_file_i/rf_reg_73_ ;
 wire \register_file_i/rf_reg_740_ ;
 wire \register_file_i/rf_reg_741_ ;
 wire \register_file_i/rf_reg_742_ ;
 wire \register_file_i/rf_reg_743_ ;
 wire \register_file_i/rf_reg_744_ ;
 wire \register_file_i/rf_reg_745_ ;
 wire \register_file_i/rf_reg_746_ ;
 wire \register_file_i/rf_reg_747_ ;
 wire \register_file_i/rf_reg_748_ ;
 wire \register_file_i/rf_reg_749_ ;
 wire \register_file_i/rf_reg_74_ ;
 wire \register_file_i/rf_reg_750_ ;
 wire \register_file_i/rf_reg_751_ ;
 wire \register_file_i/rf_reg_752_ ;
 wire \register_file_i/rf_reg_753_ ;
 wire \register_file_i/rf_reg_754_ ;
 wire \register_file_i/rf_reg_755_ ;
 wire \register_file_i/rf_reg_756_ ;
 wire \register_file_i/rf_reg_757_ ;
 wire \register_file_i/rf_reg_758_ ;
 wire \register_file_i/rf_reg_759_ ;
 wire \register_file_i/rf_reg_75_ ;
 wire \register_file_i/rf_reg_760_ ;
 wire \register_file_i/rf_reg_761_ ;
 wire \register_file_i/rf_reg_762_ ;
 wire \register_file_i/rf_reg_763_ ;
 wire \register_file_i/rf_reg_764_ ;
 wire \register_file_i/rf_reg_765_ ;
 wire \register_file_i/rf_reg_766_ ;
 wire \register_file_i/rf_reg_767_ ;
 wire \register_file_i/rf_reg_768_ ;
 wire \register_file_i/rf_reg_769_ ;
 wire \register_file_i/rf_reg_76_ ;
 wire \register_file_i/rf_reg_770_ ;
 wire \register_file_i/rf_reg_771_ ;
 wire \register_file_i/rf_reg_772_ ;
 wire \register_file_i/rf_reg_773_ ;
 wire \register_file_i/rf_reg_774_ ;
 wire \register_file_i/rf_reg_775_ ;
 wire \register_file_i/rf_reg_776_ ;
 wire \register_file_i/rf_reg_777_ ;
 wire \register_file_i/rf_reg_778_ ;
 wire \register_file_i/rf_reg_779_ ;
 wire \register_file_i/rf_reg_77_ ;
 wire \register_file_i/rf_reg_780_ ;
 wire \register_file_i/rf_reg_781_ ;
 wire \register_file_i/rf_reg_782_ ;
 wire \register_file_i/rf_reg_783_ ;
 wire \register_file_i/rf_reg_784_ ;
 wire \register_file_i/rf_reg_785_ ;
 wire \register_file_i/rf_reg_786_ ;
 wire \register_file_i/rf_reg_787_ ;
 wire \register_file_i/rf_reg_788_ ;
 wire \register_file_i/rf_reg_789_ ;
 wire \register_file_i/rf_reg_78_ ;
 wire \register_file_i/rf_reg_790_ ;
 wire \register_file_i/rf_reg_791_ ;
 wire \register_file_i/rf_reg_792_ ;
 wire \register_file_i/rf_reg_793_ ;
 wire \register_file_i/rf_reg_794_ ;
 wire \register_file_i/rf_reg_795_ ;
 wire \register_file_i/rf_reg_796_ ;
 wire \register_file_i/rf_reg_797_ ;
 wire \register_file_i/rf_reg_798_ ;
 wire \register_file_i/rf_reg_799_ ;
 wire \register_file_i/rf_reg_79_ ;
 wire \register_file_i/rf_reg_800_ ;
 wire \register_file_i/rf_reg_801_ ;
 wire \register_file_i/rf_reg_802_ ;
 wire \register_file_i/rf_reg_803_ ;
 wire \register_file_i/rf_reg_804_ ;
 wire \register_file_i/rf_reg_805_ ;
 wire \register_file_i/rf_reg_806_ ;
 wire \register_file_i/rf_reg_807_ ;
 wire \register_file_i/rf_reg_808_ ;
 wire \register_file_i/rf_reg_809_ ;
 wire \register_file_i/rf_reg_80_ ;
 wire \register_file_i/rf_reg_810_ ;
 wire \register_file_i/rf_reg_811_ ;
 wire \register_file_i/rf_reg_812_ ;
 wire \register_file_i/rf_reg_813_ ;
 wire \register_file_i/rf_reg_814_ ;
 wire \register_file_i/rf_reg_815_ ;
 wire \register_file_i/rf_reg_816_ ;
 wire \register_file_i/rf_reg_817_ ;
 wire \register_file_i/rf_reg_818_ ;
 wire \register_file_i/rf_reg_819_ ;
 wire \register_file_i/rf_reg_81_ ;
 wire \register_file_i/rf_reg_820_ ;
 wire \register_file_i/rf_reg_821_ ;
 wire \register_file_i/rf_reg_822_ ;
 wire \register_file_i/rf_reg_823_ ;
 wire \register_file_i/rf_reg_824_ ;
 wire \register_file_i/rf_reg_825_ ;
 wire \register_file_i/rf_reg_826_ ;
 wire \register_file_i/rf_reg_827_ ;
 wire \register_file_i/rf_reg_828_ ;
 wire \register_file_i/rf_reg_829_ ;
 wire \register_file_i/rf_reg_82_ ;
 wire \register_file_i/rf_reg_830_ ;
 wire \register_file_i/rf_reg_831_ ;
 wire \register_file_i/rf_reg_832_ ;
 wire \register_file_i/rf_reg_833_ ;
 wire \register_file_i/rf_reg_834_ ;
 wire \register_file_i/rf_reg_835_ ;
 wire \register_file_i/rf_reg_836_ ;
 wire \register_file_i/rf_reg_837_ ;
 wire \register_file_i/rf_reg_838_ ;
 wire \register_file_i/rf_reg_839_ ;
 wire \register_file_i/rf_reg_83_ ;
 wire \register_file_i/rf_reg_840_ ;
 wire \register_file_i/rf_reg_841_ ;
 wire \register_file_i/rf_reg_842_ ;
 wire \register_file_i/rf_reg_843_ ;
 wire \register_file_i/rf_reg_844_ ;
 wire \register_file_i/rf_reg_845_ ;
 wire \register_file_i/rf_reg_846_ ;
 wire \register_file_i/rf_reg_847_ ;
 wire \register_file_i/rf_reg_848_ ;
 wire \register_file_i/rf_reg_849_ ;
 wire \register_file_i/rf_reg_84_ ;
 wire \register_file_i/rf_reg_850_ ;
 wire \register_file_i/rf_reg_851_ ;
 wire \register_file_i/rf_reg_852_ ;
 wire \register_file_i/rf_reg_853_ ;
 wire \register_file_i/rf_reg_854_ ;
 wire \register_file_i/rf_reg_855_ ;
 wire \register_file_i/rf_reg_856_ ;
 wire \register_file_i/rf_reg_857_ ;
 wire \register_file_i/rf_reg_858_ ;
 wire \register_file_i/rf_reg_859_ ;
 wire \register_file_i/rf_reg_85_ ;
 wire \register_file_i/rf_reg_860_ ;
 wire \register_file_i/rf_reg_861_ ;
 wire \register_file_i/rf_reg_862_ ;
 wire \register_file_i/rf_reg_863_ ;
 wire \register_file_i/rf_reg_864_ ;
 wire \register_file_i/rf_reg_865_ ;
 wire \register_file_i/rf_reg_866_ ;
 wire \register_file_i/rf_reg_867_ ;
 wire \register_file_i/rf_reg_868_ ;
 wire \register_file_i/rf_reg_869_ ;
 wire \register_file_i/rf_reg_86_ ;
 wire \register_file_i/rf_reg_870_ ;
 wire \register_file_i/rf_reg_871_ ;
 wire \register_file_i/rf_reg_872_ ;
 wire \register_file_i/rf_reg_873_ ;
 wire \register_file_i/rf_reg_874_ ;
 wire \register_file_i/rf_reg_875_ ;
 wire \register_file_i/rf_reg_876_ ;
 wire \register_file_i/rf_reg_877_ ;
 wire \register_file_i/rf_reg_878_ ;
 wire \register_file_i/rf_reg_879_ ;
 wire \register_file_i/rf_reg_87_ ;
 wire \register_file_i/rf_reg_880_ ;
 wire \register_file_i/rf_reg_881_ ;
 wire \register_file_i/rf_reg_882_ ;
 wire \register_file_i/rf_reg_883_ ;
 wire \register_file_i/rf_reg_884_ ;
 wire \register_file_i/rf_reg_885_ ;
 wire \register_file_i/rf_reg_886_ ;
 wire \register_file_i/rf_reg_887_ ;
 wire \register_file_i/rf_reg_888_ ;
 wire \register_file_i/rf_reg_889_ ;
 wire \register_file_i/rf_reg_88_ ;
 wire \register_file_i/rf_reg_890_ ;
 wire \register_file_i/rf_reg_891_ ;
 wire \register_file_i/rf_reg_892_ ;
 wire \register_file_i/rf_reg_893_ ;
 wire \register_file_i/rf_reg_894_ ;
 wire \register_file_i/rf_reg_895_ ;
 wire \register_file_i/rf_reg_896_ ;
 wire \register_file_i/rf_reg_897_ ;
 wire \register_file_i/rf_reg_898_ ;
 wire \register_file_i/rf_reg_899_ ;
 wire \register_file_i/rf_reg_89_ ;
 wire \register_file_i/rf_reg_900_ ;
 wire \register_file_i/rf_reg_901_ ;
 wire \register_file_i/rf_reg_902_ ;
 wire \register_file_i/rf_reg_903_ ;
 wire \register_file_i/rf_reg_904_ ;
 wire \register_file_i/rf_reg_905_ ;
 wire \register_file_i/rf_reg_906_ ;
 wire \register_file_i/rf_reg_907_ ;
 wire \register_file_i/rf_reg_908_ ;
 wire \register_file_i/rf_reg_909_ ;
 wire \register_file_i/rf_reg_90_ ;
 wire \register_file_i/rf_reg_910_ ;
 wire \register_file_i/rf_reg_911_ ;
 wire \register_file_i/rf_reg_912_ ;
 wire \register_file_i/rf_reg_913_ ;
 wire \register_file_i/rf_reg_914_ ;
 wire \register_file_i/rf_reg_915_ ;
 wire \register_file_i/rf_reg_916_ ;
 wire \register_file_i/rf_reg_917_ ;
 wire \register_file_i/rf_reg_918_ ;
 wire \register_file_i/rf_reg_919_ ;
 wire \register_file_i/rf_reg_91_ ;
 wire \register_file_i/rf_reg_920_ ;
 wire \register_file_i/rf_reg_921_ ;
 wire \register_file_i/rf_reg_922_ ;
 wire \register_file_i/rf_reg_923_ ;
 wire \register_file_i/rf_reg_924_ ;
 wire \register_file_i/rf_reg_925_ ;
 wire \register_file_i/rf_reg_926_ ;
 wire \register_file_i/rf_reg_927_ ;
 wire \register_file_i/rf_reg_928_ ;
 wire \register_file_i/rf_reg_929_ ;
 wire \register_file_i/rf_reg_92_ ;
 wire \register_file_i/rf_reg_930_ ;
 wire \register_file_i/rf_reg_931_ ;
 wire \register_file_i/rf_reg_932_ ;
 wire \register_file_i/rf_reg_933_ ;
 wire \register_file_i/rf_reg_934_ ;
 wire \register_file_i/rf_reg_935_ ;
 wire \register_file_i/rf_reg_936_ ;
 wire \register_file_i/rf_reg_937_ ;
 wire \register_file_i/rf_reg_938_ ;
 wire \register_file_i/rf_reg_939_ ;
 wire \register_file_i/rf_reg_93_ ;
 wire \register_file_i/rf_reg_940_ ;
 wire \register_file_i/rf_reg_941_ ;
 wire \register_file_i/rf_reg_942_ ;
 wire \register_file_i/rf_reg_943_ ;
 wire \register_file_i/rf_reg_944_ ;
 wire \register_file_i/rf_reg_945_ ;
 wire \register_file_i/rf_reg_946_ ;
 wire \register_file_i/rf_reg_947_ ;
 wire \register_file_i/rf_reg_948_ ;
 wire \register_file_i/rf_reg_949_ ;
 wire \register_file_i/rf_reg_94_ ;
 wire \register_file_i/rf_reg_950_ ;
 wire \register_file_i/rf_reg_951_ ;
 wire \register_file_i/rf_reg_952_ ;
 wire \register_file_i/rf_reg_953_ ;
 wire \register_file_i/rf_reg_954_ ;
 wire \register_file_i/rf_reg_955_ ;
 wire \register_file_i/rf_reg_956_ ;
 wire \register_file_i/rf_reg_957_ ;
 wire \register_file_i/rf_reg_958_ ;
 wire \register_file_i/rf_reg_959_ ;
 wire \register_file_i/rf_reg_95_ ;
 wire \register_file_i/rf_reg_960_ ;
 wire \register_file_i/rf_reg_961_ ;
 wire \register_file_i/rf_reg_962_ ;
 wire \register_file_i/rf_reg_963_ ;
 wire \register_file_i/rf_reg_964_ ;
 wire \register_file_i/rf_reg_965_ ;
 wire \register_file_i/rf_reg_966_ ;
 wire \register_file_i/rf_reg_967_ ;
 wire \register_file_i/rf_reg_968_ ;
 wire \register_file_i/rf_reg_969_ ;
 wire \register_file_i/rf_reg_96_ ;
 wire \register_file_i/rf_reg_970_ ;
 wire \register_file_i/rf_reg_971_ ;
 wire \register_file_i/rf_reg_972_ ;
 wire \register_file_i/rf_reg_973_ ;
 wire \register_file_i/rf_reg_974_ ;
 wire \register_file_i/rf_reg_975_ ;
 wire \register_file_i/rf_reg_976_ ;
 wire \register_file_i/rf_reg_977_ ;
 wire \register_file_i/rf_reg_978_ ;
 wire \register_file_i/rf_reg_979_ ;
 wire \register_file_i/rf_reg_97_ ;
 wire \register_file_i/rf_reg_980_ ;
 wire \register_file_i/rf_reg_981_ ;
 wire \register_file_i/rf_reg_982_ ;
 wire \register_file_i/rf_reg_983_ ;
 wire \register_file_i/rf_reg_984_ ;
 wire \register_file_i/rf_reg_985_ ;
 wire \register_file_i/rf_reg_986_ ;
 wire \register_file_i/rf_reg_987_ ;
 wire \register_file_i/rf_reg_988_ ;
 wire \register_file_i/rf_reg_989_ ;
 wire \register_file_i/rf_reg_98_ ;
 wire \register_file_i/rf_reg_990_ ;
 wire \register_file_i/rf_reg_991_ ;
 wire \register_file_i/rf_reg_992_ ;
 wire \register_file_i/rf_reg_993_ ;
 wire \register_file_i/rf_reg_994_ ;
 wire \register_file_i/rf_reg_995_ ;
 wire \register_file_i/rf_reg_996_ ;
 wire \register_file_i/rf_reg_997_ ;
 wire \register_file_i/rf_reg_998_ ;
 wire \register_file_i/rf_reg_999_ ;
 wire \register_file_i/rf_reg_99_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net8;
 wire net9;
 wire net10;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2470;
 wire net2487;
 wire net2488;
 wire net2489;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_38_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_55_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_80_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_leaf_105_clk_i;
 wire clknet_leaf_106_clk_i;
 wire clknet_leaf_107_clk_i;
 wire clknet_leaf_108_clk_i;
 wire clknet_leaf_109_clk_i;
 wire clknet_leaf_110_clk_i;
 wire clknet_leaf_111_clk_i;
 wire clknet_leaf_112_clk_i;
 wire clknet_leaf_113_clk_i;
 wire clknet_leaf_114_clk_i;
 wire clknet_leaf_115_clk_i;
 wire clknet_leaf_116_clk_i;
 wire clknet_leaf_117_clk_i;
 wire clknet_leaf_118_clk_i;
 wire clknet_leaf_119_clk_i;
 wire clknet_leaf_120_clk_i;
 wire clknet_leaf_121_clk_i;
 wire clknet_leaf_122_clk_i;
 wire clknet_leaf_123_clk_i;
 wire clknet_leaf_124_clk_i;
 wire clknet_leaf_125_clk_i;
 wire clknet_leaf_126_clk_i;
 wire clknet_leaf_127_clk_i;
 wire clknet_leaf_128_clk_i;
 wire clknet_leaf_129_clk_i;
 wire clknet_leaf_130_clk_i;
 wire clknet_leaf_131_clk_i;
 wire clknet_leaf_132_clk_i;
 wire clknet_leaf_133_clk_i;
 wire clknet_leaf_134_clk_i;
 wire clknet_leaf_135_clk_i;
 wire clknet_leaf_136_clk_i;
 wire clknet_leaf_137_clk_i;
 wire clknet_leaf_138_clk_i;
 wire clknet_leaf_139_clk_i;
 wire clknet_leaf_140_clk_i;
 wire clknet_leaf_141_clk_i;
 wire clknet_leaf_142_clk_i;
 wire clknet_leaf_143_clk_i;
 wire clknet_leaf_144_clk_i;
 wire clknet_leaf_145_clk_i;
 wire clknet_leaf_146_clk_i;
 wire clknet_leaf_147_clk_i;
 wire clknet_leaf_148_clk_i;
 wire clknet_leaf_149_clk_i;
 wire clknet_leaf_151_clk_i;
 wire clknet_leaf_152_clk_i;
 wire clknet_leaf_153_clk_i;
 wire clknet_leaf_154_clk_i;
 wire clknet_leaf_155_clk_i;
 wire clknet_leaf_156_clk_i;
 wire clknet_leaf_157_clk_i;
 wire clknet_leaf_158_clk_i;
 wire clknet_leaf_159_clk_i;
 wire clknet_leaf_160_clk_i;
 wire clknet_leaf_161_clk_i;
 wire clknet_leaf_162_clk_i;
 wire clknet_leaf_163_clk_i;
 wire clknet_leaf_164_clk_i;
 wire clknet_leaf_165_clk_i;
 wire clknet_leaf_166_clk_i;
 wire clknet_leaf_167_clk_i;
 wire clknet_leaf_168_clk_i;
 wire clknet_leaf_169_clk_i;
 wire clknet_leaf_170_clk_i;
 wire clknet_leaf_171_clk_i;
 wire clknet_leaf_172_clk_i;
 wire clknet_leaf_173_clk_i;
 wire clknet_leaf_174_clk_i;
 wire clknet_leaf_175_clk_i;
 wire clknet_leaf_176_clk_i;
 wire clknet_leaf_177_clk_i;
 wire clknet_leaf_178_clk_i;
 wire clknet_leaf_179_clk_i;
 wire clknet_leaf_180_clk_i;
 wire clknet_leaf_181_clk_i;
 wire clknet_leaf_183_clk_i;
 wire clknet_leaf_184_clk_i;
 wire clknet_leaf_185_clk_i;
 wire clknet_leaf_186_clk_i;
 wire clknet_leaf_187_clk_i;
 wire clknet_leaf_188_clk_i;
 wire clknet_leaf_189_clk_i;
 wire clknet_leaf_190_clk_i;
 wire clknet_leaf_191_clk_i;
 wire clknet_leaf_192_clk_i;
 wire clknet_leaf_193_clk_i;
 wire clknet_leaf_194_clk_i;
 wire clknet_leaf_195_clk_i;
 wire clknet_leaf_196_clk_i;
 wire clknet_leaf_197_clk_i;
 wire clknet_leaf_198_clk_i;
 wire clknet_leaf_199_clk_i;
 wire clknet_leaf_200_clk_i;
 wire clknet_leaf_201_clk_i;
 wire clknet_leaf_202_clk_i;
 wire clknet_leaf_203_clk_i;
 wire clknet_leaf_204_clk_i;
 wire clknet_leaf_205_clk_i;
 wire clknet_leaf_206_clk_i;
 wire clknet_leaf_207_clk_i;
 wire clknet_leaf_208_clk_i;
 wire clknet_leaf_209_clk_i;
 wire clknet_leaf_210_clk_i;
 wire clknet_leaf_211_clk_i;
 wire clknet_leaf_212_clk_i;
 wire clknet_leaf_213_clk_i;
 wire clknet_leaf_214_clk_i;
 wire clknet_leaf_215_clk_i;
 wire clknet_leaf_216_clk_i;
 wire clknet_leaf_217_clk_i;
 wire clknet_leaf_218_clk_i;
 wire clknet_leaf_219_clk_i;
 wire clknet_leaf_220_clk_i;
 wire clknet_leaf_221_clk_i;
 wire clknet_leaf_222_clk_i;
 wire clknet_leaf_223_clk_i;
 wire clknet_leaf_224_clk_i;
 wire clknet_leaf_225_clk_i;
 wire clknet_leaf_226_clk_i;
 wire clknet_leaf_228_clk_i;
 wire clknet_leaf_230_clk_i;
 wire clknet_leaf_231_clk_i;
 wire clknet_leaf_232_clk_i;
 wire clknet_leaf_233_clk_i;
 wire clknet_leaf_234_clk_i;
 wire clknet_leaf_235_clk_i;
 wire clknet_leaf_236_clk_i;
 wire clknet_leaf_237_clk_i;
 wire clknet_leaf_238_clk_i;
 wire clknet_leaf_239_clk_i;
 wire clknet_leaf_240_clk_i;
 wire clknet_leaf_241_clk_i;
 wire clknet_leaf_242_clk_i;
 wire clknet_leaf_243_clk_i;
 wire clknet_leaf_244_clk_i;
 wire clknet_leaf_245_clk_i;
 wire clknet_leaf_246_clk_i;
 wire clknet_leaf_247_clk_i;
 wire clknet_leaf_248_clk_i;
 wire clknet_leaf_249_clk_i;
 wire clknet_leaf_250_clk_i;
 wire clknet_leaf_251_clk_i;
 wire clknet_leaf_252_clk_i;
 wire clknet_leaf_253_clk_i;
 wire clknet_leaf_254_clk_i;
 wire clknet_leaf_255_clk_i;
 wire clknet_leaf_256_clk_i;
 wire clknet_leaf_257_clk_i;
 wire clknet_leaf_258_clk_i;
 wire clknet_leaf_259_clk_i;
 wire clknet_leaf_260_clk_i;
 wire clknet_leaf_261_clk_i;
 wire clknet_leaf_262_clk_i;
 wire clknet_leaf_263_clk_i;
 wire clknet_leaf_264_clk_i;
 wire clknet_leaf_265_clk_i;
 wire clknet_leaf_266_clk_i;
 wire clknet_leaf_267_clk_i;
 wire clknet_leaf_268_clk_i;
 wire clknet_leaf_269_clk_i;
 wire clknet_leaf_270_clk_i;
 wire clknet_leaf_271_clk_i;
 wire clknet_leaf_272_clk_i;
 wire clknet_leaf_273_clk_i;
 wire clknet_leaf_274_clk_i;
 wire clknet_leaf_275_clk_i;
 wire clknet_leaf_276_clk_i;
 wire clknet_leaf_277_clk_i;
 wire clknet_leaf_278_clk_i;
 wire clknet_leaf_279_clk_i;
 wire clknet_leaf_280_clk_i;
 wire clknet_leaf_281_clk_i;
 wire clknet_leaf_282_clk_i;
 wire clknet_leaf_283_clk_i;
 wire clknet_leaf_284_clk_i;
 wire clknet_leaf_285_clk_i;
 wire clknet_leaf_286_clk_i;
 wire clknet_leaf_287_clk_i;
 wire clknet_leaf_288_clk_i;
 wire clknet_leaf_289_clk_i;
 wire clknet_leaf_290_clk_i;
 wire clknet_leaf_291_clk_i;
 wire clknet_leaf_292_clk_i;
 wire clknet_leaf_293_clk_i;
 wire clknet_leaf_294_clk_i;
 wire clknet_leaf_295_clk_i;
 wire clknet_leaf_296_clk_i;
 wire clknet_leaf_297_clk_i;
 wire clknet_leaf_298_clk_i;
 wire clknet_leaf_299_clk_i;
 wire clknet_leaf_300_clk_i;
 wire clknet_leaf_301_clk_i;
 wire clknet_leaf_302_clk_i;
 wire clknet_leaf_303_clk_i;
 wire clknet_leaf_304_clk_i;
 wire clknet_leaf_305_clk_i;
 wire clknet_leaf_306_clk_i;
 wire clknet_leaf_307_clk_i;
 wire clknet_leaf_308_clk_i;
 wire clknet_leaf_309_clk_i;
 wire clknet_leaf_310_clk_i;
 wire clknet_leaf_311_clk_i;
 wire clknet_leaf_312_clk_i;
 wire clknet_leaf_313_clk_i;
 wire clknet_leaf_314_clk_i;
 wire clknet_leaf_315_clk_i;
 wire clknet_leaf_316_clk_i;
 wire clknet_leaf_317_clk_i;
 wire clknet_leaf_318_clk_i;
 wire clknet_leaf_319_clk_i;
 wire clknet_leaf_320_clk_i;
 wire clknet_leaf_321_clk_i;
 wire clknet_leaf_322_clk_i;
 wire clknet_leaf_323_clk_i;
 wire clknet_leaf_324_clk_i;
 wire clknet_leaf_325_clk_i;
 wire clknet_leaf_326_clk_i;
 wire clknet_leaf_327_clk_i;
 wire clknet_leaf_328_clk_i;
 wire clknet_leaf_329_clk_i;
 wire clknet_leaf_330_clk_i;
 wire clknet_leaf_331_clk_i;
 wire clknet_leaf_332_clk_i;
 wire clknet_leaf_333_clk_i;
 wire clknet_leaf_334_clk_i;
 wire clknet_leaf_335_clk_i;
 wire clknet_leaf_336_clk_i;
 wire clknet_leaf_337_clk_i;
 wire clknet_leaf_338_clk_i;
 wire clknet_leaf_339_clk_i;
 wire clknet_leaf_340_clk_i;
 wire clknet_leaf_341_clk_i;
 wire clknet_leaf_342_clk_i;
 wire clknet_0_clk_i;
 wire clknet_2_0_0_clk_i;
 wire clknet_2_1_0_clk_i;
 wire clknet_2_2_0_clk_i;
 wire clknet_2_3_0_clk_i;
 wire clknet_6_0_0_clk_i;
 wire clknet_6_1_0_clk_i;
 wire clknet_6_2_0_clk_i;
 wire clknet_6_3_0_clk_i;
 wire clknet_6_4_0_clk_i;
 wire clknet_6_5_0_clk_i;
 wire clknet_6_6_0_clk_i;
 wire clknet_6_7_0_clk_i;
 wire clknet_6_8_0_clk_i;
 wire clknet_6_9_0_clk_i;
 wire clknet_6_10_0_clk_i;
 wire clknet_6_11_0_clk_i;
 wire clknet_6_12_0_clk_i;
 wire clknet_6_13_0_clk_i;
 wire clknet_6_14_0_clk_i;
 wire clknet_6_15_0_clk_i;
 wire clknet_6_16_0_clk_i;
 wire clknet_6_17_0_clk_i;
 wire clknet_6_18_0_clk_i;
 wire clknet_6_19_0_clk_i;
 wire clknet_6_20_0_clk_i;
 wire clknet_6_21_0_clk_i;
 wire clknet_6_22_0_clk_i;
 wire clknet_6_23_0_clk_i;
 wire clknet_6_24_0_clk_i;
 wire clknet_6_25_0_clk_i;
 wire clknet_6_26_0_clk_i;
 wire clknet_6_27_0_clk_i;
 wire clknet_6_28_0_clk_i;
 wire clknet_6_29_0_clk_i;
 wire clknet_6_30_0_clk_i;
 wire clknet_6_31_0_clk_i;
 wire clknet_6_32_0_clk_i;
 wire clknet_6_33_0_clk_i;
 wire clknet_6_34_0_clk_i;
 wire clknet_6_35_0_clk_i;
 wire clknet_6_36_0_clk_i;
 wire clknet_6_37_0_clk_i;
 wire clknet_6_38_0_clk_i;
 wire clknet_6_39_0_clk_i;
 wire clknet_6_40_0_clk_i;
 wire clknet_6_41_0_clk_i;
 wire clknet_6_42_0_clk_i;
 wire clknet_6_43_0_clk_i;
 wire clknet_6_44_0_clk_i;
 wire clknet_6_45_0_clk_i;
 wire clknet_6_46_0_clk_i;
 wire clknet_6_47_0_clk_i;
 wire clknet_6_48_0_clk_i;
 wire clknet_6_49_0_clk_i;
 wire clknet_6_50_0_clk_i;
 wire clknet_6_51_0_clk_i;
 wire clknet_6_52_0_clk_i;
 wire clknet_6_53_0_clk_i;
 wire clknet_6_54_0_clk_i;
 wire clknet_6_55_0_clk_i;
 wire clknet_6_56_0_clk_i;
 wire clknet_6_57_0_clk_i;
 wire clknet_6_58_0_clk_i;
 wire clknet_6_59_0_clk_i;
 wire clknet_6_60_0_clk_i;
 wire clknet_6_61_0_clk_i;
 wire clknet_6_62_0_clk_i;
 wire clknet_6_63_0_clk_i;
 wire net2490;
 wire net2491;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;

 sg13g2_buf_2 fanout1333 (.A(_05234_),
    .X(net1333));
 sg13g2_buf_2 fanout1332 (.A(net1333),
    .X(net1332));
 sg13g2_nand2_2 _09107_ (.Y(_01130_),
    .A(net2094),
    .B(net2098));
 sg13g2_buf_2 fanout1331 (.A(net1333),
    .X(net1331));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(_05289_));
 sg13g2_nor2_2 _09110_ (.A(net2091),
    .B(net549),
    .Y(_01133_));
 sg13g2_nand2_1 _09111_ (.Y(_01134_),
    .A(_01130_),
    .B(_01133_));
 sg13g2_nor4_2 _09112_ (.A(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .B(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .C(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ),
    .Y(_01135_),
    .D(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(net1330));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(net1329));
 sg13g2_buf_2 fanout1327 (.A(_05568_),
    .X(net1327));
 sg13g2_nor3_2 _09116_ (.A(net1995),
    .B(\id_stage_i.controller_i.instr_i_4_ ),
    .C(net1996),
    .Y(_01139_));
 sg13g2_and2_1 _09117_ (.A(_01135_),
    .B(_01139_),
    .X(_01140_));
 sg13g2_or2_1 _09118_ (.X(_01141_),
    .B(\load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ),
    .A(\load_store_unit_i.ls_fsm_cs_2_ ));
 sg13g2_buf_2 fanout1326 (.A(net1327),
    .X(net1326));
 sg13g2_buf_1 fanout1325 (.A(_05568_),
    .X(net1325));
 sg13g2_or3_2 _09121_ (.A(\load_store_unit_i.busy_o_$_OR__Y_A_$_OR__A_B ),
    .B(net1977),
    .C(\load_store_unit_i.ls_fsm_cs_1_ ),
    .X(_01144_));
 sg13g2_nand2b_1 _09122_ (.Y(_01145_),
    .B(\load_store_unit_i.handle_misaligned_q ),
    .A_N(\load_store_unit_i.ls_fsm_cs_0__$_NOT__A_Y ));
 sg13g2_a22oi_1 _09123_ (.Y(_01146_),
    .B1(_01145_),
    .B2(net1977),
    .A2(_01144_),
    .A1(_01141_));
 sg13g2_a21o_1 _09124_ (.A2(_01140_),
    .A1(_01134_),
    .B1(net1718),
    .X(_01147_));
 sg13g2_buf_2 fanout1324 (.A(_05568_),
    .X(net1324));
 sg13g2_buf_2 fanout1323 (.A(_05660_),
    .X(net1323));
 sg13g2_buf_2 fanout1322 (.A(net1323),
    .X(net1322));
 sg13g2_buf_2 fanout1321 (.A(_05683_),
    .X(net1321));
 sg13g2_or4_2 _09129_ (.A(\id_stage_i.controller_i.instr_i_2_ ),
    .B(\id_stage_i.controller_i.instr_i_3_ ),
    .C(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .D(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .X(_01152_));
 sg13g2_nor4_2 _09130_ (.A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .B(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .C(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .Y(_01153_),
    .D(_01152_));
 sg13g2_inv_1 _09131_ (.Y(_01154_),
    .A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ));
 sg13g2_nor4_1 _09132_ (.A(\id_stage_i.controller_i.instr_i_2_ ),
    .B(net1998),
    .C(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .D(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .Y(_01155_));
 sg13g2_buf_2 fanout1320 (.A(_05683_),
    .X(net1320));
 sg13g2_o21ai_1 _09134_ (.B1(\id_stage_i.controller_i.instr_i_6_ ),
    .Y(_01157_),
    .A1(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .A2(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_and3_1 _09135_ (.X(_01158_),
    .A(_01154_),
    .B(net1906),
    .C(_01157_));
 sg13g2_nand2_2 _09136_ (.Y(_01159_),
    .A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .B(\id_stage_i.controller_i.instr_i_5_ ));
 sg13g2_o21ai_1 _09137_ (.B1(_01159_),
    .Y(_01160_),
    .A1(_01140_),
    .A2(_01158_));
 sg13g2_nor2_1 _09138_ (.A(\id_stage_i.controller_i.instr_i_6_ ),
    .B(net1997),
    .Y(_01161_));
 sg13g2_nand3_1 _09139_ (.B(net1906),
    .C(_01159_),
    .A(_01161_),
    .Y(_01162_));
 sg13g2_nor4_2 _09140_ (.A(net1998),
    .B(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .C(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .Y(_01163_),
    .D(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ));
 sg13g2_nor3_2 _09141_ (.A(\id_stage_i.controller_i.instr_i_6_ ),
    .B(net1996),
    .C(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .Y(_01164_));
 sg13g2_nand2_1 _09142_ (.Y(_01165_),
    .A(_01163_),
    .B(_01164_));
 sg13g2_nor2_1 _09143_ (.A(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .B(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .Y(_01166_));
 sg13g2_nor3_1 _09144_ (.A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .B(net1997),
    .C(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .Y(_01167_));
 sg13g2_nand2_1 _09145_ (.Y(_01168_),
    .A(net1998),
    .B(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ));
 sg13g2_o21ai_1 _09146_ (.B1(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ),
    .Y(_01169_),
    .A1(\id_stage_i.controller_i.instr_i_2_ ),
    .A2(net1998));
 sg13g2_nand4_1 _09147_ (.B(net429),
    .C(_01168_),
    .A(_01166_),
    .Y(_01170_),
    .D(_01169_));
 sg13g2_and3_1 _09148_ (.X(_01171_),
    .A(_01162_),
    .B(_01165_),
    .C(_01170_));
 sg13g2_a22oi_1 _09149_ (.Y(_01172_),
    .B1(_01160_),
    .B2(_01171_),
    .A2(net412),
    .A1(net2092));
 sg13g2_nand2b_1 _09150_ (.Y(_01173_),
    .B(_01172_),
    .A_N(_01147_));
 sg13g2_buf_2 fanout1319 (.A(_08425_),
    .X(net1319));
 sg13g2_buf_2 fanout1318 (.A(net1319),
    .X(net1318));
 sg13g2_a221oi_1 _09153_ (.B2(_01171_),
    .C1(_01147_),
    .B1(_01160_),
    .A1(net2092),
    .Y(_01176_),
    .A2(net412));
 sg13g2_and2_1 _09154_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .B(net1619),
    .X(_01177_));
 sg13g2_a21oi_1 _09155_ (.A1(crash_dump_o_32_),
    .A2(net1598),
    .Y(_01178_),
    .B1(_01177_));
 sg13g2_buf_2 fanout1317 (.A(net1318),
    .X(net1317));
 sg13g2_buf_2 fanout1316 (.A(net1319),
    .X(net1316));
 sg13g2_nor3_1 _09158_ (.A(net2089),
    .B(net549),
    .C(\id_stage_i.controller_i.instr_i_12_ ),
    .Y(_01181_));
 sg13g2_nand2_1 _09159_ (.Y(_01182_),
    .A(net2096),
    .B(_01181_));
 sg13g2_buf_2 fanout1315 (.A(net1316),
    .X(net1315));
 sg13g2_a21o_1 _09161_ (.A2(_01182_),
    .A1(_01139_),
    .B1(net429),
    .X(_01184_));
 sg13g2_nor2_1 _09162_ (.A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .B(net1997),
    .Y(_01185_));
 sg13g2_nand2b_1 _09163_ (.Y(_01186_),
    .B(_01185_),
    .A_N(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_and2_2 _09164_ (.A(net436),
    .B(\ex_block_i.alu_i.instr_first_cycle_i_$_AND__Y_B ),
    .X(_01187_));
 sg13g2_nor2_1 _09165_ (.A(_01186_),
    .B(_01187_),
    .Y(_01188_));
 sg13g2_inv_1 _09166_ (.Y(_01189_),
    .A(_01163_));
 sg13g2_nand2_2 _09167_ (.Y(_01190_),
    .A(net436),
    .B(\ex_block_i.alu_i.instr_first_cycle_i_$_AND__Y_B ));
 sg13g2_a21oi_1 _09168_ (.A1(net429),
    .A2(_01190_),
    .Y(_01191_),
    .B1(_01164_));
 sg13g2_nor2_1 _09169_ (.A(_01189_),
    .B(_01191_),
    .Y(_01192_));
 sg13g2_a221oi_1 _09170_ (.B2(net1905),
    .C1(_01192_),
    .B1(_01188_),
    .A1(_01135_),
    .Y(_01193_),
    .A2(_01184_));
 sg13g2_a21o_1 _09171_ (.A2(_01193_),
    .A1(_01172_),
    .B1(net1718),
    .X(_01194_));
 sg13g2_buf_2 fanout1314 (.A(\cs_registers_i/_0583_ ),
    .X(net1314));
 sg13g2_buf_4 fanout1313 (.X(net1313),
    .A(net1314));
 sg13g2_buf_4 fanout1312 (.X(net1312),
    .A(net1314));
 sg13g2_nand2b_2 _09175_ (.Y(_01198_),
    .B(_01133_),
    .A_N(net2098));
 sg13g2_nand2_1 _09176_ (.Y(_01199_),
    .A(net412),
    .B(net1716));
 sg13g2_nor2_1 _09177_ (.A(net1620),
    .B(net397),
    .Y(_01200_));
 sg13g2_buf_4 fanout1311 (.X(net1311),
    .A(net1312));
 sg13g2_a221oi_1 _09179_ (.B2(net2083),
    .C1(net1591),
    .B1(_01200_),
    .A1(crash_dump_o_96_),
    .Y(_01202_),
    .A2(net1620));
 sg13g2_a21oi_1 _09180_ (.A1(_01178_),
    .A2(net1589),
    .Y(alu_operand_a_ex_0_),
    .B1(_01202_));
 sg13g2_buf_2 fanout1310 (.A(net1311),
    .X(net1310));
 sg13g2_buf_4 fanout1309 (.X(net1309),
    .A(net1311));
 sg13g2_mux2_1 _09183_ (.A0(crash_dump_o_106_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ),
    .S(net1589),
    .X(_01205_));
 sg13g2_inv_1 _09184_ (.Y(_01206_),
    .A(_01205_));
 sg13g2_buf_4 fanout1308 (.X(net1308),
    .A(net1312));
 sg13g2_buf_2 fanout1307 (.A(\cs_registers_i/_1400_ ),
    .X(net1307));
 sg13g2_nand3_1 _09187_ (.B(net1594),
    .C(net1582),
    .A(crash_dump_o_42_),
    .Y(_01209_));
 sg13g2_o21ai_1 _09188_ (.B1(_01209_),
    .Y(_01210_),
    .A1(net1593),
    .A2(_01206_));
 sg13g2_buf_2 fanout1306 (.A(net1307),
    .X(net1306));
 sg13g2_mux2_1 _09190_ (.A0(crash_dump_o_43_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ),
    .S(net1619),
    .X(_01211_));
 sg13g2_inv_1 _09191_ (.Y(_01212_),
    .A(crash_dump_o_107_));
 sg13g2_nor3_1 _09192_ (.A(_01212_),
    .B(net1599),
    .C(net1589),
    .Y(_01213_));
 sg13g2_a21o_2 _09193_ (.A2(_01211_),
    .A1(net1589),
    .B1(_01213_),
    .X(_01214_));
 sg13g2_buf_2 fanout1305 (.A(net1306),
    .X(net1305));
 sg13g2_mux2_1 _09195_ (.A0(crash_dump_o_108_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ),
    .S(net1582),
    .X(_01215_));
 sg13g2_and3_1 _09196_ (.X(_01216_),
    .A(crash_dump_o_44_),
    .B(net1593),
    .C(net1582));
 sg13g2_a21o_2 _09197_ (.A2(_01215_),
    .A1(net1617),
    .B1(_01216_),
    .X(_01217_));
 sg13g2_buf_1 fanout1304 (.A(\cs_registers_i/_1400_ ),
    .X(net1304));
 sg13g2_mux2_1 _09199_ (.A0(crash_dump_o_109_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ),
    .S(net1584),
    .X(_01218_));
 sg13g2_inv_1 _09200_ (.Y(_01219_),
    .A(_01218_));
 sg13g2_nand3_1 _09201_ (.B(net1595),
    .C(net1586),
    .A(crash_dump_o_45_),
    .Y(_01220_));
 sg13g2_o21ai_1 _09202_ (.B1(_01220_),
    .Y(alu_operand_a_ex_13_),
    .A1(net1595),
    .A2(_01219_));
 sg13g2_mux2_1 _09203_ (.A0(crash_dump_o_110_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ),
    .S(net1584),
    .X(_01221_));
 sg13g2_nand2_1 _09204_ (.Y(_01222_),
    .A(net1617),
    .B(_01221_));
 sg13g2_nand3_1 _09205_ (.B(net1593),
    .C(net1584),
    .A(crash_dump_o_46_),
    .Y(_01223_));
 sg13g2_and2_2 _09206_ (.A(_01222_),
    .B(_01223_),
    .X(_01224_));
 sg13g2_inv_2 _09207_ (.Y(alu_operand_a_ex_14_),
    .A(_01224_));
 sg13g2_mux2_1 _09208_ (.A0(crash_dump_o_47_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ),
    .S(net1618),
    .X(_01225_));
 sg13g2_inv_2 _09209_ (.Y(_01226_),
    .A(crash_dump_o_111_));
 sg13g2_nor3_1 _09210_ (.A(_01226_),
    .B(net1595),
    .C(net1587),
    .Y(_01227_));
 sg13g2_a21oi_2 _09211_ (.B1(_01227_),
    .Y(_01228_),
    .A2(_01225_),
    .A1(net1586));
 sg13g2_inv_2 _09212_ (.Y(alu_operand_a_ex_15_),
    .A(_01228_));
 sg13g2_buf_1 fanout1303 (.A(net1304),
    .X(net1303));
 sg13g2_buf_2 fanout1302 (.A(net1304),
    .X(net1302));
 sg13g2_mux2_1 _09215_ (.A0(crash_dump_o_112_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .S(net1586),
    .X(_01231_));
 sg13g2_nand2_1 _09216_ (.Y(_01232_),
    .A(net1618),
    .B(_01231_));
 sg13g2_nand3_1 _09217_ (.B(net1596),
    .C(net1587),
    .A(crash_dump_o_48_),
    .Y(_01233_));
 sg13g2_and2_2 _09218_ (.A(_01232_),
    .B(_01233_),
    .X(_01234_));
 sg13g2_inv_2 _09219_ (.Y(alu_operand_a_ex_16_),
    .A(_01234_));
 sg13g2_buf_4 fanout1301 (.X(net1301),
    .A(net1304));
 sg13g2_mux2_1 _09221_ (.A0(crash_dump_o_113_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ),
    .S(net1587),
    .X(_01236_));
 sg13g2_inv_1 _09222_ (.Y(_01237_),
    .A(_01236_));
 sg13g2_buf_1 fanout1300 (.A(\cs_registers_i/_1400_ ),
    .X(net1300));
 sg13g2_nand3_1 _09224_ (.B(net1597),
    .C(net1588),
    .A(crash_dump_o_49_),
    .Y(_01239_));
 sg13g2_o21ai_1 _09225_ (.B1(_01239_),
    .Y(alu_operand_a_ex_17_),
    .A1(net1596),
    .A2(_01237_));
 sg13g2_inv_2 _09226_ (.Y(_01240_),
    .A(crash_dump_o_114_));
 sg13g2_nand2_1 _09227_ (.Y(_01241_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ),
    .B(net1587));
 sg13g2_o21ai_1 _09228_ (.B1(_01241_),
    .Y(_01242_),
    .A1(_01240_),
    .A2(net1587));
 sg13g2_inv_1 _09229_ (.Y(_01243_),
    .A(_01242_));
 sg13g2_nand3_1 _09230_ (.B(net1596),
    .C(net1588),
    .A(crash_dump_o_50_),
    .Y(_01244_));
 sg13g2_o21ai_1 _09231_ (.B1(_01244_),
    .Y(alu_operand_a_ex_18_),
    .A1(net1596),
    .A2(_01243_));
 sg13g2_mux2_1 _09232_ (.A0(crash_dump_o_115_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ),
    .S(net1583),
    .X(_01245_));
 sg13g2_inv_1 _09233_ (.Y(_01246_),
    .A(_01245_));
 sg13g2_nand3_1 _09234_ (.B(net1593),
    .C(net1583),
    .A(crash_dump_o_51_),
    .Y(_01247_));
 sg13g2_o21ai_1 _09235_ (.B1(_01247_),
    .Y(_01248_),
    .A1(net1593),
    .A2(_01246_));
 sg13g2_buf_2 fanout1299 (.A(net1300),
    .X(net1299));
 sg13g2_and2_1 _09237_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ),
    .B(net1620),
    .X(_01249_));
 sg13g2_a21oi_2 _09238_ (.B1(_01249_),
    .Y(_01250_),
    .A2(net1598),
    .A1(crash_dump_o_33_));
 sg13g2_a221oi_1 _09239_ (.B2(net531),
    .C1(net1591),
    .B1(_01200_),
    .A1(crash_dump_o_97_),
    .Y(_01251_),
    .A2(net1620));
 sg13g2_a21oi_2 _09240_ (.B1(_01251_),
    .Y(alu_operand_a_ex_1_),
    .A2(_01250_),
    .A1(net1591));
 sg13g2_mux2_1 _09241_ (.A0(crash_dump_o_116_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ),
    .S(net1586),
    .X(_01252_));
 sg13g2_inv_1 _09242_ (.Y(_01253_),
    .A(_01252_));
 sg13g2_nand3_1 _09243_ (.B(net1596),
    .C(net1586),
    .A(crash_dump_o_52_),
    .Y(_01254_));
 sg13g2_o21ai_1 _09244_ (.B1(_01254_),
    .Y(alu_operand_a_ex_20_),
    .A1(net1595),
    .A2(_01253_));
 sg13g2_inv_2 _09245_ (.Y(_01255_),
    .A(crash_dump_o_117_));
 sg13g2_nand2_1 _09246_ (.Y(_01256_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ),
    .B(net1590));
 sg13g2_o21ai_1 _09247_ (.B1(_01256_),
    .Y(_01257_),
    .A1(_01255_),
    .A2(net1590));
 sg13g2_inv_1 _09248_ (.Y(_01258_),
    .A(_01257_));
 sg13g2_nand3_1 _09249_ (.B(net1598),
    .C(net1590),
    .A(crash_dump_o_53_),
    .Y(_01259_));
 sg13g2_o21ai_1 _09250_ (.B1(_01259_),
    .Y(alu_operand_a_ex_21_),
    .A1(net1598),
    .A2(_01258_));
 sg13g2_mux2_1 _09251_ (.A0(crash_dump_o_118_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ),
    .S(net1586),
    .X(_01260_));
 sg13g2_inv_1 _09252_ (.Y(_01261_),
    .A(_01260_));
 sg13g2_nand3_1 _09253_ (.B(net1596),
    .C(net1587),
    .A(crash_dump_o_54_),
    .Y(_01262_));
 sg13g2_o21ai_1 _09254_ (.B1(_01262_),
    .Y(alu_operand_a_ex_22_),
    .A1(net1596),
    .A2(_01261_));
 sg13g2_nand2_1 _09255_ (.Y(_01263_),
    .A(crash_dump_o_119_),
    .B(net1618));
 sg13g2_mux2_1 _09256_ (.A0(crash_dump_o_55_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ),
    .S(net1618),
    .X(_01264_));
 sg13g2_nand2_1 _09257_ (.Y(_01265_),
    .A(net1586),
    .B(_01264_));
 sg13g2_o21ai_1 _09258_ (.B1(_01265_),
    .Y(alu_operand_a_ex_23_),
    .A1(net1587),
    .A2(_01263_));
 sg13g2_mux2_1 _09259_ (.A0(crash_dump_o_120_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ),
    .S(net1590),
    .X(_01266_));
 sg13g2_inv_1 _09260_ (.Y(_01267_),
    .A(_01266_));
 sg13g2_nand3_1 _09261_ (.B(net1598),
    .C(net1590),
    .A(crash_dump_o_56_),
    .Y(_01268_));
 sg13g2_o21ai_1 _09262_ (.B1(_01268_),
    .Y(alu_operand_a_ex_24_),
    .A1(net1598),
    .A2(_01267_));
 sg13g2_buf_2 fanout1298 (.A(net1299),
    .X(net1298));
 sg13g2_mux2_1 _09264_ (.A0(crash_dump_o_121_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ),
    .S(net1583),
    .X(_01270_));
 sg13g2_inv_1 _09265_ (.Y(_01271_),
    .A(_01270_));
 sg13g2_buf_2 fanout1297 (.A(net1298),
    .X(net1297));
 sg13g2_nand3_1 _09267_ (.B(net1597),
    .C(net1588),
    .A(crash_dump_o_57_),
    .Y(_01273_));
 sg13g2_o21ai_1 _09268_ (.B1(_01273_),
    .Y(alu_operand_a_ex_25_),
    .A1(net1597),
    .A2(_01271_));
 sg13g2_mux2_1 _09269_ (.A0(crash_dump_o_122_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ),
    .S(net1584),
    .X(_01274_));
 sg13g2_inv_1 _09270_ (.Y(_01275_),
    .A(_01274_));
 sg13g2_nand3_1 _09271_ (.B(net1594),
    .C(net1585),
    .A(crash_dump_o_58_),
    .Y(_01276_));
 sg13g2_o21ai_1 _09272_ (.B1(_01276_),
    .Y(alu_operand_a_ex_26_),
    .A1(net1594),
    .A2(_01275_));
 sg13g2_nand2_1 _09273_ (.Y(_01277_),
    .A(crash_dump_o_123_),
    .B(net1621));
 sg13g2_mux2_1 _09274_ (.A0(crash_dump_o_59_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ),
    .S(net1621),
    .X(_01278_));
 sg13g2_nand2_1 _09275_ (.Y(_01279_),
    .A(net1592),
    .B(_01278_));
 sg13g2_o21ai_1 _09276_ (.B1(_01279_),
    .Y(_01280_),
    .A1(net1590),
    .A2(_01277_));
 sg13g2_buf_2 fanout1296 (.A(net1298),
    .X(net1296));
 sg13g2_inv_2 _09278_ (.Y(_01281_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_28_ ));
 sg13g2_nand2_1 _09279_ (.Y(_01282_),
    .A(crash_dump_o_60_),
    .B(net1594));
 sg13g2_o21ai_1 _09280_ (.B1(_01282_),
    .Y(_01283_),
    .A1(_01281_),
    .A2(net1594));
 sg13g2_inv_2 _09281_ (.Y(_01284_),
    .A(crash_dump_o_124_));
 sg13g2_nor3_1 _09282_ (.A(_01284_),
    .B(net1594),
    .C(net1585),
    .Y(_01285_));
 sg13g2_a21o_2 _09283_ (.A2(_01283_),
    .A1(net1585),
    .B1(_01285_),
    .X(_01286_));
 sg13g2_buf_2 fanout1295 (.A(net1300),
    .X(net1295));
 sg13g2_nand2_1 _09285_ (.Y(_01287_),
    .A(crash_dump_o_125_),
    .B(net1617));
 sg13g2_mux2_1 _09286_ (.A0(crash_dump_o_61_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ),
    .S(net1617),
    .X(_01288_));
 sg13g2_nand2_1 _09287_ (.Y(_01289_),
    .A(net1585),
    .B(_01288_));
 sg13g2_o21ai_1 _09288_ (.B1(_01289_),
    .Y(_01290_),
    .A1(net1585),
    .A2(_01287_));
 sg13g2_buf_2 fanout1294 (.A(net1300),
    .X(net1294));
 sg13g2_and2_1 _09290_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ),
    .B(net1620),
    .X(_01291_));
 sg13g2_a21oi_1 _09291_ (.A1(crash_dump_o_34_),
    .A2(net1598),
    .Y(_01292_),
    .B1(_01291_));
 sg13g2_a221oi_1 _09292_ (.B2(net529),
    .C1(net1591),
    .B1(_01200_),
    .A1(crash_dump_o_98_),
    .Y(_01293_),
    .A2(net1620));
 sg13g2_a21oi_2 _09293_ (.B1(_01293_),
    .Y(alu_operand_a_ex_2_),
    .A2(_01292_),
    .A1(net1591));
 sg13g2_mux2_1 _09294_ (.A0(crash_dump_o_126_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ),
    .S(net1584),
    .X(_01294_));
 sg13g2_inv_1 _09295_ (.Y(_01295_),
    .A(_01294_));
 sg13g2_nand3_1 _09296_ (.B(net1595),
    .C(net1584),
    .A(crash_dump_o_62_),
    .Y(_01296_));
 sg13g2_o21ai_1 _09297_ (.B1(_01296_),
    .Y(alu_operand_a_ex_30_),
    .A1(net1595),
    .A2(_01295_));
 sg13g2_buf_2 fanout1293 (.A(net1294),
    .X(net1293));
 sg13g2_mux2_1 _09299_ (.A0(crash_dump_o_127_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .S(net1590),
    .X(_01298_));
 sg13g2_inv_1 _09300_ (.Y(_01299_),
    .A(_01298_));
 sg13g2_nand3_1 _09301_ (.B(net1599),
    .C(net1590),
    .A(crash_dump_o_63_),
    .Y(_01300_));
 sg13g2_o21ai_1 _09302_ (.B1(_01300_),
    .Y(alu_operand_a_ex_31_),
    .A1(net1599),
    .A2(_01299_));
 sg13g2_mux2_1 _09303_ (.A0(crash_dump_o_35_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .S(net1620),
    .X(_01301_));
 sg13g2_nor2b_1 _09304_ (.A(_01301_),
    .B_N(net1591),
    .Y(_01302_));
 sg13g2_a221oi_1 _09305_ (.B2(net2009),
    .C1(net1591),
    .B1(_01200_),
    .A1(crash_dump_o_99_),
    .Y(_01303_),
    .A2(net1620));
 sg13g2_nor2_2 _09306_ (.A(_01302_),
    .B(_01303_),
    .Y(alu_operand_a_ex_3_));
 sg13g2_and2_1 _09307_ (.A(net412),
    .B(net1716),
    .X(_01304_));
 sg13g2_buf_2 fanout1292 (.A(net1294),
    .X(net1292));
 sg13g2_and2_1 _09309_ (.A(\id_stage_i.controller_i.instr_i_19_ ),
    .B(net1676),
    .X(_01306_));
 sg13g2_mux4_1 _09310_ (.S0(net1598),
    .A0(crash_dump_o_100_),
    .A1(_01306_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ),
    .A3(crash_dump_o_36_),
    .S1(net1591),
    .X(_01307_));
 sg13g2_buf_4 fanout1291 (.X(net1291),
    .A(net1292));
 sg13g2_mux2_1 _09312_ (.A0(crash_dump_o_101_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ),
    .S(net1582),
    .X(_01308_));
 sg13g2_nand2_1 _09313_ (.Y(_01309_),
    .A(net1617),
    .B(_01308_));
 sg13g2_nand3_1 _09314_ (.B(net1593),
    .C(net1582),
    .A(crash_dump_o_37_),
    .Y(_01310_));
 sg13g2_nand2_2 _09315_ (.Y(alu_operand_a_ex_5_),
    .A(_01309_),
    .B(_01310_));
 sg13g2_mux2_1 _09316_ (.A0(crash_dump_o_102_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ),
    .S(net1582),
    .X(_01311_));
 sg13g2_nand2_1 _09317_ (.Y(_01312_),
    .A(net1617),
    .B(_01311_));
 sg13g2_nand3_1 _09318_ (.B(net1593),
    .C(net1582),
    .A(crash_dump_o_38_),
    .Y(_01313_));
 sg13g2_nand2_2 _09319_ (.Y(_01314_),
    .A(_01312_),
    .B(_01313_));
 sg13g2_buf_4 fanout1290 (.X(net1290),
    .A(\cs_registers_i/_1578_ ));
 sg13g2_mux2_1 _09321_ (.A0(crash_dump_o_103_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ),
    .S(net1582),
    .X(_01315_));
 sg13g2_nand2_1 _09322_ (.Y(_01316_),
    .A(net1617),
    .B(_01315_));
 sg13g2_nand3_1 _09323_ (.B(net1593),
    .C(net1583),
    .A(crash_dump_o_39_),
    .Y(_01317_));
 sg13g2_and2_2 _09324_ (.A(_01316_),
    .B(_01317_),
    .X(_01318_));
 sg13g2_inv_4 _09325_ (.A(_01318_),
    .Y(alu_operand_a_ex_7_));
 sg13g2_mux2_1 _09326_ (.A0(crash_dump_o_104_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ),
    .S(net1585),
    .X(_01319_));
 sg13g2_nand2_1 _09327_ (.Y(_01320_),
    .A(net1617),
    .B(_01319_));
 sg13g2_nand3_1 _09328_ (.B(net1594),
    .C(net1585),
    .A(crash_dump_o_40_),
    .Y(_01321_));
 sg13g2_and2_1 _09329_ (.A(_01320_),
    .B(_01321_),
    .X(_01322_));
 sg13g2_inv_2 _09330_ (.Y(alu_operand_a_ex_8_),
    .A(_01322_));
 sg13g2_mux2_1 _09331_ (.A0(crash_dump_o_105_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ),
    .S(net1589),
    .X(_01323_));
 sg13g2_inv_1 _09332_ (.Y(_01324_),
    .A(_01323_));
 sg13g2_nand3_1 _09333_ (.B(net1595),
    .C(net1586),
    .A(crash_dump_o_41_),
    .Y(_01325_));
 sg13g2_o21ai_1 _09334_ (.B1(_01325_),
    .Y(_01326_),
    .A1(net1595),
    .A2(_01324_));
 sg13g2_buf_4 fanout1289 (.X(net1289),
    .A(net1290));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1289));
 sg13g2_buf_4 fanout1287 (.X(net1287),
    .A(net1288));
 sg13g2_nor4_2 _09338_ (.A(net2103),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .Y(_01329_),
    .D(\id_stage_i.controller_i.ctrl_fsm_cs_2__$_NOT__A_Y ));
 sg13g2_buf_4 fanout1286 (.X(net1286),
    .A(net1290));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(net1290));
 sg13g2_buf_4 fanout1284 (.X(net1284),
    .A(net1285));
 sg13g2_a21oi_1 _09342_ (.A1(net548),
    .A2(net551),
    .Y(_01333_),
    .B1(net2088));
 sg13g2_o21ai_1 _09343_ (.B1(_01130_),
    .Y(_01334_),
    .A1(_01133_),
    .A2(_01333_));
 sg13g2_a22oi_1 _09344_ (.Y(_01335_),
    .B1(_01334_),
    .B2(net1905),
    .A2(net1716),
    .A1(_01163_));
 sg13g2_nor3_2 _09345_ (.A(net1998),
    .B(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .C(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .Y(_01336_));
 sg13g2_nor2_2 _09346_ (.A(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .B(\id_stage_i.controller_i.instr_i_2_ ),
    .Y(_01337_));
 sg13g2_a21oi_1 _09347_ (.A1(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .A2(net1995),
    .Y(_01338_),
    .B1(net1997));
 sg13g2_nand3_1 _09348_ (.B(_01337_),
    .C(_01338_),
    .A(_01336_),
    .Y(_01339_));
 sg13g2_nor2_2 _09349_ (.A(net1995),
    .B(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .Y(_01340_));
 sg13g2_nand3_1 _09350_ (.B(_01163_),
    .C(_01340_),
    .A(_01159_),
    .Y(_01341_));
 sg13g2_and2_1 _09351_ (.A(_01339_),
    .B(_01341_),
    .X(_01342_));
 sg13g2_nand2_1 _09352_ (.Y(_01343_),
    .A(_01139_),
    .B(net1905));
 sg13g2_o21ai_1 _09353_ (.B1(net429),
    .Y(_01344_),
    .A1(_01135_),
    .A2(_01163_));
 sg13g2_nand4_1 _09354_ (.B(_01342_),
    .C(_01343_),
    .A(_01160_),
    .Y(_01345_),
    .D(_01344_));
 sg13g2_o21ai_1 _09355_ (.B1(_01345_),
    .Y(_01346_),
    .A1(_01186_),
    .A2(_01335_));
 sg13g2_buf_4 fanout1283 (.X(net1283),
    .A(alu_operand_a_ex_14_));
 sg13g2_nor2_1 _09357_ (.A(net2003),
    .B(net2004),
    .Y(_01348_));
 sg13g2_buf_2 fanout1282 (.A(alu_operand_a_ex_20_),
    .X(net1282));
 sg13g2_buf_4 fanout1281 (.X(net1281),
    .A(alu_operand_a_ex_20_));
 sg13g2_buf_1 fanout1280 (.A(alu_operand_a_ex_8_),
    .X(net1280));
 sg13g2_buf_4 fanout1279 (.X(net1279),
    .A(alu_operand_a_ex_8_));
 sg13g2_buf_2 fanout1278 (.A(_02004_),
    .X(net1278));
 sg13g2_or4_1 _09363_ (.A(net2001),
    .B(\id_stage_i.controller_i.instr_i_27_ ),
    .C(\id_stage_i.controller_i.instr_i_28_ ),
    .D(\id_stage_i.controller_i.instr_i_29_ ),
    .X(_01354_));
 sg13g2_nor2_1 _09364_ (.A(net441),
    .B(_01354_),
    .Y(_01355_));
 sg13g2_buf_2 fanout1277 (.A(csr_addr_11_),
    .X(net1277));
 sg13g2_or3_2 _09366_ (.A(net2092),
    .B(net2096),
    .C(net550),
    .X(_01357_));
 sg13g2_a21oi_1 _09367_ (.A1(_01348_),
    .A2(_01355_),
    .Y(_01358_),
    .B1(_01357_));
 sg13g2_and2_1 _09368_ (.A(net441),
    .B(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .X(_01359_));
 sg13g2_nor2_1 _09369_ (.A(_01354_),
    .B(_01359_),
    .Y(_01360_));
 sg13g2_inv_2 _09370_ (.Y(_01361_),
    .A(net549));
 sg13g2_nor2_1 _09371_ (.A(net2086),
    .B(net2094),
    .Y(_01362_));
 sg13g2_nand2_1 _09372_ (.Y(_01363_),
    .A(_01361_),
    .B(_01362_));
 sg13g2_a21oi_1 _09373_ (.A1(_01348_),
    .A2(_01360_),
    .Y(_01364_),
    .B1(_01363_));
 sg13g2_nand2_2 _09374_ (.Y(_01365_),
    .A(net1905),
    .B(_01164_));
 sg13g2_inv_1 _09375_ (.Y(_01366_),
    .A(_01365_));
 sg13g2_o21ai_1 _09376_ (.B1(_01366_),
    .Y(_01367_),
    .A1(_01358_),
    .A2(_01364_));
 sg13g2_inv_1 _09377_ (.Y(_01368_),
    .A(net548));
 sg13g2_mux2_1 _09378_ (.A0(_01368_),
    .A1(net2096),
    .S(net2098),
    .X(_01369_));
 sg13g2_nor2_1 _09379_ (.A(net550),
    .B(_01369_),
    .Y(_01370_));
 sg13g2_o21ai_1 _09380_ (.B1(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .Y(_01371_),
    .A1(net1996),
    .A2(_01370_));
 sg13g2_or2_1 _09381_ (.X(_01372_),
    .B(net1997),
    .A(net1995));
 sg13g2_or2_2 _09382_ (.X(_01373_),
    .B(net549),
    .A(net2095));
 sg13g2_buf_2 fanout1276 (.A(csr_addr_3_),
    .X(net1276));
 sg13g2_a21o_1 _09384_ (.A2(net551),
    .A1(net548),
    .B1(net2097),
    .X(_01375_));
 sg13g2_a21oi_1 _09385_ (.A1(_01373_),
    .A2(_01375_),
    .Y(_01376_),
    .B1(net2090));
 sg13g2_nor3_1 _09386_ (.A(_01372_),
    .B(_01152_),
    .C(_01376_),
    .Y(_01377_));
 sg13g2_a221oi_1 _09387_ (.B2(_01377_),
    .C1(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .B1(_01371_),
    .A1(_01134_),
    .Y(_01378_),
    .A2(_01140_));
 sg13g2_nor4_2 _09388_ (.A(net2003),
    .B(net2002),
    .C(\id_stage_i.controller_i.instr_i_27_ ),
    .Y(_01379_),
    .D(\id_stage_i.controller_i.instr_i_30_ ));
 sg13g2_nor2_2 _09389_ (.A(\id_stage_i.controller_i.instr_i_28_ ),
    .B(\id_stage_i.controller_i.instr_i_29_ ),
    .Y(_01380_));
 sg13g2_and2_1 _09390_ (.A(_01379_),
    .B(_01380_),
    .X(_01381_));
 sg13g2_buf_2 fanout1275 (.A(net1276),
    .X(net1275));
 sg13g2_buf_2 fanout1274 (.A(csr_addr_4_),
    .X(net1274));
 sg13g2_o21ai_1 _09393_ (.B1(_01130_),
    .Y(_01384_),
    .A1(_01368_),
    .A2(_01361_));
 sg13g2_a221oi_1 _09394_ (.B2(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .C1(_01384_),
    .B1(net2005),
    .A1(net2089),
    .Y(_01385_),
    .A2(net2087));
 sg13g2_nor3_1 _09395_ (.A(net2003),
    .B(net2001),
    .C(\id_stage_i.controller_i.instr_i_27_ ),
    .Y(_01386_));
 sg13g2_nor3_1 _09396_ (.A(\id_stage_i.controller_i.instr_i_28_ ),
    .B(\id_stage_i.controller_i.instr_i_29_ ),
    .C(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .Y(_01387_));
 sg13g2_nand2_1 _09397_ (.Y(_01388_),
    .A(_01386_),
    .B(_01387_));
 sg13g2_nor2_1 _09398_ (.A(net2089),
    .B(net2098),
    .Y(_01389_));
 sg13g2_o21ai_1 _09399_ (.B1(_01361_),
    .Y(_01390_),
    .A1(_01362_),
    .A2(_01389_));
 sg13g2_nor3_1 _09400_ (.A(net2004),
    .B(_01388_),
    .C(_01390_),
    .Y(_01391_));
 sg13g2_a21oi_1 _09401_ (.A1(_01381_),
    .A2(_01385_),
    .Y(_01392_),
    .B1(_01391_));
 sg13g2_nor2_1 _09402_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.operator_i_0__$_MUX__Y_A_$_MUX__Y_S_$_OR__Y_B ),
    .B(_01373_),
    .Y(_01393_));
 sg13g2_and3_1 _09403_ (.X(_01394_),
    .A(_01336_),
    .B(_01340_),
    .C(_01337_));
 sg13g2_buf_2 fanout1273 (.A(csr_addr_4_),
    .X(net1273));
 sg13g2_o21ai_1 _09405_ (.B1(net411),
    .Y(_01396_),
    .A1(_01392_),
    .A2(_01393_));
 sg13g2_or2_2 _09406_ (.X(_01397_),
    .B(net2097),
    .A(net547));
 sg13g2_a22oi_1 _09407_ (.Y(_01398_),
    .B1(_01397_),
    .B2(net2096),
    .A2(net552),
    .A1(net548));
 sg13g2_nand2_1 _09408_ (.Y(_01399_),
    .A(net1716),
    .B(_01398_));
 sg13g2_nor2_1 _09409_ (.A(\id_stage_i.controller_i.instr_i_24_ ),
    .B(net2005),
    .Y(_01400_));
 sg13g2_nand2_2 _09410_ (.Y(_01401_),
    .A(_01400_),
    .B(_01379_));
 sg13g2_or4_1 _09411_ (.A(net2003),
    .B(net2002),
    .C(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .D(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .X(_01402_));
 sg13g2_or3_2 _09412_ (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__B_A ),
    .C(_01402_),
    .X(_01403_));
 sg13g2_nand2_1 _09413_ (.Y(_01404_),
    .A(_01401_),
    .B(_01403_));
 sg13g2_nor2_1 _09414_ (.A(\id_stage_i.controller_i.instr_i_19_ ),
    .B(net2083),
    .Y(_01405_));
 sg13g2_nor3_1 _09415_ (.A(net531),
    .B(net529),
    .C(net2009),
    .Y(_01406_));
 sg13g2_nand2_2 _09416_ (.Y(_01407_),
    .A(_01405_),
    .B(_01406_));
 sg13g2_inv_1 _09417_ (.Y(_01408_),
    .A(_01407_));
 sg13g2_nor2_2 _09418_ (.A(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .Y(_01409_));
 sg13g2_buf_2 fanout1272 (.A(csr_addr_5_),
    .X(net1272));
 sg13g2_buf_1 fanout1271 (.A(net1272),
    .X(net1271));
 sg13g2_nor4_2 _09421_ (.A(net464),
    .B(net442),
    .C(net2008),
    .Y(_01412_),
    .D(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_and2_1 _09422_ (.A(_01409_),
    .B(_01412_),
    .X(_01413_));
 sg13g2_nor2_1 _09423_ (.A(net448),
    .B(net2008),
    .Y(_01414_));
 sg13g2_nor4_1 _09424_ (.A(\id_stage_i.controller_i.instr_i_29_ ),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .C(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .D(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .Y(_01415_));
 sg13g2_nand2_1 _09425_ (.Y(_01416_),
    .A(_01414_),
    .B(_01415_));
 sg13g2_and2_1 _09426_ (.A(net464),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .X(_01417_));
 sg13g2_nor3_1 _09427_ (.A(net442),
    .B(net2007),
    .C(_01417_),
    .Y(_01418_));
 sg13g2_nand3b_1 _09428_ (.B(_01380_),
    .C(_01418_),
    .Y(_01419_),
    .A_N(net448));
 sg13g2_a21oi_1 _09429_ (.A1(_01416_),
    .A2(_01419_),
    .Y(_01420_),
    .B1(_01401_));
 sg13g2_or2_1 _09430_ (.X(_01421_),
    .B(_01420_),
    .A(_01413_));
 sg13g2_or3_1 _09431_ (.A(net1993),
    .B(net1992),
    .C(\id_stage_i.controller_i.instr_i_10_ ),
    .X(_01422_));
 sg13g2_nor4_1 _09432_ (.A(net553),
    .B(\id_stage_i.controller_i.instr_i_8_ ),
    .C(net1716),
    .D(_01422_),
    .Y(_01423_));
 sg13g2_nand4_1 _09433_ (.B(_01408_),
    .C(_01421_),
    .A(_01404_),
    .Y(_01424_),
    .D(_01423_));
 sg13g2_nand3_1 _09434_ (.B(_01399_),
    .C(_01424_),
    .A(net412),
    .Y(_01425_));
 sg13g2_nand4_1 _09435_ (.B(_01378_),
    .C(_01396_),
    .A(_01367_),
    .Y(_01426_),
    .D(_01425_));
 sg13g2_or2_1 _09436_ (.X(_01427_),
    .B(_01426_),
    .A(_01346_));
 sg13g2_buf_2 fanout1270 (.A(net1272),
    .X(net1270));
 sg13g2_inv_1 _09438_ (.Y(_01429_),
    .A(\id_stage_i.id_fsm_q ));
 sg13g2_and2_1 _09439_ (.A(net428),
    .B(_01168_),
    .X(_01430_));
 sg13g2_nor4_1 _09440_ (.A(net1996),
    .B(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ),
    .C(_01372_),
    .D(_01357_),
    .Y(_01431_));
 sg13g2_nor3_2 _09441_ (.A(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .B(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .C(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ),
    .Y(_01432_));
 sg13g2_o21ai_1 _09442_ (.B1(_01432_),
    .Y(_01433_),
    .A1(_01430_),
    .A2(_01431_));
 sg13g2_nand3_1 _09443_ (.B(\id_stage_i.instr_perf_count_id_o_$_AND__Y_B ),
    .C(net1904),
    .A(net436),
    .Y(_01434_));
 sg13g2_nor3_1 _09444_ (.A(_01190_),
    .B(_01433_),
    .C(_01434_),
    .Y(_01435_));
 sg13g2_nand3b_1 _09445_ (.B(_01429_),
    .C(_01435_),
    .Y(_01436_),
    .A_N(_01427_));
 sg13g2_nand2b_1 _09446_ (.Y(_01437_),
    .B(_01436_),
    .A_N(\id_stage_i.branch_set_raw ));
 sg13g2_nand3_1 _09447_ (.B(net1904),
    .C(_01437_),
    .A(\id_stage_i.branch_set_$_AND__Y_B ),
    .Y(_01438_));
 sg13g2_buf_1 fanout1269 (.A(csr_addr_6_),
    .X(net1269));
 sg13g2_buf_2 fanout1268 (.A(csr_addr_6_),
    .X(net1268));
 sg13g2_a21oi_1 _09450_ (.A1(net2103),
    .A2(net2104),
    .Y(_01441_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ));
 sg13g2_a21oi_1 _09451_ (.A1(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .A2(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .Y(_01442_),
    .B1(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ));
 sg13g2_nor3_2 _09452_ (.A(\id_stage_i.controller_i.exc_req_q ),
    .B(\id_stage_i.controller_i.store_err_q ),
    .C(\id_stage_i.controller_i.load_err_q ),
    .Y(_01443_));
 sg13g2_inv_2 _09453_ (.Y(_01444_),
    .A(debug_ebreaku));
 sg13g2_nor3_1 _09454_ (.A(_01444_),
    .B(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .C(net2116),
    .Y(_01445_));
 sg13g2_nand3_1 _09455_ (.B(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .C(net2116),
    .A(debug_ebreakm),
    .Y(_01446_));
 sg13g2_inv_1 _09456_ (.Y(_01447_),
    .A(_01446_));
 sg13g2_nor3_2 _09457_ (.A(debug_mode),
    .B(_01445_),
    .C(_01447_),
    .Y(_01448_));
 sg13g2_inv_1 _09458_ (.Y(_01449_),
    .A(_01401_));
 sg13g2_and2_2 _09459_ (.A(net412),
    .B(_01181_),
    .X(_01450_));
 sg13g2_and3_1 _09460_ (.X(_01451_),
    .A(net436),
    .B(_01449_),
    .C(_01450_));
 sg13g2_nor3_1 _09461_ (.A(net442),
    .B(\id_stage_i.controller_i.illegal_insn_q ),
    .C(\id_stage_i.controller_i.instr_fetch_err_i ),
    .Y(_01452_));
 sg13g2_and4_1 _09462_ (.A(_01451_),
    .B(_01380_),
    .C(_01414_),
    .D(_01452_),
    .X(_01453_));
 sg13g2_buf_2 fanout1267 (.A(net1269),
    .X(net1267));
 sg13g2_nand3b_1 _09464_ (.B(_01453_),
    .C(net513),
    .Y(_01455_),
    .A_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ));
 sg13g2_or2_1 _09465_ (.X(_01456_),
    .B(_01455_),
    .A(_01448_));
 sg13g2_or2_1 _09466_ (.X(_01457_),
    .B(_01456_),
    .A(_01443_));
 sg13g2_nand3_1 _09467_ (.B(_01450_),
    .C(_01413_),
    .A(net437),
    .Y(_01458_));
 sg13g2_nand2b_1 _09468_ (.Y(_01459_),
    .B(_01404_),
    .A_N(_01458_));
 sg13g2_inv_2 _09469_ (.Y(_01460_),
    .A(net2104));
 sg13g2_inv_1 _09470_ (.Y(_01461_),
    .A(\id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_nor2_2 _09471_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_2__$_NOT__A_Y ),
    .Y(_01462_));
 sg13g2_nand3_1 _09472_ (.B(_01461_),
    .C(_01462_),
    .A(_01460_),
    .Y(_01463_));
 sg13g2_a21oi_1 _09473_ (.A1(_01443_),
    .A2(_01459_),
    .Y(_01464_),
    .B1(_01463_));
 sg13g2_a21o_1 _09474_ (.A2(csr_mstatus_mie),
    .A1(irq_pending_o),
    .B1(irq_nm_i),
    .X(_01465_));
 sg13g2_nand3_1 _09475_ (.B(\id_stage_i.controller_i.handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .C(_01465_),
    .A(\debug_single_step_$_AND__B_A ),
    .Y(_01466_));
 sg13g2_nand2_2 _09476_ (.Y(_01467_),
    .A(_01461_),
    .B(_01462_));
 sg13g2_nor3_2 _09477_ (.A(net2103),
    .B(_01466_),
    .C(_01467_),
    .Y(exc_cause_6_));
 sg13g2_a221oi_1 _09478_ (.B2(_01464_),
    .C1(exc_cause_6_),
    .B1(_01457_),
    .A1(_01441_),
    .Y(_01468_),
    .A2(_01442_));
 sg13g2_and2_2 _09479_ (.A(_01438_),
    .B(_01468_),
    .X(_01469_));
 sg13g2_buf_2 fanout1266 (.A(_04123_),
    .X(net1266));
 sg13g2_inv_1 _09481_ (.Y(_01471_),
    .A(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ));
 sg13g2_inv_4 _09482_ (.A(net430),
    .Y(_01472_));
 sg13g2_buf_1 fanout1265 (.A(net1266),
    .X(net1265));
 sg13g2_nor2_1 _09484_ (.A(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .B(\if_stage_i.prefetch_buffer_i.fifo_busy_1_ ),
    .Y(_01474_));
 sg13g2_a21oi_2 _09485_ (.B1(_01474_),
    .Y(_01475_),
    .A2(_01472_),
    .A1(_01471_));
 sg13g2_inv_1 _09486_ (.Y(_01476_),
    .A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ));
 sg13g2_nand3b_1 _09487_ (.B(_01476_),
    .C(_01462_),
    .Y(_01477_),
    .A_N(net2102));
 sg13g2_buf_2 fanout1264 (.A(net1265),
    .X(net1264));
 sg13g2_nor2_1 _09489_ (.A(net2103),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .Y(_01479_));
 sg13g2_nor2_1 _09490_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_0_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_2__$_NOT__A_Y ),
    .Y(_01480_));
 sg13g2_nor2_1 _09491_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .Y(_01481_));
 sg13g2_o21ai_1 _09492_ (.B1(_01481_),
    .Y(_01482_),
    .A1(_01479_),
    .A2(_01480_));
 sg13g2_nand2_1 _09493_ (.Y(_01483_),
    .A(net2102),
    .B(net2104));
 sg13g2_nor3_2 _09494_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .C(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .Y(_01484_));
 sg13g2_and2_1 _09495_ (.A(_01483_),
    .B(_01484_),
    .X(_01485_));
 sg13g2_nor2_1 _09496_ (.A(net2102),
    .B(_01467_),
    .Y(_01486_));
 sg13g2_nor2_1 _09497_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 sg13g2_nand4_1 _09498_ (.B(_01477_),
    .C(_01482_),
    .A(_01463_),
    .Y(_01488_),
    .D(_01487_));
 sg13g2_nand2_1 _09499_ (.Y(_01489_),
    .A(\if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__Y_B ),
    .B(_01488_));
 sg13g2_a21oi_1 _09500_ (.A1(net113),
    .A2(_01475_),
    .Y(_01490_),
    .B1(_01489_));
 sg13g2_or2_2 _09501_ (.X(instr_req_o),
    .B(_01490_),
    .A(\if_stage_i.prefetch_buffer_i.valid_req_q ));
 sg13g2_nor2_1 _09502_ (.A(debug_single_step),
    .B(irq_nm_i),
    .Y(_01491_));
 sg13g2_nor4_1 _09503_ (.A(irq_pending_o),
    .B(net2103),
    .C(debug_req_i),
    .D(debug_mode),
    .Y(_01492_));
 sg13g2_nand2_1 _09504_ (.Y(_01493_),
    .A(_01491_),
    .B(_01492_));
 sg13g2_nand2_1 _09505_ (.Y(_01494_),
    .A(net2102),
    .B(_01460_));
 sg13g2_nor3_2 _09506_ (.A(\load_store_unit_i.ls_fsm_cs_2_ ),
    .B(\load_store_unit_i.ls_fsm_cs_0_ ),
    .C(\load_store_unit_i.ls_fsm_cs_1_ ),
    .Y(_01495_));
 sg13g2_nor3_2 _09507_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .C(\id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ),
    .Y(_01496_));
 sg13g2_nor2_2 _09508_ (.A(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .B(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ),
    .Y(_01497_));
 sg13g2_nand3_1 _09509_ (.B(_01496_),
    .C(_01497_),
    .A(_01495_),
    .Y(_01498_));
 sg13g2_a21oi_2 _09510_ (.B1(_01498_),
    .Y(_01499_),
    .A2(_01494_),
    .A1(_01493_));
 sg13g2_nand2b_2 _09511_ (.Y(core_busy_o),
    .B(_01499_),
    .A_N(instr_req_o));
 sg13g2_buf_2 fanout1263 (.A(net1265),
    .X(net1263));
 sg13g2_buf_2 fanout1262 (.A(net1265),
    .X(net1262));
 sg13g2_buf_2 fanout1261 (.A(net1265),
    .X(net1261));
 sg13g2_buf_2 fanout1260 (.A(net1266),
    .X(net1260));
 sg13g2_buf_2 fanout1259 (.A(_05526_),
    .X(net1259));
 sg13g2_buf_2 fanout1258 (.A(net1259),
    .X(net1258));
 sg13g2_and2_1 _09518_ (.A(instr_rvalid_i),
    .B(\if_stage_i.prefetch_buffer_i.fifo_i.in_valid_i_$_AND__Y_B ),
    .X(_01506_));
 sg13g2_buf_2 fanout1257 (.A(_05686_),
    .X(net1257));
 sg13g2_a21oi_1 _09520_ (.A1(net1983),
    .A2(_01506_),
    .Y(_01508_),
    .B1(net431));
 sg13g2_nor2_1 _09521_ (.A(net1984),
    .B(_01506_),
    .Y(_01509_));
 sg13g2_buf_1 fanout1256 (.A(_07262_),
    .X(net1256));
 sg13g2_buf_2 fanout1255 (.A(net1256),
    .X(net1255));
 sg13g2_inv_2 _09524_ (.Y(_01512_),
    .A(net1983));
 sg13g2_and2_1 _09525_ (.A(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ),
    .B(net1983),
    .X(_01513_));
 sg13g2_a21o_1 _09526_ (.A2(_01512_),
    .A1(instr_err_i),
    .B1(_01513_),
    .X(_01514_));
 sg13g2_nand3_1 _09527_ (.B(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16_ ),
    .C(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17_ ),
    .A(net1984),
    .Y(_01515_));
 sg13g2_nand3_1 _09528_ (.B(instr_rdata_i_16_),
    .C(instr_rdata_i_17_),
    .A(_01512_),
    .Y(_01516_));
 sg13g2_nand3b_1 _09529_ (.B(_01515_),
    .C(_01516_),
    .Y(_01517_),
    .A_N(_01514_));
 sg13g2_nand2_1 _09530_ (.Y(_01518_),
    .A(net558),
    .B(_01517_));
 sg13g2_mux2_2 _09531_ (.A0(_01508_),
    .A1(_01509_),
    .S(_01518_),
    .X(_01519_));
 sg13g2_nand2_1 _09532_ (.Y(_01520_),
    .A(_01483_),
    .B(_01496_));
 sg13g2_buf_2 fanout1254 (.A(net1255),
    .X(net1254));
 sg13g2_buf_2 fanout1253 (.A(net1256),
    .X(net1253));
 sg13g2_inv_1 _09535_ (.Y(_01523_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ));
 sg13g2_inv_2 _09536_ (.Y(_01524_),
    .A(net2088));
 sg13g2_a21oi_1 _09537_ (.A1(net2094),
    .A2(net548),
    .Y(_01525_),
    .B1(net2091));
 sg13g2_a22oi_1 _09538_ (.Y(_01526_),
    .B1(net2097),
    .B2(net2094),
    .A2(net551),
    .A1(net547));
 sg13g2_o21ai_1 _09539_ (.B1(_01526_),
    .Y(_01527_),
    .A1(_01524_),
    .A2(_01525_));
 sg13g2_nand2_2 _09540_ (.Y(_01528_),
    .A(_01379_),
    .B(_01380_));
 sg13g2_nor3_2 _09541_ (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .B(_01528_),
    .C(_01393_),
    .Y(_01529_));
 sg13g2_nand2_2 _09542_ (.Y(_01530_),
    .A(net411),
    .B(_01529_));
 sg13g2_nor2_2 _09543_ (.A(_01527_),
    .B(_01530_),
    .Y(_01531_));
 sg13g2_buf_2 fanout1252 (.A(net1253),
    .X(net1252));
 sg13g2_o21ai_1 _09545_ (.B1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .Y(_01533_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ),
    .A2(_01531_));
 sg13g2_buf_1 fanout1251 (.A(alu_operand_a_ex_17_),
    .X(net1251));
 sg13g2_nor2_2 _09547_ (.A(net2111),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(_01535_));
 sg13g2_inv_1 _09548_ (.Y(_01536_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(alu_operand_a_ex_17_));
 sg13g2_buf_4 fanout1249 (.X(net1249),
    .A(_01248_));
 sg13g2_buf_2 fanout1248 (.A(net1249),
    .X(net1248));
 sg13g2_nand2_2 _09552_ (.Y(_01540_),
    .A(net2091),
    .B(net2088));
 sg13g2_nor4_2 _09553_ (.A(net2003),
    .B(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .C(_01528_),
    .Y(_01541_),
    .D(_01384_));
 sg13g2_nand3_1 _09554_ (.B(_01540_),
    .C(_01541_),
    .A(net411),
    .Y(_01542_));
 sg13g2_buf_4 fanout1247 (.X(net1247),
    .A(_03061_));
 sg13g2_buf_2 fanout1246 (.A(csr_addr_0_),
    .X(net1246));
 sg13g2_buf_2 fanout1245 (.A(net1246),
    .X(net1245));
 sg13g2_buf_2 fanout1244 (.A(net1245),
    .X(net1244));
 sg13g2_buf_4 fanout1243 (.X(net1243),
    .A(net1244));
 sg13g2_buf_2 fanout1242 (.A(net1245),
    .X(net1242));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(net1242));
 sg13g2_buf_2 fanout1240 (.A(net1241),
    .X(net1240));
 sg13g2_buf_2 fanout1239 (.A(net1241),
    .X(net1239));
 sg13g2_a221oi_1 _09564_ (.B2(net1975),
    .C1(net368),
    .B1(_01535_),
    .A1(_01523_),
    .Y(_01552_),
    .A2(_01533_));
 sg13g2_and3_1 _09565_ (.X(_01553_),
    .A(net410),
    .B(_01540_),
    .C(_01541_));
 sg13g2_buf_2 fanout1238 (.A(net1242),
    .X(net1238));
 sg13g2_buf_4 fanout1237 (.X(net1237),
    .A(net1245));
 sg13g2_buf_1 fanout1236 (.A(net1237),
    .X(net1236));
 sg13g2_buf_4 fanout1235 (.X(net1235),
    .A(net1237));
 sg13g2_buf_4 fanout1234 (.X(net1234),
    .A(net1246));
 sg13g2_buf_2 fanout1233 (.A(net1246),
    .X(net1233));
 sg13g2_buf_4 fanout1232 (.X(net1232),
    .A(net1233));
 sg13g2_o21ai_1 _09573_ (.B1(net358),
    .Y(_01561_),
    .A1(\id_stage_i.id_fsm_q ),
    .A2(_01552_));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1232));
 sg13g2_buf_4 fanout1230 (.X(net1230),
    .A(_03959_));
 sg13g2_nor2_2 _09576_ (.A(net2466),
    .B(net1976),
    .Y(_01564_));
 sg13g2_nand2b_2 _09577_ (.Y(_01565_),
    .B(_01495_),
    .A_N(_01564_));
 sg13g2_nor2_2 _09578_ (.A(_01162_),
    .B(net1490),
    .Y(_01566_));
 sg13g2_mux2_1 _09579_ (.A0(_01552_),
    .A1(_01565_),
    .S(_01566_),
    .X(_01567_));
 sg13g2_or2_2 _09580_ (.X(_01568_),
    .B(net1490),
    .A(_01434_));
 sg13g2_inv_2 _09581_ (.Y(_01569_),
    .A(_01568_));
 sg13g2_o21ai_1 _09582_ (.B1(_01569_),
    .Y(_01570_),
    .A1(_01429_),
    .A2(_01567_));
 sg13g2_a21oi_2 _09583_ (.B1(_01570_),
    .Y(_01571_),
    .A2(_01561_),
    .A1(_01433_));
 sg13g2_or4_1 _09584_ (.A(_01460_),
    .B(net437),
    .C(\id_in_ready_$_AND__Y_A_$_AND__Y_A_$_AND__A_Y_$_AND__A_B ),
    .D(_01571_),
    .X(_01572_));
 sg13g2_inv_1 _09585_ (.Y(_01573_),
    .A(\debug_single_step_$_AND__B_A ));
 sg13g2_inv_1 _09586_ (.Y(_01574_),
    .A(\id_stage_i.controller_i.do_single_step_q ));
 sg13g2_nand3_1 _09587_ (.B(debug_single_step),
    .C(net436),
    .A(\debug_single_step_$_AND__B_A ),
    .Y(_01575_));
 sg13g2_o21ai_1 _09588_ (.B1(_01575_),
    .Y(\id_stage_i.controller_i.do_single_step_d ),
    .A1(net436),
    .A2(_01574_));
 sg13g2_nor2_1 _09589_ (.A(debug_req_i),
    .B(\id_stage_i.controller_i.do_single_step_d ),
    .Y(_01576_));
 sg13g2_nor2_1 _09590_ (.A(_01573_),
    .B(_01576_),
    .Y(\id_stage_i.controller_i.enter_debug_mode_prio_d ));
 sg13g2_a21oi_2 _09591_ (.B1(\id_stage_i.controller_i.enter_debug_mode_prio_d ),
    .Y(_01577_),
    .A2(net7),
    .A1(\debug_single_step_$_AND__B_A ));
 sg13g2_nand2_1 _09592_ (.Y(_01578_),
    .A(_01466_),
    .B(_01577_));
 sg13g2_nand4_1 _09593_ (.B(_01441_),
    .C(_01572_),
    .A(_01462_),
    .Y(_01579_),
    .D(_01578_));
 sg13g2_nand3_1 _09594_ (.B(_01520_),
    .C(_01579_),
    .A(_01463_),
    .Y(_01580_));
 sg13g2_nor2_1 _09595_ (.A(_01403_),
    .B(_01458_),
    .Y(_01581_));
 sg13g2_nor2_1 _09596_ (.A(net2104),
    .B(_01467_),
    .Y(_01582_));
 sg13g2_o21ai_1 _09597_ (.B1(net437),
    .Y(_01583_),
    .A1(\id_stage_i.illegal_csr_insn_i ),
    .A2(net1490));
 sg13g2_nand2_2 _09598_ (.Y(_01584_),
    .A(_01409_),
    .B(_01412_));
 sg13g2_and2_1 _09599_ (.A(_01414_),
    .B(_01415_),
    .X(_01585_));
 sg13g2_nand2_1 _09600_ (.Y(_01586_),
    .A(csr_mstatus_tw),
    .B(_01585_));
 sg13g2_a22oi_1 _09601_ (.Y(_01587_),
    .B1(_01584_),
    .B2(_01586_),
    .A2(net2116),
    .A1(\id_stage_i.controller_i.priv_mode_i_0_ ));
 sg13g2_a22oi_1 _09602_ (.Y(_01588_),
    .B1(_01587_),
    .B2(_01451_),
    .A2(_01581_),
    .A1(\debug_single_step_$_AND__B_A ));
 sg13g2_nand2_1 _09603_ (.Y(_01589_),
    .A(_01583_),
    .B(_01588_));
 sg13g2_and2_1 _09604_ (.A(net436),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ),
    .X(_01590_));
 sg13g2_nand3_1 _09605_ (.B(_01449_),
    .C(_01450_),
    .A(net437),
    .Y(_01591_));
 sg13g2_nor2_1 _09606_ (.A(_01591_),
    .B(_01419_),
    .Y(_01592_));
 sg13g2_nor3_1 _09607_ (.A(_01589_),
    .B(net1897),
    .C(_01592_),
    .Y(_01593_));
 sg13g2_nor2_1 _09608_ (.A(net395),
    .B(_01593_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 sg13g2_a21oi_1 _09609_ (.A1(_01584_),
    .A2(_01416_),
    .Y(_01594_),
    .B1(_01591_));
 sg13g2_or2_1 _09610_ (.X(_01595_),
    .B(net1976),
    .A(data_err_i));
 sg13g2_nor2_1 _09611_ (.A(\load_store_unit_i.lsu_err_q ),
    .B(_01595_),
    .Y(_01596_));
 sg13g2_nor2_1 _09612_ (.A(_01565_),
    .B(_01596_),
    .Y(_01597_));
 sg13g2_and2_1 _09613_ (.A(\load_store_unit_i.data_we_q ),
    .B(_01597_),
    .X(\id_stage_i.controller_i.store_err_i ));
 sg13g2_and2_1 _09614_ (.A(\load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ),
    .B(_01597_),
    .X(\id_stage_i.controller_i.load_err_i ));
 sg13g2_nor2_1 _09615_ (.A(\id_stage_i.controller_i.store_err_i ),
    .B(\id_stage_i.controller_i.load_err_i ),
    .Y(_01598_));
 sg13g2_inv_1 _09616_ (.Y(_01599_),
    .A(_01598_));
 sg13g2_or4_1 _09617_ (.A(_01581_),
    .B(\id_stage_i.controller_i.exc_req_d ),
    .C(_01594_),
    .D(_01599_),
    .X(_01600_));
 sg13g2_inv_1 _09618_ (.Y(_01601_),
    .A(_01600_));
 sg13g2_nand4_1 _09619_ (.B(_01130_),
    .C(net1676),
    .A(_01368_),
    .Y(_01602_),
    .D(_01407_));
 sg13g2_nor2_1 _09620_ (.A(net548),
    .B(_01407_),
    .Y(_01603_));
 sg13g2_a21o_1 _09621_ (.A2(net551),
    .A1(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .B1(net2095),
    .X(_01604_));
 sg13g2_or3_2 _09622_ (.A(net397),
    .B(_01603_),
    .C(_01604_),
    .X(_01605_));
 sg13g2_xnor2_1 _09623_ (.Y(_01606_),
    .A(_01602_),
    .B(_01605_));
 sg13g2_inv_1 _09624_ (.Y(_01607_),
    .A(_01414_));
 sg13g2_and2_1 _09625_ (.A(net442),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .X(_01608_));
 sg13g2_nor4_1 _09626_ (.A(net464),
    .B(_01401_),
    .C(_01607_),
    .D(_01608_),
    .Y(_01609_));
 sg13g2_nor2_1 _09627_ (.A(net2007),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(_01610_));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(net1230));
 sg13g2_nor2_1 _09629_ (.A(net2002),
    .B(\id_stage_i.controller_i.instr_i_27_ ),
    .Y(_01612_));
 sg13g2_nor4_1 _09630_ (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.operator_i_0__$_MUX__Y_A_$_MUX__Y_S_$_OR__Y_B ),
    .C(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .D(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .Y(_01613_));
 sg13g2_nand4_1 _09631_ (.B(_01610_),
    .C(_01612_),
    .A(_01400_),
    .Y(_01614_),
    .D(_01613_));
 sg13g2_o21ai_1 _09632_ (.B1(_01614_),
    .Y(_01615_),
    .A1(net441),
    .A2(_01402_));
 sg13g2_o21ai_1 _09633_ (.B1(_01409_),
    .Y(_01616_),
    .A1(_01609_),
    .A2(_01615_));
 sg13g2_nand2_1 _09634_ (.Y(_01617_),
    .A(net448),
    .B(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_nand3_1 _09635_ (.B(_01418_),
    .C(_01617_),
    .A(_01409_),
    .Y(_01618_));
 sg13g2_or4_1 _09636_ (.A(_01403_),
    .B(_01602_),
    .C(_01605_),
    .D(_01618_),
    .X(_01619_));
 sg13g2_o21ai_1 _09637_ (.B1(_01619_),
    .Y(_01620_),
    .A1(_01606_),
    .A2(_01616_));
 sg13g2_o21ai_1 _09638_ (.B1(net437),
    .Y(_01621_),
    .A1(\ex_block_i.alu_i.instr_first_cycle_i_$_AND__Y_B ),
    .A2(_01565_));
 sg13g2_inv_1 _09639_ (.Y(_01622_),
    .A(_01621_));
 sg13g2_a21oi_1 _09640_ (.A1(_01566_),
    .A2(_01622_),
    .Y(_01623_),
    .B1(_01571_));
 sg13g2_nand2_2 _09641_ (.Y(_01624_),
    .A(net1905),
    .B(net428));
 sg13g2_or3_2 _09642_ (.A(\load_store_unit_i.ls_fsm_cs_2_ ),
    .B(net1977),
    .C(\load_store_unit_i.ls_fsm_cs_1_ ),
    .X(_01625_));
 sg13g2_nor2_2 _09643_ (.A(_01625_),
    .B(_01564_),
    .Y(_01626_));
 sg13g2_nor2_1 _09644_ (.A(_01162_),
    .B(_01626_),
    .Y(_01627_));
 sg13g2_a21oi_1 _09645_ (.A1(_01162_),
    .A2(_01552_),
    .Y(_01628_),
    .B1(_01627_));
 sg13g2_nor4_1 _09646_ (.A(_01429_),
    .B(net1490),
    .C(_01624_),
    .D(_01628_),
    .Y(_01629_));
 sg13g2_or2_1 _09647_ (.X(_01630_),
    .B(net1490),
    .A(net396));
 sg13g2_nand2_2 _09648_ (.Y(_01631_),
    .A(_01483_),
    .B(_01484_));
 sg13g2_nand2_1 _09649_ (.Y(_01632_),
    .A(_01457_),
    .B(net395));
 sg13g2_nand3_1 _09650_ (.B(_01520_),
    .C(_01632_),
    .A(_01631_),
    .Y(_01633_));
 sg13g2_nor4_1 _09651_ (.A(_01434_),
    .B(_01629_),
    .C(net1403),
    .D(_01633_),
    .Y(_01634_));
 sg13g2_and2_1 _09652_ (.A(_01623_),
    .B(_01634_),
    .X(_01635_));
 sg13g2_nand3_1 _09653_ (.B(_01620_),
    .C(_01635_),
    .A(net437),
    .Y(_01636_));
 sg13g2_nand3_1 _09654_ (.B(_01165_),
    .C(_01170_),
    .A(_01162_),
    .Y(_01637_));
 sg13g2_and2_1 _09655_ (.A(_01336_),
    .B(_01340_),
    .X(_01638_));
 sg13g2_a21o_1 _09656_ (.A2(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ),
    .A1(\id_stage_i.controller_i.instr_i_2_ ),
    .B1(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .X(_01639_));
 sg13g2_o21ai_1 _09657_ (.B1(_01639_),
    .Y(_01640_),
    .A1(\id_stage_i.controller_i.instr_i_2_ ),
    .A2(net1996));
 sg13g2_a21o_1 _09658_ (.A2(_01640_),
    .A1(_01638_),
    .B1(_01140_),
    .X(_01641_));
 sg13g2_nor2_2 _09659_ (.A(_01637_),
    .B(_01641_),
    .Y(_01642_));
 sg13g2_a22oi_1 _09660_ (.Y(_01643_),
    .B1(_01387_),
    .B2(_01386_),
    .A2(_01380_),
    .A1(_01379_));
 sg13g2_nand3b_1 _09661_ (.B(_01379_),
    .C(_01380_),
    .Y(_01644_),
    .A_N(net2089));
 sg13g2_o21ai_1 _09662_ (.B1(_01644_),
    .Y(_01645_),
    .A1(net2086),
    .A2(_01643_));
 sg13g2_nor2_1 _09663_ (.A(net2004),
    .B(_01373_),
    .Y(_01646_));
 sg13g2_or3_1 _09664_ (.A(net2090),
    .B(net547),
    .C(net2097),
    .X(_01647_));
 sg13g2_or2_1 _09665_ (.X(_01648_),
    .B(net547),
    .A(net2094));
 sg13g2_a221oi_1 _09666_ (.B2(_01375_),
    .C1(net2004),
    .B1(_01648_),
    .A1(net2086),
    .Y(_01649_),
    .A2(_01647_));
 sg13g2_nor4_1 _09667_ (.A(net2090),
    .B(net2004),
    .C(net549),
    .D(net2097),
    .Y(_01650_));
 sg13g2_a221oi_1 _09668_ (.B2(net2094),
    .C1(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .B1(net2097),
    .A1(net548),
    .Y(_01651_),
    .A2(net551));
 sg13g2_o21ai_1 _09669_ (.B1(_01540_),
    .Y(_01652_),
    .A1(_01650_),
    .A2(_01651_));
 sg13g2_nand2b_1 _09670_ (.Y(_01653_),
    .B(_01652_),
    .A_N(_01649_));
 sg13g2_nor3_1 _09671_ (.A(net2004),
    .B(net1716),
    .C(_01388_),
    .Y(_01654_));
 sg13g2_a221oi_1 _09672_ (.B2(_01381_),
    .C1(_01654_),
    .B1(_01653_),
    .A1(_01645_),
    .Y(_01655_),
    .A2(_01646_));
 sg13g2_and2_1 _09673_ (.A(_01373_),
    .B(_01397_),
    .X(_01656_));
 sg13g2_nand2b_1 _09674_ (.Y(_01657_),
    .B(_01524_),
    .A_N(_01375_));
 sg13g2_o21ai_1 _09675_ (.B1(_01657_),
    .Y(_01658_),
    .A1(net2091),
    .A2(_01656_));
 sg13g2_nand3_1 _09676_ (.B(_01340_),
    .C(_01337_),
    .A(_01336_),
    .Y(_01659_));
 sg13g2_nor4_1 _09677_ (.A(net2003),
    .B(net2004),
    .C(_01659_),
    .D(_01528_),
    .Y(_01660_));
 sg13g2_nand2_1 _09678_ (.Y(_01661_),
    .A(_01658_),
    .B(_01660_));
 sg13g2_nand3_1 _09679_ (.B(net428),
    .C(_01187_),
    .A(net1905),
    .Y(_01662_));
 sg13g2_nor2_2 _09680_ (.A(_01334_),
    .B(_01662_),
    .Y(_01663_));
 sg13g2_nor2_2 _09681_ (.A(net2095),
    .B(net550),
    .Y(_01664_));
 sg13g2_nand2b_1 _09682_ (.Y(_01665_),
    .B(_01664_),
    .A_N(net2091));
 sg13g2_o21ai_1 _09683_ (.B1(_01665_),
    .Y(_01666_),
    .A1(net2086),
    .A2(_01656_));
 sg13g2_nor2_2 _09684_ (.A(_01365_),
    .B(_01527_),
    .Y(_01667_));
 sg13g2_a22oi_1 _09685_ (.Y(_01668_),
    .B1(_01667_),
    .B2(_01658_),
    .A2(_01666_),
    .A1(_01663_));
 sg13g2_o21ai_1 _09686_ (.B1(_01668_),
    .Y(_01669_),
    .A1(_01655_),
    .A2(_01661_));
 sg13g2_buf_2 fanout1228 (.A(net1229),
    .X(net1228));
 sg13g2_a22oi_1 _09688_ (.Y(_01671_),
    .B1(_01653_),
    .B2(_01381_),
    .A2(_01646_),
    .A1(_01645_));
 sg13g2_o21ai_1 _09689_ (.B1(net2086),
    .Y(_01672_),
    .A1(net2091),
    .A2(_01397_));
 sg13g2_nand3b_1 _09690_ (.B(_01660_),
    .C(_01672_),
    .Y(_01673_),
    .A_N(_01656_));
 sg13g2_nor3_1 _09691_ (.A(net2086),
    .B(net2095),
    .C(net551),
    .Y(_01674_));
 sg13g2_nor2b_1 _09692_ (.A(_01397_),
    .B_N(_01540_),
    .Y(_01675_));
 sg13g2_a21o_1 _09693_ (.A2(_01674_),
    .A1(_01355_),
    .B1(_01675_),
    .X(_01676_));
 sg13g2_nor2_1 _09694_ (.A(net1716),
    .B(_01388_),
    .Y(_01677_));
 sg13g2_and2_1 _09695_ (.A(_01348_),
    .B(net410),
    .X(_01678_));
 sg13g2_a21oi_1 _09696_ (.A1(_01524_),
    .A2(_01130_),
    .Y(_01679_),
    .B1(_01389_));
 sg13g2_nor3_1 _09697_ (.A(net550),
    .B(_01662_),
    .C(_01679_),
    .Y(_01680_));
 sg13g2_a221oi_1 _09698_ (.B2(_01678_),
    .C1(_01680_),
    .B1(_01677_),
    .A1(_01667_),
    .Y(_01681_),
    .A2(_01676_));
 sg13g2_o21ai_1 _09699_ (.B1(_01681_),
    .Y(_01682_),
    .A1(_01671_),
    .A2(_01673_));
 sg13g2_buf_2 fanout1227 (.A(_03959_),
    .X(net1227));
 sg13g2_xnor2_1 _09701_ (.Y(_01684_),
    .A(net1581),
    .B(net1580));
 sg13g2_nor2_1 _09702_ (.A(_01642_),
    .B(_01684_),
    .Y(_01685_));
 sg13g2_a221oi_1 _09703_ (.B2(_01655_),
    .C1(_01642_),
    .B1(net411),
    .A1(_01134_),
    .Y(_01686_),
    .A2(_01140_));
 sg13g2_inv_1 _09704_ (.Y(_01687_),
    .A(net2003));
 sg13g2_nor2_1 _09705_ (.A(net2004),
    .B(net548),
    .Y(_01688_));
 sg13g2_nand4_1 _09706_ (.B(_01380_),
    .C(_01389_),
    .A(_01379_),
    .Y(_01689_),
    .D(_01688_));
 sg13g2_nand2_1 _09707_ (.Y(_01690_),
    .A(_01687_),
    .B(_01689_));
 sg13g2_a21o_1 _09708_ (.A2(_01646_),
    .A1(_01645_),
    .B1(_01690_),
    .X(_01691_));
 sg13g2_a21oi_1 _09709_ (.A1(_01397_),
    .A2(_01604_),
    .Y(_01692_),
    .B1(net2089));
 sg13g2_nor2_1 _09710_ (.A(net2086),
    .B(_01373_),
    .Y(_01693_));
 sg13g2_o21ai_1 _09711_ (.B1(_01164_),
    .Y(_01694_),
    .A1(_01692_),
    .A2(_01693_));
 sg13g2_nand2_1 _09712_ (.Y(_01695_),
    .A(net429),
    .B(_01187_));
 sg13g2_a21oi_2 _09713_ (.B1(_01152_),
    .Y(_01696_),
    .A2(_01695_),
    .A1(_01694_));
 sg13g2_a21oi_2 _09714_ (.B1(_01696_),
    .Y(_01697_),
    .A2(_01691_),
    .A1(net410));
 sg13g2_or2_1 _09715_ (.X(_01698_),
    .B(net547),
    .A(net2091));
 sg13g2_nand2b_1 _09716_ (.Y(_01699_),
    .B(_01130_),
    .A_N(_01698_));
 sg13g2_o21ai_1 _09717_ (.B1(_01699_),
    .Y(_01700_),
    .A1(_01363_),
    .A2(_01360_));
 sg13g2_a22oi_1 _09718_ (.Y(_01701_),
    .B1(_01700_),
    .B2(_01667_),
    .A2(_01690_),
    .A1(net410));
 sg13g2_nand2_2 _09719_ (.Y(_01702_),
    .A(_01662_),
    .B(_01701_));
 sg13g2_or2_1 _09720_ (.X(_01703_),
    .B(_01662_),
    .A(_01334_));
 sg13g2_nor2_1 _09721_ (.A(_01190_),
    .B(_01624_),
    .Y(_01704_));
 sg13g2_nand2b_1 _09722_ (.Y(_01705_),
    .B(net547),
    .A_N(net2094));
 sg13g2_nand2b_1 _09723_ (.Y(_01706_),
    .B(net2094),
    .A_N(net2097));
 sg13g2_nand2b_1 _09724_ (.Y(_01707_),
    .B(net2091),
    .A_N(net549));
 sg13g2_a21oi_1 _09725_ (.A1(_01705_),
    .A2(_01706_),
    .Y(_01708_),
    .B1(_01707_));
 sg13g2_nor3_1 _09726_ (.A(net547),
    .B(_01361_),
    .C(_01706_),
    .Y(_01709_));
 sg13g2_o21ai_1 _09727_ (.B1(_01524_),
    .Y(_01710_),
    .A1(_01708_),
    .A2(_01709_));
 sg13g2_o21ai_1 _09728_ (.B1(_01361_),
    .Y(_01711_),
    .A1(_01354_),
    .A2(_01359_));
 sg13g2_a221oi_1 _09729_ (.B2(net547),
    .C1(net2095),
    .B1(_01711_),
    .A1(net2086),
    .Y(_01712_),
    .A2(_01698_));
 sg13g2_nand4_1 _09730_ (.B(_01380_),
    .C(_01362_),
    .A(_01379_),
    .Y(_01713_),
    .D(_01688_));
 sg13g2_a21oi_1 _09731_ (.A1(_01687_),
    .A2(_01713_),
    .Y(_01714_),
    .B1(_01659_));
 sg13g2_a221oi_1 _09732_ (.B2(_01667_),
    .C1(_01714_),
    .B1(_01712_),
    .A1(_01704_),
    .Y(_01715_),
    .A2(_01710_));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_and2_1 _09734_ (.A(_01703_),
    .B(_01715_),
    .X(_01717_));
 sg13g2_and4_1 _09735_ (.A(_01686_),
    .B(_01697_),
    .C(_01702_),
    .D(_01717_),
    .X(_01718_));
 sg13g2_or2_2 _09736_ (.X(_01719_),
    .B(_01641_),
    .A(_01637_));
 sg13g2_buf_2 fanout1225 (.A(net1226),
    .X(net1225));
 sg13g2_nand2_1 _09738_ (.Y(_01721_),
    .A(_01719_),
    .B(net1580));
 sg13g2_and2_2 _09739_ (.A(_01686_),
    .B(_01715_),
    .X(_01722_));
 sg13g2_inv_1 _09740_ (.Y(_01723_),
    .A(_01722_));
 sg13g2_nand2_2 _09741_ (.Y(_01724_),
    .A(_01719_),
    .B(_01669_));
 sg13g2_nand3_1 _09742_ (.B(_01723_),
    .C(_01724_),
    .A(net1562),
    .Y(_01725_));
 sg13g2_nand4_1 _09743_ (.B(net1581),
    .C(net1580),
    .A(_01719_),
    .Y(_01726_),
    .D(_01722_));
 sg13g2_nand2_1 _09744_ (.Y(_01727_),
    .A(_01725_),
    .B(_01726_));
 sg13g2_inv_1 _09745_ (.Y(_01728_),
    .A(_01686_));
 sg13g2_nand2_1 _09746_ (.Y(_01729_),
    .A(_01663_),
    .B(_01701_));
 sg13g2_nor3_1 _09747_ (.A(_01728_),
    .B(_01697_),
    .C(_01729_),
    .Y(_01730_));
 sg13g2_a22oi_1 _09748_ (.Y(_01731_),
    .B1(_01727_),
    .B2(_01730_),
    .A2(_01718_),
    .A1(_01685_));
 sg13g2_a21o_1 _09749_ (.A2(_01691_),
    .A1(net411),
    .B1(_01696_),
    .X(_01732_));
 sg13g2_and4_1 _09750_ (.A(_01703_),
    .B(net1580),
    .C(_01732_),
    .D(_01702_),
    .X(_01733_));
 sg13g2_nor3_1 _09751_ (.A(_01642_),
    .B(net1580),
    .C(_01729_),
    .Y(_01734_));
 sg13g2_o21ai_1 _09752_ (.B1(net1581),
    .Y(_01735_),
    .A1(_01733_),
    .A2(_01734_));
 sg13g2_or3_1 _09753_ (.A(net1581),
    .B(net1562),
    .C(_01729_),
    .X(_01736_));
 sg13g2_a21oi_2 _09754_ (.B1(_01723_),
    .Y(_01737_),
    .A2(_01736_),
    .A1(_01735_));
 sg13g2_inv_1 _09755_ (.Y(_01738_),
    .A(_01715_));
 sg13g2_nand2_1 _09756_ (.Y(_01739_),
    .A(_01738_),
    .B(_01702_));
 sg13g2_o21ai_1 _09757_ (.B1(_01686_),
    .Y(_01740_),
    .A1(_01697_),
    .A2(_01739_));
 sg13g2_nand4_1 _09758_ (.B(net1562),
    .C(_01724_),
    .A(_01703_),
    .Y(_01741_),
    .D(_01740_));
 sg13g2_nand2b_1 _09759_ (.Y(_01742_),
    .B(_01741_),
    .A_N(_01737_));
 sg13g2_inv_1 _09760_ (.Y(_01743_),
    .A(net1581));
 sg13g2_nor2_1 _09761_ (.A(_01642_),
    .B(_01743_),
    .Y(_01744_));
 sg13g2_nor2_1 _09762_ (.A(_01728_),
    .B(_01729_),
    .Y(_01745_));
 sg13g2_nand3_1 _09763_ (.B(_01744_),
    .C(_01745_),
    .A(_01738_),
    .Y(_01746_));
 sg13g2_nand3_1 _09764_ (.B(net1562),
    .C(_01724_),
    .A(_01718_),
    .Y(_01747_));
 sg13g2_o21ai_1 _09765_ (.B1(_01747_),
    .Y(_01748_),
    .A1(net1562),
    .A2(_01746_));
 sg13g2_nor2_2 _09766_ (.A(_01742_),
    .B(_01748_),
    .Y(_01749_));
 sg13g2_nand2b_1 _09767_ (.Y(_01750_),
    .B(net1562),
    .A_N(_01746_));
 sg13g2_and3_2 _09768_ (.X(_01751_),
    .A(_01731_),
    .B(_01749_),
    .C(_01750_));
 sg13g2_o21ai_1 _09769_ (.B1(_01715_),
    .Y(_01752_),
    .A1(_01743_),
    .A2(net1562));
 sg13g2_nand2b_1 _09770_ (.Y(_01753_),
    .B(_01697_),
    .A_N(_01669_));
 sg13g2_nand4_1 _09771_ (.B(_01682_),
    .C(_01686_),
    .A(_01703_),
    .Y(_01754_),
    .D(_01715_));
 sg13g2_nor2_1 _09772_ (.A(_01753_),
    .B(_01754_),
    .Y(_01755_));
 sg13g2_a21o_2 _09773_ (.A2(_01752_),
    .A1(_01745_),
    .B1(_01755_),
    .X(_01756_));
 sg13g2_inv_1 _09774_ (.Y(_01757_),
    .A(net1580));
 sg13g2_o21ai_1 _09775_ (.B1(_01719_),
    .Y(_01758_),
    .A1(net1581),
    .A2(net1580));
 sg13g2_a21oi_1 _09776_ (.A1(_01757_),
    .A2(_01718_),
    .Y(_01759_),
    .B1(_01758_));
 sg13g2_xnor2_1 _09777_ (.Y(_01760_),
    .A(_01715_),
    .B(_01697_));
 sg13g2_a21oi_1 _09778_ (.A1(_01702_),
    .A2(_01760_),
    .Y(_01761_),
    .B1(_01728_));
 sg13g2_nor3_2 _09779_ (.A(_01663_),
    .B(_01759_),
    .C(_01761_),
    .Y(_01762_));
 sg13g2_or3_1 _09780_ (.A(_01737_),
    .B(_01756_),
    .C(_01762_),
    .X(_01763_));
 sg13g2_buf_1 fanout1224 (.A(net1225),
    .X(net1224));
 sg13g2_buf_2 fanout1223 (.A(net1225),
    .X(net1223));
 sg13g2_buf_2 fanout1222 (.A(_04526_),
    .X(net1222));
 sg13g2_buf_2 fanout1221 (.A(_04767_),
    .X(net1221));
 sg13g2_buf_2 fanout1220 (.A(net1221),
    .X(net1220));
 sg13g2_buf_1 fanout1219 (.A(net1221),
    .X(net1219));
 sg13g2_nor2_1 _09787_ (.A(\load_store_unit_i.ls_fsm_cs_2_ ),
    .B(\load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ),
    .Y(_01770_));
 sg13g2_nor3_2 _09788_ (.A(\load_store_unit_i.busy_o_$_OR__Y_A_$_OR__A_B ),
    .B(net1977),
    .C(\load_store_unit_i.ls_fsm_cs_1_ ),
    .Y(_01771_));
 sg13g2_nand2_1 _09789_ (.Y(_01772_),
    .A(net1977),
    .B(_01145_));
 sg13g2_o21ai_1 _09790_ (.B1(_01772_),
    .Y(_01773_),
    .A1(_01770_),
    .A2(_01771_));
 sg13g2_nand2_1 _09791_ (.Y(_01774_),
    .A(_01336_),
    .B(_01337_));
 sg13g2_mux2_1 _09792_ (.A0(net2087),
    .A1(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .S(net1997),
    .X(_01775_));
 sg13g2_nor2_1 _09793_ (.A(net1995),
    .B(_01775_),
    .Y(_01776_));
 sg13g2_a21oi_1 _09794_ (.A1(net1995),
    .A2(_01185_),
    .Y(_01777_),
    .B1(_01776_));
 sg13g2_nor3_2 _09795_ (.A(_01188_),
    .B(_01774_),
    .C(_01777_),
    .Y(_01778_));
 sg13g2_and2_1 _09796_ (.A(_01773_),
    .B(net1613),
    .X(_01779_));
 sg13g2_buf_2 fanout1218 (.A(net1221),
    .X(net1218));
 sg13g2_buf_2 fanout1217 (.A(_07276_),
    .X(net1217));
 sg13g2_buf_1 fanout1216 (.A(net1217),
    .X(net1216));
 sg13g2_buf_1 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_nor4_2 _09801_ (.A(net2089),
    .B(net2095),
    .C(net550),
    .Y(_01784_),
    .D(net1996));
 sg13g2_a21oi_1 _09802_ (.A1(_01161_),
    .A2(_01784_),
    .Y(_01785_),
    .B1(net428));
 sg13g2_nand3b_1 _09803_ (.B(net429),
    .C(_01190_),
    .Y(_01786_),
    .A_N(net1998));
 sg13g2_o21ai_1 _09804_ (.B1(_01786_),
    .Y(_01787_),
    .A1(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ),
    .A2(_01785_));
 sg13g2_inv_1 _09805_ (.Y(_01788_),
    .A(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ));
 sg13g2_a22oi_1 _09806_ (.Y(_01789_),
    .B1(net428),
    .B2(_01168_),
    .A2(_01139_),
    .A1(_01788_));
 sg13g2_nand3_1 _09807_ (.B(_01341_),
    .C(_01789_),
    .A(_01339_),
    .Y(_01790_));
 sg13g2_and3_2 _09808_ (.X(_01791_),
    .A(_01432_),
    .B(_01787_),
    .C(_01790_));
 sg13g2_buf_2 fanout1214 (.A(net1216),
    .X(net1214));
 sg13g2_nor2_2 _09810_ (.A(net1718),
    .B(_01791_),
    .Y(_01793_));
 sg13g2_nand3_1 _09811_ (.B(net428),
    .C(_01190_),
    .A(_01135_),
    .Y(_01794_));
 sg13g2_a22oi_1 _09812_ (.Y(_01795_),
    .B1(net428),
    .B2(_01190_),
    .A2(_01340_),
    .A1(_01159_));
 sg13g2_a21o_1 _09813_ (.A2(_01794_),
    .A1(_01189_),
    .B1(_01795_),
    .X(_01796_));
 sg13g2_nand3_1 _09814_ (.B(_01336_),
    .C(_01337_),
    .A(net2087),
    .Y(_01797_));
 sg13g2_nand2_1 _09815_ (.Y(_01798_),
    .A(_01135_),
    .B(_01784_));
 sg13g2_a21o_1 _09816_ (.A2(_01798_),
    .A1(_01797_),
    .B1(_01372_),
    .X(_01799_));
 sg13g2_nand2b_1 _09817_ (.Y(_01800_),
    .B(_01432_),
    .A_N(_01789_));
 sg13g2_a221oi_1 _09818_ (.B2(_01342_),
    .C1(net1718),
    .B1(_01800_),
    .A1(_01796_),
    .Y(_01801_),
    .A2(_01799_));
 sg13g2_nand3_1 _09819_ (.B(net428),
    .C(_01190_),
    .A(net1905),
    .Y(_01802_));
 sg13g2_nand2_2 _09820_ (.Y(_01803_),
    .A(_01341_),
    .B(_01802_));
 sg13g2_nor2_2 _09821_ (.A(net1717),
    .B(net387),
    .Y(_01804_));
 sg13g2_nor2b_2 _09822_ (.A(net348),
    .B_N(_01804_),
    .Y(_01805_));
 sg13g2_o21ai_1 _09823_ (.B1(net2000),
    .Y(_01806_),
    .A1(_01793_),
    .A2(_01805_));
 sg13g2_nor2_1 _09824_ (.A(_01806_),
    .B(net332),
    .Y(_01807_));
 sg13g2_a21oi_2 _09825_ (.B1(_01807_),
    .Y(_01808_),
    .A2(net329),
    .A1(net288));
 sg13g2_nor2_2 _09826_ (.A(net81),
    .B(_01808_),
    .Y(_01809_));
 sg13g2_and2_1 _09827_ (.A(net81),
    .B(_01808_),
    .X(_01810_));
 sg13g2_nor2_1 _09828_ (.A(_01809_),
    .B(_01810_),
    .Y(_01811_));
 sg13g2_xnor2_1 _09829_ (.Y(_01812_),
    .A(net189),
    .B(_01811_));
 sg13g2_a21o_1 _09830_ (.A2(net331),
    .A1(net289),
    .B1(_01807_),
    .X(_01813_));
 sg13g2_nor3_2 _09831_ (.A(_01737_),
    .B(_01756_),
    .C(_01762_),
    .Y(_01814_));
 sg13g2_buf_1 fanout1213 (.A(net1216),
    .X(net1213));
 sg13g2_buf_2 fanout1212 (.A(net1216),
    .X(net1212));
 sg13g2_buf_1 fanout1211 (.A(_07369_),
    .X(net1211));
 sg13g2_buf_2 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sg13g2_buf_2 fanout1208 (.A(net1211),
    .X(net1208));
 sg13g2_buf_2 fanout1207 (.A(net1211),
    .X(net1207));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(\cs_registers_i/_1452_ ));
 sg13g2_nand2_1 _09840_ (.Y(_01823_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_32__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1974));
 sg13g2_o21ai_1 _09841_ (.B1(_01823_),
    .Y(_01824_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .A2(net2108));
 sg13g2_buf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sg13g2_nor2_1 _09843_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ),
    .B(net2110),
    .Y(_01826_));
 sg13g2_buf_2 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_4 fanout1203 (.X(net1203),
    .A(alu_operand_a_ex_18_));
 sg13g2_buf_4 fanout1202 (.X(net1202),
    .A(alu_operand_a_ex_25_));
 sg13g2_nor3_1 _09847_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0_ ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_1_ ),
    .Y(_01830_));
 sg13g2_nor3_2 _09848_ (.A(net2105),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ),
    .Y(_01831_));
 sg13g2_or2_1 _09849_ (.X(_01832_),
    .B(net1882),
    .A(net1888));
 sg13g2_buf_2 fanout1201 (.A(_01286_),
    .X(net1201));
 sg13g2_buf_4 fanout1200 (.X(net1200),
    .A(_01286_));
 sg13g2_buf_1 fanout1199 (.A(_01290_),
    .X(net1199));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(_01290_));
 sg13g2_buf_2 fanout1197 (.A(_08547_),
    .X(net1197));
 sg13g2_buf_2 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_or2_2 _09856_ (.X(_01839_),
    .B(net2110),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ));
 sg13g2_a21oi_2 _09857_ (.B1(_01839_),
    .Y(_01840_),
    .A2(net2107),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ));
 sg13g2_buf_2 fanout1195 (.A(_08547_),
    .X(net1195));
 sg13g2_buf_2 fanout1194 (.A(_08547_),
    .X(net1194));
 sg13g2_nor3_1 _09860_ (.A(net288),
    .B(net1712),
    .C(net403),
    .Y(_01843_));
 sg13g2_a221oi_1 _09861_ (.B2(\ex_block_i.alu_i.imd_val_q_i_31__$_NOT__A_Y ),
    .C1(_01843_),
    .B1(net403),
    .A1(_01824_),
    .Y(_01844_),
    .A2(net1894));
 sg13g2_o21ai_1 _09862_ (.B1(_01844_),
    .Y(_01845_),
    .A1(_01813_),
    .A2(net173));
 sg13g2_inv_2 _09863_ (.Y(_01846_),
    .A(\ex_block_i.alu_i.imd_val_q_i_63_ ));
 sg13g2_buf_2 fanout1193 (.A(\cs_registers_i/_0472_ ),
    .X(net1193));
 sg13g2_nor2_1 _09865_ (.A(net1888),
    .B(net1882),
    .Y(_01848_));
 sg13g2_buf_2 fanout1192 (.A(\cs_registers_i/_0472_ ),
    .X(net1192));
 sg13g2_nor3_1 _09867_ (.A(_01846_),
    .B(net367),
    .C(net1675),
    .Y(_01850_));
 sg13g2_nor3_1 _09868_ (.A(net367),
    .B(_01845_),
    .C(_01850_),
    .Y(_01851_));
 sg13g2_a21oi_1 _09869_ (.A1(_01845_),
    .A2(_01850_),
    .Y(_01852_),
    .B1(_01851_));
 sg13g2_o21ai_1 _09870_ (.B1(_01852_),
    .Y(_01853_),
    .A1(net353),
    .A2(_01812_));
 sg13g2_and3_1 _09871_ (.X(_01854_),
    .A(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .B(net357),
    .C(net403));
 sg13g2_a21oi_2 _09872_ (.B1(_01854_),
    .Y(_01855_),
    .A2(net379),
    .A1(net1190));
 sg13g2_inv_2 _09873_ (.Y(_01856_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ));
 sg13g2_a21o_1 _09874_ (.A2(_01803_),
    .A1(net348),
    .B1(_01791_),
    .X(_01857_));
 sg13g2_and2_2 _09875_ (.A(_01341_),
    .B(_01802_),
    .X(_01858_));
 sg13g2_nand2b_2 _09876_ (.Y(_01859_),
    .B(_01858_),
    .A_N(net347));
 sg13g2_nand2_2 _09877_ (.Y(_01860_),
    .A(_01857_),
    .B(_01859_));
 sg13g2_nand2_1 _09878_ (.Y(_01861_),
    .A(net2000),
    .B(_01860_));
 sg13g2_nor2_1 _09879_ (.A(net1718),
    .B(_01861_),
    .Y(_01862_));
 sg13g2_nor2_1 _09880_ (.A(net332),
    .B(_01862_),
    .Y(_01863_));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(\cs_registers_i/_0550_ ));
 sg13g2_and2_2 _09882_ (.A(net348),
    .B(net387),
    .X(_01865_));
 sg13g2_nand3_1 _09883_ (.B(_01793_),
    .C(_01865_),
    .A(net441),
    .Y(_01866_));
 sg13g2_a22oi_1 _09884_ (.Y(_01867_),
    .B1(_01863_),
    .B2(_01866_),
    .A2(net331),
    .A1(_01856_));
 sg13g2_nor2_2 _09885_ (.A(net350),
    .B(net187),
    .Y(_01868_));
 sg13g2_buf_4 fanout1190 (.X(net1190),
    .A(alu_operand_a_ex_30_));
 sg13g2_nand2_1 _09887_ (.Y(_01870_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_31__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _09888_ (.B1(_01870_),
    .Y(_01871_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ),
    .A2(net2108));
 sg13g2_nor3_1 _09889_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ),
    .B(net1712),
    .C(net403),
    .Y(_01872_));
 sg13g2_a221oi_1 _09890_ (.B2(net1894),
    .C1(_01872_),
    .B1(_01871_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_30__$_NOT__A_Y ),
    .Y(_01873_),
    .A2(net407));
 sg13g2_nand2b_1 _09891_ (.Y(_01874_),
    .B(net352),
    .A_N(_01873_));
 sg13g2_o21ai_1 _09892_ (.B1(_01874_),
    .Y(_01875_),
    .A1(net174),
    .A2(_01867_));
 sg13g2_a21oi_2 _09893_ (.B1(_01875_),
    .Y(_01876_),
    .A2(net110),
    .A1(_01867_));
 sg13g2_xnor2_1 _09894_ (.Y(_01877_),
    .A(_01855_),
    .B(_01876_));
 sg13g2_buf_1 fanout1189 (.A(_04036_),
    .X(net1189));
 sg13g2_buf_2 fanout1188 (.A(_04036_),
    .X(net1188));
 sg13g2_nand3_1 _09897_ (.B(_01787_),
    .C(_01790_),
    .A(_01432_),
    .Y(_01880_));
 sg13g2_buf_2 fanout1187 (.A(_04036_),
    .X(net1187));
 sg13g2_nor2_2 _09899_ (.A(net1717),
    .B(net1613),
    .Y(_01882_));
 sg13g2_nand2_2 _09900_ (.Y(_01883_),
    .A(net1612),
    .B(_01882_));
 sg13g2_inv_1 _09901_ (.Y(_01884_),
    .A(net1999));
 sg13g2_nor2_1 _09902_ (.A(_01884_),
    .B(net387),
    .Y(_01885_));
 sg13g2_a21oi_1 _09903_ (.A1(\id_stage_i.controller_i.instr_i_27_ ),
    .A2(_01865_),
    .Y(_01886_),
    .B1(_01885_));
 sg13g2_nor2_1 _09904_ (.A(_01883_),
    .B(_01886_),
    .Y(_01887_));
 sg13g2_buf_2 fanout1186 (.A(net1187),
    .X(net1186));
 sg13g2_nand2_1 _09906_ (.Y(_01889_),
    .A(_01791_),
    .B(net387));
 sg13g2_nand2_1 _09907_ (.Y(_01890_),
    .A(net2000),
    .B(_01882_));
 sg13g2_nor2_1 _09908_ (.A(net348),
    .B(_01890_),
    .Y(_01891_));
 sg13g2_a22oi_1 _09909_ (.Y(_01892_),
    .B1(_01889_),
    .B2(_01891_),
    .A2(net331),
    .A1(net1499));
 sg13g2_nor2b_2 _09910_ (.A(_01887_),
    .B_N(_01892_),
    .Y(_01893_));
 sg13g2_xnor2_1 _09911_ (.Y(_01894_),
    .A(net122),
    .B(_01893_));
 sg13g2_buf_2 fanout1185 (.A(net1187),
    .X(net1185));
 sg13g2_nand2b_2 _09913_ (.Y(_01896_),
    .B(_01892_),
    .A_N(_01887_));
 sg13g2_and3_1 _09914_ (.X(_01897_),
    .A(net122),
    .B(net186),
    .C(_01896_));
 sg13g2_a21oi_1 _09915_ (.A1(net181),
    .A2(_01894_),
    .Y(_01898_),
    .B1(_01897_));
 sg13g2_inv_2 _09916_ (.Y(_01899_),
    .A(\ex_block_i.alu_i.imd_val_q_i_59_ ));
 sg13g2_nor3_2 _09917_ (.A(_01899_),
    .B(net364),
    .C(net1674),
    .Y(_01900_));
 sg13g2_buf_2 fanout1184 (.A(_04401_),
    .X(net1184));
 sg13g2_buf_1 fanout1183 (.A(net1184),
    .X(net1183));
 sg13g2_buf_2 fanout1182 (.A(net1183),
    .X(net1182));
 sg13g2_buf_2 fanout1181 (.A(_05153_),
    .X(net1181));
 sg13g2_a21oi_1 _09922_ (.A1(net122),
    .A2(net381),
    .Y(_01905_),
    .B1(_01900_));
 sg13g2_inv_2 _09923_ (.Y(_01906_),
    .A(net2107));
 sg13g2_inv_1 _09924_ (.Y(_01907_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_a22oi_1 _09925_ (.Y(_01908_),
    .B1(net1881),
    .B2(_01907_),
    .A2(net1971),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_28__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nand2b_1 _09926_ (.Y(_01909_),
    .B(net1893),
    .A_N(_01908_));
 sg13g2_buf_2 fanout1180 (.A(_08434_),
    .X(net1180));
 sg13g2_buf_2 fanout1179 (.A(net1180),
    .X(net1179));
 sg13g2_buf_2 fanout1178 (.A(net1179),
    .X(net1178));
 sg13g2_nor3_1 _09930_ (.A(net1499),
    .B(net1709),
    .C(net405),
    .Y(_01913_));
 sg13g2_a21oi_1 _09931_ (.A1(\ex_block_i.alu_i.imd_val_q_i_27__$_NOT__A_Y ),
    .A2(net402),
    .Y(_01914_),
    .B1(_01913_));
 sg13g2_a21o_2 _09932_ (.A2(_01914_),
    .A1(_01909_),
    .B1(net380),
    .X(_01915_));
 sg13g2_nand2_1 _09933_ (.Y(_01916_),
    .A(_01915_),
    .B(_01896_));
 sg13g2_mux2_1 _09934_ (.A0(_01900_),
    .A1(_01905_),
    .S(_01916_),
    .X(_01917_));
 sg13g2_nor2_1 _09935_ (.A(net361),
    .B(net1674),
    .Y(_01918_));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(net1178));
 sg13g2_nand2_1 _09937_ (.Y(_01920_),
    .A(\ex_block_i.alu_i.imd_val_q_i_59_ ),
    .B(net1558));
 sg13g2_nand2_2 _09938_ (.Y(_01921_),
    .A(net123),
    .B(net371));
 sg13g2_nand2_2 _09939_ (.Y(_01922_),
    .A(_01920_),
    .B(_01921_));
 sg13g2_mux2_1 _09940_ (.A0(_01922_),
    .A1(_01920_),
    .S(_01915_),
    .X(_01923_));
 sg13g2_nand2_1 _09941_ (.Y(_01924_),
    .A(net181),
    .B(_01923_));
 sg13g2_o21ai_1 _09942_ (.B1(_01924_),
    .Y(_01925_),
    .A1(net173),
    .A2(_01917_));
 sg13g2_o21ai_1 _09943_ (.B1(_01925_),
    .Y(_01926_),
    .A1(net352),
    .A2(_01898_));
 sg13g2_buf_2 fanout1176 (.A(net1180),
    .X(net1176));
 sg13g2_buf_4 fanout1175 (.X(net1175),
    .A(net1180));
 sg13g2_a22oi_1 _09946_ (.Y(_01929_),
    .B1(net1557),
    .B2(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .A2(net380),
    .A1(net1200));
 sg13g2_inv_1 _09947_ (.Y(_01930_),
    .A(_01929_));
 sg13g2_nand2b_2 _09948_ (.Y(_01931_),
    .B(_01860_),
    .A_N(_01890_));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(\cs_registers_i/_0492_ ));
 sg13g2_nand2_2 _09950_ (.Y(_01933_),
    .A(net348),
    .B(net387));
 sg13g2_nor2_1 _09951_ (.A(_01933_),
    .B(_01883_),
    .Y(_01934_));
 sg13g2_a22oi_1 _09952_ (.Y(_01935_),
    .B1(_01934_),
    .B2(\id_stage_i.controller_i.instr_i_28_ ),
    .A2(net331),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ));
 sg13g2_nand2_1 _09953_ (.Y(_01936_),
    .A(_01931_),
    .B(_01935_));
 sg13g2_a22oi_1 _09954_ (.Y(_01937_),
    .B1(net1881),
    .B2(_01281_),
    .A2(net1971),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_29__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nand2b_1 _09955_ (.Y(_01938_),
    .B(net1893),
    .A_N(_01937_));
 sg13g2_nor3_1 _09956_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .B(net1709),
    .C(net402),
    .Y(_01939_));
 sg13g2_a21oi_1 _09957_ (.A1(\ex_block_i.alu_i.imd_val_q_i_28__$_NOT__A_Y ),
    .A2(net402),
    .Y(_01940_),
    .B1(_01939_));
 sg13g2_a21oi_2 _09958_ (.B1(net370),
    .Y(_01941_),
    .A2(_01940_),
    .A1(_01938_));
 sg13g2_inv_1 _09959_ (.Y(_01942_),
    .A(_01941_));
 sg13g2_o21ai_1 _09960_ (.B1(_01942_),
    .Y(_01943_),
    .A1(net175),
    .A2(net1346));
 sg13g2_xnor2_1 _09961_ (.Y(_01944_),
    .A(net1200),
    .B(net1346));
 sg13g2_o21ai_1 _09962_ (.B1(net180),
    .Y(_01945_),
    .A1(net352),
    .A2(_01944_));
 sg13g2_nand2_1 _09963_ (.Y(_01946_),
    .A(net1200),
    .B(net371));
 sg13g2_nand3_1 _09964_ (.B(_01946_),
    .C(net1346),
    .A(net189),
    .Y(_01947_));
 sg13g2_nand2_1 _09965_ (.Y(_01948_),
    .A(_01945_),
    .B(_01947_));
 sg13g2_a21oi_1 _09966_ (.A1(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .A2(net1557),
    .Y(_01949_),
    .B1(_01941_));
 sg13g2_a22oi_1 _09967_ (.Y(_01950_),
    .B1(_01948_),
    .B2(_01949_),
    .A2(_01943_),
    .A1(_01930_));
 sg13g2_nand2_1 _09968_ (.Y(_01951_),
    .A(_01926_),
    .B(_01950_));
 sg13g2_buf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sg13g2_nand2_1 _09970_ (.Y(_01953_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_30__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _09971_ (.B1(_01953_),
    .Y(_01954_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ),
    .A2(net2106));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(\cs_registers_i/_0542_ ));
 sg13g2_nor3_1 _09973_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .B(net1709),
    .C(net405),
    .Y(_01956_));
 sg13g2_a221oi_1 _09974_ (.B2(net1892),
    .C1(_01956_),
    .B1(_01954_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_29__$_NOT__A_Y ),
    .Y(_01957_),
    .A2(net409));
 sg13g2_nor2_2 _09975_ (.A(net373),
    .B(_01957_),
    .Y(_01958_));
 sg13g2_inv_4 _09976_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .Y(_01959_));
 sg13g2_buf_2 fanout1171 (.A(_08050_),
    .X(net1171));
 sg13g2_nor2_1 _09978_ (.A(_01791_),
    .B(_01933_),
    .Y(_01961_));
 sg13g2_nand2_1 _09979_ (.Y(_01962_),
    .A(\id_stage_i.controller_i.instr_i_29_ ),
    .B(_01961_));
 sg13g2_a21oi_2 _09980_ (.B1(_01778_),
    .Y(_01963_),
    .A2(_01860_),
    .A1(net2000));
 sg13g2_a221oi_1 _09981_ (.B2(_01963_),
    .C1(net1717),
    .B1(_01962_),
    .A1(_01959_),
    .Y(_01964_),
    .A2(net1614));
 sg13g2_buf_2 fanout1170 (.A(net1171),
    .X(net1170));
 sg13g2_nor2_1 _09983_ (.A(net174),
    .B(net1345),
    .Y(_01966_));
 sg13g2_o21ai_1 _09984_ (.B1(net1198),
    .Y(_01967_),
    .A1(_01958_),
    .A2(_01966_));
 sg13g2_nor2_1 _09985_ (.A(_01958_),
    .B(net1345),
    .Y(_01968_));
 sg13g2_mux2_1 _09986_ (.A0(_01968_),
    .A1(net1345),
    .S(net1198),
    .X(_01969_));
 sg13g2_nand2b_1 _09987_ (.Y(_01970_),
    .B(net1345),
    .A_N(_01958_));
 sg13g2_nor3_1 _09988_ (.A(net1198),
    .B(net179),
    .C(_01970_),
    .Y(_01971_));
 sg13g2_a21oi_1 _09989_ (.A1(net179),
    .A2(_01969_),
    .Y(_01972_),
    .B1(_01971_));
 sg13g2_and2_1 _09990_ (.A(net361),
    .B(_01972_),
    .X(_01973_));
 sg13g2_nand2_1 _09991_ (.Y(_01974_),
    .A(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .B(net398));
 sg13g2_and2_1 _09992_ (.A(net351),
    .B(_01974_),
    .X(_01975_));
 sg13g2_xor2_1 _09993_ (.B(_01974_),
    .A(_01958_),
    .X(_01976_));
 sg13g2_nor3_1 _09994_ (.A(net367),
    .B(_01966_),
    .C(_01976_),
    .Y(_01977_));
 sg13g2_a221oi_1 _09995_ (.B2(_01966_),
    .C1(_01977_),
    .B1(_01975_),
    .A1(_01967_),
    .Y(_01978_),
    .A2(_01973_));
 sg13g2_nor3_1 _09996_ (.A(_01877_),
    .B(_01951_),
    .C(_01978_),
    .Y(_01979_));
 sg13g2_buf_1 fanout1169 (.A(_08429_),
    .X(net1169));
 sg13g2_buf_1 fanout1168 (.A(net1169),
    .X(net1168));
 sg13g2_and3_1 _09999_ (.X(_01982_),
    .A(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .B(net359),
    .C(net402));
 sg13g2_a21oi_2 _10000_ (.B1(_01982_),
    .Y(_01983_),
    .A2(net379),
    .A1(net1202));
 sg13g2_nand2_1 _10001_ (.Y(_01984_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_26__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _10002_ (.B1(_01984_),
    .Y(_01985_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ),
    .A2(net2106));
 sg13g2_buf_2 fanout1167 (.A(net1168),
    .X(net1167));
 sg13g2_nor3_1 _10004_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_25_ ),
    .B(net1710),
    .C(net402),
    .Y(_01987_));
 sg13g2_a221oi_1 _10005_ (.B2(net1892),
    .C1(_01987_),
    .B1(_01985_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_25__$_NOT__A_Y ),
    .Y(_01988_),
    .A2(net406));
 sg13g2_nor2_1 _10006_ (.A(net365),
    .B(_01988_),
    .Y(_01989_));
 sg13g2_inv_4 _10007_ (.A(net1496),
    .Y(_01990_));
 sg13g2_nand3_1 _10008_ (.B(_01793_),
    .C(_01865_),
    .A(net2006),
    .Y(_01991_));
 sg13g2_o21ai_1 _10009_ (.B1(_01773_),
    .Y(_01992_),
    .A1(net1614),
    .A2(_01889_));
 sg13g2_a221oi_1 _10010_ (.B2(_01991_),
    .C1(_01992_),
    .B1(_01863_),
    .A1(_01990_),
    .Y(_01993_),
    .A2(net1614));
 sg13g2_nand2b_1 _10011_ (.Y(_01994_),
    .B(_01993_),
    .A_N(_01989_));
 sg13g2_a21oi_1 _10012_ (.A1(net365),
    .A2(_01993_),
    .Y(_01995_),
    .B1(_01989_));
 sg13g2_nand2_1 _10013_ (.Y(_01996_),
    .A(net179),
    .B(_01995_));
 sg13g2_o21ai_1 _10014_ (.B1(_01996_),
    .Y(_01997_),
    .A1(net174),
    .A2(_01994_));
 sg13g2_nor2_1 _10015_ (.A(_01983_),
    .B(_01997_),
    .Y(_01998_));
 sg13g2_nand2_1 _10016_ (.Y(_01999_),
    .A(_01983_),
    .B(_01997_));
 sg13g2_nor2b_2 _10017_ (.A(_01998_),
    .B_N(_01999_),
    .Y(_02000_));
 sg13g2_buf_2 fanout1166 (.A(net1167),
    .X(net1166));
 sg13g2_inv_1 _10019_ (.Y(_02002_),
    .A(net1497));
 sg13g2_nand3_1 _10020_ (.B(_01793_),
    .C(_01865_),
    .A(\id_stage_i.controller_i.instr_i_26_ ),
    .Y(_02003_));
 sg13g2_a221oi_1 _10021_ (.B2(_02003_),
    .C1(_01992_),
    .B1(_01863_),
    .A1(_02002_),
    .Y(_02004_),
    .A2(net1614));
 sg13g2_buf_2 fanout1165 (.A(net1168),
    .X(net1165));
 sg13g2_xor2_1 _10023_ (.B(net1278),
    .A(net87),
    .X(_02006_));
 sg13g2_buf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_nand2_1 _10025_ (.Y(_02008_),
    .A(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .B(net1558));
 sg13g2_nand2_1 _10026_ (.Y(_02009_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_27__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1972));
 sg13g2_o21ai_1 _10027_ (.B1(_02009_),
    .Y(_02010_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2_ ));
 sg13g2_nor3_1 _10028_ (.A(net1497),
    .B(net1709),
    .C(net402),
    .Y(_02011_));
 sg13g2_a221oi_1 _10029_ (.B2(net1896),
    .C1(_02011_),
    .B1(_02010_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_26__$_NOT__A_Y ),
    .Y(_02012_),
    .A2(net406));
 sg13g2_xnor2_1 _10030_ (.Y(_02013_),
    .A(_02008_),
    .B(_02012_));
 sg13g2_nand2_1 _10031_ (.Y(_02014_),
    .A(net357),
    .B(_02013_));
 sg13g2_o21ai_1 _10032_ (.B1(_02014_),
    .Y(_02015_),
    .A1(net352),
    .A2(_02006_));
 sg13g2_and2_1 _10033_ (.A(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .B(net1558),
    .X(_02016_));
 sg13g2_nor2_1 _10034_ (.A(net365),
    .B(_02012_),
    .Y(_02017_));
 sg13g2_nand2b_1 _10035_ (.Y(_02018_),
    .B(net1278),
    .A_N(_02017_));
 sg13g2_and3_1 _10036_ (.X(_02019_),
    .A(net351),
    .B(_02008_),
    .C(_02012_));
 sg13g2_a22oi_1 _10037_ (.Y(_02020_),
    .B1(_02019_),
    .B2(net1278),
    .A2(_02018_),
    .A1(_02016_));
 sg13g2_nand2_1 _10038_ (.Y(_02021_),
    .A(net367),
    .B(_02006_));
 sg13g2_nand3_1 _10039_ (.B(_02020_),
    .C(_02021_),
    .A(net189),
    .Y(_02022_));
 sg13g2_o21ai_1 _10040_ (.B1(_02022_),
    .Y(_02023_),
    .A1(net185),
    .A2(_02015_));
 sg13g2_buf_2 fanout1163 (.A(net1169),
    .X(net1163));
 sg13g2_nand2_2 _10042_ (.Y(_02025_),
    .A(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .B(net1558));
 sg13g2_nand2_1 _10043_ (.Y(_02026_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_24__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _10044_ (.B1(_02026_),
    .Y(_02027_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ),
    .A2(net2106));
 sg13g2_buf_2 fanout1162 (.A(net1163),
    .X(net1162));
 sg13g2_buf_2 fanout1161 (.A(\cs_registers_i/_0604_ ),
    .X(net1161));
 sg13g2_nor3_1 _10047_ (.A(net1494),
    .B(net1709),
    .C(net404),
    .Y(_02030_));
 sg13g2_a221oi_1 _10048_ (.B2(net1892),
    .C1(_02030_),
    .B1(_02027_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_23__$_NOT__A_Y ),
    .Y(_02031_),
    .A2(net409));
 sg13g2_nand2b_1 _10049_ (.Y(_02032_),
    .B(net351),
    .A_N(_02031_));
 sg13g2_and2_1 _10050_ (.A(net351),
    .B(_02031_),
    .X(_02033_));
 sg13g2_nand2_1 _10051_ (.Y(_02034_),
    .A(net1612),
    .B(net348));
 sg13g2_nor2_1 _10052_ (.A(_01858_),
    .B(_02034_),
    .Y(_02035_));
 sg13g2_nand2_1 _10053_ (.Y(_02036_),
    .A(net2008),
    .B(_02035_));
 sg13g2_inv_1 _10054_ (.Y(_02037_),
    .A(net1613));
 sg13g2_o21ai_1 _10055_ (.B1(_01773_),
    .Y(_02038_),
    .A1(net1494),
    .A2(_02037_));
 sg13g2_a21oi_1 _10056_ (.A1(_01963_),
    .A2(_02036_),
    .Y(_02039_),
    .B1(_02038_));
 sg13g2_a22oi_1 _10057_ (.Y(_02040_),
    .B1(_02033_),
    .B2(net1344),
    .A2(_02032_),
    .A1(net173));
 sg13g2_a21o_2 _10058_ (.A2(_02036_),
    .A1(_01963_),
    .B1(_02038_),
    .X(_02041_));
 sg13g2_and2_1 _10059_ (.A(net149),
    .B(net370),
    .X(_02042_));
 sg13g2_nand3_1 _10060_ (.B(_02041_),
    .C(_02042_),
    .A(net181),
    .Y(_02043_));
 sg13g2_o21ai_1 _10061_ (.B1(_02043_),
    .Y(_02044_),
    .A1(_02025_),
    .A2(_02040_));
 sg13g2_nor2_1 _10062_ (.A(net365),
    .B(net1344),
    .Y(_02045_));
 sg13g2_a21oi_1 _10063_ (.A1(net1344),
    .A2(_02042_),
    .Y(_02046_),
    .B1(_02045_));
 sg13g2_o21ai_1 _10064_ (.B1(_02032_),
    .Y(_02047_),
    .A1(net173),
    .A2(_02046_));
 sg13g2_nand3_1 _10065_ (.B(net172),
    .C(net1344),
    .A(net380),
    .Y(_02048_));
 sg13g2_nand3_1 _10066_ (.B(_02025_),
    .C(_02041_),
    .A(net188),
    .Y(_02049_));
 sg13g2_a21oi_1 _10067_ (.A1(_02048_),
    .A2(_02049_),
    .Y(_02050_),
    .B1(net149));
 sg13g2_a21oi_1 _10068_ (.A1(_02025_),
    .A2(_02047_),
    .Y(_02051_),
    .B1(_02050_));
 sg13g2_nand2b_2 _10069_ (.Y(_02052_),
    .B(_02051_),
    .A_N(_02044_));
 sg13g2_and2_1 _10070_ (.A(net125),
    .B(net364),
    .X(_02053_));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_and2_1 _10072_ (.A(net556),
    .B(net1558),
    .X(_02055_));
 sg13g2_nor2_2 _10073_ (.A(_02053_),
    .B(_02055_),
    .Y(_02056_));
 sg13g2_buf_1 fanout1159 (.A(\cs_registers_i/_0627_ ),
    .X(net1159));
 sg13g2_inv_4 _10075_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .Y(_02058_));
 sg13g2_nand2_1 _10076_ (.Y(_02059_),
    .A(\id_stage_i.controller_i.instr_i_24_ ),
    .B(_01961_));
 sg13g2_a221oi_1 _10077_ (.B2(_02059_),
    .C1(net1717),
    .B1(_01963_),
    .A1(_02058_),
    .Y(_02060_),
    .A2(net1614));
 sg13g2_nand2_2 _10078_ (.Y(_02061_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_25__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10079_ (.B1(_02061_),
    .Y(_02062_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ),
    .A2(net2106));
 sg13g2_nor3_1 _10080_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .B(net1709),
    .C(net402),
    .Y(_02063_));
 sg13g2_a221oi_1 _10081_ (.B2(net1892),
    .C1(_02063_),
    .B1(_02062_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_24__$_NOT__A_Y ),
    .Y(_02064_),
    .A2(net407));
 sg13g2_nor2_1 _10082_ (.A(net372),
    .B(_02064_),
    .Y(_02065_));
 sg13g2_a21oi_1 _10083_ (.A1(net110),
    .A2(_02060_),
    .Y(_02066_),
    .B1(_02065_));
 sg13g2_o21ai_1 _10084_ (.B1(_02066_),
    .Y(_02067_),
    .A1(net172),
    .A2(_02060_));
 sg13g2_xor2_1 _10085_ (.B(_02067_),
    .A(_02056_),
    .X(_02068_));
 sg13g2_inv_1 _10086_ (.Y(_02069_),
    .A(_02068_));
 sg13g2_and4_2 _10087_ (.A(_02000_),
    .B(_02023_),
    .C(_02052_),
    .D(_02069_),
    .X(_02070_));
 sg13g2_and2_1 _10088_ (.A(_01979_),
    .B(_02070_),
    .X(_02071_));
 sg13g2_inv_1 _10089_ (.Y(_02072_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ));
 sg13g2_a22oi_1 _10090_ (.Y(_02073_),
    .B1(net1881),
    .B2(_02072_),
    .A2(net1972),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_15__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_buf_2 fanout1158 (.A(\cs_registers_i/_0627_ ),
    .X(net1158));
 sg13g2_buf_1 fanout1157 (.A(\cs_registers_i/_0630_ ),
    .X(net1157));
 sg13g2_nor3_1 _10093_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .B(net1714),
    .C(net401),
    .Y(_02076_));
 sg13g2_a21oi_1 _10094_ (.A1(\ex_block_i.alu_i.imd_val_q_i_14__$_NOT__A_Y ),
    .A2(net401),
    .Y(_02077_),
    .B1(_02076_));
 sg13g2_o21ai_1 _10095_ (.B1(_02077_),
    .Y(_02078_),
    .A1(_01839_),
    .A2(_02073_));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(\cs_registers_i/_0630_ ));
 sg13g2_and2_1 _10097_ (.A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(net1559),
    .X(_02080_));
 sg13g2_or2_2 _10098_ (.X(_02081_),
    .B(net1613),
    .A(net1717));
 sg13g2_mux2_1 _10099_ (.A0(_01933_),
    .A1(_01859_),
    .S(_01791_),
    .X(_02082_));
 sg13g2_nor2_1 _10100_ (.A(_02081_),
    .B(_02082_),
    .Y(_02083_));
 sg13g2_nand4_1 _10101_ (.B(net1612),
    .C(_01933_),
    .A(net1999),
    .Y(_02084_),
    .D(_01882_));
 sg13g2_inv_1 _10102_ (.Y(_02085_),
    .A(_02084_));
 sg13g2_a221oi_1 _10103_ (.B2(net2093),
    .C1(_02085_),
    .B1(_02083_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .Y(_02086_),
    .A2(net330));
 sg13g2_buf_4 fanout1155 (.X(net1155),
    .A(\cs_registers_i/_0636_ ));
 sg13g2_nand2_1 _10105_ (.Y(_02088_),
    .A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(net1559));
 sg13g2_o21ai_1 _10106_ (.B1(_02088_),
    .Y(_02089_),
    .A1(_01224_),
    .A2(net353));
 sg13g2_and2_1 _10107_ (.A(net241),
    .B(_02089_),
    .X(_02090_));
 sg13g2_nand2_1 _10108_ (.Y(_02091_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_14__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1974));
 sg13g2_o21ai_1 _10109_ (.B1(_02091_),
    .Y(_02092_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ),
    .A2(net2109));
 sg13g2_buf_1 fanout1154 (.A(\cs_registers_i/_0645_ ),
    .X(net1154));
 sg13g2_nor3_1 _10111_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .B(net1714),
    .C(net404),
    .Y(_02094_));
 sg13g2_a221oi_1 _10112_ (.B2(net1895),
    .C1(_02094_),
    .B1(_02092_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_13__$_NOT__A_Y ),
    .Y(_02095_),
    .A2(net406));
 sg13g2_nor2_2 _10113_ (.A(net362),
    .B(_02095_),
    .Y(_02096_));
 sg13g2_inv_4 _10114_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .Y(_02097_));
 sg13g2_nor2_2 _10115_ (.A(net1612),
    .B(net387),
    .Y(_02098_));
 sg13g2_a22oi_1 _10116_ (.Y(_02099_),
    .B1(_02098_),
    .B2(net551),
    .A2(_01880_),
    .A1(net1999));
 sg13g2_or2_1 _10117_ (.X(_02100_),
    .B(_02099_),
    .A(net347));
 sg13g2_nand2_1 _10118_ (.Y(_02101_),
    .A(net1999),
    .B(_01858_));
 sg13g2_o21ai_1 _10119_ (.B1(_02101_),
    .Y(_02102_),
    .A1(_01361_),
    .A2(_01933_));
 sg13g2_a21oi_1 _10120_ (.A1(net1612),
    .A2(_02102_),
    .Y(_02103_),
    .B1(net1613));
 sg13g2_a221oi_1 _10121_ (.B2(_02103_),
    .C1(net1717),
    .B1(_02100_),
    .A1(_02097_),
    .Y(_02104_),
    .A2(net1613));
 sg13g2_nand2b_1 _10122_ (.Y(_02105_),
    .B(_02104_),
    .A_N(_02096_));
 sg13g2_a21oi_1 _10123_ (.A1(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .A2(net401),
    .Y(_02106_),
    .B1(_02078_));
 sg13g2_nor2_1 _10124_ (.A(net369),
    .B(_02106_),
    .Y(_02107_));
 sg13g2_a21oi_1 _10125_ (.A1(net1283),
    .A2(net379),
    .Y(_02108_),
    .B1(_02107_));
 sg13g2_nand2b_1 _10126_ (.Y(_02109_),
    .B(_02108_),
    .A_N(net241));
 sg13g2_nor4_2 _10127_ (.A(net350),
    .B(_01737_),
    .C(_01756_),
    .Y(_02110_),
    .D(_01762_));
 sg13g2_a21oi_1 _10128_ (.A1(_02105_),
    .A2(_02109_),
    .Y(_02111_),
    .B1(_02110_));
 sg13g2_nor2_1 _10129_ (.A(_01224_),
    .B(net241),
    .Y(_02112_));
 sg13g2_nand2_1 _10130_ (.Y(_02113_),
    .A(net241),
    .B(_02108_));
 sg13g2_o21ai_1 _10131_ (.B1(_02113_),
    .Y(_02114_),
    .A1(_02096_),
    .A2(_02104_));
 sg13g2_inv_1 _10132_ (.Y(_02115_),
    .A(\ex_block_i.alu_i.imd_val_q_i_45_ ));
 sg13g2_nor3_2 _10133_ (.A(_02115_),
    .B(net361),
    .C(net1675),
    .Y(_02116_));
 sg13g2_a21oi_2 _10134_ (.B1(_02116_),
    .Y(_02117_),
    .A2(net378),
    .A1(net1352));
 sg13g2_a21oi_1 _10135_ (.A1(net178),
    .A2(_02114_),
    .Y(_02118_),
    .B1(_02117_));
 sg13g2_a21oi_1 _10136_ (.A1(net110),
    .A2(_02112_),
    .Y(_02119_),
    .B1(_02118_));
 sg13g2_nor2_1 _10137_ (.A(_02111_),
    .B(_02119_),
    .Y(_02120_));
 sg13g2_a221oi_1 _10138_ (.B2(net186),
    .C1(_02120_),
    .B1(_02090_),
    .A1(_02078_),
    .Y(_02121_),
    .A2(_02080_));
 sg13g2_nor2_1 _10139_ (.A(net152),
    .B(net356),
    .Y(_02122_));
 sg13g2_inv_1 _10140_ (.Y(_02123_),
    .A(_02122_));
 sg13g2_nand2_1 _10141_ (.Y(_02124_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_11__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _10142_ (.B1(_02124_),
    .Y(_02125_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ),
    .A2(net2106));
 sg13g2_buf_1 fanout1153 (.A(net1154),
    .X(net1153));
 sg13g2_nor3_1 _10144_ (.A(net258),
    .B(net1710),
    .C(net404),
    .Y(_02127_));
 sg13g2_a221oi_1 _10145_ (.B2(net1892),
    .C1(_02127_),
    .B1(_02125_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_10__$_NOT__A_Y ),
    .Y(_02128_),
    .A2(net407));
 sg13g2_buf_2 fanout1152 (.A(net1154),
    .X(net1152));
 sg13g2_nand2_2 _10147_ (.Y(_02130_),
    .A(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .B(net399));
 sg13g2_and2_1 _10148_ (.A(net350),
    .B(_02130_),
    .X(_02131_));
 sg13g2_nand2_1 _10149_ (.Y(_02132_),
    .A(_02128_),
    .B(_02131_));
 sg13g2_a21oi_2 _10150_ (.B1(_02081_),
    .Y(_02133_),
    .A2(_01859_),
    .A1(_01857_));
 sg13g2_a22oi_1 _10151_ (.Y(_02134_),
    .B1(_02133_),
    .B2(net441),
    .A2(net331),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_10_ ));
 sg13g2_a21oi_1 _10152_ (.A1(_02123_),
    .A2(_02132_),
    .Y(_02135_),
    .B1(_02134_));
 sg13g2_nand2_1 _10153_ (.Y(_02136_),
    .A(_02134_),
    .B(_02122_));
 sg13g2_nand3_1 _10154_ (.B(_02132_),
    .C(_02136_),
    .A(net180),
    .Y(_02137_));
 sg13g2_o21ai_1 _10155_ (.B1(_02137_),
    .Y(_02138_),
    .A1(net175),
    .A2(_02135_));
 sg13g2_nand2_1 _10156_ (.Y(_02139_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_10__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _10157_ (.B1(_02139_),
    .Y(_02140_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ),
    .A2(net2106));
 sg13g2_buf_1 fanout1151 (.A(\cs_registers_i/_0645_ ),
    .X(net1151));
 sg13g2_nor3_1 _10159_ (.A(net1466),
    .B(net1710),
    .C(net400),
    .Y(_02142_));
 sg13g2_a221oi_1 _10160_ (.B2(net1892),
    .C1(_02142_),
    .B1(_02140_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_9__$_NOT__A_Y ),
    .Y(_02143_),
    .A2(net407));
 sg13g2_buf_2 fanout1150 (.A(\cs_registers_i/_0645_ ),
    .X(net1150));
 sg13g2_nand2b_2 _10162_ (.Y(_02145_),
    .B(net354),
    .A_N(_02143_));
 sg13g2_inv_1 _10163_ (.Y(_02146_),
    .A(_02145_));
 sg13g2_buf_2 fanout1149 (.A(\cs_registers_i/_0827_ ),
    .X(net1149));
 sg13g2_a22oi_1 _10165_ (.Y(_02148_),
    .B1(_02133_),
    .B2(\id_stage_i.controller_i.instr_i_29_ ),
    .A2(net330),
    .A1(net1466));
 sg13g2_buf_2 fanout1148 (.A(\cs_registers_i/_0827_ ),
    .X(net1148));
 sg13g2_and2_2 _10167_ (.A(net192),
    .B(net374),
    .X(_02150_));
 sg13g2_a22oi_1 _10168_ (.Y(_02151_),
    .B1(_02148_),
    .B2(_02150_),
    .A2(net1557),
    .A1(net2115));
 sg13g2_or2_1 _10169_ (.X(_02152_),
    .B(_02148_),
    .A(net354));
 sg13g2_a21oi_1 _10170_ (.A1(_02145_),
    .A2(_02152_),
    .Y(_02153_),
    .B1(net192));
 sg13g2_nor2_1 _10171_ (.A(net364),
    .B(_02143_),
    .Y(_02154_));
 sg13g2_nand2_1 _10172_ (.Y(_02155_),
    .A(net2115),
    .B(net1557));
 sg13g2_o21ai_1 _10173_ (.B1(_02155_),
    .Y(_02156_),
    .A1(_02153_),
    .A2(_02154_));
 sg13g2_o21ai_1 _10174_ (.B1(_02156_),
    .Y(_02157_),
    .A1(_02146_),
    .A2(_02151_));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(_03059_));
 sg13g2_a22oi_1 _10176_ (.Y(_02159_),
    .B1(_02133_),
    .B2(\id_stage_i.controller_i.instr_i_28_ ),
    .A2(net331),
    .A1(net1463));
 sg13g2_and3_1 _10177_ (.X(_02160_),
    .A(_01322_),
    .B(net369),
    .C(net1401));
 sg13g2_buf_2 fanout1146 (.A(_03059_),
    .X(net1146));
 sg13g2_buf_4 fanout1145 (.X(net1145),
    .A(_03059_));
 sg13g2_buf_1 fanout1144 (.A(_08312_),
    .X(net1144));
 sg13g2_a22oi_1 _10181_ (.Y(_02164_),
    .B1(_02133_),
    .B2(\id_stage_i.controller_i.instr_i_27_ ),
    .A2(net330),
    .A1(net282));
 sg13g2_buf_4 fanout1143 (.X(net1143),
    .A(net1144));
 sg13g2_nor2_1 _10183_ (.A(_01318_),
    .B(net1400),
    .Y(_02166_));
 sg13g2_nor2_1 _10184_ (.A(_01322_),
    .B(net1401),
    .Y(_02167_));
 sg13g2_nor3_1 _10185_ (.A(net355),
    .B(_02166_),
    .C(_02167_),
    .Y(_02168_));
 sg13g2_nand2_1 _10186_ (.Y(_02169_),
    .A(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .B(net1559));
 sg13g2_nand2_1 _10187_ (.Y(_02170_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_8__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10188_ (.B1(_02170_),
    .Y(_02171_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ),
    .A2(net2109));
 sg13g2_nor3_1 _10189_ (.A(net282),
    .B(net1712),
    .C(net403),
    .Y(_02172_));
 sg13g2_a221oi_1 _10190_ (.B2(net1894),
    .C1(_02172_),
    .B1(_02171_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_7__$_NOT__A_Y ),
    .Y(_02173_),
    .A2(net406));
 sg13g2_nor2_1 _10191_ (.A(_02169_),
    .B(_02173_),
    .Y(_02174_));
 sg13g2_inv_2 _10192_ (.Y(_02175_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_a22oi_1 _10193_ (.Y(_02176_),
    .B1(net1881),
    .B2(_02175_),
    .A2(net1972),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_9__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nand2b_1 _10194_ (.Y(_02177_),
    .B(net1893),
    .A_N(_02176_));
 sg13g2_nor3_1 _10195_ (.A(net1463),
    .B(net1711),
    .C(net400),
    .Y(_02178_));
 sg13g2_a21oi_2 _10196_ (.B1(_02178_),
    .Y(_02179_),
    .A2(net403),
    .A1(\ex_block_i.alu_i.imd_val_q_i_8__$_NOT__A_Y ));
 sg13g2_nand2_2 _10197_ (.Y(_02180_),
    .A(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .B(net399));
 sg13g2_nand3_1 _10198_ (.B(_02179_),
    .C(_02180_),
    .A(_02177_),
    .Y(_02181_));
 sg13g2_nand2_1 _10199_ (.Y(_02182_),
    .A(_02177_),
    .B(_02179_));
 sg13g2_nand2b_1 _10200_ (.Y(_02183_),
    .B(_02182_),
    .A_N(_02180_));
 sg13g2_nand2_1 _10201_ (.Y(_02184_),
    .A(net356),
    .B(_02183_));
 sg13g2_a21oi_1 _10202_ (.A1(_02174_),
    .A2(_02181_),
    .Y(_02185_),
    .B1(_02184_));
 sg13g2_nor3_2 _10203_ (.A(_02160_),
    .B(_02168_),
    .C(_02185_),
    .Y(_02186_));
 sg13g2_nand2_1 _10204_ (.Y(_02187_),
    .A(_02157_),
    .B(_02186_));
 sg13g2_a21oi_2 _10205_ (.B1(_02150_),
    .Y(_02188_),
    .A2(net1557),
    .A1(net2115));
 sg13g2_inv_1 _10206_ (.Y(_02189_),
    .A(_02188_));
 sg13g2_inv_2 _10207_ (.Y(_02190_),
    .A(net258));
 sg13g2_nand2_2 _10208_ (.Y(_02191_),
    .A(_01773_),
    .B(net1613));
 sg13g2_nand2_1 _10209_ (.Y(_02192_),
    .A(net441),
    .B(_02133_));
 sg13g2_o21ai_1 _10210_ (.B1(_02192_),
    .Y(_02193_),
    .A1(_02190_),
    .A2(_02191_));
 sg13g2_inv_2 _10211_ (.Y(_02194_),
    .A(_02148_));
 sg13g2_a22oi_1 _10212_ (.Y(_02195_),
    .B1(_02194_),
    .B2(net193),
    .A2(_02193_),
    .A1(net152));
 sg13g2_inv_1 _10213_ (.Y(_02196_),
    .A(_02195_));
 sg13g2_nor3_1 _10214_ (.A(net372),
    .B(_02128_),
    .C(_02130_),
    .Y(_02197_));
 sg13g2_a221oi_1 _10215_ (.B2(net370),
    .C1(_02197_),
    .B1(_02196_),
    .A1(_02146_),
    .Y(_02198_),
    .A2(_02189_));
 sg13g2_nand2_1 _10216_ (.Y(_02199_),
    .A(_02187_),
    .B(_02198_));
 sg13g2_nand2_1 _10217_ (.Y(_02200_),
    .A(_02145_),
    .B(_02194_));
 sg13g2_nor2_1 _10218_ (.A(net362),
    .B(_02180_),
    .Y(_02201_));
 sg13g2_a21o_1 _10219_ (.A2(net378),
    .A1(net1279),
    .B1(_02201_),
    .X(_02202_));
 sg13g2_a22oi_1 _10220_ (.Y(_02203_),
    .B1(_02202_),
    .B2(net1401),
    .A2(_02201_),
    .A1(_02182_));
 sg13g2_inv_4 _10221_ (.A(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .Y(_02204_));
 sg13g2_nor3_2 _10222_ (.A(_02204_),
    .B(net363),
    .C(net1674),
    .Y(_02205_));
 sg13g2_nand2b_1 _10223_ (.Y(_02206_),
    .B(_02173_),
    .A_N(net1400));
 sg13g2_nor2_1 _10224_ (.A(_01318_),
    .B(net356),
    .Y(_02207_));
 sg13g2_a22oi_1 _10225_ (.Y(_02208_),
    .B1(_02207_),
    .B2(net1400),
    .A2(_02206_),
    .A1(_02205_));
 sg13g2_nor2_1 _10226_ (.A(net369),
    .B(_02181_),
    .Y(_02209_));
 sg13g2_a21oi_1 _10227_ (.A1(_01322_),
    .A2(net380),
    .Y(_02210_),
    .B1(_02209_));
 sg13g2_nor2_1 _10228_ (.A(net1401),
    .B(_02210_),
    .Y(_02211_));
 sg13g2_a21oi_2 _10229_ (.B1(_02211_),
    .Y(_02212_),
    .A2(_02208_),
    .A1(_02203_));
 sg13g2_o21ai_1 _10230_ (.B1(_02212_),
    .Y(_02213_),
    .A1(_02189_),
    .A2(_02200_));
 sg13g2_a21oi_1 _10231_ (.A1(_02193_),
    .A2(_02128_),
    .Y(_02214_),
    .B1(_02130_));
 sg13g2_and3_1 _10232_ (.X(_02215_),
    .A(net152),
    .B(net372),
    .C(_02134_));
 sg13g2_a221oi_1 _10233_ (.B2(net350),
    .C1(_02215_),
    .B1(_02214_),
    .A1(_02189_),
    .Y(_02216_),
    .A2(_02200_));
 sg13g2_nand2_1 _10234_ (.Y(_02217_),
    .A(_02213_),
    .B(_02216_));
 sg13g2_mux2_1 _10235_ (.A0(_02199_),
    .A1(_02217_),
    .S(net184),
    .X(_02218_));
 sg13g2_a21oi_1 _10236_ (.A1(_02205_),
    .A2(_02173_),
    .Y(_02219_),
    .B1(_02207_));
 sg13g2_nand2_2 _10237_ (.Y(_02220_),
    .A(net148),
    .B(net364));
 sg13g2_nand2_2 _10238_ (.Y(_02221_),
    .A(net1400),
    .B(_02220_));
 sg13g2_o21ai_1 _10239_ (.B1(_02221_),
    .Y(_02222_),
    .A1(net364),
    .A2(_02173_));
 sg13g2_nand2_1 _10240_ (.Y(_02223_),
    .A(_02169_),
    .B(_02222_));
 sg13g2_o21ai_1 _10241_ (.B1(_02223_),
    .Y(_02224_),
    .A1(net1400),
    .A2(_02219_));
 sg13g2_o21ai_1 _10242_ (.B1(_02134_),
    .Y(_02225_),
    .A1(_02122_),
    .A2(_02131_));
 sg13g2_inv_1 _10243_ (.Y(_02226_),
    .A(_02128_));
 sg13g2_nand3_1 _10244_ (.B(net399),
    .C(_02128_),
    .A(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .Y(_02227_));
 sg13g2_nand2_1 _10245_ (.Y(_02228_),
    .A(net152),
    .B(net372));
 sg13g2_o21ai_1 _10246_ (.B1(_02228_),
    .Y(_02229_),
    .A1(net364),
    .A2(_02227_));
 sg13g2_a22oi_1 _10247_ (.Y(_02230_),
    .B1(_02229_),
    .B2(_02193_),
    .A2(_02131_),
    .A1(_02226_));
 sg13g2_nand2_1 _10248_ (.Y(_02231_),
    .A(_02225_),
    .B(_02230_));
 sg13g2_inv_1 _10249_ (.Y(_02232_),
    .A(_02203_));
 sg13g2_xor2_1 _10250_ (.B(_02200_),
    .A(_02188_),
    .X(_02233_));
 sg13g2_nor3_1 _10251_ (.A(_02211_),
    .B(_02232_),
    .C(_02233_),
    .Y(_02234_));
 sg13g2_nand3_1 _10252_ (.B(_02231_),
    .C(_02234_),
    .A(_02224_),
    .Y(_02235_));
 sg13g2_xnor2_1 _10253_ (.Y(_02236_),
    .A(_01318_),
    .B(net1400));
 sg13g2_nor2_1 _10254_ (.A(_02204_),
    .B(net1674),
    .Y(_02237_));
 sg13g2_xnor2_1 _10255_ (.Y(_02238_),
    .A(_02173_),
    .B(_02237_));
 sg13g2_nor2_1 _10256_ (.A(net370),
    .B(_02238_),
    .Y(_02239_));
 sg13g2_a21oi_2 _10257_ (.B1(_02239_),
    .Y(_02240_),
    .A2(_02236_),
    .A1(net365));
 sg13g2_nand2_1 _10258_ (.Y(_02241_),
    .A(net2115),
    .B(net398));
 sg13g2_xnor2_1 _10259_ (.Y(_02242_),
    .A(_02145_),
    .B(_02241_));
 sg13g2_xor2_1 _10260_ (.B(_02130_),
    .A(_02128_),
    .X(_02243_));
 sg13g2_nand4_1 _10261_ (.B(_02181_),
    .C(_02183_),
    .A(net359),
    .Y(_02244_),
    .D(_02243_));
 sg13g2_xnor2_1 _10262_ (.Y(_02245_),
    .A(net1279),
    .B(net1401));
 sg13g2_xnor2_1 _10263_ (.Y(_02246_),
    .A(net151),
    .B(_02134_));
 sg13g2_nand2_1 _10264_ (.Y(_02247_),
    .A(_02145_),
    .B(_02148_));
 sg13g2_xor2_1 _10265_ (.B(_02247_),
    .A(net192),
    .X(_02248_));
 sg13g2_nand4_1 _10266_ (.B(_02245_),
    .C(_02246_),
    .A(net380),
    .Y(_02249_),
    .D(_02248_));
 sg13g2_o21ai_1 _10267_ (.B1(_02249_),
    .Y(_02250_),
    .A1(_02242_),
    .A2(_02244_));
 sg13g2_nand3_1 _10268_ (.B(_02240_),
    .C(_02250_),
    .A(net179),
    .Y(_02251_));
 sg13g2_o21ai_1 _10269_ (.B1(_02251_),
    .Y(_02252_),
    .A1(net173),
    .A2(_02235_));
 sg13g2_nand2_1 _10270_ (.Y(_02253_),
    .A(_01773_),
    .B(_01880_));
 sg13g2_nor2b_1 _10271_ (.A(_01804_),
    .B_N(net347),
    .Y(_02254_));
 sg13g2_nor3_1 _10272_ (.A(_02253_),
    .B(_01805_),
    .C(_02254_),
    .Y(_02255_));
 sg13g2_a22oi_1 _10273_ (.Y(_02256_),
    .B1(_02255_),
    .B2(net553),
    .A2(_01805_),
    .A1(\id_stage_i.controller_i.instr_i_24_ ));
 sg13g2_buf_4 fanout1142 (.X(net1142),
    .A(net1144));
 sg13g2_nor2_1 _10275_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ),
    .B(_02191_),
    .Y(_02258_));
 sg13g2_a21oi_2 _10276_ (.B1(_02258_),
    .Y(_02259_),
    .A2(_02256_),
    .A1(_02191_));
 sg13g2_nand3_1 _10277_ (.B(net171),
    .C(net1399),
    .A(net378),
    .Y(_02260_));
 sg13g2_a21o_2 _10278_ (.A2(_02256_),
    .A1(_02191_),
    .B1(_02258_),
    .X(_02261_));
 sg13g2_nand2_1 _10279_ (.Y(_02262_),
    .A(net187),
    .B(_02261_));
 sg13g2_inv_1 _10280_ (.Y(_02263_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_a22oi_1 _10281_ (.Y(_02264_),
    .B1(net1881),
    .B2(_02263_),
    .A2(net1972),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_5__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nand2b_1 _10282_ (.Y(_02265_),
    .B(net1896),
    .A_N(_02264_));
 sg13g2_or2_1 _10283_ (.X(_02266_),
    .B(\ex_block_i.alu_i.imd_val_q_i_4__$_NOT__A_Y ),
    .A(\ex_block_i.alu_i.imd_val_q_i_36_ ));
 sg13g2_o21ai_1 _10284_ (.B1(net1674),
    .Y(_02267_),
    .A1(net1507),
    .A2(net1711));
 sg13g2_o21ai_1 _10285_ (.B1(_02267_),
    .Y(_02268_),
    .A1(net1674),
    .A2(_02266_));
 sg13g2_a21o_1 _10286_ (.A2(_02268_),
    .A1(_02265_),
    .B1(net381),
    .X(_02269_));
 sg13g2_nand2_2 _10287_ (.Y(_02270_),
    .A(net1406),
    .B(net363));
 sg13g2_and2_1 _10288_ (.A(_02269_),
    .B(_02270_),
    .X(_02271_));
 sg13g2_nand3_1 _10289_ (.B(_02262_),
    .C(_02271_),
    .A(_02260_),
    .Y(_02272_));
 sg13g2_nand2_1 _10290_ (.Y(_02273_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_4__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1974));
 sg13g2_o21ai_1 _10291_ (.B1(_02273_),
    .Y(_02274_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .A2(net2109));
 sg13g2_buf_2 fanout1141 (.A(net1144),
    .X(net1141));
 sg13g2_nor3_1 _10293_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_3_ ),
    .B(net1714),
    .C(net400),
    .Y(_02276_));
 sg13g2_a221oi_1 _10294_ (.B2(net1895),
    .C1(_02276_),
    .B1(_02274_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_3__$_NOT__A_Y ),
    .Y(_02277_),
    .A2(net405));
 sg13g2_nand2b_2 _10295_ (.Y(_02278_),
    .B(net349),
    .A_N(_02277_));
 sg13g2_nand2_1 _10296_ (.Y(_02279_),
    .A(net178),
    .B(_02278_));
 sg13g2_inv_1 _10297_ (.Y(_02280_),
    .A(\ex_block_i.alu_i.imd_val_q_i_35_ ));
 sg13g2_nor2_1 _10298_ (.A(_02280_),
    .B(net1674),
    .Y(_02281_));
 sg13g2_mux2_2 _10299_ (.A0(net1408),
    .A1(_02281_),
    .S(net349),
    .X(_02282_));
 sg13g2_inv_4 _10300_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_3_ ),
    .Y(_02283_));
 sg13g2_inv_1 _10301_ (.Y(_02284_),
    .A(\id_stage_i.controller_i.instr_i_10_ ));
 sg13g2_or4_1 _10302_ (.A(_02284_),
    .B(_02253_),
    .C(_01805_),
    .D(_02254_),
    .X(_02285_));
 sg13g2_a21oi_1 _10303_ (.A1(net2008),
    .A2(_01805_),
    .Y(_02286_),
    .B1(net332));
 sg13g2_a22oi_1 _10304_ (.Y(_02287_),
    .B1(_02285_),
    .B2(_02286_),
    .A2(net329),
    .A1(_02283_));
 sg13g2_nand2_2 _10305_ (.Y(_02288_),
    .A(_02278_),
    .B(_02287_));
 sg13g2_nand3_1 _10306_ (.B(_02282_),
    .C(_02288_),
    .A(_02279_),
    .Y(_02289_));
 sg13g2_inv_2 _10307_ (.Y(_02290_),
    .A(_02282_));
 sg13g2_nand2_1 _10308_ (.Y(_02291_),
    .A(net361),
    .B(_02287_));
 sg13g2_nor2_1 _10309_ (.A(_02290_),
    .B(_02291_),
    .Y(_02292_));
 sg13g2_inv_1 _10310_ (.Y(_02293_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_a22oi_1 _10311_ (.Y(_02294_),
    .B1(net1881),
    .B2(_02293_),
    .A2(net1974),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1144));
 sg13g2_buf_2 fanout1139 (.A(_08460_),
    .X(net1139));
 sg13g2_buf_1 fanout1138 (.A(_08460_),
    .X(net1138));
 sg13g2_nor3_1 _10315_ (.A(net1503),
    .B(net1712),
    .C(net400),
    .Y(_02298_));
 sg13g2_a21oi_1 _10316_ (.A1(\ex_block_i.alu_i.imd_val_q_i_1__$_NOT__A_Y ),
    .A2(net400),
    .Y(_02299_),
    .B1(_02298_));
 sg13g2_o21ai_1 _10317_ (.B1(_02299_),
    .Y(_02300_),
    .A1(_01839_),
    .A2(_02294_));
 sg13g2_nand2_1 _10318_ (.Y(_02301_),
    .A(\ex_block_i.alu_i.imd_val_q_i_33_ ),
    .B(net398));
 sg13g2_buf_2 fanout1137 (.A(_08460_),
    .X(net1137));
 sg13g2_o21ai_1 _10320_ (.B1(net1674),
    .Y(_02303_),
    .A1(net280),
    .A2(net1712));
 sg13g2_inv_1 _10321_ (.Y(_02304_),
    .A(\ex_block_i.alu_i.imd_val_q_i_32_ ));
 sg13g2_nand3b_1 _10322_ (.B(_02304_),
    .C(net399),
    .Y(_02305_),
    .A_N(\ex_block_i.alu_i.imd_val_q_i_0__$_NOT__A_Y ));
 sg13g2_inv_1 _10323_ (.Y(_02306_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ));
 sg13g2_a22oi_1 _10324_ (.Y(_02307_),
    .B1(_01906_),
    .B2(_02306_),
    .A2(net1974),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_1__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nor2_1 _10325_ (.A(_01839_),
    .B(_02307_),
    .Y(_02308_));
 sg13g2_a21oi_2 _10326_ (.B1(_02308_),
    .Y(_02309_),
    .A2(_02305_),
    .A1(_02303_));
 sg13g2_nand2_1 _10327_ (.Y(_02310_),
    .A(_02301_),
    .B(_02309_));
 sg13g2_nor2_1 _10328_ (.A(_02301_),
    .B(_02309_),
    .Y(_02311_));
 sg13g2_a21oi_1 _10329_ (.A1(_02300_),
    .A2(_02310_),
    .Y(_02312_),
    .B1(_02311_));
 sg13g2_nand2_1 _10330_ (.Y(_02313_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_3__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1974));
 sg13g2_o21ai_1 _10331_ (.B1(_02313_),
    .Y(_02314_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ),
    .A2(net2108));
 sg13g2_buf_2 fanout1136 (.A(net1138),
    .X(net1136));
 sg13g2_nor3_1 _10333_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ),
    .B(net1713),
    .C(net400),
    .Y(_02316_));
 sg13g2_a221oi_1 _10334_ (.B2(net1894),
    .C1(_02316_),
    .B1(_02314_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_2__$_NOT__A_Y ),
    .Y(_02317_),
    .A2(net405));
 sg13g2_nor2_1 _10335_ (.A(net363),
    .B(_02317_),
    .Y(_02318_));
 sg13g2_nand2b_1 _10336_ (.Y(_02319_),
    .B(_02318_),
    .A_N(_02312_));
 sg13g2_inv_4 _10337_ (.A(net1504),
    .Y(_02320_));
 sg13g2_nor2_1 _10338_ (.A(net348),
    .B(_01804_),
    .Y(_02321_));
 sg13g2_nor3_1 _10339_ (.A(net1717),
    .B(_01803_),
    .C(_02034_),
    .Y(_02322_));
 sg13g2_o21ai_1 _10340_ (.B1(net1992),
    .Y(_02323_),
    .A1(_02321_),
    .A2(_02322_));
 sg13g2_inv_1 _10341_ (.Y(_02324_),
    .A(\id_stage_i.imm_b_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_inv_1 _10342_ (.Y(_02325_),
    .A(net347));
 sg13g2_o21ai_1 _10343_ (.B1(_01804_),
    .Y(_02326_),
    .A1(_02324_),
    .A2(_02325_));
 sg13g2_a221oi_1 _10344_ (.B2(_02253_),
    .C1(net332),
    .B1(_02326_),
    .A1(\id_stage_i.controller_i.instr_i_22_ ),
    .Y(_02327_),
    .A2(_01805_));
 sg13g2_a22oi_1 _10345_ (.Y(_02328_),
    .B1(_02323_),
    .B2(_02327_),
    .A2(net330),
    .A1(_02320_));
 sg13g2_buf_2 fanout1135 (.A(_08475_),
    .X(net1135));
 sg13g2_nand2_1 _10347_ (.Y(_02330_),
    .A(net369),
    .B(net1398));
 sg13g2_inv_8 _10348_ (.Y(_02331_),
    .A(net1411));
 sg13g2_nand2_1 _10349_ (.Y(_02332_),
    .A(net1503),
    .B(net1614));
 sg13g2_inv_1 _10350_ (.Y(_02333_),
    .A(\id_stage_i.controller_i.instr_i_8_ ));
 sg13g2_buf_2 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_nand2_1 _10352_ (.Y(_02335_),
    .A(net440),
    .B(_01858_));
 sg13g2_mux2_1 _10353_ (.A0(_02333_),
    .A1(_02335_),
    .S(_01791_),
    .X(_02336_));
 sg13g2_nor3_1 _10354_ (.A(_02325_),
    .B(_02081_),
    .C(_02336_),
    .Y(_02337_));
 sg13g2_and3_1 _10355_ (.X(_02338_),
    .A(net448),
    .B(_02325_),
    .C(_02037_));
 sg13g2_o21ai_1 _10356_ (.B1(_01858_),
    .Y(_02339_),
    .A1(_02337_),
    .A2(_02338_));
 sg13g2_a21o_2 _10357_ (.A2(_02339_),
    .A1(_02332_),
    .B1(net1717),
    .X(_02340_));
 sg13g2_nand3b_1 _10358_ (.B(_02321_),
    .C(_01882_),
    .Y(_02341_),
    .A_N(_02336_));
 sg13g2_nand3_1 _10359_ (.B(_02340_),
    .C(_02341_),
    .A(_02331_),
    .Y(_02342_));
 sg13g2_mux2_1 _10360_ (.A0(net513),
    .A1(net1994),
    .S(net348),
    .X(_02343_));
 sg13g2_nor2_1 _10361_ (.A(net387),
    .B(_01883_),
    .Y(_02344_));
 sg13g2_a22oi_1 _10362_ (.Y(_02345_),
    .B1(_02343_),
    .B2(_02344_),
    .A2(net329),
    .A1(net280));
 sg13g2_nor2b_2 _10363_ (.A(net1457),
    .B_N(net197),
    .Y(_02346_));
 sg13g2_a21oi_2 _10364_ (.B1(_02331_),
    .Y(_02347_),
    .A2(_02341_),
    .A1(_02340_));
 sg13g2_a21oi_2 _10365_ (.B1(_02347_),
    .Y(_02348_),
    .A2(_02346_),
    .A1(_02342_));
 sg13g2_and2_1 _10366_ (.A(_02278_),
    .B(_02291_),
    .X(_02349_));
 sg13g2_and2_1 _10367_ (.A(_02290_),
    .B(_02349_),
    .X(_02350_));
 sg13g2_a221oi_1 _10368_ (.B2(net370),
    .C1(_02350_),
    .B1(_02348_),
    .A1(_02319_),
    .Y(_02351_),
    .A2(_02330_));
 sg13g2_o21ai_1 _10369_ (.B1(net178),
    .Y(_02352_),
    .A1(_02292_),
    .A2(_02351_));
 sg13g2_nand2_1 _10370_ (.Y(_02353_),
    .A(_02289_),
    .B(_02352_));
 sg13g2_nand2_1 _10371_ (.Y(_02354_),
    .A(_02272_),
    .B(_02353_));
 sg13g2_nand2_1 _10372_ (.Y(_02355_),
    .A(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .B(net1559));
 sg13g2_nor3_1 _10373_ (.A(net1507),
    .B(net1711),
    .C(net401),
    .Y(_02356_));
 sg13g2_a21oi_1 _10374_ (.A1(\ex_block_i.alu_i.imd_val_q_i_4__$_NOT__A_Y ),
    .A2(net401),
    .Y(_02357_),
    .B1(_02356_));
 sg13g2_a21oi_2 _10375_ (.B1(net363),
    .Y(_02358_),
    .A2(_02357_),
    .A1(_02265_));
 sg13g2_nor2_1 _10376_ (.A(_02261_),
    .B(_02358_),
    .Y(_02359_));
 sg13g2_or2_1 _10377_ (.X(_02360_),
    .B(_02359_),
    .A(_02355_));
 sg13g2_xnor2_1 _10378_ (.Y(_02361_),
    .A(net188),
    .B(net1399));
 sg13g2_inv_1 _10379_ (.Y(_02362_),
    .A(_02358_));
 sg13g2_a22oi_1 _10380_ (.Y(_02363_),
    .B1(_02361_),
    .B2(_02362_),
    .A2(_02360_),
    .A1(_02270_));
 sg13g2_a22oi_1 _10381_ (.Y(_02364_),
    .B1(net1559),
    .B2(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .A2(net380),
    .A1(net1349));
 sg13g2_buf_2 fanout1133 (.A(_08565_),
    .X(net1133));
 sg13g2_buf_2 fanout1132 (.A(\cs_registers_i/_0545_ ),
    .X(net1132));
 sg13g2_a22oi_1 _10384_ (.Y(_02367_),
    .B1(_02133_),
    .B2(net2006),
    .A2(net330),
    .A1(net1511));
 sg13g2_nand2_2 _10385_ (.Y(_02368_),
    .A(net187),
    .B(_02367_));
 sg13g2_nand2_1 _10386_ (.Y(_02369_),
    .A(\ex_block_i.alu_i.imd_val_q_i_37_ ),
    .B(net398));
 sg13g2_nand2_1 _10387_ (.Y(_02370_),
    .A(net1404),
    .B(net374));
 sg13g2_o21ai_1 _10388_ (.B1(_02370_),
    .Y(_02371_),
    .A1(net363),
    .A2(_02369_));
 sg13g2_nand2b_1 _10389_ (.Y(_02372_),
    .B(_02371_),
    .A_N(_02368_));
 sg13g2_nand2_1 _10390_ (.Y(_02373_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_6__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1972));
 sg13g2_o21ai_1 _10391_ (.B1(_02373_),
    .Y(_02374_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ),
    .A2(net2107));
 sg13g2_nor3_1 _10392_ (.A(net1511),
    .B(net1709),
    .C(net400),
    .Y(_02375_));
 sg13g2_a221oi_1 _10393_ (.B2(net1893),
    .C1(_02375_),
    .B1(_02374_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_5__$_NOT__A_Y ),
    .Y(_02376_),
    .A2(net405));
 sg13g2_nor3_1 _10394_ (.A(net362),
    .B(_02376_),
    .C(_02369_),
    .Y(_02377_));
 sg13g2_nor3_1 _10395_ (.A(net183),
    .B(_02370_),
    .C(_02367_),
    .Y(_02378_));
 sg13g2_nor2_1 _10396_ (.A(_02377_),
    .B(_02378_),
    .Y(_02379_));
 sg13g2_and2_1 _10397_ (.A(_02372_),
    .B(_02379_),
    .X(_02380_));
 sg13g2_nand2_1 _10398_ (.Y(_02381_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_7__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1972));
 sg13g2_o21ai_1 _10399_ (.B1(_02381_),
    .Y(_02382_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ),
    .A2(net2107));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(\cs_registers_i/_0545_ ));
 sg13g2_nor3_1 _10401_ (.A(net1513),
    .B(net1711),
    .C(net401),
    .Y(_02384_));
 sg13g2_a221oi_1 _10402_ (.B2(net1896),
    .C1(_02384_),
    .B1(_02382_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_6__$_NOT__A_Y ),
    .Y(_02385_),
    .A2(net407));
 sg13g2_nor2_2 _10403_ (.A(net368),
    .B(_02385_),
    .Y(_02386_));
 sg13g2_a22oi_1 _10404_ (.Y(_02387_),
    .B1(_02133_),
    .B2(\id_stage_i.controller_i.instr_i_26_ ),
    .A2(net330),
    .A1(net1513));
 sg13g2_inv_1 _10405_ (.Y(_02388_),
    .A(_02387_));
 sg13g2_nor2_1 _10406_ (.A(net171),
    .B(_02388_),
    .Y(_02389_));
 sg13g2_nor3_1 _10407_ (.A(net350),
    .B(net187),
    .C(_02387_),
    .Y(_02390_));
 sg13g2_or3_2 _10408_ (.A(_02386_),
    .B(_02389_),
    .C(_02390_),
    .X(_02391_));
 sg13g2_inv_1 _10409_ (.Y(_02392_),
    .A(_02391_));
 sg13g2_a21oi_1 _10410_ (.A1(_02364_),
    .A2(_02380_),
    .Y(_02393_),
    .B1(_02392_));
 sg13g2_nor2_1 _10411_ (.A(_02364_),
    .B(_02380_),
    .Y(_02394_));
 sg13g2_o21ai_1 _10412_ (.B1(_02310_),
    .Y(_02395_),
    .A1(_02300_),
    .A2(_02311_));
 sg13g2_nand3_1 _10413_ (.B(_02317_),
    .C(_02395_),
    .A(net356),
    .Y(_02396_));
 sg13g2_o21ai_1 _10414_ (.B1(_02396_),
    .Y(_02397_),
    .A1(net349),
    .A2(net1398));
 sg13g2_o21ai_1 _10415_ (.B1(_02397_),
    .Y(_02398_),
    .A1(net355),
    .A2(_02348_));
 sg13g2_nand2_2 _10416_ (.Y(_02399_),
    .A(\ex_block_i.alu_i.imd_val_q_i_34_ ),
    .B(net399));
 sg13g2_nand2_1 _10417_ (.Y(_02400_),
    .A(net1409),
    .B(net362));
 sg13g2_o21ai_1 _10418_ (.B1(_02400_),
    .Y(_02401_),
    .A1(net373),
    .A2(_02399_));
 sg13g2_and2_1 _10419_ (.A(net171),
    .B(_02401_),
    .X(_02402_));
 sg13g2_nor2_1 _10420_ (.A(net361),
    .B(_02301_),
    .Y(_02403_));
 sg13g2_a21oi_2 _10421_ (.B1(_02403_),
    .Y(_02404_),
    .A2(net378),
    .A1(net1411));
 sg13g2_a22oi_1 _10422_ (.Y(_02405_),
    .B1(_02340_),
    .B2(_02341_),
    .A2(_02300_),
    .A1(net349));
 sg13g2_nand2b_1 _10423_ (.Y(_02406_),
    .B(net362),
    .A_N(net197));
 sg13g2_nand2_1 _10424_ (.Y(_02407_),
    .A(net356),
    .B(_02309_));
 sg13g2_a21oi_2 _10425_ (.B1(net1457),
    .Y(_02408_),
    .A2(_02407_),
    .A1(_02406_));
 sg13g2_a21o_1 _10426_ (.A2(_02405_),
    .A1(_02404_),
    .B1(_02408_),
    .X(_02409_));
 sg13g2_or2_1 _10427_ (.X(_02410_),
    .B(_02405_),
    .A(_02404_));
 sg13g2_inv_1 _10428_ (.Y(_02411_),
    .A(_02399_));
 sg13g2_inv_4 _10429_ (.A(_02328_),
    .Y(_02412_));
 sg13g2_a22oi_1 _10430_ (.Y(_02413_),
    .B1(_02401_),
    .B2(_02412_),
    .A2(_02411_),
    .A1(_02318_));
 sg13g2_nand3_1 _10431_ (.B(_02410_),
    .C(_02413_),
    .A(_02409_),
    .Y(_02414_));
 sg13g2_nand3_1 _10432_ (.B(_02317_),
    .C(_02399_),
    .A(net359),
    .Y(_02415_));
 sg13g2_o21ai_1 _10433_ (.B1(_02415_),
    .Y(_02416_),
    .A1(net1409),
    .A2(net354));
 sg13g2_nand2_1 _10434_ (.Y(_02417_),
    .A(net1398),
    .B(_02416_));
 sg13g2_and2_1 _10435_ (.A(net183),
    .B(_02417_),
    .X(_02418_));
 sg13g2_a22oi_1 _10436_ (.Y(_02419_),
    .B1(_02414_),
    .B2(_02418_),
    .A2(_02402_),
    .A1(_02398_));
 sg13g2_nand2_1 _10437_ (.Y(_02420_),
    .A(net178),
    .B(_02350_));
 sg13g2_nor2_1 _10438_ (.A(_02282_),
    .B(_02288_),
    .Y(_02421_));
 sg13g2_nand2_1 _10439_ (.Y(_02422_),
    .A(net187),
    .B(_02421_));
 sg13g2_nand3_1 _10440_ (.B(_02420_),
    .C(_02422_),
    .A(_02272_),
    .Y(_02423_));
 sg13g2_nor2_2 _10441_ (.A(_02419_),
    .B(_02423_),
    .Y(_02424_));
 sg13g2_nor4_2 _10442_ (.A(_02363_),
    .B(_02393_),
    .C(_02394_),
    .Y(_02425_),
    .D(_02424_));
 sg13g2_nand2_1 _10443_ (.Y(_02426_),
    .A(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .B(net1559));
 sg13g2_nand3_1 _10444_ (.B(net1349),
    .C(net373),
    .A(net1404),
    .Y(_02427_));
 sg13g2_and2_1 _10445_ (.A(_02376_),
    .B(_02369_),
    .X(_02428_));
 sg13g2_and2_1 _10446_ (.A(net354),
    .B(_02428_),
    .X(_02429_));
 sg13g2_a21oi_1 _10447_ (.A1(_02426_),
    .A2(_02427_),
    .Y(_02430_),
    .B1(_02429_));
 sg13g2_nor4_1 _10448_ (.A(net110),
    .B(_02387_),
    .C(_02386_),
    .D(_02430_),
    .Y(_02431_));
 sg13g2_nor4_1 _10449_ (.A(net183),
    .B(_02388_),
    .C(_02386_),
    .D(_02430_),
    .Y(_02432_));
 sg13g2_or2_1 _10450_ (.X(_02433_),
    .B(_02432_),
    .A(_02431_));
 sg13g2_nand2_1 _10451_ (.Y(_02434_),
    .A(net356),
    .B(_02428_));
 sg13g2_inv_2 _10452_ (.Y(_02435_),
    .A(_02367_));
 sg13g2_nand3_1 _10453_ (.B(_02434_),
    .C(_02435_),
    .A(net178),
    .Y(_02436_));
 sg13g2_a22oi_1 _10454_ (.Y(_02437_),
    .B1(_02368_),
    .B2(_02436_),
    .A2(_02433_),
    .A1(_02364_));
 sg13g2_nand3_1 _10455_ (.B(_01310_),
    .C(net372),
    .A(_01309_),
    .Y(_02438_));
 sg13g2_inv_1 _10456_ (.Y(_02439_),
    .A(net1349));
 sg13g2_o21ai_1 _10457_ (.B1(_02426_),
    .Y(_02440_),
    .A1(_02439_),
    .A2(net355));
 sg13g2_a21oi_1 _10458_ (.A1(_02434_),
    .A2(_02438_),
    .Y(_02441_),
    .B1(_02440_));
 sg13g2_nor2_1 _10459_ (.A(_02433_),
    .B(_02441_),
    .Y(_02442_));
 sg13g2_nor2_1 _10460_ (.A(_02437_),
    .B(_02442_),
    .Y(_02443_));
 sg13g2_a21oi_2 _10461_ (.B1(_02443_),
    .Y(_02444_),
    .A2(_02425_),
    .A1(_02354_));
 sg13g2_a22oi_1 _10462_ (.Y(_02445_),
    .B1(_02252_),
    .B2(_02444_),
    .A2(_02218_),
    .A1(_02138_));
 sg13g2_nand2_1 _10463_ (.Y(_02446_),
    .A(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .B(net1559));
 sg13g2_nand2_1 _10464_ (.Y(_02447_),
    .A(_02104_),
    .B(_02446_));
 sg13g2_nor4_1 _10465_ (.A(_01737_),
    .B(_01756_),
    .C(_01762_),
    .D(_02447_),
    .Y(_02448_));
 sg13g2_nor2_1 _10466_ (.A(net1352),
    .B(net360),
    .Y(_02449_));
 sg13g2_nor2_1 _10467_ (.A(net171),
    .B(_02104_),
    .Y(_02450_));
 sg13g2_nor4_1 _10468_ (.A(_02096_),
    .B(_02117_),
    .C(_02448_),
    .D(_02450_),
    .Y(_02451_));
 sg13g2_a21o_1 _10469_ (.A2(_02450_),
    .A1(_02117_),
    .B1(_02451_),
    .X(_02452_));
 sg13g2_a221oi_1 _10470_ (.B2(_02449_),
    .C1(_02452_),
    .B1(_02448_),
    .A1(_02096_),
    .Y(_02453_),
    .A2(_02117_));
 sg13g2_nor3_1 _10471_ (.A(net368),
    .B(_02078_),
    .C(_02086_),
    .Y(_02454_));
 sg13g2_nand3_1 _10472_ (.B(_02088_),
    .C(net241),
    .A(_01224_),
    .Y(_02455_));
 sg13g2_nand2_1 _10473_ (.Y(_02456_),
    .A(net187),
    .B(_02455_));
 sg13g2_o21ai_1 _10474_ (.B1(net359),
    .Y(_02457_),
    .A1(_02078_),
    .A2(_02088_));
 sg13g2_a21o_1 _10475_ (.A2(_02086_),
    .A1(net1283),
    .B1(_02080_),
    .X(_02458_));
 sg13g2_nor2_1 _10476_ (.A(net349),
    .B(net241),
    .Y(_02459_));
 sg13g2_a22oi_1 _10477_ (.Y(_02460_),
    .B1(_02459_),
    .B2(_01224_),
    .A2(_02458_),
    .A1(_02457_));
 sg13g2_nand2_1 _10478_ (.Y(_02461_),
    .A(net178),
    .B(_02460_));
 sg13g2_nor2_1 _10479_ (.A(net349),
    .B(_02112_),
    .Y(_02462_));
 sg13g2_a21oi_1 _10480_ (.A1(net356),
    .A2(_02078_),
    .Y(_02463_),
    .B1(net183));
 sg13g2_nor4_1 _10481_ (.A(_02080_),
    .B(_02454_),
    .C(_02462_),
    .D(_02463_),
    .Y(_02464_));
 sg13g2_a221oi_1 _10482_ (.B2(_02461_),
    .C1(_02464_),
    .B1(_02456_),
    .A1(_02080_),
    .Y(_02465_),
    .A2(_02454_));
 sg13g2_or2_1 _10483_ (.X(_02466_),
    .B(_02465_),
    .A(_02453_));
 sg13g2_inv_1 _10484_ (.Y(_02467_),
    .A(net1412));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(\cs_registers_i/_0631_ ));
 sg13g2_a221oi_1 _10486_ (.B2(\id_stage_i.controller_i.instr_i_12_ ),
    .C1(_02085_),
    .B1(_02083_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .Y(_02469_),
    .A2(net329));
 sg13g2_nor2_1 _10487_ (.A(_02467_),
    .B(_02469_),
    .Y(_02470_));
 sg13g2_nand2_2 _10488_ (.Y(_02471_),
    .A(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .B(net398));
 sg13g2_nand2_1 _10489_ (.Y(_02472_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_12__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10490_ (.B1(_02472_),
    .Y(_02473_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ),
    .A2(net2108));
 sg13g2_buf_2 fanout1129 (.A(net1130),
    .X(net1129));
 sg13g2_nor3_1 _10492_ (.A(net1468),
    .B(net1712),
    .C(net403),
    .Y(_02475_));
 sg13g2_a221oi_1 _10493_ (.B2(net1894),
    .C1(_02475_),
    .B1(_02473_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_11__$_NOT__A_Y ),
    .Y(_02476_),
    .A2(net405));
 sg13g2_nor3_1 _10494_ (.A(net362),
    .B(_02471_),
    .C(_02476_),
    .Y(_02477_));
 sg13g2_inv_2 _10495_ (.Y(_02478_),
    .A(net1467));
 sg13g2_a22oi_1 _10496_ (.Y(_02479_),
    .B1(_02321_),
    .B2(net1994),
    .A2(_01804_),
    .A1(net1999));
 sg13g2_nand2b_1 _10497_ (.Y(_02480_),
    .B(_01793_),
    .A_N(_02479_));
 sg13g2_nand3_1 _10498_ (.B(_02253_),
    .C(_01805_),
    .A(net513),
    .Y(_02481_));
 sg13g2_and2_1 _10499_ (.A(_02191_),
    .B(_02481_),
    .X(_02482_));
 sg13g2_a22oi_1 _10500_ (.Y(_02483_),
    .B1(_02480_),
    .B2(_02482_),
    .A2(net330),
    .A1(_02478_));
 sg13g2_nand3_1 _10501_ (.B(net368),
    .C(_02483_),
    .A(net1414),
    .Y(_02484_));
 sg13g2_nand2b_1 _10502_ (.Y(_02485_),
    .B(_02484_),
    .A_N(_02477_));
 sg13g2_nand2_1 _10503_ (.Y(_02486_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_13__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1972));
 sg13g2_o21ai_1 _10504_ (.B1(_02486_),
    .Y(_02487_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ),
    .A2(net2107));
 sg13g2_nor3_1 _10505_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .B(net1711),
    .C(net400),
    .Y(_02488_));
 sg13g2_a221oi_1 _10506_ (.B2(net1893),
    .C1(_02488_),
    .B1(_02487_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_12__$_NOT__A_Y ),
    .Y(_02489_),
    .A2(net405));
 sg13g2_buf_4 fanout1128 (.X(net1128),
    .A(_03060_));
 sg13g2_nand2_2 _10508_ (.Y(_02491_),
    .A(net2114),
    .B(net398));
 sg13g2_nand3_1 _10509_ (.B(_02489_),
    .C(_02491_),
    .A(net355),
    .Y(_02492_));
 sg13g2_nand3_1 _10510_ (.B(net373),
    .C(_02469_),
    .A(_02467_),
    .Y(_02493_));
 sg13g2_and2_1 _10511_ (.A(_02492_),
    .B(_02493_),
    .X(_02494_));
 sg13g2_nor3_1 _10512_ (.A(net362),
    .B(_02489_),
    .C(_02491_),
    .Y(_02495_));
 sg13g2_a221oi_1 _10513_ (.B2(_02494_),
    .C1(_02495_),
    .B1(_02485_),
    .A1(net378),
    .Y(_02496_),
    .A2(_02470_));
 sg13g2_nor2_1 _10514_ (.A(net361),
    .B(_02491_),
    .Y(_02497_));
 sg13g2_a21oi_1 _10515_ (.A1(net1412),
    .A2(net378),
    .Y(_02498_),
    .B1(_02497_));
 sg13g2_nor2b_1 _10516_ (.A(_02498_),
    .B_N(_02469_),
    .Y(_02499_));
 sg13g2_o21ai_1 _10517_ (.B1(_02492_),
    .Y(_02500_),
    .A1(net1412),
    .A2(net349));
 sg13g2_nand2b_1 _10518_ (.Y(_02501_),
    .B(_02500_),
    .A_N(_02469_));
 sg13g2_nand2_1 _10519_ (.Y(_02502_),
    .A(net1414),
    .B(net373));
 sg13g2_o21ai_1 _10520_ (.B1(_02502_),
    .Y(_02503_),
    .A1(net373),
    .A2(_02471_));
 sg13g2_nor2_1 _10521_ (.A(net362),
    .B(_02476_),
    .Y(_02504_));
 sg13g2_nand2b_1 _10522_ (.Y(_02505_),
    .B(_02483_),
    .A_N(_02504_));
 sg13g2_and3_1 _10523_ (.X(_02506_),
    .A(_02501_),
    .B(_02503_),
    .C(_02505_));
 sg13g2_nor3_1 _10524_ (.A(_02495_),
    .B(_02499_),
    .C(_02506_),
    .Y(_02507_));
 sg13g2_mux2_1 _10525_ (.A0(_02496_),
    .A1(_02507_),
    .S(net184),
    .X(_02508_));
 sg13g2_or2_1 _10526_ (.X(_02509_),
    .B(_02508_),
    .A(_02466_));
 sg13g2_nand3_1 _10527_ (.B(_02445_),
    .C(_02509_),
    .A(_02121_),
    .Y(_02510_));
 sg13g2_nand2_2 _10528_ (.Y(_02511_),
    .A(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .B(net1557));
 sg13g2_nand2_2 _10529_ (.Y(_02512_),
    .A(net1351),
    .B(net373));
 sg13g2_inv_1 _10530_ (.Y(_02513_),
    .A(_02512_));
 sg13g2_nand2_1 _10531_ (.Y(_02514_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_16__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1971));
 sg13g2_o21ai_1 _10532_ (.B1(_02514_),
    .Y(_02515_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ),
    .A2(net2106));
 sg13g2_buf_2 fanout1127 (.A(net1128),
    .X(net1127));
 sg13g2_nor3_1 _10534_ (.A(net1469),
    .B(net1709),
    .C(net403),
    .Y(_02517_));
 sg13g2_a221oi_1 _10535_ (.B2(net1892),
    .C1(_02517_),
    .B1(_02515_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_15__$_NOT__A_Y ),
    .Y(_02518_),
    .A2(net407));
 sg13g2_nor2_2 _10536_ (.A(net361),
    .B(_02518_),
    .Y(_02519_));
 sg13g2_a21oi_1 _10537_ (.A1(net2083),
    .A2(_01865_),
    .Y(_02520_),
    .B1(_01885_));
 sg13g2_nand2_1 _10538_ (.Y(_02521_),
    .A(net1999),
    .B(net1612));
 sg13g2_nand2_1 _10539_ (.Y(_02522_),
    .A(net2083),
    .B(_02098_));
 sg13g2_nand2_1 _10540_ (.Y(_02523_),
    .A(_02521_),
    .B(_02522_));
 sg13g2_nor2_1 _10541_ (.A(net347),
    .B(_02081_),
    .Y(_02524_));
 sg13g2_a22oi_1 _10542_ (.Y(_02525_),
    .B1(_02523_),
    .B2(_02524_),
    .A2(net329),
    .A1(net1469));
 sg13g2_o21ai_1 _10543_ (.B1(_02525_),
    .Y(_02526_),
    .A1(_01883_),
    .A2(_02520_));
 sg13g2_buf_2 fanout1126 (.A(net1127),
    .X(net1126));
 sg13g2_nor2_1 _10545_ (.A(net172),
    .B(net1343),
    .Y(_02528_));
 sg13g2_nor2_1 _10546_ (.A(_02519_),
    .B(_02528_),
    .Y(_02529_));
 sg13g2_nand3_1 _10547_ (.B(net110),
    .C(net1343),
    .A(_01228_),
    .Y(_02530_));
 sg13g2_o21ai_1 _10548_ (.B1(_02530_),
    .Y(_02531_),
    .A1(_02513_),
    .A2(_02529_));
 sg13g2_o21ai_1 _10549_ (.B1(_02511_),
    .Y(_02532_),
    .A1(net1343),
    .A2(_02512_));
 sg13g2_o21ai_1 _10550_ (.B1(_02511_),
    .Y(_02533_),
    .A1(net171),
    .A2(_02512_));
 sg13g2_a22oi_1 _10551_ (.Y(_02534_),
    .B1(_02533_),
    .B2(net1343),
    .A2(_02532_),
    .A1(net174));
 sg13g2_nor2_1 _10552_ (.A(_02519_),
    .B(_02534_),
    .Y(_02535_));
 sg13g2_a21oi_2 _10553_ (.B1(_02535_),
    .Y(_02536_),
    .A2(_02531_),
    .A1(_02511_));
 sg13g2_nand3_1 _10554_ (.B(net349),
    .C(net399),
    .A(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .Y(_02537_));
 sg13g2_o21ai_1 _10555_ (.B1(_02537_),
    .Y(_02538_),
    .A1(_01234_),
    .A2(net354));
 sg13g2_nand2_1 _10556_ (.Y(_02539_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_17__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10557_ (.B1(_02539_),
    .Y(_02540_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .A2(net2108));
 sg13g2_buf_4 fanout1125 (.X(net1125),
    .A(net1126));
 sg13g2_nor3_1 _10559_ (.A(net1471),
    .B(net1713),
    .C(net401),
    .Y(_02542_));
 sg13g2_a221oi_1 _10560_ (.B2(net1894),
    .C1(_02542_),
    .B1(_02540_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_16__$_NOT__A_Y ),
    .Y(_02543_),
    .A2(net405));
 sg13g2_nor2_1 _10561_ (.A(net373),
    .B(_02543_),
    .Y(_02544_));
 sg13g2_nand2_1 _10562_ (.Y(_02545_),
    .A(net531),
    .B(_02098_));
 sg13g2_a21oi_1 _10563_ (.A1(_02521_),
    .A2(_02545_),
    .Y(_02546_),
    .B1(net347));
 sg13g2_a21oi_1 _10564_ (.A1(net531),
    .A2(_01865_),
    .Y(_02547_),
    .B1(_01885_));
 sg13g2_nor2_1 _10565_ (.A(_01791_),
    .B(_02547_),
    .Y(_02548_));
 sg13g2_nor3_1 _10566_ (.A(net1613),
    .B(_02546_),
    .C(_02548_),
    .Y(_02549_));
 sg13g2_o21ai_1 _10567_ (.B1(_01773_),
    .Y(_02550_),
    .A1(net1471),
    .A2(_02037_));
 sg13g2_nor2_2 _10568_ (.A(_02549_),
    .B(_02550_),
    .Y(_02551_));
 sg13g2_nand2b_2 _10569_ (.Y(_02552_),
    .B(_02551_),
    .A_N(_02544_));
 sg13g2_nor2_1 _10570_ (.A(net171),
    .B(_02552_),
    .Y(_02553_));
 sg13g2_a21o_2 _10571_ (.A2(_02551_),
    .A1(net378),
    .B1(_02544_),
    .X(_02554_));
 sg13g2_or2_1 _10572_ (.X(_02555_),
    .B(_02554_),
    .A(net183));
 sg13g2_nor2b_1 _10573_ (.A(_02553_),
    .B_N(_02555_),
    .Y(_02556_));
 sg13g2_xor2_1 _10574_ (.B(_02556_),
    .A(_02538_),
    .X(_02557_));
 sg13g2_inv_1 _10575_ (.Y(_02558_),
    .A(_02524_));
 sg13g2_a22oi_1 _10576_ (.Y(_02559_),
    .B1(_02098_),
    .B2(\id_stage_i.controller_i.instr_i_18_ ),
    .A2(net1612),
    .A1(net1999));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(net1125));
 sg13g2_a21oi_1 _10578_ (.A1(\id_stage_i.controller_i.instr_i_18_ ),
    .A2(_01865_),
    .Y(_02561_),
    .B1(_01885_));
 sg13g2_nor2_1 _10579_ (.A(_01883_),
    .B(_02561_),
    .Y(_02562_));
 sg13g2_a21oi_1 _10580_ (.A1(net1516),
    .A2(net329),
    .Y(_02563_),
    .B1(_02562_));
 sg13g2_o21ai_1 _10581_ (.B1(_02563_),
    .Y(_02564_),
    .A1(_02558_),
    .A2(_02559_));
 sg13g2_nand2_1 _10582_ (.Y(_02565_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_19__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1974));
 sg13g2_o21ai_1 _10583_ (.B1(_02565_),
    .Y(_02566_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ),
    .A2(net2108));
 sg13g2_nor3_1 _10584_ (.A(net1516),
    .B(net1713),
    .C(net401),
    .Y(_02567_));
 sg13g2_a221oi_1 _10585_ (.B2(net1895),
    .C1(_02567_),
    .B1(_02566_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_18__$_NOT__A_Y ),
    .Y(_02568_),
    .A2(net406));
 sg13g2_nand2b_1 _10586_ (.Y(_02569_),
    .B(net354),
    .A_N(_02568_));
 sg13g2_o21ai_1 _10587_ (.B1(_02569_),
    .Y(_02570_),
    .A1(net171),
    .A2(_02564_));
 sg13g2_a21o_2 _10588_ (.A2(_02564_),
    .A1(net110),
    .B1(_02570_),
    .X(_02571_));
 sg13g2_inv_2 _10589_ (.Y(_02572_),
    .A(\ex_block_i.alu_i.imd_val_q_i_50_ ));
 sg13g2_nor3_1 _10590_ (.A(_02572_),
    .B(net372),
    .C(net1675),
    .Y(_02573_));
 sg13g2_a21oi_2 _10591_ (.B1(_02573_),
    .Y(_02574_),
    .A2(net379),
    .A1(net1203));
 sg13g2_xnor2_1 _10592_ (.Y(_02575_),
    .A(_02571_),
    .B(_02574_));
 sg13g2_inv_2 _10593_ (.Y(_02576_),
    .A(\ex_block_i.alu_i.imd_val_q_i_49_ ));
 sg13g2_nor3_1 _10594_ (.A(_02576_),
    .B(net372),
    .C(net1675),
    .Y(_02577_));
 sg13g2_a21oi_2 _10595_ (.B1(_02577_),
    .Y(_02578_),
    .A2(net379),
    .A1(net1250));
 sg13g2_nand2_1 _10596_ (.Y(_02579_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_18__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10597_ (.B1(_02579_),
    .Y(_02580_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ),
    .A2(net2109));
 sg13g2_buf_2 fanout1123 (.A(_04624_),
    .X(net1123));
 sg13g2_buf_2 fanout1122 (.A(_08071_),
    .X(net1122));
 sg13g2_buf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sg13g2_nor3_1 _10601_ (.A(net284),
    .B(net1713),
    .C(net404),
    .Y(_02584_));
 sg13g2_a221oi_1 _10602_ (.B2(net1894),
    .C1(_02584_),
    .B1(_02580_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_17__$_NOT__A_Y ),
    .Y(_02585_),
    .A2(net406));
 sg13g2_nand3_1 _10603_ (.B(net347),
    .C(net387),
    .A(net530),
    .Y(_02586_));
 sg13g2_o21ai_1 _10604_ (.B1(_02586_),
    .Y(_02587_),
    .A1(_01884_),
    .A2(net347));
 sg13g2_nor2b_1 _10605_ (.A(_01801_),
    .B_N(net525),
    .Y(_02588_));
 sg13g2_a22oi_1 _10606_ (.Y(_02589_),
    .B1(_02588_),
    .B2(_02098_),
    .A2(_02587_),
    .A1(net1612));
 sg13g2_and4_1 _10607_ (.A(net1999),
    .B(_01880_),
    .C(_01804_),
    .D(_02191_),
    .X(_02590_));
 sg13g2_a21oi_1 _10608_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ),
    .A2(net329),
    .Y(_02591_),
    .B1(_02590_));
 sg13g2_o21ai_1 _10609_ (.B1(_02591_),
    .Y(_02592_),
    .A1(_02081_),
    .A2(_02589_));
 sg13g2_o21ai_1 _10610_ (.B1(_02592_),
    .Y(_02593_),
    .A1(net370),
    .A2(_02585_));
 sg13g2_nand2_1 _10611_ (.Y(_02594_),
    .A(net360),
    .B(_02585_));
 sg13g2_o21ai_1 _10612_ (.B1(_02594_),
    .Y(_02595_),
    .A1(net354),
    .A2(_02592_));
 sg13g2_nor2_1 _10613_ (.A(net183),
    .B(_02595_),
    .Y(_02596_));
 sg13g2_a21oi_2 _10614_ (.B1(_02596_),
    .Y(_02597_),
    .A2(_02593_),
    .A1(net187));
 sg13g2_xor2_1 _10615_ (.B(_02597_),
    .A(_02578_),
    .X(_02598_));
 sg13g2_nand2_1 _10616_ (.Y(_02599_),
    .A(_02575_),
    .B(_02598_));
 sg13g2_inv_1 _10617_ (.Y(_02600_),
    .A(_02599_));
 sg13g2_nand2_1 _10618_ (.Y(_02601_),
    .A(_02557_),
    .B(_02600_));
 sg13g2_xnor2_1 _10619_ (.Y(_02602_),
    .A(net1412),
    .B(_02469_));
 sg13g2_xnor2_1 _10620_ (.Y(_02603_),
    .A(_02489_),
    .B(_02491_));
 sg13g2_nand2_1 _10621_ (.Y(_02604_),
    .A(net359),
    .B(_02603_));
 sg13g2_o21ai_1 _10622_ (.B1(_02604_),
    .Y(_02605_),
    .A1(net354),
    .A2(_02602_));
 sg13g2_nand2b_1 _10623_ (.Y(_02606_),
    .B(_02469_),
    .A_N(_02498_));
 sg13g2_nand3b_1 _10624_ (.B(_02606_),
    .C(_02501_),
    .Y(_02607_),
    .A_N(_02495_));
 sg13g2_mux2_2 _10625_ (.A0(_02605_),
    .A1(_02607_),
    .S(net183),
    .X(_02608_));
 sg13g2_xnor2_1 _10626_ (.Y(_02609_),
    .A(_02503_),
    .B(_02505_));
 sg13g2_o21ai_1 _10627_ (.B1(_02507_),
    .Y(_02610_),
    .A1(_02608_),
    .A2(_02609_));
 sg13g2_xor2_1 _10628_ (.B(_02483_),
    .A(net1414),
    .X(_02611_));
 sg13g2_xnor2_1 _10629_ (.Y(_02612_),
    .A(_02471_),
    .B(_02476_));
 sg13g2_nor2_1 _10630_ (.A(net363),
    .B(_02612_),
    .Y(_02613_));
 sg13g2_a21oi_1 _10631_ (.A1(net369),
    .A2(_02611_),
    .Y(_02614_),
    .B1(_02613_));
 sg13g2_o21ai_1 _10632_ (.B1(_02496_),
    .Y(_02615_),
    .A1(_02608_),
    .A2(_02614_));
 sg13g2_or2_1 _10633_ (.X(_02616_),
    .B(_02615_),
    .A(net184));
 sg13g2_o21ai_1 _10634_ (.B1(_02616_),
    .Y(_02617_),
    .A1(net174),
    .A2(_02610_));
 sg13g2_or2_1 _10635_ (.X(_02618_),
    .B(_02466_),
    .A(_02617_));
 sg13g2_and2_2 _10636_ (.A(_02121_),
    .B(_02618_),
    .X(_02619_));
 sg13g2_nand2_2 _10637_ (.Y(_02620_),
    .A(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .B(net399));
 sg13g2_nand2_1 _10638_ (.Y(_02621_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_22__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10639_ (.B1(_02621_),
    .Y(_02622_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ),
    .A2(net2108));
 sg13g2_buf_2 fanout1120 (.A(_08503_),
    .X(net1120));
 sg13g2_nor3_1 _10641_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_21_ ),
    .B(net1713),
    .C(net404),
    .Y(_02624_));
 sg13g2_a221oi_1 _10642_ (.B2(net1895),
    .C1(_02624_),
    .B1(_02622_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_21__$_NOT__A_Y ),
    .Y(_02625_),
    .A2(net407));
 sg13g2_xor2_1 _10643_ (.B(_02625_),
    .A(_02620_),
    .X(_02626_));
 sg13g2_buf_2 fanout1119 (.A(\cs_registers_i/_0507_ ),
    .X(net1119));
 sg13g2_nand2_2 _10645_ (.Y(_02628_),
    .A(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .B(net398));
 sg13g2_nand2_1 _10646_ (.Y(_02629_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_23__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1973));
 sg13g2_o21ai_1 _10647_ (.B1(_02629_),
    .Y(_02630_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ),
    .A2(net2108));
 sg13g2_buf_2 fanout1118 (.A(net1119),
    .X(net1118));
 sg13g2_nor3_1 _10649_ (.A(net1491),
    .B(net1712),
    .C(net404),
    .Y(_02632_));
 sg13g2_a221oi_1 _10650_ (.B2(net1894),
    .C1(_02632_),
    .B1(_02630_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_22__$_NOT__A_Y ),
    .Y(_02633_),
    .A2(net407));
 sg13g2_xor2_1 _10651_ (.B(_02633_),
    .A(_02628_),
    .X(_02634_));
 sg13g2_nand3_1 _10652_ (.B(_02626_),
    .C(_02634_),
    .A(net357),
    .Y(_02635_));
 sg13g2_inv_4 _10653_ (.A(net1520),
    .Y(_02636_));
 sg13g2_nand2_1 _10654_ (.Y(_02637_),
    .A(net448),
    .B(_02035_));
 sg13g2_a221oi_1 _10655_ (.B2(_02637_),
    .C1(_01992_),
    .B1(_01963_),
    .A1(_02636_),
    .Y(_02638_),
    .A2(net1614));
 sg13g2_buf_2 fanout1117 (.A(\cs_registers_i/_0546_ ),
    .X(net1117));
 sg13g2_xnor2_1 _10657_ (.Y(_02640_),
    .A(net126),
    .B(_02638_));
 sg13g2_a22oi_1 _10658_ (.Y(_02641_),
    .B1(_01934_),
    .B2(net447),
    .A2(net330),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_22_ ));
 sg13g2_nand2_2 _10659_ (.Y(_02642_),
    .A(_01931_),
    .B(_02641_));
 sg13g2_buf_1 fanout1116 (.A(\cs_registers_i/_0770_ ),
    .X(net1116));
 sg13g2_xor2_1 _10661_ (.B(net1397),
    .A(net195),
    .X(_02644_));
 sg13g2_nand3b_1 _10662_ (.B(_02644_),
    .C(net365),
    .Y(_02645_),
    .A_N(_02640_));
 sg13g2_inv_1 _10663_ (.Y(_02646_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_a22oi_1 _10664_ (.Y(_02647_),
    .B1(_01906_),
    .B2(_02646_),
    .A2(net1974),
    .A1(\ex_block_i.alu_i.multdiv_operand_b_i_21__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ));
 sg13g2_nor2_1 _10665_ (.A(_01839_),
    .B(_02647_),
    .Y(_02648_));
 sg13g2_buf_2 fanout1115 (.A(\cs_registers_i/_0770_ ),
    .X(net1115));
 sg13g2_nor3_1 _10667_ (.A(net287),
    .B(net1712),
    .C(net404),
    .Y(_02650_));
 sg13g2_a21o_1 _10668_ (.A2(net406),
    .A1(\ex_block_i.alu_i.imd_val_q_i_20__$_NOT__A_Y ),
    .B1(_02650_),
    .X(_02651_));
 sg13g2_o21ai_1 _10669_ (.B1(net360),
    .Y(_02652_),
    .A1(_02648_),
    .A2(_02651_));
 sg13g2_and2_1 _10670_ (.A(net287),
    .B(net332),
    .X(_02653_));
 sg13g2_a221oi_1 _10671_ (.B2(net464),
    .C1(_02653_),
    .B1(_01934_),
    .A1(_02191_),
    .Y(_02654_),
    .A2(_01862_));
 sg13g2_nor2_1 _10672_ (.A(\ex_block_i.alu_i.imd_val_q_i_20__$_NOT__A_Y ),
    .B(_02648_),
    .Y(_02655_));
 sg13g2_nand2_1 _10673_ (.Y(_02656_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .B(net398));
 sg13g2_nor3_1 _10674_ (.A(net363),
    .B(_02655_),
    .C(_02656_),
    .Y(_02657_));
 sg13g2_a21oi_1 _10675_ (.A1(net1281),
    .A2(net380),
    .Y(_02658_),
    .B1(_02657_));
 sg13g2_a21o_1 _10676_ (.A2(_02654_),
    .A1(_02652_),
    .B1(_02658_),
    .X(_02659_));
 sg13g2_nor2_1 _10677_ (.A(net1281),
    .B(net360),
    .Y(_02660_));
 sg13g2_a22oi_1 _10678_ (.Y(_02661_),
    .B1(_02660_),
    .B2(_02654_),
    .A2(_02656_),
    .A1(net350));
 sg13g2_inv_1 _10679_ (.Y(_02662_),
    .A(_02661_));
 sg13g2_nand2_1 _10680_ (.Y(_02663_),
    .A(_02652_),
    .B(_02662_));
 sg13g2_nand2_1 _10681_ (.Y(_02664_),
    .A(_02659_),
    .B(_02663_));
 sg13g2_a21oi_1 _10682_ (.A1(_02635_),
    .A2(_02645_),
    .Y(_02665_),
    .B1(_02664_));
 sg13g2_nand2_1 _10683_ (.Y(_02666_),
    .A(net513),
    .B(_02035_));
 sg13g2_nand2_1 _10684_ (.Y(_02667_),
    .A(_01861_),
    .B(_02666_));
 sg13g2_mux2_1 _10685_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ),
    .A1(_02667_),
    .S(_02037_),
    .X(_02668_));
 sg13g2_nand3_1 _10686_ (.B(_02652_),
    .C(_02668_),
    .A(_01773_),
    .Y(_02669_));
 sg13g2_nand2_1 _10687_ (.Y(_02670_),
    .A(net1281),
    .B(net372));
 sg13g2_o21ai_1 _10688_ (.B1(_02670_),
    .Y(_02671_),
    .A1(net364),
    .A2(_02656_));
 sg13g2_xnor2_1 _10689_ (.Y(_02672_),
    .A(_02669_),
    .B(_02671_));
 sg13g2_nor2_1 _10690_ (.A(net353),
    .B(_02644_),
    .Y(_02673_));
 sg13g2_nand2_1 _10691_ (.Y(_02674_),
    .A(_02625_),
    .B(net240));
 sg13g2_xnor2_1 _10692_ (.Y(_02675_),
    .A(_02620_),
    .B(_02674_));
 sg13g2_nand2_1 _10693_ (.Y(_02676_),
    .A(_02633_),
    .B(net1397));
 sg13g2_xor2_1 _10694_ (.B(_02676_),
    .A(_02628_),
    .X(_02677_));
 sg13g2_nor2_1 _10695_ (.A(net365),
    .B(_02677_),
    .Y(_02678_));
 sg13g2_a22oi_1 _10696_ (.Y(_02679_),
    .B1(_02675_),
    .B2(_02678_),
    .A2(_02673_),
    .A1(_02640_));
 sg13g2_nor3_1 _10697_ (.A(net172),
    .B(_02672_),
    .C(_02679_),
    .Y(_02680_));
 sg13g2_a21oi_2 _10698_ (.B1(_02680_),
    .Y(_02681_),
    .A2(_02665_),
    .A1(net181));
 sg13g2_nand2_1 _10699_ (.Y(_02682_),
    .A(\id_stage_i.controller_i.instr_i_19_ ),
    .B(_02083_));
 sg13g2_buf_4 fanout1114 (.X(net1114),
    .A(\cs_registers_i/_0773_ ));
 sg13g2_buf_8 fanout1113 (.A(_03077_),
    .X(net1113));
 sg13g2_a21oi_1 _10702_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ),
    .A2(net329),
    .Y(_02685_),
    .B1(_02085_));
 sg13g2_nand2_2 _10703_ (.Y(_02686_),
    .A(_02682_),
    .B(_02685_));
 sg13g2_buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sg13g2_xnor2_1 _10705_ (.Y(_02688_),
    .A(net178),
    .B(net170));
 sg13g2_a21o_1 _10706_ (.A2(net169),
    .A1(net1248),
    .B1(net356),
    .X(_02689_));
 sg13g2_a22oi_1 _10707_ (.Y(_02690_),
    .B1(_02689_),
    .B2(net178),
    .A2(net170),
    .A1(net351));
 sg13g2_o21ai_1 _10708_ (.B1(_02690_),
    .Y(_02691_),
    .A1(net1248),
    .A2(_02688_));
 sg13g2_buf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sg13g2_nand2_1 _10710_ (.Y(_02693_),
    .A(\ex_block_i.alu_i.multdiv_operand_b_i_20__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .B(net1972));
 sg13g2_o21ai_1 _10711_ (.B1(_02693_),
    .Y(_02694_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ),
    .A2(net2107));
 sg13g2_nor3_1 _10712_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ),
    .B(net1711),
    .C(net404),
    .Y(_02695_));
 sg13g2_a221oi_1 _10713_ (.B2(net1893),
    .C1(_02695_),
    .B1(_02694_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_19__$_NOT__A_Y ),
    .Y(_02696_),
    .A2(net406));
 sg13g2_nor2_1 _10714_ (.A(net363),
    .B(_02696_),
    .Y(_02697_));
 sg13g2_a21oi_2 _10715_ (.B1(_02697_),
    .Y(_02698_),
    .A2(net1560),
    .A1(\ex_block_i.alu_i.imd_val_q_i_51_ ));
 sg13g2_nand2b_1 _10716_ (.Y(_02699_),
    .B(net184),
    .A_N(net169));
 sg13g2_nand2b_1 _10717_ (.Y(_02700_),
    .B(net350),
    .A_N(_02696_));
 sg13g2_a22oi_1 _10718_ (.Y(_02701_),
    .B1(net1560),
    .B2(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .A2(net379),
    .A1(net1248));
 sg13g2_a21oi_1 _10719_ (.A1(_02699_),
    .A2(_02700_),
    .Y(_02702_),
    .B1(_02701_));
 sg13g2_a21oi_2 _10720_ (.B1(_02702_),
    .Y(_02703_),
    .A2(_02698_),
    .A1(_02691_));
 sg13g2_nand2b_1 _10721_ (.Y(_02704_),
    .B(_02703_),
    .A_N(_02681_));
 sg13g2_nor4_2 _10722_ (.A(_02536_),
    .B(_02601_),
    .C(_02619_),
    .Y(_02705_),
    .D(_02704_));
 sg13g2_o21ai_1 _10723_ (.B1(net408),
    .Y(_02706_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .A2(\ex_block_i.alu_i.imd_val_q_i_50_ ));
 sg13g2_nor3_1 _10724_ (.A(net1250),
    .B(net1203),
    .C(net359),
    .Y(_02707_));
 sg13g2_a21oi_2 _10725_ (.B1(_02707_),
    .Y(_02708_),
    .A2(_02706_),
    .A1(net359));
 sg13g2_inv_1 _10726_ (.Y(_02709_),
    .A(_02708_));
 sg13g2_a21oi_1 _10727_ (.A1(_02578_),
    .A2(_02709_),
    .Y(_02710_),
    .B1(_02574_));
 sg13g2_nand2b_1 _10728_ (.Y(_02711_),
    .B(_02574_),
    .A_N(_02571_));
 sg13g2_nand2_1 _10729_ (.Y(_02712_),
    .A(_02578_),
    .B(_02597_));
 sg13g2_inv_1 _10730_ (.Y(_02713_),
    .A(_02519_));
 sg13g2_a22oi_1 _10731_ (.Y(_02714_),
    .B1(_02512_),
    .B2(_02511_),
    .A2(net1343),
    .A1(_02713_));
 sg13g2_o21ai_1 _10732_ (.B1(_02714_),
    .Y(_02715_),
    .A1(_02538_),
    .A2(_02552_));
 sg13g2_nand2_1 _10733_ (.Y(_02716_),
    .A(_02538_),
    .B(_02552_));
 sg13g2_and2_1 _10734_ (.A(_02715_),
    .B(_02716_),
    .X(_02717_));
 sg13g2_inv_1 _10735_ (.Y(_02718_),
    .A(_02717_));
 sg13g2_a21o_1 _10736_ (.A2(_02515_),
    .A1(net1892),
    .B1(\ex_block_i.alu_i.imd_val_q_i_15__$_NOT__A_Y ),
    .X(_02719_));
 sg13g2_nand3_1 _10737_ (.B(net1558),
    .C(_02719_),
    .A(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .Y(_02720_));
 sg13g2_nor2_1 _10738_ (.A(_02519_),
    .B(net1343),
    .Y(_02721_));
 sg13g2_a21oi_1 _10739_ (.A1(_02512_),
    .A2(_02720_),
    .Y(_02722_),
    .B1(_02721_));
 sg13g2_o21ai_1 _10740_ (.B1(_02538_),
    .Y(_02723_),
    .A1(_02554_),
    .A2(_02722_));
 sg13g2_nand2_1 _10741_ (.Y(_02724_),
    .A(_02554_),
    .B(_02722_));
 sg13g2_nand2_1 _10742_ (.Y(_02725_),
    .A(_02723_),
    .B(_02724_));
 sg13g2_mux2_1 _10743_ (.A0(_02718_),
    .A1(_02725_),
    .S(net171),
    .X(_02726_));
 sg13g2_and2_1 _10744_ (.A(_02712_),
    .B(_02726_),
    .X(_02727_));
 sg13g2_nor2_1 _10745_ (.A(_02574_),
    .B(_02578_),
    .Y(_02728_));
 sg13g2_a21oi_1 _10746_ (.A1(_02571_),
    .A2(_02708_),
    .Y(_02729_),
    .B1(_02728_));
 sg13g2_nor2_1 _10747_ (.A(_02597_),
    .B(_02729_),
    .Y(_02730_));
 sg13g2_a221oi_1 _10748_ (.B2(_02727_),
    .C1(_02730_),
    .B1(_02711_),
    .A1(_02571_),
    .Y(_02731_),
    .A2(_02710_));
 sg13g2_nand2b_1 _10749_ (.Y(_02732_),
    .B(net369),
    .A_N(net195));
 sg13g2_nand3_1 _10750_ (.B(_02628_),
    .C(_02633_),
    .A(net360),
    .Y(_02733_));
 sg13g2_and2_1 _10751_ (.A(_02732_),
    .B(_02733_),
    .X(_02734_));
 sg13g2_inv_1 _10752_ (.Y(_02735_),
    .A(_02734_));
 sg13g2_and2_1 _10753_ (.A(net126),
    .B(net240),
    .X(_02736_));
 sg13g2_nor3_1 _10754_ (.A(net370),
    .B(_02620_),
    .C(_02625_),
    .Y(_02737_));
 sg13g2_a21oi_2 _10755_ (.B1(_02737_),
    .Y(_02738_),
    .A2(_02736_),
    .A1(_02110_));
 sg13g2_nor2_1 _10756_ (.A(net370),
    .B(_02620_),
    .Y(_02739_));
 sg13g2_a21oi_1 _10757_ (.A1(net126),
    .A2(net380),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_or2_1 _10758_ (.X(_02741_),
    .B(_02740_),
    .A(net240));
 sg13g2_a22oi_1 _10759_ (.Y(_02742_),
    .B1(_02738_),
    .B2(_02741_),
    .A2(_02735_),
    .A1(net1397));
 sg13g2_a21oi_1 _10760_ (.A1(net371),
    .A2(net1397),
    .Y(_02743_),
    .B1(_02734_));
 sg13g2_nor3_1 _10761_ (.A(net186),
    .B(_02738_),
    .C(_02743_),
    .Y(_02744_));
 sg13g2_a21oi_1 _10762_ (.A1(net188),
    .A2(_02742_),
    .Y(_02745_),
    .B1(_02744_));
 sg13g2_nand3_1 _10763_ (.B(net369),
    .C(net169),
    .A(net1248),
    .Y(_02746_));
 sg13g2_nand3_1 _10764_ (.B(net1560),
    .C(_02697_),
    .A(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .Y(_02747_));
 sg13g2_and2_1 _10765_ (.A(_02746_),
    .B(_02747_),
    .X(_02748_));
 sg13g2_nand2_2 _10766_ (.Y(_02749_),
    .A(_02659_),
    .B(_02748_));
 sg13g2_or2_1 _10767_ (.X(_02750_),
    .B(_02732_),
    .A(net1397));
 sg13g2_nand4_1 _10768_ (.B(_02733_),
    .C(_02749_),
    .A(_02663_),
    .Y(_02751_),
    .D(_02750_));
 sg13g2_nor2_1 _10769_ (.A(net186),
    .B(_02751_),
    .Y(_02752_));
 sg13g2_a21oi_1 _10770_ (.A1(net169),
    .A2(_02700_),
    .Y(_02753_),
    .B1(_02701_));
 sg13g2_a21oi_2 _10771_ (.B1(_02753_),
    .Y(_02754_),
    .A2(_02671_),
    .A1(_02669_));
 sg13g2_nand2_1 _10772_ (.Y(_02755_),
    .A(net1397),
    .B(_02735_));
 sg13g2_o21ai_1 _10773_ (.B1(_02755_),
    .Y(_02756_),
    .A1(_02669_),
    .A2(_02671_));
 sg13g2_nor3_1 _10774_ (.A(net172),
    .B(_02754_),
    .C(_02756_),
    .Y(_02757_));
 sg13g2_nand3_1 _10775_ (.B(_02620_),
    .C(_02625_),
    .A(net359),
    .Y(_02758_));
 sg13g2_o21ai_1 _10776_ (.B1(_02758_),
    .Y(_02759_),
    .A1(net126),
    .A2(net353));
 sg13g2_o21ai_1 _10777_ (.B1(_02759_),
    .Y(_02760_),
    .A1(net174),
    .A2(net240));
 sg13g2_a21o_1 _10778_ (.A2(net240),
    .A1(_01868_),
    .B1(_02760_),
    .X(_02761_));
 sg13g2_o21ai_1 _10779_ (.B1(_02761_),
    .Y(_02762_),
    .A1(_02752_),
    .A2(_02757_));
 sg13g2_nand2_1 _10780_ (.Y(_02763_),
    .A(net195),
    .B(net371));
 sg13g2_o21ai_1 _10781_ (.B1(_02763_),
    .Y(_02764_),
    .A1(net371),
    .A2(_02628_));
 sg13g2_nor2_1 _10782_ (.A(net172),
    .B(net1397),
    .Y(_02765_));
 sg13g2_and2_1 _10783_ (.A(net195),
    .B(_02642_),
    .X(_02766_));
 sg13g2_nor3_1 _10784_ (.A(net366),
    .B(_02628_),
    .C(_02633_),
    .Y(_02767_));
 sg13g2_a221oi_1 _10785_ (.B2(net110),
    .C1(_02767_),
    .B1(_02766_),
    .A1(_02764_),
    .Y(_02768_),
    .A2(_02765_));
 sg13g2_and3_1 _10786_ (.X(_02769_),
    .A(_02745_),
    .B(_02762_),
    .C(_02768_));
 sg13g2_o21ai_1 _10787_ (.B1(_02769_),
    .Y(_02770_),
    .A1(_02704_),
    .A2(_02731_));
 sg13g2_a21o_2 _10788_ (.A2(_02705_),
    .A1(_02510_),
    .B1(_02770_),
    .X(_02771_));
 sg13g2_buf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sg13g2_a21oi_1 _10790_ (.A1(net179),
    .A2(net1278),
    .Y(_02773_),
    .B1(net87));
 sg13g2_nor2_1 _10791_ (.A(net352),
    .B(_02773_),
    .Y(_02774_));
 sg13g2_buf_4 fanout1109 (.X(net1109),
    .A(net1110));
 sg13g2_nor2_1 _10793_ (.A(net176),
    .B(net1278),
    .Y(_02776_));
 sg13g2_nor4_1 _10794_ (.A(_02016_),
    .B(_02774_),
    .C(_02017_),
    .D(_02776_),
    .Y(_02777_));
 sg13g2_inv_1 _10795_ (.Y(_02778_),
    .A(_01983_));
 sg13g2_or2_1 _10796_ (.X(_02779_),
    .B(_02031_),
    .A(_02025_));
 sg13g2_a21oi_1 _10797_ (.A1(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .A2(net1558),
    .Y(_02780_),
    .B1(_02042_));
 sg13g2_a21oi_1 _10798_ (.A1(_02779_),
    .A2(net1344),
    .Y(_02781_),
    .B1(_02780_));
 sg13g2_inv_1 _10799_ (.Y(_02782_),
    .A(_02065_));
 sg13g2_nand2_1 _10800_ (.Y(_02783_),
    .A(_02060_),
    .B(_02782_));
 sg13g2_nor2_1 _10801_ (.A(_02781_),
    .B(_02783_),
    .Y(_02784_));
 sg13g2_nand2_1 _10802_ (.Y(_02785_),
    .A(_02781_),
    .B(_02783_));
 sg13g2_o21ai_1 _10803_ (.B1(_02785_),
    .Y(_02786_),
    .A1(_02056_),
    .A2(_02784_));
 sg13g2_o21ai_1 _10804_ (.B1(_02786_),
    .Y(_02787_),
    .A1(_02778_),
    .A2(_01994_));
 sg13g2_a21oi_1 _10805_ (.A1(net556),
    .A2(net402),
    .Y(_02788_),
    .B1(net364));
 sg13g2_nand2_1 _10806_ (.Y(_02789_),
    .A(net1344),
    .B(_02042_));
 sg13g2_a22oi_1 _10807_ (.Y(_02790_),
    .B1(_02779_),
    .B2(_02789_),
    .A2(_02788_),
    .A1(_02782_));
 sg13g2_o21ai_1 _10808_ (.B1(_02060_),
    .Y(_02791_),
    .A1(_02053_),
    .A2(_02790_));
 sg13g2_o21ai_1 _10809_ (.B1(_02065_),
    .Y(_02792_),
    .A1(_02790_),
    .A2(_02055_));
 sg13g2_o21ai_1 _10810_ (.B1(_02790_),
    .Y(_02793_),
    .A1(net125),
    .A2(net351));
 sg13g2_nand3_1 _10811_ (.B(_02792_),
    .C(_02793_),
    .A(_02791_),
    .Y(_02794_));
 sg13g2_nand2_1 _10812_ (.Y(_02795_),
    .A(_01995_),
    .B(_01983_));
 sg13g2_nand3_1 _10813_ (.B(_02794_),
    .C(_02795_),
    .A(net179),
    .Y(_02796_));
 sg13g2_o21ai_1 _10814_ (.B1(_02796_),
    .Y(_02797_),
    .A1(net173),
    .A2(_02787_));
 sg13g2_a21oi_1 _10815_ (.A1(net87),
    .A2(net379),
    .Y(_02798_),
    .B1(_02016_));
 sg13g2_nor3_1 _10816_ (.A(net176),
    .B(net1278),
    .C(_02798_),
    .Y(_02799_));
 sg13g2_and2_1 _10817_ (.A(net87),
    .B(_02004_),
    .X(_02800_));
 sg13g2_a22oi_1 _10818_ (.Y(_02801_),
    .B1(_02110_),
    .B2(_02800_),
    .A2(_02017_),
    .A1(_02016_));
 sg13g2_inv_1 _10819_ (.Y(_02802_),
    .A(_02801_));
 sg13g2_nor4_1 _10820_ (.A(_02797_),
    .B(_01998_),
    .C(_02799_),
    .D(_02802_),
    .Y(_02803_));
 sg13g2_nor2_2 _10821_ (.A(_02777_),
    .B(_02803_),
    .Y(_02804_));
 sg13g2_nand2_1 _10822_ (.Y(_02805_),
    .A(_01868_),
    .B(net1345));
 sg13g2_nand2_1 _10823_ (.Y(_02806_),
    .A(net1198),
    .B(net371));
 sg13g2_o21ai_1 _10824_ (.B1(_02806_),
    .Y(_02807_),
    .A1(net366),
    .A2(_01974_));
 sg13g2_nor2_1 _10825_ (.A(_01958_),
    .B(_02807_),
    .Y(_02808_));
 sg13g2_nand3b_1 _10826_ (.B(_02805_),
    .C(_02808_),
    .Y(_02809_),
    .A_N(_01966_));
 sg13g2_nand3_1 _10827_ (.B(_01926_),
    .C(_01950_),
    .A(_02809_),
    .Y(_02810_));
 sg13g2_nand2_1 _10828_ (.Y(_02811_),
    .A(_01855_),
    .B(_01876_));
 sg13g2_nor2b_1 _10829_ (.A(_02810_),
    .B_N(_02811_),
    .Y(_02812_));
 sg13g2_buf_2 fanout1108 (.A(net1109),
    .X(net1108));
 sg13g2_nand2_2 _10831_ (.Y(_02814_),
    .A(_01922_),
    .B(_01916_));
 sg13g2_a21oi_1 _10832_ (.A1(_01931_),
    .A2(_01935_),
    .Y(_02815_),
    .B1(_01941_));
 sg13g2_o21ai_1 _10833_ (.B1(_02815_),
    .Y(_02816_),
    .A1(_01929_),
    .A2(_02814_));
 sg13g2_nand2_1 _10834_ (.Y(_02817_),
    .A(_01929_),
    .B(_02814_));
 sg13g2_a22oi_1 _10835_ (.Y(_02818_),
    .B1(_02816_),
    .B2(_02817_),
    .A2(_01970_),
    .A1(_02807_));
 sg13g2_a21oi_1 _10836_ (.A1(_02808_),
    .A2(net1345),
    .Y(_02819_),
    .B1(_02818_));
 sg13g2_nand2_1 _10837_ (.Y(_02820_),
    .A(net367),
    .B(net1345));
 sg13g2_nand4_1 _10838_ (.B(net357),
    .C(net399),
    .A(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .Y(_02821_),
    .D(_01958_));
 sg13g2_a21o_1 _10839_ (.A2(_02821_),
    .A1(_02806_),
    .B1(_01968_),
    .X(_02822_));
 sg13g2_inv_1 _10840_ (.Y(_02823_),
    .A(_01909_));
 sg13g2_o21ai_1 _10841_ (.B1(_01900_),
    .Y(_02824_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_27__$_NOT__A_Y ),
    .A2(_02823_));
 sg13g2_a22oi_1 _10842_ (.Y(_02825_),
    .B1(_02824_),
    .B2(_01921_),
    .A2(_01893_),
    .A1(_01915_));
 sg13g2_nand2b_1 _10843_ (.Y(_02826_),
    .B(_01938_),
    .A_N(\ex_block_i.alu_i.imd_val_q_i_28__$_NOT__A_Y ));
 sg13g2_nand3_1 _10844_ (.B(net1558),
    .C(_02826_),
    .A(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .Y(_02827_));
 sg13g2_nor2_1 _10845_ (.A(_01941_),
    .B(net1346),
    .Y(_02828_));
 sg13g2_a21oi_1 _10846_ (.A1(_01946_),
    .A2(_02827_),
    .Y(_02829_),
    .B1(_02828_));
 sg13g2_a21oi_1 _10847_ (.A1(net371),
    .A2(net1346),
    .Y(_02830_),
    .B1(_01941_));
 sg13g2_o21ai_1 _10848_ (.B1(_01929_),
    .Y(_02831_),
    .A1(_01905_),
    .A2(_02830_));
 sg13g2_o21ai_1 _10849_ (.B1(_02831_),
    .Y(_02832_),
    .A1(_02825_),
    .A2(_02829_));
 sg13g2_a221oi_1 _10850_ (.B2(_02832_),
    .C1(net185),
    .B1(_02822_),
    .A1(_02808_),
    .Y(_02833_),
    .A2(_02820_));
 sg13g2_a21oi_2 _10851_ (.B1(_02833_),
    .Y(_02834_),
    .A2(_02819_),
    .A1(net190));
 sg13g2_o21ai_1 _10852_ (.B1(_02834_),
    .Y(_02835_),
    .A1(_01855_),
    .A2(_01876_));
 sg13g2_a22oi_1 _10853_ (.Y(_02836_),
    .B1(_02835_),
    .B2(_02811_),
    .A2(_02812_),
    .A1(_02804_));
 sg13g2_inv_1 _10854_ (.Y(_02837_),
    .A(_02836_));
 sg13g2_a21oi_1 _10855_ (.A1(_02071_),
    .A2(_02771_),
    .Y(_02838_),
    .B1(_02837_));
 sg13g2_xor2_1 _10856_ (.B(_02838_),
    .A(_01853_),
    .X(data_addr_o_31_));
 sg13g2_and2_1 _10857_ (.A(_01686_),
    .B(_01701_),
    .X(_02840_));
 sg13g2_nand2_1 _10858_ (.Y(_02841_),
    .A(_01686_),
    .B(_01697_));
 sg13g2_nand3_1 _10859_ (.B(_01669_),
    .C(_02841_),
    .A(_01719_),
    .Y(_02842_));
 sg13g2_a221oi_1 _10860_ (.B2(_02842_),
    .C1(_01754_),
    .B1(_01753_),
    .A1(_01662_),
    .Y(_02843_),
    .A2(_02840_));
 sg13g2_o21ai_1 _10861_ (.B1(_01724_),
    .Y(_02844_),
    .A1(net1581),
    .A2(_01738_));
 sg13g2_nand3_1 _10862_ (.B(_01730_),
    .C(_02844_),
    .A(net1580),
    .Y(_02845_));
 sg13g2_nor2b_2 _10863_ (.A(_02843_),
    .B_N(_02845_),
    .Y(_02846_));
 sg13g2_nand3b_1 _10864_ (.B(_02846_),
    .C(_01731_),
    .Y(_02847_),
    .A_N(net37));
 sg13g2_nand3b_1 _10865_ (.B(net37),
    .C(_01749_),
    .Y(_02848_),
    .A_N(_02846_));
 sg13g2_a21oi_1 _10866_ (.A1(_02847_),
    .A2(_02848_),
    .Y(_02849_),
    .B1(_01809_));
 sg13g2_nor2b_1 _10867_ (.A(_02846_),
    .B_N(_01731_),
    .Y(_02850_));
 sg13g2_nand2b_1 _10868_ (.Y(_02851_),
    .B(_02850_),
    .A_N(net36));
 sg13g2_nand3_1 _10869_ (.B(_02846_),
    .C(net36),
    .A(_01749_),
    .Y(_02852_));
 sg13g2_a21oi_1 _10870_ (.A1(_02851_),
    .A2(_02852_),
    .Y(_02853_),
    .B1(_01810_));
 sg13g2_a22oi_1 _10871_ (.Y(_02854_),
    .B1(_01810_),
    .B2(_01731_),
    .A2(_01809_),
    .A1(_01749_));
 sg13g2_a221oi_1 _10872_ (.B2(_01749_),
    .C1(_02846_),
    .B1(_01810_),
    .A1(_01731_),
    .Y(_02855_),
    .A2(_01809_));
 sg13g2_a21oi_1 _10873_ (.A1(_02846_),
    .A2(_02854_),
    .Y(_02856_),
    .B1(_02855_));
 sg13g2_nor3_2 _10874_ (.A(_02849_),
    .B(_02853_),
    .C(_02856_),
    .Y(_02857_));
 sg13g2_nor3_1 _10875_ (.A(\id_stage_i.id_fsm_q ),
    .B(net1490),
    .C(_01624_),
    .Y(_02858_));
 sg13g2_o21ai_1 _10876_ (.B1(_02858_),
    .Y(_02859_),
    .A1(_01751_),
    .A2(_02857_));
 sg13g2_nand2b_1 _10877_ (.Y(_02860_),
    .B(_02859_),
    .A_N(_01636_));
 sg13g2_a21oi_1 _10878_ (.A1(_01601_),
    .A2(_02860_),
    .Y(_02861_),
    .B1(net1715));
 sg13g2_nor2_1 _10879_ (.A(\id_stage_i.id_fsm_q ),
    .B(net1490),
    .Y(_02862_));
 sg13g2_nand2b_2 _10880_ (.Y(_02863_),
    .B(_02862_),
    .A_N(_01624_));
 sg13g2_nor2_1 _10881_ (.A(_02863_),
    .B(_01751_),
    .Y(_02864_));
 sg13g2_a21oi_1 _10882_ (.A1(_02857_),
    .A2(_02864_),
    .Y(_02865_),
    .B1(_01636_));
 sg13g2_o21ai_1 _10883_ (.B1(_02865_),
    .Y(_02866_),
    .A1(_02863_),
    .A2(_01750_));
 sg13g2_a21oi_1 _10884_ (.A1(_01601_),
    .A2(_02866_),
    .Y(_02867_),
    .B1(net1715));
 sg13g2_a21oi_2 _10885_ (.B1(_02804_),
    .Y(_02868_),
    .A2(_02771_),
    .A1(_02070_));
 sg13g2_o21ai_1 _10886_ (.B1(_02834_),
    .Y(_02869_),
    .A1(_02810_),
    .A2(_02868_));
 sg13g2_xnor2_1 _10887_ (.Y(data_addr_o_30_),
    .A(_01877_),
    .B(_02869_));
 sg13g2_xnor2_1 _10888_ (.Y(data_addr_o_27_),
    .A(_01926_),
    .B(_02868_));
 sg13g2_buf_2 fanout1107 (.A(net1108),
    .X(net1107));
 sg13g2_buf_2 fanout1106 (.A(net1108),
    .X(net1106));
 sg13g2_o21ai_1 _10891_ (.B1(_02128_),
    .Y(_02872_),
    .A1(net177),
    .A2(_02193_));
 sg13g2_xnor2_1 _10892_ (.Y(_02873_),
    .A(_02130_),
    .B(_02872_));
 sg13g2_xnor2_1 _10893_ (.Y(_02874_),
    .A(net190),
    .B(_02246_));
 sg13g2_nor2_1 _10894_ (.A(net353),
    .B(_02874_),
    .Y(_02875_));
 sg13g2_a21oi_1 _10895_ (.A1(net358),
    .A2(_02873_),
    .Y(_02876_),
    .B1(_02875_));
 sg13g2_nor2_1 _10896_ (.A(net186),
    .B(_02152_),
    .Y(_02877_));
 sg13g2_o21ai_1 _10897_ (.B1(_02145_),
    .Y(_02878_),
    .A1(net174),
    .A2(_02194_));
 sg13g2_nor2_1 _10898_ (.A(_02877_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_mux2_1 _10899_ (.A0(_02186_),
    .A1(_02212_),
    .S(net185),
    .X(_02880_));
 sg13g2_xnor2_1 _10900_ (.Y(_02881_),
    .A(net180),
    .B(_02245_));
 sg13g2_a21oi_1 _10901_ (.A1(net188),
    .A2(net1401),
    .Y(_02882_),
    .B1(_02181_));
 sg13g2_a21oi_1 _10902_ (.A1(net189),
    .A2(net1401),
    .Y(_02883_),
    .B1(_02182_));
 sg13g2_nor2_1 _10903_ (.A(_02180_),
    .B(_02883_),
    .Y(_02884_));
 sg13g2_nor3_1 _10904_ (.A(net367),
    .B(_02882_),
    .C(_02884_),
    .Y(_02885_));
 sg13g2_a21oi_2 _10905_ (.B1(_02885_),
    .Y(_02886_),
    .A2(_02881_),
    .A1(net366));
 sg13g2_nand2b_1 _10906_ (.Y(_02887_),
    .B(net176),
    .A_N(_02240_));
 sg13g2_o21ai_1 _10907_ (.B1(_02887_),
    .Y(_02888_),
    .A1(net175),
    .A2(_02224_));
 sg13g2_inv_1 _10908_ (.Y(_02889_),
    .A(_02888_));
 sg13g2_and2_1 _10909_ (.A(_02444_),
    .B(_02889_),
    .X(_02890_));
 sg13g2_nor2b_1 _10910_ (.A(_02886_),
    .B_N(_02890_),
    .Y(_02891_));
 sg13g2_nand2_1 _10911_ (.Y(_02892_),
    .A(_02188_),
    .B(_02879_));
 sg13g2_o21ai_1 _10912_ (.B1(_02892_),
    .Y(_02893_),
    .A1(_02880_),
    .A2(_02891_));
 sg13g2_o21ai_1 _10913_ (.B1(_02893_),
    .Y(_02894_),
    .A1(_02188_),
    .A2(_02879_));
 sg13g2_xor2_1 _10914_ (.B(_02894_),
    .A(_02876_),
    .X(_02895_));
 sg13g2_nand2_1 _10915_ (.Y(_02896_),
    .A(net1248),
    .B(net366));
 sg13g2_nand3_1 _10916_ (.B(_02698_),
    .C(_02896_),
    .A(net170),
    .Y(_02897_));
 sg13g2_a21o_1 _10917_ (.A2(_02897_),
    .A1(_02671_),
    .B1(_02669_),
    .X(_02898_));
 sg13g2_o21ai_1 _10918_ (.B1(_02898_),
    .Y(_02899_),
    .A1(_02671_),
    .A2(_02897_));
 sg13g2_o21ai_1 _10919_ (.B1(net368),
    .Y(_02900_),
    .A1(net1248),
    .A2(net169));
 sg13g2_nand3_1 _10920_ (.B(_02659_),
    .C(_02900_),
    .A(_02698_),
    .Y(_02901_));
 sg13g2_nand3_1 _10921_ (.B(_02663_),
    .C(_02901_),
    .A(net182),
    .Y(_02902_));
 sg13g2_o21ai_1 _10922_ (.B1(_02902_),
    .Y(_02903_),
    .A1(net177),
    .A2(_02899_));
 sg13g2_nor2_1 _10923_ (.A(_02536_),
    .B(_02601_),
    .Y(_02904_));
 sg13g2_nand2_1 _10924_ (.Y(_02905_),
    .A(_02138_),
    .B(_02218_));
 sg13g2_nor3_1 _10925_ (.A(net183),
    .B(_02605_),
    .C(_02614_),
    .Y(_02906_));
 sg13g2_nor3_1 _10926_ (.A(net174),
    .B(_02607_),
    .C(_02609_),
    .Y(_02907_));
 sg13g2_nor2_1 _10927_ (.A(_02906_),
    .B(_02907_),
    .Y(_02908_));
 sg13g2_o21ai_1 _10928_ (.B1(_02508_),
    .Y(_02909_),
    .A1(_02905_),
    .A2(_02908_));
 sg13g2_nand2b_1 _10929_ (.Y(_02910_),
    .B(_02909_),
    .A_N(_02466_));
 sg13g2_nor2_1 _10930_ (.A(_02466_),
    .B(_02908_),
    .Y(_02911_));
 sg13g2_nand3_1 _10931_ (.B(_02444_),
    .C(_02911_),
    .A(_02252_),
    .Y(_02912_));
 sg13g2_nand3_1 _10932_ (.B(_02910_),
    .C(_02912_),
    .A(_02121_),
    .Y(_02913_));
 sg13g2_nand2_1 _10933_ (.Y(_02914_),
    .A(_02904_),
    .B(_02913_));
 sg13g2_a21oi_1 _10934_ (.A1(_02728_),
    .A2(_02725_),
    .Y(_02915_),
    .B1(_02749_));
 sg13g2_nand2_1 _10935_ (.Y(_02916_),
    .A(net181),
    .B(_02915_));
 sg13g2_nand2_1 _10936_ (.Y(_02917_),
    .A(_02728_),
    .B(_02718_));
 sg13g2_nand3_1 _10937_ (.B(_02754_),
    .C(_02917_),
    .A(net190),
    .Y(_02918_));
 sg13g2_nor2_1 _10938_ (.A(_02597_),
    .B(_02709_),
    .Y(_02919_));
 sg13g2_or3_1 _10939_ (.A(_02710_),
    .B(_02727_),
    .C(_02919_),
    .X(_02920_));
 sg13g2_nor2b_1 _10940_ (.A(_02726_),
    .B_N(_02578_),
    .Y(_02921_));
 sg13g2_nor3_1 _10941_ (.A(_02574_),
    .B(_02597_),
    .C(_02921_),
    .Y(_02922_));
 sg13g2_a221oi_1 _10942_ (.B2(_02571_),
    .C1(_02922_),
    .B1(_02920_),
    .A1(_02916_),
    .Y(_02923_),
    .A2(_02918_));
 sg13g2_nand2_2 _10943_ (.Y(_02924_),
    .A(_02914_),
    .B(_02923_));
 sg13g2_nand2_2 _10944_ (.Y(_02925_),
    .A(_02903_),
    .B(_02924_));
 sg13g2_o21ai_1 _10945_ (.B1(_02625_),
    .Y(_02926_),
    .A1(net177),
    .A2(net240));
 sg13g2_xnor2_1 _10946_ (.Y(_02927_),
    .A(_02620_),
    .B(_02926_));
 sg13g2_xnor2_1 _10947_ (.Y(_02928_),
    .A(net182),
    .B(_02640_));
 sg13g2_nor2_1 _10948_ (.A(net352),
    .B(_02928_),
    .Y(_02929_));
 sg13g2_a21oi_1 _10949_ (.A1(net358),
    .A2(_02927_),
    .Y(_02930_),
    .B1(_02929_));
 sg13g2_xor2_1 _10950_ (.B(_02930_),
    .A(_02925_),
    .X(data_addr_o_21_));
 sg13g2_inv_2 _10951_ (.Y(_02931_),
    .A(data_addr_o_21_));
 sg13g2_o21ai_1 _10952_ (.B1(_01915_),
    .Y(_02932_),
    .A1(net177),
    .A2(_01896_));
 sg13g2_nor3_1 _10953_ (.A(net186),
    .B(_01921_),
    .C(_01893_),
    .Y(_02933_));
 sg13g2_o21ai_1 _10954_ (.B1(_01922_),
    .Y(_02934_),
    .A1(_02932_),
    .A2(_02933_));
 sg13g2_xor2_1 _10955_ (.B(_02934_),
    .A(_01950_),
    .X(_02935_));
 sg13g2_or2_1 _10956_ (.X(_02936_),
    .B(_02794_),
    .A(net185));
 sg13g2_o21ai_1 _10957_ (.B1(_02936_),
    .Y(_02937_),
    .A1(net177),
    .A2(_02786_));
 sg13g2_xnor2_1 _10958_ (.Y(_02938_),
    .A(_02000_),
    .B(_02937_));
 sg13g2_nand2_1 _10959_ (.Y(_02939_),
    .A(net188),
    .B(_02041_));
 sg13g2_nor2_1 _10960_ (.A(net186),
    .B(_02041_),
    .Y(_02940_));
 sg13g2_inv_1 _10961_ (.Y(_02941_),
    .A(_02779_));
 sg13g2_a21oi_1 _10962_ (.A1(_02042_),
    .A2(_02940_),
    .Y(_02942_),
    .B1(_02941_));
 sg13g2_o21ai_1 _10963_ (.B1(_02942_),
    .Y(_02943_),
    .A1(_02780_),
    .A2(_02939_));
 sg13g2_xnor2_1 _10964_ (.Y(_02944_),
    .A(_02068_),
    .B(_02943_));
 sg13g2_nor3_1 _10965_ (.A(_02052_),
    .B(_02938_),
    .C(_02944_),
    .Y(_02945_));
 sg13g2_o21ai_1 _10966_ (.B1(_02945_),
    .Y(_02946_),
    .A1(_02804_),
    .A2(_02935_));
 sg13g2_nand2_1 _10967_ (.Y(_02947_),
    .A(net366),
    .B(net175));
 sg13g2_nor2_1 _10968_ (.A(_02947_),
    .B(_01893_),
    .Y(_02948_));
 sg13g2_nor3_1 _10969_ (.A(_01922_),
    .B(_02948_),
    .C(_02932_),
    .Y(_02949_));
 sg13g2_xnor2_1 _10970_ (.Y(_02950_),
    .A(_01950_),
    .B(_02949_));
 sg13g2_nand2_1 _10971_ (.Y(_02951_),
    .A(_02804_),
    .B(_02950_));
 sg13g2_nor2b_1 _10972_ (.A(_02946_),
    .B_N(_02951_),
    .Y(_02952_));
 sg13g2_a21o_1 _10973_ (.A2(_01979_),
    .A1(_01853_),
    .B1(_02950_),
    .X(_02953_));
 sg13g2_o21ai_1 _10974_ (.B1(net368),
    .Y(_02954_),
    .A1(net122),
    .A2(_01896_));
 sg13g2_o21ai_1 _10975_ (.B1(net368),
    .Y(_02955_),
    .A1(net122),
    .A2(net176));
 sg13g2_a22oi_1 _10976_ (.Y(_02956_),
    .B1(_02955_),
    .B2(_01896_),
    .A2(_02954_),
    .A1(net176));
 sg13g2_inv_1 _10977_ (.Y(_02957_),
    .A(_02956_));
 sg13g2_nor2b_1 _10978_ (.A(_01900_),
    .B_N(_01915_),
    .Y(_02958_));
 sg13g2_a221oi_1 _10979_ (.B2(_02958_),
    .C1(_02933_),
    .B1(_02957_),
    .A1(_01922_),
    .Y(_02959_),
    .A2(_02932_));
 sg13g2_nand2_1 _10980_ (.Y(_02960_),
    .A(_02070_),
    .B(_02959_));
 sg13g2_a21oi_1 _10981_ (.A1(_02804_),
    .A2(_02959_),
    .Y(_02961_),
    .B1(_02935_));
 sg13g2_o21ai_1 _10982_ (.B1(net366),
    .Y(_02962_),
    .A1(net149),
    .A2(_02940_));
 sg13g2_and4_1 _10983_ (.A(_02025_),
    .B(_02032_),
    .C(_02962_),
    .D(_02939_),
    .X(_02963_));
 sg13g2_xnor2_1 _10984_ (.Y(_02964_),
    .A(_02068_),
    .B(_02963_));
 sg13g2_nand2_1 _10985_ (.Y(_02965_),
    .A(_02056_),
    .B(_02963_));
 sg13g2_nand2_1 _10986_ (.Y(_02966_),
    .A(_02067_),
    .B(_02965_));
 sg13g2_o21ai_1 _10987_ (.B1(_02966_),
    .Y(_02967_),
    .A1(_02056_),
    .A2(_02963_));
 sg13g2_xnor2_1 _10988_ (.Y(_02968_),
    .A(_02000_),
    .B(_02967_));
 sg13g2_nand3_1 _10989_ (.B(_02951_),
    .C(_02968_),
    .A(_02964_),
    .Y(_02969_));
 sg13g2_a221oi_1 _10990_ (.B2(_02961_),
    .C1(_02969_),
    .B1(_02960_),
    .A1(_02070_),
    .Y(_02970_),
    .A2(_02953_));
 sg13g2_mux2_1 _10991_ (.A0(_02952_),
    .A1(_02970_),
    .S(_02771_),
    .X(_02971_));
 sg13g2_a21oi_1 _10992_ (.A1(net180),
    .A2(net1343),
    .Y(_02972_),
    .B1(net1351));
 sg13g2_or2_1 _10993_ (.X(_02973_),
    .B(_02972_),
    .A(net351));
 sg13g2_nand3_1 _10994_ (.B(_02529_),
    .C(_02973_),
    .A(_02511_),
    .Y(_02974_));
 sg13g2_o21ai_1 _10995_ (.B1(_02703_),
    .Y(_02975_),
    .A1(_02052_),
    .A2(_02681_));
 sg13g2_nand2_1 _10996_ (.Y(_02976_),
    .A(_02600_),
    .B(_02975_));
 sg13g2_nand3_1 _10997_ (.B(_02974_),
    .C(_02976_),
    .A(_02557_),
    .Y(_02977_));
 sg13g2_or2_1 _10998_ (.X(_02978_),
    .B(_02974_),
    .A(_02557_));
 sg13g2_a21oi_1 _10999_ (.A1(_02977_),
    .A2(_02978_),
    .Y(_02979_),
    .B1(_02536_));
 sg13g2_nand2b_1 _11000_ (.Y(_02980_),
    .B(_02555_),
    .A_N(_02553_));
 sg13g2_or2_1 _11001_ (.X(_02981_),
    .B(_02597_),
    .A(_02578_));
 sg13g2_mux2_1 _11002_ (.A0(_02712_),
    .A1(_02981_),
    .S(_02575_),
    .X(_02982_));
 sg13g2_nand2_1 _11003_ (.Y(_02983_),
    .A(_02980_),
    .B(_02982_));
 sg13g2_mux2_2 _11004_ (.A0(_02714_),
    .A1(_02722_),
    .S(net176),
    .X(_02984_));
 sg13g2_nand2_1 _11005_ (.Y(_02985_),
    .A(_02974_),
    .B(_02984_));
 sg13g2_o21ai_1 _11006_ (.B1(_02985_),
    .Y(_02986_),
    .A1(_02983_),
    .A2(_02984_));
 sg13g2_nand3_1 _11007_ (.B(_02974_),
    .C(_02984_),
    .A(_02557_),
    .Y(_02987_));
 sg13g2_o21ai_1 _11008_ (.B1(_02987_),
    .Y(_02988_),
    .A1(_02557_),
    .A2(_02986_));
 sg13g2_nand2_1 _11009_ (.Y(_02989_),
    .A(_02536_),
    .B(_02988_));
 sg13g2_nor2_1 _11010_ (.A(_02913_),
    .B(_02989_),
    .Y(_02990_));
 sg13g2_a21oi_1 _11011_ (.A1(_02913_),
    .A2(_02979_),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_and2_1 _11012_ (.A(_02704_),
    .B(_02769_),
    .X(_02992_));
 sg13g2_nand3b_1 _11013_ (.B(_02964_),
    .C(_02071_),
    .Y(_02993_),
    .A_N(_02992_));
 sg13g2_nor2_1 _11014_ (.A(_01853_),
    .B(_02837_),
    .Y(_02994_));
 sg13g2_nand2_1 _11015_ (.Y(_02995_),
    .A(_02993_),
    .B(_02994_));
 sg13g2_nor2b_1 _11016_ (.A(_02608_),
    .B_N(_02503_),
    .Y(_02996_));
 sg13g2_nand2_1 _11017_ (.Y(_02997_),
    .A(_02480_),
    .B(_02482_));
 sg13g2_o21ai_1 _11018_ (.B1(_02997_),
    .Y(_02998_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ),
    .A2(_02191_));
 sg13g2_a21oi_1 _11019_ (.A1(net189),
    .A2(_02998_),
    .Y(_02999_),
    .B1(_02504_));
 sg13g2_o21ai_1 _11020_ (.B1(_02999_),
    .Y(_03000_),
    .A1(_02947_),
    .A2(_02998_));
 sg13g2_inv_1 _11021_ (.Y(_03001_),
    .A(_02608_));
 sg13g2_nor3_1 _11022_ (.A(_03001_),
    .B(_02503_),
    .C(_03000_),
    .Y(_03002_));
 sg13g2_a21o_1 _11023_ (.A2(_03000_),
    .A1(_02996_),
    .B1(_03002_),
    .X(_03003_));
 sg13g2_xnor2_1 _11024_ (.Y(_03004_),
    .A(_02503_),
    .B(_03000_));
 sg13g2_nor3_1 _11025_ (.A(_02608_),
    .B(_02445_),
    .C(_03004_),
    .Y(_03005_));
 sg13g2_a21o_1 _11026_ (.A2(_03003_),
    .A1(_02445_),
    .B1(_03005_),
    .X(_03006_));
 sg13g2_a22oi_1 _11027_ (.Y(_03007_),
    .B1(_02348_),
    .B2(net379),
    .A2(_02330_),
    .A1(_02319_));
 sg13g2_o21ai_1 _11028_ (.B1(_02398_),
    .Y(_03008_),
    .A1(_03007_),
    .A2(_02401_));
 sg13g2_xnor2_1 _11029_ (.Y(_03009_),
    .A(_02349_),
    .B(_03008_));
 sg13g2_nand2_1 _11030_ (.Y(_03010_),
    .A(_02404_),
    .B(_02405_));
 sg13g2_o21ai_1 _11031_ (.B1(_02408_),
    .Y(_03011_),
    .A1(_02404_),
    .A2(_02405_));
 sg13g2_nand3_1 _11032_ (.B(_03010_),
    .C(_03011_),
    .A(_02417_),
    .Y(_03012_));
 sg13g2_nand2_2 _11033_ (.Y(_03013_),
    .A(_02413_),
    .B(_03012_));
 sg13g2_xor2_1 _11034_ (.B(_03013_),
    .A(_02288_),
    .X(_03014_));
 sg13g2_nor2_1 _11035_ (.A(net173),
    .B(_03014_),
    .Y(_03015_));
 sg13g2_a21oi_2 _11036_ (.B1(_03015_),
    .Y(_03016_),
    .A2(_03009_),
    .A1(net181));
 sg13g2_xnor2_1 _11037_ (.Y(data_addr_o_3_),
    .A(_02290_),
    .B(_03016_));
 sg13g2_a21o_1 _11038_ (.A2(_02814_),
    .A1(_02815_),
    .B1(_01929_),
    .X(_03017_));
 sg13g2_o21ai_1 _11039_ (.B1(_03017_),
    .Y(_03018_),
    .A1(_02815_),
    .A2(_02814_));
 sg13g2_o21ai_1 _11040_ (.B1(net1346),
    .Y(_03019_),
    .A1(net1200),
    .A2(_02825_));
 sg13g2_o21ai_1 _11041_ (.B1(net1200),
    .Y(_03020_),
    .A1(_01941_),
    .A2(_02825_));
 sg13g2_a21o_1 _11042_ (.A2(_03020_),
    .A1(_03019_),
    .B1(net358),
    .X(_03021_));
 sg13g2_nand2b_1 _11043_ (.Y(_03022_),
    .B(_02825_),
    .A_N(_01949_));
 sg13g2_nand3_1 _11044_ (.B(net1557),
    .C(_01941_),
    .A(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .Y(_03023_));
 sg13g2_nand4_1 _11045_ (.B(_03021_),
    .C(_03022_),
    .A(net181),
    .Y(_03024_),
    .D(_03023_));
 sg13g2_o21ai_1 _11046_ (.B1(_03024_),
    .Y(_03025_),
    .A1(net176),
    .A2(_03018_));
 sg13g2_nand2_1 _11047_ (.Y(_03026_),
    .A(_01951_),
    .B(_03025_));
 sg13g2_xor2_1 _11048_ (.B(_03026_),
    .A(_01978_),
    .X(_03027_));
 sg13g2_a21oi_1 _11049_ (.A1(_01876_),
    .A2(_02834_),
    .Y(_03028_),
    .B1(_01855_));
 sg13g2_nor2_1 _11050_ (.A(_01876_),
    .B(_02834_),
    .Y(_03029_));
 sg13g2_o21ai_1 _11051_ (.B1(_01853_),
    .Y(_03030_),
    .A1(_03028_),
    .A2(_03029_));
 sg13g2_nand2_1 _11052_ (.Y(_03031_),
    .A(_02538_),
    .B(_02974_));
 sg13g2_nor2_1 _11053_ (.A(_02538_),
    .B(_02974_),
    .Y(_03032_));
 sg13g2_a21o_1 _11054_ (.A2(_03031_),
    .A1(_02980_),
    .B1(_03032_),
    .X(_03033_));
 sg13g2_nor2_1 _11055_ (.A(_02703_),
    .B(_02731_),
    .Y(_03034_));
 sg13g2_a21oi_1 _11056_ (.A1(_02982_),
    .A2(_03033_),
    .Y(_03035_),
    .B1(_03034_));
 sg13g2_and2_1 _11057_ (.A(net110),
    .B(_02104_),
    .X(_03036_));
 sg13g2_nor3_1 _11058_ (.A(_02096_),
    .B(_02450_),
    .C(_03036_),
    .Y(_03037_));
 sg13g2_nor2_1 _11059_ (.A(_02117_),
    .B(_03037_),
    .Y(_03038_));
 sg13g2_xor2_1 _11060_ (.B(_03038_),
    .A(_02465_),
    .X(_03039_));
 sg13g2_nand3_1 _11061_ (.B(_02453_),
    .C(_03039_),
    .A(_02617_),
    .Y(_03040_));
 sg13g2_mux2_1 _11062_ (.A0(_02348_),
    .A1(_02395_),
    .S(net353),
    .X(_03041_));
 sg13g2_xnor2_1 _11063_ (.Y(_03042_),
    .A(_02317_),
    .B(_02399_));
 sg13g2_xor2_1 _11064_ (.B(net1398),
    .A(net1409),
    .X(_03043_));
 sg13g2_nor2_1 _11065_ (.A(net353),
    .B(_03043_),
    .Y(_03044_));
 sg13g2_a21oi_1 _11066_ (.A1(net357),
    .A2(_03042_),
    .Y(_03045_),
    .B1(_03044_));
 sg13g2_xnor2_1 _11067_ (.Y(_03046_),
    .A(_03041_),
    .B(_03045_));
 sg13g2_nand2_1 _11068_ (.Y(_03047_),
    .A(_02409_),
    .B(_02410_));
 sg13g2_nand2_1 _11069_ (.Y(_03048_),
    .A(_02317_),
    .B(net1398));
 sg13g2_xnor2_1 _11070_ (.Y(_03049_),
    .A(_02399_),
    .B(_03048_));
 sg13g2_a21oi_1 _11071_ (.A1(net357),
    .A2(_03049_),
    .Y(_03050_),
    .B1(_03044_));
 sg13g2_xnor2_1 _11072_ (.Y(_03051_),
    .A(_03047_),
    .B(_03050_));
 sg13g2_mux2_2 _11073_ (.A0(_03046_),
    .A1(_03051_),
    .S(net185),
    .X(data_addr_o_2_));
 sg13g2_buf_1 fanout1105 (.A(net1110),
    .X(net1105));
 sg13g2_and3_1 _11075_ (.X(_03053_),
    .A(net197),
    .B(net371),
    .C(net1457));
 sg13g2_nor2_1 _11076_ (.A(_02304_),
    .B(net1675),
    .Y(_03054_));
 sg13g2_o21ai_1 _11077_ (.B1(_03054_),
    .Y(_03055_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_0__$_NOT__A_Y ),
    .A2(_02308_));
 sg13g2_nand2_1 _11078_ (.Y(_03056_),
    .A(net180),
    .B(_02309_));
 sg13g2_a21oi_1 _11079_ (.A1(_03055_),
    .A2(_03056_),
    .Y(_03057_),
    .B1(net366));
 sg13g2_and4_1 _11080_ (.A(\ex_block_i.alu_i.imd_val_q_i_32_ ),
    .B(net187),
    .C(net1559),
    .D(net1457),
    .X(_03058_));
 sg13g2_nor4_2 _11081_ (.A(_02408_),
    .B(_03053_),
    .C(_03057_),
    .Y(_03059_),
    .D(_03058_));
 sg13g2_inv_1 _11082_ (.Y(_03060_),
    .A(net1145));
 sg13g2_and2_2 _11083_ (.A(_02340_),
    .B(_02341_),
    .X(_03061_));
 sg13g2_buf_1 fanout1104 (.A(net1105),
    .X(net1104));
 sg13g2_xor2_1 _11085_ (.B(_02346_),
    .A(net1247),
    .X(_03063_));
 sg13g2_xnor2_1 _11086_ (.Y(_03064_),
    .A(_02300_),
    .B(_02309_));
 sg13g2_nand2_1 _11087_ (.Y(_03065_),
    .A(net357),
    .B(_03064_));
 sg13g2_o21ai_1 _11088_ (.B1(_03065_),
    .Y(_03066_),
    .A1(net350),
    .A2(_03063_));
 sg13g2_inv_4 _11089_ (.A(net1457),
    .Y(_03067_));
 sg13g2_nor2_1 _11090_ (.A(_03067_),
    .B(_02405_),
    .Y(_03068_));
 sg13g2_o21ai_1 _11091_ (.B1(_02406_),
    .Y(_03069_),
    .A1(_02300_),
    .A2(_02407_));
 sg13g2_nand2_1 _11092_ (.Y(_03070_),
    .A(_03067_),
    .B(_03069_));
 sg13g2_nor2_1 _11093_ (.A(net369),
    .B(_02309_),
    .Y(_03071_));
 sg13g2_a21o_1 _11094_ (.A2(net378),
    .A1(net198),
    .B1(_03071_),
    .X(_03072_));
 sg13g2_a22oi_1 _11095_ (.Y(_03073_),
    .B1(_03072_),
    .B2(net1247),
    .A2(_03071_),
    .A1(_02300_));
 sg13g2_o21ai_1 _11096_ (.B1(_03073_),
    .Y(_03074_),
    .A1(net1247),
    .A2(_03070_));
 sg13g2_o21ai_1 _11097_ (.B1(net188),
    .Y(_03075_),
    .A1(_03068_),
    .A2(_03074_));
 sg13g2_o21ai_1 _11098_ (.B1(_03075_),
    .Y(_03076_),
    .A1(net185),
    .A2(_03066_));
 sg13g2_xor2_1 _11099_ (.B(_03076_),
    .A(_02404_),
    .X(_03077_));
 sg13g2_nor2_2 _11100_ (.A(net1128),
    .B(net1113),
    .Y(_03078_));
 sg13g2_xnor2_1 _11101_ (.Y(_03079_),
    .A(_02440_),
    .B(_02391_));
 sg13g2_a21oi_1 _11102_ (.A1(net180),
    .A2(_02435_),
    .Y(_03080_),
    .B1(_02438_));
 sg13g2_or2_1 _11103_ (.X(_03081_),
    .B(_03080_),
    .A(_02429_));
 sg13g2_nand2_1 _11104_ (.Y(_03082_),
    .A(_02368_),
    .B(_03081_));
 sg13g2_mux2_1 _11105_ (.A0(_02664_),
    .A1(_02672_),
    .S(net184),
    .X(_03083_));
 sg13g2_a21oi_1 _11106_ (.A1(net179),
    .A2(net170),
    .Y(_03084_),
    .B1(net1248));
 sg13g2_or2_1 _11107_ (.X(_03085_),
    .B(_03084_),
    .A(net351));
 sg13g2_nand3_1 _11108_ (.B(_02698_),
    .C(_03085_),
    .A(_02699_),
    .Y(_03086_));
 sg13g2_xnor2_1 _11109_ (.Y(_03087_),
    .A(_03083_),
    .B(_03086_));
 sg13g2_a21oi_1 _11110_ (.A1(_03079_),
    .A2(_03082_),
    .Y(_03088_),
    .B1(_03087_));
 sg13g2_nand3b_1 _11111_ (.B(_03078_),
    .C(_03088_),
    .Y(_03089_),
    .A_N(data_addr_o_2_));
 sg13g2_a21oi_2 _11112_ (.B1(_03089_),
    .Y(_03090_),
    .A2(_03040_),
    .A1(_02618_));
 sg13g2_nand4_1 _11113_ (.B(_03030_),
    .C(_03035_),
    .A(_03027_),
    .Y(_03091_),
    .D(_03090_));
 sg13g2_nand2b_1 _11114_ (.Y(_03092_),
    .B(_02770_),
    .A_N(_02052_));
 sg13g2_nand3_1 _11115_ (.B(_02804_),
    .C(_02812_),
    .A(_01853_),
    .Y(_03093_));
 sg13g2_nand3_1 _11116_ (.B(_02355_),
    .C(_02359_),
    .A(net179),
    .Y(_03094_));
 sg13g2_o21ai_1 _11117_ (.B1(_03094_),
    .Y(_03095_),
    .A1(net352),
    .A2(_02262_));
 sg13g2_o21ai_1 _11118_ (.B1(net366),
    .Y(_03096_),
    .A1(net1406),
    .A2(net1399));
 sg13g2_o21ai_1 _11119_ (.B1(net365),
    .Y(_03097_),
    .A1(net1406),
    .A2(net173));
 sg13g2_a22oi_1 _11120_ (.Y(_03098_),
    .B1(_03097_),
    .B2(net1399),
    .A2(_03096_),
    .A1(net175));
 sg13g2_o21ai_1 _11121_ (.B1(_02355_),
    .Y(_03099_),
    .A1(_02358_),
    .A2(_03098_));
 sg13g2_nand4_1 _11122_ (.B(net1560),
    .C(_02262_),
    .A(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .Y(_03100_),
    .D(_02362_));
 sg13g2_a22oi_1 _11123_ (.Y(_03101_),
    .B1(_03099_),
    .B2(_03100_),
    .A2(_03095_),
    .A1(net1406));
 sg13g2_nand2_1 _11124_ (.Y(_03102_),
    .A(net180),
    .B(_02349_));
 sg13g2_o21ai_1 _11125_ (.B1(_03102_),
    .Y(_03103_),
    .A1(net172),
    .A2(_02288_));
 sg13g2_a21oi_1 _11126_ (.A1(_02290_),
    .A2(_03103_),
    .Y(_03104_),
    .B1(_02419_));
 sg13g2_nor2_1 _11127_ (.A(_02353_),
    .B(_03104_),
    .Y(_03105_));
 sg13g2_xnor2_1 _11128_ (.Y(data_addr_o_4_),
    .A(_03101_),
    .B(_03105_));
 sg13g2_a21oi_1 _11129_ (.A1(_02376_),
    .A2(_02368_),
    .Y(_03106_),
    .B1(_02369_));
 sg13g2_a21oi_1 _11130_ (.A1(_02428_),
    .A2(_02368_),
    .Y(_03107_),
    .B1(_03106_));
 sg13g2_xnor2_1 _11131_ (.Y(_03108_),
    .A(net1404),
    .B(_02435_));
 sg13g2_xnor2_1 _11132_ (.Y(_03109_),
    .A(net180),
    .B(_03108_));
 sg13g2_nor2_1 _11133_ (.A(net352),
    .B(_03109_),
    .Y(_03110_));
 sg13g2_a21oi_2 _11134_ (.B1(_03110_),
    .Y(_03111_),
    .A2(_03107_),
    .A1(net357));
 sg13g2_nand2_1 _11135_ (.Y(_03112_),
    .A(_02372_),
    .B(_02379_));
 sg13g2_nor2_1 _11136_ (.A(_03112_),
    .B(_03079_),
    .Y(_03113_));
 sg13g2_a21oi_1 _11137_ (.A1(_02282_),
    .A2(_02288_),
    .Y(_03114_),
    .B1(_03013_));
 sg13g2_nor2_1 _11138_ (.A(_02421_),
    .B(_03114_),
    .Y(_03115_));
 sg13g2_a21oi_1 _11139_ (.A1(net1399),
    .A2(_02271_),
    .Y(_03116_),
    .B1(net172));
 sg13g2_or2_1 _11140_ (.X(_03117_),
    .B(_02349_),
    .A(_02290_));
 sg13g2_nand2_1 _11141_ (.Y(_03118_),
    .A(_03008_),
    .B(_03117_));
 sg13g2_a221oi_1 _11142_ (.B2(_02269_),
    .C1(net184),
    .B1(_03096_),
    .A1(_02290_),
    .Y(_03119_),
    .A2(_02349_));
 sg13g2_a221oi_1 _11143_ (.B2(_03119_),
    .C1(_02363_),
    .B1(_03118_),
    .A1(_03115_),
    .Y(_03120_),
    .A2(_03116_));
 sg13g2_mux2_1 _11144_ (.A0(_03111_),
    .A1(_03113_),
    .S(_03120_),
    .X(_03121_));
 sg13g2_nor2_1 _11145_ (.A(data_addr_o_4_),
    .B(_03121_),
    .Y(_03122_));
 sg13g2_nand3_1 _11146_ (.B(_03093_),
    .C(_03122_),
    .A(_03092_),
    .Y(_03123_));
 sg13g2_nor3_1 _11147_ (.A(data_addr_o_3_),
    .B(_03091_),
    .C(_03123_),
    .Y(_03124_));
 sg13g2_xor2_1 _11148_ (.B(_02233_),
    .A(_02212_),
    .X(_03125_));
 sg13g2_or2_1 _11149_ (.X(_03126_),
    .B(_02186_),
    .A(_02157_));
 sg13g2_nand3_1 _11150_ (.B(_02187_),
    .C(_03126_),
    .A(net182),
    .Y(_03127_));
 sg13g2_o21ai_1 _11151_ (.B1(_03127_),
    .Y(_03128_),
    .A1(net177),
    .A2(_03125_));
 sg13g2_o21ai_1 _11152_ (.B1(net1400),
    .Y(_03129_),
    .A1(_02205_),
    .A2(_02207_));
 sg13g2_nor3_1 _11153_ (.A(net184),
    .B(net1400),
    .C(_02220_),
    .Y(_03130_));
 sg13g2_nor2_1 _11154_ (.A(_02174_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_o21ai_1 _11155_ (.B1(_03131_),
    .Y(_03132_),
    .A1(net175),
    .A2(_03129_));
 sg13g2_xnor2_1 _11156_ (.Y(_03133_),
    .A(_02886_),
    .B(_03132_));
 sg13g2_or3_1 _11157_ (.A(_02444_),
    .B(_03128_),
    .C(_03133_),
    .X(_03134_));
 sg13g2_a22oi_1 _11158_ (.Y(_03135_),
    .B1(_02150_),
    .B2(net189),
    .A2(net1557),
    .A1(net2115));
 sg13g2_or2_1 _11159_ (.X(_03136_),
    .B(_03135_),
    .A(_02148_));
 sg13g2_o21ai_1 _11160_ (.B1(_03136_),
    .Y(_03137_),
    .A1(net185),
    .A2(_02151_));
 sg13g2_nor2b_1 _11161_ (.A(_02150_),
    .B_N(_02878_),
    .Y(_03138_));
 sg13g2_nor3_1 _11162_ (.A(net192),
    .B(net188),
    .C(_02152_),
    .Y(_03139_));
 sg13g2_or2_1 _11163_ (.X(_03140_),
    .B(_03139_),
    .A(_03138_));
 sg13g2_a22oi_1 _11164_ (.Y(_03141_),
    .B1(_03140_),
    .B2(_02155_),
    .A2(_03137_),
    .A1(_02145_));
 sg13g2_nor3_1 _11165_ (.A(net185),
    .B(_02186_),
    .C(_02240_),
    .Y(_03142_));
 sg13g2_nor3_1 _11166_ (.A(net175),
    .B(_02212_),
    .C(_02224_),
    .Y(_03143_));
 sg13g2_nor2_1 _11167_ (.A(_03142_),
    .B(_03143_),
    .Y(_03144_));
 sg13g2_nor2b_1 _11168_ (.A(_02886_),
    .B_N(_03144_),
    .Y(_03145_));
 sg13g2_or3_1 _11169_ (.A(_02880_),
    .B(_03141_),
    .C(_03145_),
    .X(_03146_));
 sg13g2_nand2b_1 _11170_ (.Y(_03147_),
    .B(_02888_),
    .A_N(_03132_));
 sg13g2_nand2_1 _11171_ (.Y(_03148_),
    .A(_03141_),
    .B(_03144_));
 sg13g2_a21o_1 _11172_ (.A2(_03148_),
    .A1(_03147_),
    .B1(_02886_),
    .X(_03149_));
 sg13g2_and2_1 _11173_ (.A(_03141_),
    .B(_03144_),
    .X(_03150_));
 sg13g2_a22oi_1 _11174_ (.Y(_03151_),
    .B1(_03150_),
    .B2(_02880_),
    .A2(_03147_),
    .A1(_02886_));
 sg13g2_nand4_1 _11175_ (.B(_03146_),
    .C(_03149_),
    .A(_02444_),
    .Y(_03152_),
    .D(_03151_));
 sg13g2_a21oi_1 _11176_ (.A1(_02440_),
    .A2(_02391_),
    .Y(_03153_),
    .B1(_03112_));
 sg13g2_o21ai_1 _11177_ (.B1(_03153_),
    .Y(_03154_),
    .A1(_03111_),
    .A2(_03120_));
 sg13g2_o21ai_1 _11178_ (.B1(_03154_),
    .Y(_03155_),
    .A1(_02440_),
    .A2(_02391_));
 sg13g2_mux2_2 _11179_ (.A0(_02444_),
    .A1(_03155_),
    .S(_02889_),
    .X(data_addr_o_7_));
 sg13g2_a21oi_2 _11180_ (.B1(data_addr_o_7_),
    .Y(_03156_),
    .A2(_03152_),
    .A1(_03134_));
 sg13g2_nand4_1 _11181_ (.B(_03006_),
    .C(_03124_),
    .A(_02995_),
    .Y(_03157_),
    .D(_03156_));
 sg13g2_a22oi_1 _11182_ (.Y(_03158_),
    .B1(_02992_),
    .B2(_02994_),
    .A2(_02731_),
    .A1(_02703_));
 sg13g2_nor2_1 _11183_ (.A(_02914_),
    .B(_02975_),
    .Y(_03159_));
 sg13g2_a21o_1 _11184_ (.A2(_02556_),
    .A1(_02538_),
    .B1(_02984_),
    .X(_03160_));
 sg13g2_o21ai_1 _11185_ (.B1(_03031_),
    .Y(_03161_),
    .A1(_02980_),
    .A2(_03032_));
 sg13g2_o21ai_1 _11186_ (.B1(_03161_),
    .Y(_03162_),
    .A1(_02913_),
    .A2(_03160_));
 sg13g2_nand2b_1 _11187_ (.Y(_03163_),
    .B(_02599_),
    .A_N(_03162_));
 sg13g2_o21ai_1 _11188_ (.B1(_03163_),
    .Y(_03164_),
    .A1(_03158_),
    .A2(_03159_));
 sg13g2_nor3_1 _11189_ (.A(_02991_),
    .B(_03157_),
    .C(_03164_),
    .Y(_03165_));
 sg13g2_nand4_1 _11190_ (.B(_02931_),
    .C(_02971_),
    .A(_02895_),
    .Y(_03166_),
    .D(_03165_));
 sg13g2_xnor2_1 _11191_ (.Y(_03167_),
    .A(net190),
    .B(_02644_));
 sg13g2_o21ai_1 _11192_ (.B1(_02633_),
    .Y(_03168_),
    .A1(net177),
    .A2(net1397));
 sg13g2_xnor2_1 _11193_ (.Y(_03169_),
    .A(_02628_),
    .B(_03168_));
 sg13g2_nand2_1 _11194_ (.Y(_03170_),
    .A(net358),
    .B(_03169_));
 sg13g2_o21ai_1 _11195_ (.B1(_03170_),
    .Y(_03171_),
    .A1(net353),
    .A2(_03167_));
 sg13g2_o21ai_1 _11196_ (.B1(_02738_),
    .Y(_03172_),
    .A1(net177),
    .A2(_02741_));
 sg13g2_mux2_1 _11197_ (.A0(_02761_),
    .A1(_03172_),
    .S(_02925_),
    .X(_03173_));
 sg13g2_xnor2_1 _11198_ (.Y(_03174_),
    .A(_03171_),
    .B(_03173_));
 sg13g2_and3_1 _11199_ (.X(_03175_),
    .A(_02052_),
    .B(_02069_),
    .C(_02771_));
 sg13g2_nand2b_1 _11200_ (.Y(_03176_),
    .B(_02937_),
    .A_N(_01998_));
 sg13g2_o21ai_1 _11201_ (.B1(_01999_),
    .Y(_03177_),
    .A1(_03175_),
    .A2(_03176_));
 sg13g2_xnor2_1 _11202_ (.Y(_03178_),
    .A(net190),
    .B(_02006_));
 sg13g2_nand2_1 _11203_ (.Y(_03179_),
    .A(net182),
    .B(_02014_));
 sg13g2_nand2_1 _11204_ (.Y(_03180_),
    .A(net189),
    .B(_02020_));
 sg13g2_a22oi_1 _11205_ (.Y(_03181_),
    .B1(_03179_),
    .B2(_03180_),
    .A2(_03178_),
    .A1(net361));
 sg13g2_xor2_1 _11206_ (.B(_03181_),
    .A(_03177_),
    .X(_03182_));
 sg13g2_nand2_1 _11207_ (.Y(_03183_),
    .A(_03174_),
    .B(_03182_));
 sg13g2_or4_2 _11208_ (.A(data_addr_o_30_),
    .B(data_addr_o_27_),
    .C(_03166_),
    .D(_03183_),
    .X(_03184_));
 sg13g2_buf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sg13g2_mux2_1 _11210_ (.A0(_02861_),
    .A1(_02867_),
    .S(_03184_),
    .X(_03186_));
 sg13g2_a21oi_1 _11211_ (.A1(_02858_),
    .A2(_02857_),
    .Y(_03187_),
    .B1(_01629_));
 sg13g2_o21ai_1 _11212_ (.B1(_01623_),
    .Y(_03188_),
    .A1(_01434_),
    .A2(_03187_));
 sg13g2_nor2b_2 _11213_ (.A(_01746_),
    .B_N(_01721_),
    .Y(_03189_));
 sg13g2_nor2_1 _11214_ (.A(_01434_),
    .B(_02863_),
    .Y(\id_stage_i.perf_branch_o ));
 sg13g2_nand3_1 _11215_ (.B(_03184_),
    .C(\id_stage_i.perf_branch_o ),
    .A(_03189_),
    .Y(_03190_));
 sg13g2_nand2_1 _11216_ (.Y(_03191_),
    .A(_01751_),
    .B(\id_stage_i.perf_branch_o ));
 sg13g2_or2_1 _11217_ (.X(_03192_),
    .B(_03191_),
    .A(_03184_));
 sg13g2_nand3b_1 _11218_ (.B(_03190_),
    .C(_03192_),
    .Y(_03193_),
    .A_N(_03188_));
 sg13g2_or2_1 _11219_ (.X(_03194_),
    .B(_03193_),
    .A(_03186_));
 sg13g2_or2_2 _11220_ (.X(_03195_),
    .B(_03194_),
    .A(_01580_));
 sg13g2_nor2_2 _11221_ (.A(_01519_),
    .B(_03195_),
    .Y(_03196_));
 sg13g2_buf_2 fanout1102 (.A(net1103),
    .X(net1102));
 sg13g2_buf_1 fanout1101 (.A(\cs_registers_i/_0640_ ),
    .X(net1101));
 sg13g2_buf_2 fanout1100 (.A(\cs_registers_i/_0640_ ),
    .X(net1100));
 sg13g2_mux2_1 _11225_ (.A0(crash_dump_o_100_),
    .A1(crash_dump_o_68_),
    .S(net771),
    .X(_00000_));
 sg13g2_mux2_1 _11226_ (.A0(crash_dump_o_101_),
    .A1(crash_dump_o_69_),
    .S(net771),
    .X(_00001_));
 sg13g2_mux2_1 _11227_ (.A0(crash_dump_o_102_),
    .A1(crash_dump_o_70_),
    .S(net771),
    .X(_00002_));
 sg13g2_mux2_1 _11228_ (.A0(crash_dump_o_103_),
    .A1(crash_dump_o_71_),
    .S(net771),
    .X(_00003_));
 sg13g2_inv_2 _11229_ (.Y(_03200_),
    .A(crash_dump_o_104_));
 sg13g2_buf_2 fanout1099 (.A(_03368_),
    .X(net1099));
 sg13g2_buf_2 fanout1098 (.A(\cs_registers_i/_0715_ ),
    .X(net1098));
 sg13g2_buf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sg13g2_nand2_2 _11233_ (.Y(_03204_),
    .A(crash_dump_o_72_),
    .B(net779));
 sg13g2_o21ai_1 _11234_ (.B1(_03204_),
    .Y(_00004_),
    .A1(_03200_),
    .A2(net779));
 sg13g2_mux2_1 _11235_ (.A0(crash_dump_o_105_),
    .A1(crash_dump_o_73_),
    .S(net771),
    .X(_00005_));
 sg13g2_mux2_1 _11236_ (.A0(crash_dump_o_106_),
    .A1(crash_dump_o_74_),
    .S(net771),
    .X(_00006_));
 sg13g2_nand2_2 _11237_ (.Y(_03205_),
    .A(crash_dump_o_75_),
    .B(net770));
 sg13g2_o21ai_1 _11238_ (.B1(_03205_),
    .Y(_00007_),
    .A1(_01212_),
    .A2(net770));
 sg13g2_mux2_1 _11239_ (.A0(crash_dump_o_108_),
    .A1(crash_dump_o_76_),
    .S(net772),
    .X(_00008_));
 sg13g2_buf_2 fanout1096 (.A(\cs_registers_i/_0715_ ),
    .X(net1096));
 sg13g2_mux2_1 _11241_ (.A0(crash_dump_o_109_),
    .A1(crash_dump_o_77_),
    .S(net771),
    .X(_00009_));
 sg13g2_inv_2 _11242_ (.Y(_03207_),
    .A(crash_dump_o_110_));
 sg13g2_nand2_2 _11243_ (.Y(_03208_),
    .A(crash_dump_o_78_),
    .B(net779));
 sg13g2_o21ai_1 _11244_ (.B1(_03208_),
    .Y(_00010_),
    .A1(_03207_),
    .A2(net779));
 sg13g2_buf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sg13g2_nand2_2 _11246_ (.Y(_03210_),
    .A(crash_dump_o_79_),
    .B(net770));
 sg13g2_o21ai_1 _11247_ (.B1(_03210_),
    .Y(_00011_),
    .A1(_01226_),
    .A2(net770));
 sg13g2_mux2_1 _11248_ (.A0(crash_dump_o_112_),
    .A1(crash_dump_o_80_),
    .S(net772),
    .X(_00012_));
 sg13g2_mux2_1 _11249_ (.A0(crash_dump_o_113_),
    .A1(crash_dump_o_81_),
    .S(net773),
    .X(_00013_));
 sg13g2_nand2_2 _11250_ (.Y(_03211_),
    .A(crash_dump_o_82_),
    .B(net773));
 sg13g2_o21ai_1 _11251_ (.B1(_03211_),
    .Y(_00014_),
    .A1(_01240_),
    .A2(net773));
 sg13g2_mux2_1 _11252_ (.A0(crash_dump_o_115_),
    .A1(crash_dump_o_83_),
    .S(net773),
    .X(_00015_));
 sg13g2_mux2_1 _11253_ (.A0(crash_dump_o_116_),
    .A1(crash_dump_o_84_),
    .S(net774),
    .X(_00016_));
 sg13g2_nand2_2 _11254_ (.Y(_03212_),
    .A(crash_dump_o_85_),
    .B(net779));
 sg13g2_o21ai_1 _11255_ (.B1(_03212_),
    .Y(_00017_),
    .A1(_01255_),
    .A2(net779));
 sg13g2_mux2_1 _11256_ (.A0(crash_dump_o_118_),
    .A1(crash_dump_o_86_),
    .S(net777),
    .X(_00018_));
 sg13g2_mux2_1 _11257_ (.A0(crash_dump_o_119_),
    .A1(crash_dump_o_87_),
    .S(net772),
    .X(_00019_));
 sg13g2_mux2_1 _11258_ (.A0(crash_dump_o_120_),
    .A1(crash_dump_o_88_),
    .S(net772),
    .X(_00020_));
 sg13g2_mux2_1 _11259_ (.A0(crash_dump_o_121_),
    .A1(crash_dump_o_89_),
    .S(net772),
    .X(_00021_));
 sg13g2_mux2_1 _11260_ (.A0(crash_dump_o_122_),
    .A1(crash_dump_o_90_),
    .S(net773),
    .X(_00022_));
 sg13g2_buf_2 fanout1094 (.A(\cs_registers_i/_0814_ ),
    .X(net1094));
 sg13g2_mux2_1 _11262_ (.A0(crash_dump_o_123_),
    .A1(crash_dump_o_91_),
    .S(net773),
    .X(_00023_));
 sg13g2_nand2_2 _11263_ (.Y(_03214_),
    .A(crash_dump_o_92_),
    .B(net779));
 sg13g2_o21ai_1 _11264_ (.B1(_03214_),
    .Y(_00024_),
    .A1(_01284_),
    .A2(net779));
 sg13g2_mux2_1 _11265_ (.A0(crash_dump_o_125_),
    .A1(crash_dump_o_93_),
    .S(net774),
    .X(_00025_));
 sg13g2_mux2_1 _11266_ (.A0(crash_dump_o_126_),
    .A1(crash_dump_o_94_),
    .S(net774),
    .X(_00026_));
 sg13g2_mux2_1 _11267_ (.A0(crash_dump_o_127_),
    .A1(crash_dump_o_95_),
    .S(net774),
    .X(_00027_));
 sg13g2_buf_2 fanout1093 (.A(\cs_registers_i/_0596_ ),
    .X(net1093));
 sg13g2_inv_1 _11269_ (.Y(_03216_),
    .A(_01566_));
 sg13g2_nor3_2 _11270_ (.A(_01190_),
    .B(_01434_),
    .C(_03216_),
    .Y(_03217_));
 sg13g2_and2_1 _11271_ (.A(_01495_),
    .B(_03217_),
    .X(_03218_));
 sg13g2_nor2_2 _11272_ (.A(net1977),
    .B(_01141_),
    .Y(_03219_));
 sg13g2_or2_1 _11273_ (.X(_03220_),
    .B(\load_store_unit_i.ls_fsm_cs_0__$_NOT__A_Y ),
    .A(\load_store_unit_i.ls_fsm_cs_2_ ));
 sg13g2_a21oi_1 _11274_ (.A1(\load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ),
    .A2(\load_store_unit_i.ls_fsm_cs_1_ ),
    .Y(_03221_),
    .B1(_03220_));
 sg13g2_nor2_2 _11275_ (.A(_03219_),
    .B(_03221_),
    .Y(_03222_));
 sg13g2_nor2_1 _11276_ (.A(_01771_),
    .B(_01495_),
    .Y(_03223_));
 sg13g2_inv_1 _11277_ (.Y(_03224_),
    .A(data_gnt_i));
 sg13g2_nand2b_1 _11278_ (.Y(_03225_),
    .B(_03219_),
    .A_N(net1976));
 sg13g2_o21ai_1 _11279_ (.B1(_01144_),
    .Y(_03226_),
    .A1(_03224_),
    .A2(_03225_));
 sg13g2_nor2b_1 _11280_ (.A(data_err_i),
    .B_N(net2466),
    .Y(_03227_));
 sg13g2_inv_1 _11281_ (.Y(_03228_),
    .A(\load_store_unit_i.lsu_err_q_$_NOT__A_Y ));
 sg13g2_o21ai_1 _11282_ (.B1(\load_store_unit_i.ls_fsm_cs_1_ ),
    .Y(_03229_),
    .A1(\load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ),
    .A2(_03228_));
 sg13g2_nor2_1 _11283_ (.A(net1976),
    .B(data_gnt_i),
    .Y(_03230_));
 sg13g2_nor2_1 _11284_ (.A(_03230_),
    .B(_03220_),
    .Y(_03231_));
 sg13g2_a22oi_1 _11285_ (.Y(_03232_),
    .B1(_03229_),
    .B2(_03231_),
    .A2(_03227_),
    .A1(_03226_));
 sg13g2_a21oi_1 _11286_ (.A1(_03222_),
    .A2(_03223_),
    .Y(_03233_),
    .B1(_03232_));
 sg13g2_a21oi_2 _11287_ (.B1(_03233_),
    .Y(_03234_),
    .A2(_03218_),
    .A1(data_gnt_i));
 sg13g2_buf_1 fanout1092 (.A(net1093),
    .X(net1092));
 sg13g2_buf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sg13g2_buf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_nor3_1 _11291_ (.A(net1718),
    .B(net1147),
    .C(net86),
    .Y(_03238_));
 sg13g2_a21o_1 _11292_ (.A2(_03234_),
    .A1(crash_dump_o_32_),
    .B1(_03238_),
    .X(_00028_));
 sg13g2_inv_2 _11293_ (.Y(_03239_),
    .A(net1113));
 sg13g2_nor3_1 _11294_ (.A(net1718),
    .B(_03239_),
    .C(net86),
    .Y(_03240_));
 sg13g2_a21o_1 _11295_ (.A2(net86),
    .A1(crash_dump_o_33_),
    .B1(_03240_),
    .X(_00029_));
 sg13g2_mux2_1 _11296_ (.A0(data_addr_o_2_),
    .A1(crash_dump_o_34_),
    .S(net83),
    .X(_00030_));
 sg13g2_mux2_1 _11297_ (.A0(net2490),
    .A1(crash_dump_o_35_),
    .S(net83),
    .X(_00031_));
 sg13g2_buf_2 fanout1089 (.A(net1091),
    .X(net1089));
 sg13g2_mux2_1 _11299_ (.A0(data_addr_o_4_),
    .A1(crash_dump_o_36_),
    .S(net84),
    .X(_00032_));
 sg13g2_nand2_1 _11300_ (.Y(_03242_),
    .A(net181),
    .B(_03008_));
 sg13g2_o21ai_1 _11301_ (.B1(_03242_),
    .Y(_03243_),
    .A1(net175),
    .A2(_03013_));
 sg13g2_inv_4 _11302_ (.A(_02287_),
    .Y(_03244_));
 sg13g2_nor2_1 _11303_ (.A(net184),
    .B(_02291_),
    .Y(_03245_));
 sg13g2_a21oi_1 _11304_ (.A1(net188),
    .A2(_03244_),
    .Y(_03246_),
    .B1(_03245_));
 sg13g2_nand2_1 _11305_ (.Y(_03247_),
    .A(_02278_),
    .B(_03246_));
 sg13g2_nand2_1 _11306_ (.Y(_03248_),
    .A(_02282_),
    .B(_03247_));
 sg13g2_nor2_1 _11307_ (.A(_02282_),
    .B(_03247_),
    .Y(_03249_));
 sg13g2_a21oi_1 _11308_ (.A1(_03243_),
    .A2(_03248_),
    .Y(_03250_),
    .B1(_03249_));
 sg13g2_o21ai_1 _11309_ (.B1(_02272_),
    .Y(_03251_),
    .A1(_02363_),
    .A2(_03250_));
 sg13g2_xor2_1 _11310_ (.B(_03251_),
    .A(_03111_),
    .X(data_addr_o_5_));
 sg13g2_mux2_1 _11311_ (.A0(data_addr_o_5_),
    .A1(crash_dump_o_37_),
    .S(net84),
    .X(_00033_));
 sg13g2_a22oi_1 _11312_ (.Y(_03252_),
    .B1(_03081_),
    .B2(_02368_),
    .A2(_03120_),
    .A1(_02380_));
 sg13g2_xnor2_1 _11313_ (.Y(data_addr_o_6_),
    .A(_03079_),
    .B(_03252_));
 sg13g2_mux2_1 _11314_ (.A0(data_addr_o_6_),
    .A1(crash_dump_o_38_),
    .S(net84),
    .X(_00034_));
 sg13g2_mux2_1 _11315_ (.A0(data_addr_o_7_),
    .A1(crash_dump_o_39_),
    .S(net84),
    .X(_00035_));
 sg13g2_nor2_2 _11316_ (.A(_02890_),
    .B(_03132_),
    .Y(_03253_));
 sg13g2_xor2_1 _11317_ (.B(_03253_),
    .A(_02886_),
    .X(data_addr_o_8_));
 sg13g2_mux2_1 _11318_ (.A0(data_addr_o_8_),
    .A1(crash_dump_o_40_),
    .S(net84),
    .X(_00036_));
 sg13g2_nor2_1 _11319_ (.A(_02444_),
    .B(_03128_),
    .Y(_03254_));
 sg13g2_nand2b_1 _11320_ (.Y(_03255_),
    .B(_02886_),
    .A_N(_02880_));
 sg13g2_nand3_1 _11321_ (.B(_03144_),
    .C(_03255_),
    .A(_03141_),
    .Y(_03256_));
 sg13g2_nand3_1 _11322_ (.B(_03146_),
    .C(_03256_),
    .A(_02444_),
    .Y(_03257_));
 sg13g2_nor2b_2 _11323_ (.A(_03254_),
    .B_N(_03257_),
    .Y(data_addr_o_9_));
 sg13g2_mux2_1 _11324_ (.A0(data_addr_o_9_),
    .A1(crash_dump_o_41_),
    .S(net84),
    .X(_00037_));
 sg13g2_inv_16 _11325_ (.A(_02895_),
    .Y(data_addr_o_10_));
 sg13g2_mux2_1 _11326_ (.A0(data_addr_o_10_),
    .A1(crash_dump_o_42_),
    .S(net84),
    .X(_00038_));
 sg13g2_xor2_1 _11327_ (.B(_03004_),
    .A(_02445_),
    .X(data_addr_o_11_));
 sg13g2_mux2_1 _11328_ (.A0(data_addr_o_11_),
    .A1(crash_dump_o_43_),
    .S(net83),
    .X(_00039_));
 sg13g2_nand2_1 _11329_ (.Y(_03258_),
    .A(_02503_),
    .B(_03000_));
 sg13g2_nor2_1 _11330_ (.A(_02503_),
    .B(_03000_),
    .Y(_03259_));
 sg13g2_a21oi_2 _11331_ (.B1(_03259_),
    .Y(_03260_),
    .A2(_03258_),
    .A1(_02445_));
 sg13g2_xnor2_1 _11332_ (.Y(data_addr_o_12_),
    .A(_02608_),
    .B(_03260_));
 sg13g2_mux2_1 _11333_ (.A0(data_addr_o_12_),
    .A1(crash_dump_o_44_),
    .S(net83),
    .X(_00040_));
 sg13g2_or2_1 _11334_ (.X(_03261_),
    .B(_02908_),
    .A(_02445_));
 sg13g2_and2_2 _11335_ (.A(_02508_),
    .B(_03261_),
    .X(_03262_));
 sg13g2_xor2_1 _11336_ (.B(_03262_),
    .A(_02453_),
    .X(data_addr_o_13_));
 sg13g2_mux2_1 _11337_ (.A0(data_addr_o_13_),
    .A1(crash_dump_o_45_),
    .S(net83),
    .X(_00041_));
 sg13g2_nor2_1 _11338_ (.A(_02453_),
    .B(_03262_),
    .Y(_03263_));
 sg13g2_nor2_1 _11339_ (.A(_03038_),
    .B(_03263_),
    .Y(_03264_));
 sg13g2_xnor2_1 _11340_ (.Y(_03265_),
    .A(_02465_),
    .B(_03264_));
 sg13g2_inv_16 _11341_ (.A(_03265_),
    .Y(data_addr_o_14_));
 sg13g2_buf_2 fanout1088 (.A(net1092),
    .X(net1088));
 sg13g2_mux2_1 _11343_ (.A0(data_addr_o_14_),
    .A1(crash_dump_o_46_),
    .S(net86),
    .X(_00042_));
 sg13g2_xnor2_1 _11344_ (.Y(data_addr_o_15_),
    .A(_02536_),
    .B(_02913_));
 sg13g2_mux2_1 _11345_ (.A0(data_addr_o_15_),
    .A1(crash_dump_o_47_),
    .S(net85),
    .X(_00043_));
 sg13g2_o21ai_1 _11346_ (.B1(_02974_),
    .Y(_03267_),
    .A1(_02913_),
    .A2(_02984_));
 sg13g2_xnor2_1 _11347_ (.Y(data_addr_o_16_),
    .A(_02557_),
    .B(_03267_));
 sg13g2_mux2_1 _11348_ (.A0(data_addr_o_16_),
    .A1(crash_dump_o_48_),
    .S(net85),
    .X(_00044_));
 sg13g2_xnor2_1 _11349_ (.Y(data_addr_o_17_),
    .A(_02598_),
    .B(_03162_));
 sg13g2_mux2_1 _11350_ (.A0(data_addr_o_17_),
    .A1(crash_dump_o_49_),
    .S(net85),
    .X(_00045_));
 sg13g2_inv_1 _11351_ (.Y(_03268_),
    .A(_02712_));
 sg13g2_a21oi_1 _11352_ (.A1(_02981_),
    .A2(_03162_),
    .Y(_03269_),
    .B1(_03268_));
 sg13g2_xor2_1 _11353_ (.B(_03269_),
    .A(_02575_),
    .X(data_addr_o_18_));
 sg13g2_mux2_1 _11354_ (.A0(data_addr_o_18_),
    .A1(crash_dump_o_50_),
    .S(net85),
    .X(_00046_));
 sg13g2_and2_1 _11355_ (.A(_02731_),
    .B(_02914_),
    .X(_03270_));
 sg13g2_xnor2_1 _11356_ (.Y(data_addr_o_19_),
    .A(_02703_),
    .B(_03270_));
 sg13g2_mux2_1 _11357_ (.A0(data_addr_o_19_),
    .A1(crash_dump_o_51_),
    .S(net85),
    .X(_00047_));
 sg13g2_inv_1 _11358_ (.Y(_03271_),
    .A(_03270_));
 sg13g2_nor2_1 _11359_ (.A(net186),
    .B(_02748_),
    .Y(_03272_));
 sg13g2_a221oi_1 _11360_ (.B2(_03271_),
    .C1(_03272_),
    .B1(_03086_),
    .A1(net189),
    .Y(_03273_),
    .A2(_02753_));
 sg13g2_xnor2_1 _11361_ (.Y(_03274_),
    .A(_03083_),
    .B(_03273_));
 sg13g2_inv_16 _11362_ (.A(_03274_),
    .Y(data_addr_o_20_));
 sg13g2_nand2_1 _11363_ (.Y(_03275_),
    .A(crash_dump_o_52_),
    .B(net83));
 sg13g2_o21ai_1 _11364_ (.B1(_03275_),
    .Y(_00048_),
    .A1(net83),
    .A2(_03274_));
 sg13g2_nand2_1 _11365_ (.Y(_03276_),
    .A(crash_dump_o_53_),
    .B(net83));
 sg13g2_o21ai_1 _11366_ (.B1(_03276_),
    .Y(_00049_),
    .A1(_02931_),
    .A2(net82));
 sg13g2_inv_16 _11367_ (.A(_03174_),
    .Y(data_addr_o_22_));
 sg13g2_nand2_1 _11368_ (.Y(_03277_),
    .A(crash_dump_o_54_),
    .B(net82));
 sg13g2_o21ai_1 _11369_ (.B1(_03277_),
    .Y(_00050_),
    .A1(_03174_),
    .A2(net82));
 sg13g2_xnor2_1 _11370_ (.Y(_03278_),
    .A(_02052_),
    .B(_02771_));
 sg13g2_inv_16 _11371_ (.A(_03278_),
    .Y(data_addr_o_23_));
 sg13g2_mux2_1 _11372_ (.A0(data_addr_o_23_),
    .A1(crash_dump_o_55_),
    .S(net85),
    .X(_00051_));
 sg13g2_a21oi_1 _11373_ (.A1(_02052_),
    .A2(_02771_),
    .Y(_03279_),
    .B1(_02943_));
 sg13g2_xnor2_1 _11374_ (.Y(data_addr_o_24_),
    .A(_02069_),
    .B(_03279_));
 sg13g2_mux2_1 _11375_ (.A0(data_addr_o_24_),
    .A1(crash_dump_o_56_),
    .S(net85),
    .X(_00052_));
 sg13g2_inv_1 _11376_ (.Y(_03280_),
    .A(_02968_));
 sg13g2_mux2_2 _11377_ (.A0(_02938_),
    .A1(_03280_),
    .S(_02771_),
    .X(data_addr_o_25_));
 sg13g2_mux2_1 _11378_ (.A0(data_addr_o_25_),
    .A1(crash_dump_o_57_),
    .S(net85),
    .X(_00053_));
 sg13g2_inv_16 _11379_ (.A(_03182_),
    .Y(data_addr_o_26_));
 sg13g2_mux2_1 _11380_ (.A0(data_addr_o_26_),
    .A1(crash_dump_o_58_),
    .S(net84),
    .X(_00054_));
 sg13g2_mux2_1 _11381_ (.A0(data_addr_o_27_),
    .A1(crash_dump_o_59_),
    .S(net82),
    .X(_00055_));
 sg13g2_nor2_1 _11382_ (.A(_02868_),
    .B(_02950_),
    .Y(_03281_));
 sg13g2_a21oi_2 _11383_ (.B1(_03281_),
    .Y(data_addr_o_28_),
    .A2(_02935_),
    .A1(_02868_));
 sg13g2_mux2_1 _11384_ (.A0(data_addr_o_28_),
    .A1(crash_dump_o_60_),
    .S(net82),
    .X(_00056_));
 sg13g2_o21ai_1 _11385_ (.B1(_03025_),
    .Y(_03282_),
    .A1(_01951_),
    .A2(_02868_));
 sg13g2_xnor2_1 _11386_ (.Y(data_addr_o_29_),
    .A(_01978_),
    .B(_03282_));
 sg13g2_mux2_1 _11387_ (.A0(data_addr_o_29_),
    .A1(crash_dump_o_61_),
    .S(net82),
    .X(_00057_));
 sg13g2_mux2_1 _11388_ (.A0(net2494),
    .A1(crash_dump_o_62_),
    .S(net82),
    .X(_00058_));
 sg13g2_buf_2 fanout1087 (.A(\cs_registers_i/_1178_ ),
    .X(net1087));
 sg13g2_mux2_1 _11390_ (.A0(net37),
    .A1(crash_dump_o_63_),
    .S(net82),
    .X(_00059_));
 sg13g2_nand2_2 _11391_ (.Y(_03283_),
    .A(_01438_),
    .B(_01468_));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_1 fanout1085 (.A(net1086),
    .X(net1085));
 sg13g2_buf_2 fanout1084 (.A(net1085),
    .X(net1084));
 sg13g2_buf_1 fanout1083 (.A(net1085),
    .X(net1083));
 sg13g2_buf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sg13g2_buf_2 fanout1081 (.A(_05797_),
    .X(net1081));
 sg13g2_nand2b_1 _11398_ (.Y(_03290_),
    .B(net768),
    .A_N(_01517_));
 sg13g2_nand2_1 _11399_ (.Y(_03291_),
    .A(instr_rdata_i_0_),
    .B(instr_rdata_i_1_));
 sg13g2_nand3_1 _11400_ (.B(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0_ ),
    .C(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1_ ),
    .A(net1983),
    .Y(_03292_));
 sg13g2_o21ai_1 _11401_ (.B1(_03292_),
    .Y(_03293_),
    .A1(net1983),
    .A2(_03291_));
 sg13g2_or3_2 _11402_ (.A(net557),
    .B(_01514_),
    .C(_03293_),
    .X(_03294_));
 sg13g2_inv_4 _11403_ (.A(_03294_),
    .Y(_03295_));
 sg13g2_a22oi_1 _11404_ (.Y(_03296_),
    .B1(_03295_),
    .B2(net768),
    .A2(_03290_),
    .A1(net561));
 sg13g2_buf_2 fanout1080 (.A(_06765_),
    .X(net1080));
 sg13g2_o21ai_1 _11406_ (.B1(_01631_),
    .Y(_03298_),
    .A1(net2102),
    .A2(_01467_));
 sg13g2_nor3_1 _11407_ (.A(_01464_),
    .B(net1715),
    .C(_03298_),
    .Y(_03299_));
 sg13g2_buf_2 fanout1079 (.A(\cs_registers_i/_1455_ ),
    .X(net1079));
 sg13g2_buf_1 fanout1078 (.A(net1079),
    .X(net1078));
 sg13g2_buf_2 fanout1077 (.A(net1078),
    .X(net1077));
 sg13g2_nand2_1 _11411_ (.Y(_03303_),
    .A(net1113),
    .B(net1556));
 sg13g2_nand2_2 _11412_ (.Y(_03304_),
    .A(_01401_),
    .B(_01581_));
 sg13g2_nand2_2 _11413_ (.Y(_03305_),
    .A(_01443_),
    .B(net395));
 sg13g2_nor4_1 _11414_ (.A(net1904),
    .B(_03298_),
    .C(_03304_),
    .D(_03305_),
    .Y(_03306_));
 sg13g2_buf_2 fanout1076 (.A(_06724_),
    .X(net1076));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(_08551_));
 sg13g2_buf_1 fanout1074 (.A(_08551_),
    .X(net1074));
 sg13g2_nor2_2 _11418_ (.A(_01443_),
    .B(_01463_),
    .Y(_03310_));
 sg13g2_a21oi_1 _11419_ (.A1(_01463_),
    .A2(_03298_),
    .Y(_03311_),
    .B1(_03310_));
 sg13g2_nor3_1 _11420_ (.A(_01591_),
    .B(_01584_),
    .C(_03305_),
    .Y(csr_restore_mret_id));
 sg13g2_nor2_1 _11421_ (.A(net1715),
    .B(_01487_),
    .Y(_03312_));
 sg13g2_o21ai_1 _11422_ (.B1(_03304_),
    .Y(_03313_),
    .A1(net344),
    .A2(_03312_));
 sg13g2_o21ai_1 _11423_ (.B1(_03313_),
    .Y(_03314_),
    .A1(net1715),
    .A2(_03311_));
 sg13g2_buf_1 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_2 fanout1072 (.A(net1073),
    .X(net1072));
 sg13g2_buf_2 fanout1071 (.A(\cs_registers_i/_0698_ ),
    .X(net1071));
 sg13g2_a22oi_1 _11427_ (.Y(_03318_),
    .B1(net1489),
    .B2(crash_dump_o_1_),
    .A2(net1550),
    .A1(csr_depc_1_));
 sg13g2_inv_1 _11428_ (.Y(_03319_),
    .A(_01459_));
 sg13g2_a21oi_1 _11429_ (.A1(net395),
    .A2(_03319_),
    .Y(_03320_),
    .B1(_01487_));
 sg13g2_nor2_1 _11430_ (.A(_03310_),
    .B(_03320_),
    .Y(_03321_));
 sg13g2_nor2_2 _11431_ (.A(net1904),
    .B(_03321_),
    .Y(_03322_));
 sg13g2_or4_2 _11432_ (.A(net1555),
    .B(net1545),
    .C(net1456),
    .D(net1484),
    .X(_03323_));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(\cs_registers_i/_0698_ ));
 sg13g2_nand2_2 _11434_ (.Y(_03325_),
    .A(net106),
    .B(net235));
 sg13g2_a21o_1 _11435_ (.A2(_03318_),
    .A1(_03303_),
    .B1(_03325_),
    .X(_03326_));
 sg13g2_o21ai_1 _11436_ (.B1(_03326_),
    .Y(_00060_),
    .A1(net105),
    .A2(_03296_));
 sg13g2_nand2b_1 _11437_ (.Y(_03327_),
    .B(net395),
    .A_N(_01443_));
 sg13g2_nor2_1 _11438_ (.A(\id_stage_i.controller_i.store_err_q ),
    .B(\id_stage_i.controller_i.load_err_q ),
    .Y(_03328_));
 sg13g2_inv_1 _11439_ (.Y(_03329_),
    .A(net2101));
 sg13g2_nand2_1 _11440_ (.Y(_03330_),
    .A(net437),
    .B(\id_stage_i.controller_i.instr_fetch_err_i ));
 sg13g2_nand2_1 _11441_ (.Y(_03331_),
    .A(_03329_),
    .B(net1880));
 sg13g2_nor3_1 _11442_ (.A(_03328_),
    .B(_01592_),
    .C(_03331_),
    .Y(_03332_));
 sg13g2_nand2_1 _11443_ (.Y(_03333_),
    .A(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .B(net2116));
 sg13g2_nand3b_1 _11444_ (.B(_01448_),
    .C(net513),
    .Y(_03334_),
    .A_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ));
 sg13g2_o21ai_1 _11445_ (.B1(_03334_),
    .Y(_03335_),
    .A1(net464),
    .A2(_03333_));
 sg13g2_nand2_1 _11446_ (.Y(_03336_),
    .A(_01453_),
    .B(_03335_));
 sg13g2_a21oi_1 _11447_ (.A1(_03329_),
    .A2(_01419_),
    .Y(_03337_),
    .B1(_03336_));
 sg13g2_nor3_1 _11448_ (.A(net1903),
    .B(net328),
    .C(_03337_),
    .Y(_03338_));
 sg13g2_inv_1 _11449_ (.Y(_03339_),
    .A(exc_cause_6_));
 sg13g2_a21oi_2 _11450_ (.B1(_03339_),
    .Y(_03340_),
    .A2(irq_nm_i),
    .A1(\id_stage_i.controller_i.handle_irq_$_AND__Y_A_$_AND__Y_B ));
 sg13g2_inv_1 _11451_ (.Y(_03341_),
    .A(\id_stage_i.controller_i.irqs_i_2_ ));
 sg13g2_inv_1 _11452_ (.Y(_03342_),
    .A(\id_stage_i.controller_i.irqs_i_6_ ));
 sg13g2_inv_1 _11453_ (.Y(_03343_),
    .A(\id_stage_i.controller_i.irqs_i_10_ ));
 sg13g2_inv_1 _11454_ (.Y(_03344_),
    .A(\id_stage_i.controller_i.irqs_i_14_ ));
 sg13g2_a21oi_1 _11455_ (.A1(_03344_),
    .A2(\id_stage_i.controller_i.irqs_i_15_ ),
    .Y(_03345_),
    .B1(\id_stage_i.controller_i.irqs_i_13_ ));
 sg13g2_inv_1 _11456_ (.Y(_03346_),
    .A(\id_stage_i.controller_i.irqs_i_11_ ));
 sg13g2_o21ai_1 _11457_ (.B1(_03346_),
    .Y(_03347_),
    .A1(\id_stage_i.controller_i.irqs_i_12_ ),
    .A2(_03345_));
 sg13g2_a21oi_1 _11458_ (.A1(_03343_),
    .A2(_03347_),
    .Y(_03348_),
    .B1(\id_stage_i.controller_i.irqs_i_9_ ));
 sg13g2_inv_1 _11459_ (.Y(_03349_),
    .A(\id_stage_i.controller_i.irqs_i_7_ ));
 sg13g2_o21ai_1 _11460_ (.B1(_03349_),
    .Y(_03350_),
    .A1(\id_stage_i.controller_i.irqs_i_8_ ),
    .A2(_03348_));
 sg13g2_a21oi_1 _11461_ (.A1(_03342_),
    .A2(_03350_),
    .Y(_03351_),
    .B1(\id_stage_i.controller_i.irqs_i_5_ ));
 sg13g2_inv_1 _11462_ (.Y(_03352_),
    .A(\id_stage_i.controller_i.irqs_i_3_ ));
 sg13g2_o21ai_1 _11463_ (.B1(_03352_),
    .Y(_03353_),
    .A1(\id_stage_i.controller_i.irqs_i_4_ ),
    .A2(_03351_));
 sg13g2_a21oi_1 _11464_ (.A1(_03341_),
    .A2(_03353_),
    .Y(_03354_),
    .B1(\id_stage_i.controller_i.irqs_i_1_ ));
 sg13g2_nor4_2 _11465_ (.A(\id_stage_i.controller_i.irqs_i_4_ ),
    .B(\id_stage_i.controller_i.irqs_i_5_ ),
    .C(\id_stage_i.controller_i.irqs_i_6_ ),
    .Y(_03355_),
    .D(\id_stage_i.controller_i.irqs_i_7_ ));
 sg13g2_or2_1 _11466_ (.X(_03356_),
    .B(\id_stage_i.controller_i.irqs_i_1_ ),
    .A(\id_stage_i.controller_i.irqs_i_0_ ));
 sg13g2_nor3_1 _11467_ (.A(\id_stage_i.controller_i.irqs_i_2_ ),
    .B(\id_stage_i.controller_i.irqs_i_3_ ),
    .C(_03356_),
    .Y(_03357_));
 sg13g2_nor4_2 _11468_ (.A(\id_stage_i.controller_i.irqs_i_8_ ),
    .B(\id_stage_i.controller_i.irqs_i_9_ ),
    .C(\id_stage_i.controller_i.irqs_i_10_ ),
    .Y(_03358_),
    .D(\id_stage_i.controller_i.irqs_i_11_ ));
 sg13g2_nor4_2 _11469_ (.A(\id_stage_i.controller_i.irqs_i_14_ ),
    .B(\id_stage_i.controller_i.irqs_i_15_ ),
    .C(\id_stage_i.controller_i.irqs_i_12_ ),
    .Y(_03359_),
    .D(\id_stage_i.controller_i.irqs_i_13_ ));
 sg13g2_nand4_1 _11470_ (.B(_03357_),
    .C(_03358_),
    .A(_03355_),
    .Y(_03360_),
    .D(_03359_));
 sg13g2_o21ai_1 _11471_ (.B1(_03360_),
    .Y(_03361_),
    .A1(\id_stage_i.controller_i.irqs_i_0_ ),
    .A2(_03354_));
 sg13g2_nand2_2 _11472_ (.Y(_03362_),
    .A(_03340_),
    .B(_03361_));
 sg13g2_o21ai_1 _11473_ (.B1(_03362_),
    .Y(exc_cause_0_),
    .A1(net1645),
    .A2(_03338_));
 sg13g2_inv_1 _11474_ (.Y(_03363_),
    .A(exc_cause_0_));
 sg13g2_nand4_1 _11475_ (.B(_01631_),
    .C(net1645),
    .A(net1715),
    .Y(_03364_),
    .D(_03320_));
 sg13g2_a22oi_1 _11476_ (.Y(_03365_),
    .B1(net1484),
    .B2(crash_dump_o_2_),
    .A2(net1545),
    .A1(csr_depc_2_));
 sg13g2_o21ai_1 _11477_ (.B1(_03365_),
    .Y(_03366_),
    .A1(_03363_),
    .A2(_03364_));
 sg13g2_a21oi_2 _11478_ (.B1(_03366_),
    .Y(_03367_),
    .A2(net1551),
    .A1(data_addr_o_2_));
 sg13g2_or2_1 _11479_ (.X(_03368_),
    .B(_03367_),
    .A(_03325_));
 sg13g2_buf_2 fanout1069 (.A(\cs_registers_i/_0808_ ),
    .X(net1069));
 sg13g2_nand2_1 _11481_ (.Y(_03370_),
    .A(_03295_),
    .B(net1099));
 sg13g2_buf_4 fanout1068 (.X(net1068),
    .A(\cs_registers_i/_0808_ ));
 sg13g2_buf_4 fanout1067 (.X(net1067),
    .A(\cs_registers_i/_0932_ ));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(\cs_registers_i/_1100_ ));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(\cs_registers_i/_1304_ ));
 sg13g2_o21ai_1 _11486_ (.B1(net114),
    .Y(_03375_),
    .A1(_01519_),
    .A2(_03195_));
 sg13g2_a21oi_2 _11487_ (.B1(crash_dump_o_66_),
    .Y(_03376_),
    .A2(net2488),
    .A1(_03370_));
 sg13g2_buf_4 fanout1064 (.X(net1064),
    .A(\cs_registers_i/_1322_ ));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(\cs_registers_i/_1694_ ));
 sg13g2_and3_1 _11490_ (.X(_03379_),
    .A(crash_dump_o_66_),
    .B(net778),
    .C(_03294_));
 sg13g2_o21ai_1 _11491_ (.B1(net1099),
    .Y(_03380_),
    .A1(net106),
    .A2(_03379_));
 sg13g2_nor2b_1 _11492_ (.A(_03376_),
    .B_N(_03380_),
    .Y(_00061_));
 sg13g2_xnor2_1 _11493_ (.Y(_03381_),
    .A(crash_dump_o_67_),
    .B(_03379_));
 sg13g2_nor2_1 _11494_ (.A(_01592_),
    .B(_03331_),
    .Y(_03382_));
 sg13g2_inv_1 _11495_ (.Y(_03383_),
    .A(\id_stage_i.controller_i.load_err_q ));
 sg13g2_buf_2 fanout1062 (.A(_06861_),
    .X(net1062));
 sg13g2_nand2_1 _11497_ (.Y(_03385_),
    .A(net2100),
    .B(net1879));
 sg13g2_a22oi_1 _11498_ (.Y(_03386_),
    .B1(_03336_),
    .B2(_03385_),
    .A2(_03382_),
    .A1(_03383_));
 sg13g2_a21oi_1 _11499_ (.A1(\id_stage_i.controller_i.store_err_q ),
    .A2(_03382_),
    .Y(_03387_),
    .B1(_03386_));
 sg13g2_nor2_1 _11500_ (.A(\id_stage_i.controller_i.irqs_i_14_ ),
    .B(\id_stage_i.controller_i.irqs_i_15_ ),
    .Y(_03388_));
 sg13g2_nor3_1 _11501_ (.A(\id_stage_i.controller_i.irqs_i_12_ ),
    .B(\id_stage_i.controller_i.irqs_i_13_ ),
    .C(_03388_),
    .Y(_03389_));
 sg13g2_nor3_1 _11502_ (.A(\id_stage_i.controller_i.irqs_i_10_ ),
    .B(\id_stage_i.controller_i.irqs_i_11_ ),
    .C(_03389_),
    .Y(_03390_));
 sg13g2_nor3_1 _11503_ (.A(\id_stage_i.controller_i.irqs_i_8_ ),
    .B(\id_stage_i.controller_i.irqs_i_9_ ),
    .C(_03390_),
    .Y(_03391_));
 sg13g2_nor3_1 _11504_ (.A(\id_stage_i.controller_i.irqs_i_6_ ),
    .B(\id_stage_i.controller_i.irqs_i_7_ ),
    .C(_03391_),
    .Y(_03392_));
 sg13g2_nor3_1 _11505_ (.A(\id_stage_i.controller_i.irqs_i_4_ ),
    .B(\id_stage_i.controller_i.irqs_i_5_ ),
    .C(_03392_),
    .Y(_03393_));
 sg13g2_nor3_1 _11506_ (.A(\id_stage_i.controller_i.irqs_i_2_ ),
    .B(\id_stage_i.controller_i.irqs_i_3_ ),
    .C(_03393_),
    .Y(_03394_));
 sg13g2_o21ai_1 _11507_ (.B1(_03360_),
    .Y(_03395_),
    .A1(_03356_),
    .A2(_03394_));
 sg13g2_nand2_2 _11508_ (.Y(_03396_),
    .A(_03340_),
    .B(_03395_));
 sg13g2_o21ai_1 _11509_ (.B1(_03396_),
    .Y(exc_cause_1_),
    .A1(net1645),
    .A2(_03387_));
 sg13g2_a21oi_1 _11510_ (.A1(_01443_),
    .A2(_01631_),
    .Y(_03397_),
    .B1(_01463_));
 sg13g2_o21ai_1 _11511_ (.B1(_03305_),
    .Y(_03398_),
    .A1(net395),
    .A2(_01485_));
 sg13g2_nand2_1 _11512_ (.Y(_03399_),
    .A(_03320_),
    .B(_03398_));
 sg13g2_nand2_1 _11513_ (.Y(_03400_),
    .A(debug_mode),
    .B(_03310_));
 sg13g2_a21oi_1 _11514_ (.A1(_03399_),
    .A2(_03400_),
    .Y(_03401_),
    .B1(net1904));
 sg13g2_o21ai_1 _11515_ (.B1(_03401_),
    .Y(_03402_),
    .A1(exc_cause_1_),
    .A2(_03397_));
 sg13g2_a22oi_1 _11516_ (.Y(_03403_),
    .B1(net1489),
    .B2(crash_dump_o_3_),
    .A2(net1550),
    .A1(csr_depc_3_));
 sg13g2_nand2_2 _11517_ (.Y(_03404_),
    .A(_03402_),
    .B(_03403_));
 sg13g2_a21oi_2 _11518_ (.B1(_03404_),
    .Y(_03405_),
    .A2(net1551),
    .A1(data_addr_o_3_));
 sg13g2_nor2_2 _11519_ (.A(_03325_),
    .B(_03405_),
    .Y(_03406_));
 sg13g2_inv_1 _11520_ (.Y(_03407_),
    .A(_03406_));
 sg13g2_o21ai_1 _11521_ (.B1(_03407_),
    .Y(_00062_),
    .A1(net105),
    .A2(_03381_));
 sg13g2_inv_1 _11522_ (.Y(_03408_),
    .A(crash_dump_o_68_));
 sg13g2_and3_1 _11523_ (.X(_03409_),
    .A(crash_dump_o_66_),
    .B(crash_dump_o_67_),
    .C(_03294_));
 sg13g2_o21ai_1 _11524_ (.B1(_03117_),
    .Y(_03410_),
    .A1(_02350_),
    .A2(_03008_));
 sg13g2_mux2_1 _11525_ (.A0(_03115_),
    .A1(_03410_),
    .S(net176),
    .X(_03411_));
 sg13g2_xor2_1 _11526_ (.B(_03411_),
    .A(_03101_),
    .X(_03412_));
 sg13g2_nand2_1 _11527_ (.Y(_03413_),
    .A(net1551),
    .B(_03412_));
 sg13g2_o21ai_1 _11528_ (.B1(_03359_),
    .Y(_03414_),
    .A1(\id_stage_i.controller_i.irqs_i_18_ ),
    .A2(\id_stage_i.controller_i.irqs_i_16_ ));
 sg13g2_nand2_1 _11529_ (.Y(_03415_),
    .A(_03358_),
    .B(_03414_));
 sg13g2_nand2_1 _11530_ (.Y(_03416_),
    .A(_03340_),
    .B(_03357_));
 sg13g2_a21oi_2 _11531_ (.B1(_03416_),
    .Y(_03417_),
    .A2(_03415_),
    .A1(_03355_));
 sg13g2_a21o_1 _11532_ (.A2(net325),
    .A1(_03310_),
    .B1(_03417_),
    .X(exc_cause_2_));
 sg13g2_nor2b_1 _11533_ (.A(_03364_),
    .B_N(exc_cause_2_),
    .Y(_03418_));
 sg13g2_a221oi_1 _11534_ (.B2(crash_dump_o_4_),
    .C1(_03418_),
    .B1(net1489),
    .A1(csr_depc_4_),
    .Y(_03419_),
    .A2(net1550));
 sg13g2_a21oi_2 _11535_ (.B1(_03325_),
    .Y(_03420_),
    .A2(_03419_),
    .A1(_03413_));
 sg13g2_o21ai_1 _11536_ (.B1(net2489),
    .Y(_03421_),
    .A1(_03409_),
    .A2(_03420_));
 sg13g2_buf_2 fanout1061 (.A(_00615_),
    .X(net1061));
 sg13g2_nand3_1 _11538_ (.B(net776),
    .C(_03409_),
    .A(crash_dump_o_68_),
    .Y(_03423_));
 sg13g2_a21oi_1 _11539_ (.A1(net115),
    .A2(_03423_),
    .Y(_03424_),
    .B1(_03420_));
 sg13g2_a21oi_1 _11540_ (.A1(_03408_),
    .A2(_03421_),
    .Y(_00063_),
    .B1(_03424_));
 sg13g2_buf_2 fanout1060 (.A(_00621_),
    .X(net1060));
 sg13g2_xor2_1 _11542_ (.B(_03423_),
    .A(crash_dump_o_69_),
    .X(_03426_));
 sg13g2_buf_4 fanout1059 (.X(net1059),
    .A(\cs_registers_i/_0653_ ));
 sg13g2_nor4_2 _11544_ (.A(net1555),
    .B(net1545),
    .C(net1456),
    .Y(_03428_),
    .D(net1484));
 sg13g2_nand2_1 _11545_ (.Y(_03429_),
    .A(_03358_),
    .B(_03359_));
 sg13g2_o21ai_1 _11546_ (.B1(_03355_),
    .Y(_03430_),
    .A1(\id_stage_i.controller_i.irqs_i_16_ ),
    .A2(_03429_));
 sg13g2_nand3b_1 _11547_ (.B(_01453_),
    .C(_03310_),
    .Y(_03431_),
    .A_N(net464));
 sg13g2_o21ai_1 _11548_ (.B1(_03431_),
    .Y(exc_cause_3_),
    .A1(_03416_),
    .A2(_03430_));
 sg13g2_nand2b_1 _11549_ (.Y(_03432_),
    .B(exc_cause_3_),
    .A_N(_03364_));
 sg13g2_a22oi_1 _11550_ (.Y(_03433_),
    .B1(net1489),
    .B2(crash_dump_o_5_),
    .A2(net1550),
    .A1(csr_depc_5_));
 sg13g2_nand2_2 _11551_ (.Y(_03434_),
    .A(_03432_),
    .B(_03433_));
 sg13g2_a21oi_1 _11552_ (.A1(data_addr_o_5_),
    .A2(net1551),
    .Y(_03435_),
    .B1(_03434_));
 sg13g2_nor2_1 _11553_ (.A(net1395),
    .B(_03435_),
    .Y(_03436_));
 sg13g2_nor2_1 _11554_ (.A(net113),
    .B(_03436_),
    .Y(_03437_));
 sg13g2_a21oi_1 _11555_ (.A1(net116),
    .A2(_03426_),
    .Y(_00064_),
    .B1(_03437_));
 sg13g2_nand4_1 _11556_ (.B(crash_dump_o_69_),
    .C(net777),
    .A(crash_dump_o_68_),
    .Y(_03438_),
    .D(_03409_));
 sg13g2_xor2_1 _11557_ (.B(_03438_),
    .A(crash_dump_o_70_),
    .X(_03439_));
 sg13g2_nand2_2 _11558_ (.Y(_03440_),
    .A(_03340_),
    .B(_03360_));
 sg13g2_a22oi_1 _11559_ (.Y(_03441_),
    .B1(net1484),
    .B2(crash_dump_o_6_),
    .A2(net1545),
    .A1(csr_depc_6_));
 sg13g2_o21ai_1 _11560_ (.B1(_03441_),
    .Y(_03442_),
    .A1(_03364_),
    .A2(_03440_));
 sg13g2_a21oi_2 _11561_ (.B1(_03442_),
    .Y(_03443_),
    .A2(net1551),
    .A1(data_addr_o_6_));
 sg13g2_nor2_2 _11562_ (.A(net1396),
    .B(_03443_),
    .Y(_03444_));
 sg13g2_nor2_1 _11563_ (.A(net113),
    .B(_03444_),
    .Y(_03445_));
 sg13g2_a21oi_1 _11564_ (.A1(net115),
    .A2(_03439_),
    .Y(_00065_),
    .B1(_03445_));
 sg13g2_inv_1 _11565_ (.Y(_03446_),
    .A(crash_dump_o_71_));
 sg13g2_and4_1 _11566_ (.A(crash_dump_o_68_),
    .B(crash_dump_o_69_),
    .C(crash_dump_o_70_),
    .D(_03409_),
    .X(_03447_));
 sg13g2_nand2_1 _11567_ (.Y(_03448_),
    .A(data_addr_o_7_),
    .B(net1551));
 sg13g2_and3_1 _11568_ (.X(exc_cause_5_),
    .A(\id_stage_i.controller_i.handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .B(irq_nm_i),
    .C(exc_cause_6_));
 sg13g2_nor2b_1 _11569_ (.A(_03364_),
    .B_N(exc_cause_5_),
    .Y(_03449_));
 sg13g2_a221oi_1 _11570_ (.B2(crash_dump_o_7_),
    .C1(_03449_),
    .B1(net1487),
    .A1(csr_depc_7_),
    .Y(_03450_),
    .A2(net1548));
 sg13g2_a21oi_2 _11571_ (.B1(_03325_),
    .Y(_03451_),
    .A2(_03450_),
    .A1(_03448_));
 sg13g2_o21ai_1 _11572_ (.B1(net2489),
    .Y(_03452_),
    .A1(_03447_),
    .A2(_03451_));
 sg13g2_nand3_1 _11573_ (.B(net778),
    .C(_03447_),
    .A(crash_dump_o_71_),
    .Y(_03453_));
 sg13g2_a21oi_1 _11574_ (.A1(net116),
    .A2(_03453_),
    .Y(_03454_),
    .B1(_03451_));
 sg13g2_a21oi_1 _11575_ (.A1(_03446_),
    .A2(_03452_),
    .Y(_00066_),
    .B1(_03454_));
 sg13g2_xor2_1 _11576_ (.B(_03453_),
    .A(crash_dump_o_72_),
    .X(_03455_));
 sg13g2_inv_1 _11577_ (.Y(_03456_),
    .A(boot_addr_i_8_));
 sg13g2_and3_1 _11578_ (.X(_03457_),
    .A(_01631_),
    .B(net1456),
    .C(_03400_));
 sg13g2_buf_2 fanout1058 (.A(\cs_registers_i/_0764_ ),
    .X(net1058));
 sg13g2_a22oi_1 _11580_ (.Y(_03459_),
    .B1(net1488),
    .B2(crash_dump_o_8_),
    .A2(net1549),
    .A1(csr_depc_8_));
 sg13g2_nand2_1 _11581_ (.Y(_03460_),
    .A(net237),
    .B(_03459_));
 sg13g2_a221oi_1 _11582_ (.B2(csr_mtvec_8_),
    .C1(_03460_),
    .B1(net1393),
    .A1(data_addr_o_8_),
    .Y(_03461_),
    .A2(net1555));
 sg13g2_a21oi_2 _11583_ (.B1(_03461_),
    .Y(_03462_),
    .A2(net1395),
    .A1(_03456_));
 sg13g2_nor2_1 _11584_ (.A(net113),
    .B(_03462_),
    .Y(_03463_));
 sg13g2_a21oi_1 _11585_ (.A1(net115),
    .A2(_03455_),
    .Y(_00067_),
    .B1(_03463_));
 sg13g2_nand4_1 _11586_ (.B(crash_dump_o_72_),
    .C(net778),
    .A(crash_dump_o_71_),
    .Y(_03464_),
    .D(_03447_));
 sg13g2_xnor2_1 _11587_ (.Y(_03465_),
    .A(crash_dump_o_73_),
    .B(_03464_));
 sg13g2_nor2_1 _11588_ (.A(boot_addr_i_9_),
    .B(net237),
    .Y(_03466_));
 sg13g2_a22oi_1 _11589_ (.Y(_03467_),
    .B1(net1484),
    .B2(crash_dump_o_9_),
    .A2(net1545),
    .A1(csr_depc_9_));
 sg13g2_nand2_1 _11590_ (.Y(_03468_),
    .A(net237),
    .B(_03467_));
 sg13g2_a221oi_1 _11591_ (.B2(csr_mtvec_9_),
    .C1(_03468_),
    .B1(net1394),
    .A1(data_addr_o_9_),
    .Y(_03469_),
    .A2(net1555));
 sg13g2_nor3_2 _11592_ (.A(net111),
    .B(_03466_),
    .C(_03469_),
    .Y(_03470_));
 sg13g2_a21o_1 _11593_ (.A2(_03465_),
    .A1(net119),
    .B1(_03470_),
    .X(_00068_));
 sg13g2_and4_1 _11594_ (.A(crash_dump_o_71_),
    .B(crash_dump_o_72_),
    .C(crash_dump_o_73_),
    .D(_03447_),
    .X(_03471_));
 sg13g2_nand2_2 _11595_ (.Y(_03472_),
    .A(net775),
    .B(_03471_));
 sg13g2_xor2_1 _11596_ (.B(_03472_),
    .A(crash_dump_o_74_),
    .X(_03473_));
 sg13g2_nand2_1 _11597_ (.Y(_03474_),
    .A(csr_mtvec_10_),
    .B(net1392));
 sg13g2_nand2_1 _11598_ (.Y(_03475_),
    .A(data_addr_o_10_),
    .B(net1552));
 sg13g2_a22oi_1 _11599_ (.Y(_03476_),
    .B1(net1485),
    .B2(crash_dump_o_10_),
    .A2(net1546),
    .A1(csr_depc_10_));
 sg13g2_nand4_1 _11600_ (.B(_03474_),
    .C(_03475_),
    .A(net236),
    .Y(_03477_),
    .D(_03476_));
 sg13g2_o21ai_1 _11601_ (.B1(_03477_),
    .Y(_03478_),
    .A1(boot_addr_i_10_),
    .A2(net235));
 sg13g2_and2_1 _11602_ (.A(net104),
    .B(_03478_),
    .X(_03479_));
 sg13g2_a21oi_1 _11603_ (.A1(net115),
    .A2(_03473_),
    .Y(_00069_),
    .B1(_03479_));
 sg13g2_nand3_1 _11604_ (.B(net775),
    .C(_03471_),
    .A(crash_dump_o_74_),
    .Y(_03480_));
 sg13g2_xnor2_1 _11605_ (.Y(_03481_),
    .A(crash_dump_o_75_),
    .B(_03480_));
 sg13g2_nand2_2 _11606_ (.Y(_03482_),
    .A(_01631_),
    .B(_03400_));
 sg13g2_o21ai_1 _11607_ (.B1(net1456),
    .Y(_03483_),
    .A1(csr_mtvec_11_),
    .A2(_03482_));
 sg13g2_a22oi_1 _11608_ (.Y(_03484_),
    .B1(net1484),
    .B2(crash_dump_o_11_),
    .A2(net1545),
    .A1(csr_depc_11_));
 sg13g2_nand3_1 _11609_ (.B(_03483_),
    .C(_03484_),
    .A(net236),
    .Y(_03485_));
 sg13g2_a21oi_1 _11610_ (.A1(data_addr_o_11_),
    .A2(net1551),
    .Y(_03486_),
    .B1(_03485_));
 sg13g2_o21ai_1 _11611_ (.B1(net107),
    .Y(_03487_),
    .A1(boot_addr_i_11_),
    .A2(net235));
 sg13g2_nor2_2 _11612_ (.A(_03486_),
    .B(_03487_),
    .Y(_03488_));
 sg13g2_a21o_1 _11613_ (.A2(_03481_),
    .A1(net118),
    .B1(_03488_),
    .X(_00070_));
 sg13g2_nand4_1 _11614_ (.B(crash_dump_o_75_),
    .C(net775),
    .A(crash_dump_o_74_),
    .Y(_03489_),
    .D(_03471_));
 sg13g2_xnor2_1 _11615_ (.Y(_03490_),
    .A(crash_dump_o_76_),
    .B(_03489_));
 sg13g2_buf_4 fanout1057 (.X(net1057),
    .A(\cs_registers_i/_0764_ ));
 sg13g2_nor2_1 _11617_ (.A(boot_addr_i_12_),
    .B(net238),
    .Y(_03492_));
 sg13g2_a22oi_1 _11618_ (.Y(_03493_),
    .B1(net1485),
    .B2(crash_dump_o_12_),
    .A2(net1546),
    .A1(csr_depc_12_));
 sg13g2_nand2_1 _11619_ (.Y(_03494_),
    .A(net238),
    .B(_03493_));
 sg13g2_a221oi_1 _11620_ (.B2(csr_mtvec_12_),
    .C1(_03494_),
    .B1(net1392),
    .A1(data_addr_o_12_),
    .Y(_03495_),
    .A2(net1552));
 sg13g2_nor3_2 _11621_ (.A(net112),
    .B(_03492_),
    .C(_03495_),
    .Y(_03496_));
 sg13g2_a21o_1 _11622_ (.A2(_03490_),
    .A1(net118),
    .B1(_03496_),
    .X(_00071_));
 sg13g2_and4_1 _11623_ (.A(crash_dump_o_74_),
    .B(crash_dump_o_75_),
    .C(crash_dump_o_76_),
    .D(_03471_),
    .X(_03497_));
 sg13g2_nand2_2 _11624_ (.Y(_03498_),
    .A(net777),
    .B(_03497_));
 sg13g2_xnor2_1 _11625_ (.Y(_03499_),
    .A(crash_dump_o_77_),
    .B(_03498_));
 sg13g2_nand2_1 _11626_ (.Y(_03500_),
    .A(data_addr_o_13_),
    .B(net1556));
 sg13g2_a22oi_1 _11627_ (.Y(_03501_),
    .B1(net1488),
    .B2(crash_dump_o_13_),
    .A2(net1549),
    .A1(csr_depc_13_));
 sg13g2_nand2_1 _11628_ (.Y(_03502_),
    .A(net237),
    .B(_03501_));
 sg13g2_a21oi_2 _11629_ (.B1(_03502_),
    .Y(_03503_),
    .A2(net1394),
    .A1(csr_mtvec_13_));
 sg13g2_o21ai_1 _11630_ (.B1(net108),
    .Y(_03504_),
    .A1(boot_addr_i_13_),
    .A2(net235));
 sg13g2_a21oi_2 _11631_ (.B1(_03504_),
    .Y(_03505_),
    .A2(_03503_),
    .A1(_03500_));
 sg13g2_a21o_1 _11632_ (.A2(_03499_),
    .A1(net118),
    .B1(_03505_),
    .X(_00072_));
 sg13g2_nand3_1 _11633_ (.B(net775),
    .C(_03497_),
    .A(crash_dump_o_77_),
    .Y(_03506_));
 sg13g2_xor2_1 _11634_ (.B(_03506_),
    .A(crash_dump_o_78_),
    .X(_03507_));
 sg13g2_inv_1 _11635_ (.Y(_03508_),
    .A(net1556));
 sg13g2_nand2_1 _11636_ (.Y(_03509_),
    .A(_02117_),
    .B(_03037_));
 sg13g2_xor2_1 _11637_ (.B(_03509_),
    .A(_02465_),
    .X(_03510_));
 sg13g2_nand2_1 _11638_ (.Y(_03511_),
    .A(csr_mtvec_14_),
    .B(net1394));
 sg13g2_a22oi_1 _11639_ (.Y(_03512_),
    .B1(net1489),
    .B2(crash_dump_o_14_),
    .A2(net1550),
    .A1(csr_depc_14_));
 sg13g2_and3_2 _11640_ (.X(_03513_),
    .A(net235),
    .B(_03511_),
    .C(_03512_));
 sg13g2_o21ai_1 _11641_ (.B1(_03513_),
    .Y(_03514_),
    .A1(_03508_),
    .A2(_03510_));
 sg13g2_o21ai_1 _11642_ (.B1(_03513_),
    .Y(_03515_),
    .A1(_03039_),
    .A2(_03508_));
 sg13g2_mux2_2 _11643_ (.A0(_03514_),
    .A1(_03515_),
    .S(_03262_),
    .X(_03516_));
 sg13g2_o21ai_1 _11644_ (.B1(_03516_),
    .Y(_03517_),
    .A1(boot_addr_i_14_),
    .A2(net235));
 sg13g2_and2_1 _11645_ (.A(net104),
    .B(_03517_),
    .X(_03518_));
 sg13g2_a21oi_1 _11646_ (.A1(net115),
    .A2(_03507_),
    .Y(_00073_),
    .B1(_03518_));
 sg13g2_nand4_1 _11647_ (.B(crash_dump_o_78_),
    .C(net775),
    .A(crash_dump_o_77_),
    .Y(_03519_),
    .D(_03497_));
 sg13g2_xor2_1 _11648_ (.B(_03519_),
    .A(crash_dump_o_79_),
    .X(_03520_));
 sg13g2_buf_4 fanout1056 (.X(net1056),
    .A(\cs_registers_i/_0790_ ));
 sg13g2_nand2b_1 _11650_ (.Y(_03522_),
    .B(net1395),
    .A_N(boot_addr_i_15_));
 sg13g2_nand2_1 _11651_ (.Y(_03523_),
    .A(csr_mtvec_15_),
    .B(net1394));
 sg13g2_nand2_1 _11652_ (.Y(_03524_),
    .A(data_addr_o_15_),
    .B(net1554));
 sg13g2_a22oi_1 _11653_ (.Y(_03525_),
    .B1(net1484),
    .B2(crash_dump_o_15_),
    .A2(net1545),
    .A1(csr_depc_15_));
 sg13g2_nand4_1 _11654_ (.B(_03523_),
    .C(_03524_),
    .A(net237),
    .Y(_03526_),
    .D(_03525_));
 sg13g2_nand3_1 _11655_ (.B(_03522_),
    .C(_03526_),
    .A(net107),
    .Y(_03527_));
 sg13g2_o21ai_1 _11656_ (.B1(_03527_),
    .Y(_00074_),
    .A1(net105),
    .A2(_03520_));
 sg13g2_and4_1 _11657_ (.A(crash_dump_o_77_),
    .B(crash_dump_o_78_),
    .C(crash_dump_o_79_),
    .D(_03497_),
    .X(_03528_));
 sg13g2_nand2_2 _11658_ (.Y(_03529_),
    .A(net776),
    .B(_03528_));
 sg13g2_xor2_1 _11659_ (.B(_03529_),
    .A(crash_dump_o_80_),
    .X(_03530_));
 sg13g2_nand2b_1 _11660_ (.Y(_03531_),
    .B(net1395),
    .A_N(boot_addr_i_16_));
 sg13g2_o21ai_1 _11661_ (.B1(net1456),
    .Y(_03532_),
    .A1(csr_mtvec_16_),
    .A2(_03482_));
 sg13g2_nand2_1 _11662_ (.Y(_03533_),
    .A(data_addr_o_16_),
    .B(net1554));
 sg13g2_a22oi_1 _11663_ (.Y(_03534_),
    .B1(net1484),
    .B2(crash_dump_o_16_),
    .A2(net1545),
    .A1(csr_depc_16_));
 sg13g2_nand4_1 _11664_ (.B(_03532_),
    .C(_03533_),
    .A(net237),
    .Y(_03535_),
    .D(_03534_));
 sg13g2_nand3_1 _11665_ (.B(_03531_),
    .C(_03535_),
    .A(net107),
    .Y(_03536_));
 sg13g2_o21ai_1 _11666_ (.B1(_03536_),
    .Y(_00075_),
    .A1(net105),
    .A2(_03530_));
 sg13g2_buf_4 fanout1055 (.X(net1055),
    .A(\cs_registers_i/_0834_ ));
 sg13g2_nand2_1 _11668_ (.Y(_03538_),
    .A(csr_mtvec_17_),
    .B(net1392));
 sg13g2_a22oi_1 _11669_ (.Y(_03539_),
    .B1(net1487),
    .B2(crash_dump_o_17_),
    .A2(net1548),
    .A1(csr_depc_17_));
 sg13g2_nand2_1 _11670_ (.Y(_03540_),
    .A(data_addr_o_17_),
    .B(net1551));
 sg13g2_nand3_1 _11671_ (.B(_03539_),
    .C(_03540_),
    .A(_03538_),
    .Y(_03541_));
 sg13g2_nand2b_1 _11672_ (.Y(_03542_),
    .B(net1396),
    .A_N(boot_addr_i_17_));
 sg13g2_o21ai_1 _11673_ (.B1(_03542_),
    .Y(_03543_),
    .A1(net1396),
    .A2(_03541_));
 sg13g2_nand3_1 _11674_ (.B(net776),
    .C(_03528_),
    .A(crash_dump_o_80_),
    .Y(_03544_));
 sg13g2_xnor2_1 _11675_ (.Y(_03545_),
    .A(crash_dump_o_81_),
    .B(_03544_));
 sg13g2_nor2_1 _11676_ (.A(net106),
    .B(_03545_),
    .Y(_03546_));
 sg13g2_a21oi_1 _11677_ (.A1(net109),
    .A2(_03543_),
    .Y(_00076_),
    .B1(_03546_));
 sg13g2_nand2_1 _11678_ (.Y(_03547_),
    .A(csr_mtvec_18_),
    .B(net1392));
 sg13g2_nand2_1 _11679_ (.Y(_03548_),
    .A(data_addr_o_18_),
    .B(net1552));
 sg13g2_a22oi_1 _11680_ (.Y(_03549_),
    .B1(net1485),
    .B2(crash_dump_o_18_),
    .A2(net1546),
    .A1(csr_depc_18_));
 sg13g2_nand3_1 _11681_ (.B(_03548_),
    .C(_03549_),
    .A(_03547_),
    .Y(_03550_));
 sg13g2_nand2b_1 _11682_ (.Y(_03551_),
    .B(net1396),
    .A_N(boot_addr_i_18_));
 sg13g2_o21ai_1 _11683_ (.B1(_03551_),
    .Y(_03552_),
    .A1(net1396),
    .A2(_03550_));
 sg13g2_nand4_1 _11684_ (.B(crash_dump_o_81_),
    .C(net776),
    .A(crash_dump_o_80_),
    .Y(_03553_),
    .D(_03528_));
 sg13g2_xnor2_1 _11685_ (.Y(_03554_),
    .A(crash_dump_o_82_),
    .B(_03553_));
 sg13g2_nor2_1 _11686_ (.A(net106),
    .B(_03554_),
    .Y(_03555_));
 sg13g2_a21oi_1 _11687_ (.A1(net109),
    .A2(_03552_),
    .Y(_00077_),
    .B1(_03555_));
 sg13g2_and4_1 _11688_ (.A(crash_dump_o_80_),
    .B(crash_dump_o_81_),
    .C(crash_dump_o_82_),
    .D(_03528_),
    .X(_03556_));
 sg13g2_nand2_2 _11689_ (.Y(_03557_),
    .A(net775),
    .B(_03556_));
 sg13g2_xnor2_1 _11690_ (.Y(_03558_),
    .A(crash_dump_o_83_),
    .B(_03557_));
 sg13g2_a22oi_1 _11691_ (.Y(_03559_),
    .B1(net1487),
    .B2(crash_dump_o_19_),
    .A2(net1548),
    .A1(csr_depc_19_));
 sg13g2_nand2_1 _11692_ (.Y(_03560_),
    .A(net237),
    .B(_03559_));
 sg13g2_a221oi_1 _11693_ (.B2(csr_mtvec_19_),
    .C1(_03560_),
    .B1(net1392),
    .A1(data_addr_o_19_),
    .Y(_03561_),
    .A2(net1554));
 sg13g2_buf_2 fanout1054 (.A(\cs_registers_i/_0860_ ),
    .X(net1054));
 sg13g2_o21ai_1 _11695_ (.B1(net107),
    .Y(_03563_),
    .A1(boot_addr_i_19_),
    .A2(net236));
 sg13g2_nor2_2 _11696_ (.A(_03561_),
    .B(_03563_),
    .Y(_03564_));
 sg13g2_a21o_1 _11697_ (.A2(_03558_),
    .A1(net118),
    .B1(_03564_),
    .X(_00078_));
 sg13g2_nand3_1 _11698_ (.B(net774),
    .C(_03556_),
    .A(crash_dump_o_83_),
    .Y(_03565_));
 sg13g2_xor2_1 _11699_ (.B(_03565_),
    .A(crash_dump_o_84_),
    .X(_03566_));
 sg13g2_o21ai_1 _11700_ (.B1(net1456),
    .Y(_03567_),
    .A1(csr_mtvec_20_),
    .A2(_03482_));
 sg13g2_nand2_1 _11701_ (.Y(_03568_),
    .A(data_addr_o_20_),
    .B(net1552));
 sg13g2_a22oi_1 _11702_ (.Y(_03569_),
    .B1(net1485),
    .B2(crash_dump_o_20_),
    .A2(net1546),
    .A1(csr_depc_20_));
 sg13g2_nand3_1 _11703_ (.B(_03568_),
    .C(_03569_),
    .A(_03567_),
    .Y(_03570_));
 sg13g2_buf_8 fanout1053 (.A(\cs_registers_i/_0860_ ),
    .X(net1053));
 sg13g2_mux2_1 _11705_ (.A0(boot_addr_i_20_),
    .A1(_03570_),
    .S(net236),
    .X(_03572_));
 sg13g2_nor2_2 _11706_ (.A(net113),
    .B(_03572_),
    .Y(_03573_));
 sg13g2_a21oi_1 _11707_ (.A1(net115),
    .A2(_03566_),
    .Y(_00079_),
    .B1(_03573_));
 sg13g2_nand4_1 _11708_ (.B(crash_dump_o_84_),
    .C(net774),
    .A(crash_dump_o_83_),
    .Y(_03574_),
    .D(_03556_));
 sg13g2_xnor2_1 _11709_ (.Y(_03575_),
    .A(crash_dump_o_85_),
    .B(_03574_));
 sg13g2_nand2_1 _11710_ (.Y(_03576_),
    .A(csr_mtvec_21_),
    .B(net1393));
 sg13g2_nand2_1 _11711_ (.Y(_03577_),
    .A(data_addr_o_21_),
    .B(net1552));
 sg13g2_a22oi_1 _11712_ (.Y(_03578_),
    .B1(net1486),
    .B2(crash_dump_o_21_),
    .A2(net1547),
    .A1(csr_depc_21_));
 sg13g2_nand4_1 _11713_ (.B(_03576_),
    .C(_03577_),
    .A(net238),
    .Y(_03579_),
    .D(_03578_));
 sg13g2_o21ai_1 _11714_ (.B1(_03579_),
    .Y(_03580_),
    .A1(boot_addr_i_21_),
    .A2(net236));
 sg13g2_nor2_2 _11715_ (.A(net112),
    .B(_03580_),
    .Y(_03581_));
 sg13g2_a21o_1 _11716_ (.A2(_03575_),
    .A1(net118),
    .B1(_03581_),
    .X(_00080_));
 sg13g2_and4_1 _11717_ (.A(crash_dump_o_83_),
    .B(crash_dump_o_84_),
    .C(crash_dump_o_85_),
    .D(_03556_),
    .X(_03582_));
 sg13g2_nand2_2 _11718_ (.Y(_03583_),
    .A(net772),
    .B(_03582_));
 sg13g2_xor2_1 _11719_ (.B(_03583_),
    .A(crash_dump_o_86_),
    .X(_03584_));
 sg13g2_a22oi_1 _11720_ (.Y(_03585_),
    .B1(net1485),
    .B2(crash_dump_o_22_),
    .A2(net1546),
    .A1(csr_depc_22_));
 sg13g2_inv_1 _11721_ (.Y(_03586_),
    .A(_03585_));
 sg13g2_a221oi_1 _11722_ (.B2(csr_mtvec_22_),
    .C1(_03586_),
    .B1(net1393),
    .A1(data_addr_o_22_),
    .Y(_03587_),
    .A2(net1553));
 sg13g2_nor2_1 _11723_ (.A(boot_addr_i_22_),
    .B(net237),
    .Y(_03588_));
 sg13g2_a21oi_2 _11724_ (.B1(_03588_),
    .Y(_03589_),
    .A2(_03587_),
    .A1(net238));
 sg13g2_nor2_2 _11725_ (.A(net113),
    .B(_03589_),
    .Y(_03590_));
 sg13g2_a21oi_1 _11726_ (.A1(net115),
    .A2(_03584_),
    .Y(_00081_),
    .B1(_03590_));
 sg13g2_a22oi_1 _11727_ (.Y(_03591_),
    .B1(net1488),
    .B2(crash_dump_o_23_),
    .A2(net1549),
    .A1(csr_depc_23_));
 sg13g2_nand2_1 _11728_ (.Y(_03592_),
    .A(net238),
    .B(_03591_));
 sg13g2_a221oi_1 _11729_ (.B2(csr_mtvec_23_),
    .C1(_03592_),
    .B1(net1393),
    .A1(data_addr_o_23_),
    .Y(_03593_),
    .A2(net1553));
 sg13g2_o21ai_1 _11730_ (.B1(net107),
    .Y(_03594_),
    .A1(boot_addr_i_23_),
    .A2(net235));
 sg13g2_nor2_2 _11731_ (.A(_03593_),
    .B(_03594_),
    .Y(_03595_));
 sg13g2_a21o_1 _11732_ (.A2(_03582_),
    .A1(crash_dump_o_86_),
    .B1(_03595_),
    .X(_03596_));
 sg13g2_a21oi_1 _11733_ (.A1(net2488),
    .A2(_03596_),
    .Y(_03597_),
    .B1(crash_dump_o_87_));
 sg13g2_nand4_1 _11734_ (.B(crash_dump_o_87_),
    .C(net772),
    .A(crash_dump_o_86_),
    .Y(_03598_),
    .D(_03582_));
 sg13g2_a21oi_1 _11735_ (.A1(net115),
    .A2(_03598_),
    .Y(_03599_),
    .B1(_03595_));
 sg13g2_nor2_1 _11736_ (.A(_03597_),
    .B(_03599_),
    .Y(_00082_));
 sg13g2_xnor2_1 _11737_ (.Y(_03600_),
    .A(crash_dump_o_88_),
    .B(_03598_));
 sg13g2_a22oi_1 _11738_ (.Y(_03601_),
    .B1(net1486),
    .B2(crash_dump_o_24_),
    .A2(net1547),
    .A1(csr_depc_24_));
 sg13g2_nand2_1 _11739_ (.Y(_03602_),
    .A(net238),
    .B(_03601_));
 sg13g2_a221oi_1 _11740_ (.B2(csr_mtvec_24_),
    .C1(_03602_),
    .B1(net1393),
    .A1(data_addr_o_24_),
    .Y(_03603_),
    .A2(net1553));
 sg13g2_o21ai_1 _11741_ (.B1(net108),
    .Y(_03604_),
    .A1(boot_addr_i_24_),
    .A2(net235));
 sg13g2_nor2_2 _11742_ (.A(_03603_),
    .B(_03604_),
    .Y(_03605_));
 sg13g2_a21o_1 _11743_ (.A2(_03600_),
    .A1(net118),
    .B1(_03605_),
    .X(_00083_));
 sg13g2_o21ai_1 _11744_ (.B1(net1456),
    .Y(_03606_),
    .A1(csr_mtvec_25_),
    .A2(_03482_));
 sg13g2_nand2_1 _11745_ (.Y(_03607_),
    .A(data_addr_o_25_),
    .B(net1553));
 sg13g2_a22oi_1 _11746_ (.Y(_03608_),
    .B1(net1485),
    .B2(crash_dump_o_25_),
    .A2(net1546),
    .A1(csr_depc_25_));
 sg13g2_nand4_1 _11747_ (.B(_03606_),
    .C(_03607_),
    .A(net238),
    .Y(_03609_),
    .D(_03608_));
 sg13g2_o21ai_1 _11748_ (.B1(_03609_),
    .Y(_03610_),
    .A1(boot_addr_i_25_),
    .A2(net236));
 sg13g2_and4_1 _11749_ (.A(crash_dump_o_86_),
    .B(crash_dump_o_87_),
    .C(crash_dump_o_88_),
    .D(_03582_),
    .X(_03611_));
 sg13g2_nand2_2 _11750_ (.Y(_03612_),
    .A(net776),
    .B(_03611_));
 sg13g2_xnor2_1 _11751_ (.Y(_03613_),
    .A(crash_dump_o_89_),
    .B(_03612_));
 sg13g2_nor2_1 _11752_ (.A(net106),
    .B(_03613_),
    .Y(_03614_));
 sg13g2_a21oi_1 _11753_ (.A1(_03283_),
    .A2(_03610_),
    .Y(_00084_),
    .B1(_03614_));
 sg13g2_nand3_1 _11754_ (.B(net774),
    .C(_03611_),
    .A(crash_dump_o_89_),
    .Y(_03615_));
 sg13g2_xnor2_1 _11755_ (.Y(_03616_),
    .A(crash_dump_o_90_),
    .B(_03615_));
 sg13g2_nand2_1 _11756_ (.Y(_03617_),
    .A(csr_mtvec_26_),
    .B(net1392));
 sg13g2_nand2_1 _11757_ (.Y(_03618_),
    .A(data_addr_o_26_),
    .B(net1552));
 sg13g2_a22oi_1 _11758_ (.Y(_03619_),
    .B1(net1487),
    .B2(crash_dump_o_26_),
    .A2(net1548),
    .A1(csr_depc_26_));
 sg13g2_nand4_1 _11759_ (.B(_03617_),
    .C(_03618_),
    .A(net239),
    .Y(_03620_),
    .D(_03619_));
 sg13g2_o21ai_1 _11760_ (.B1(_03620_),
    .Y(_03621_),
    .A1(boot_addr_i_26_),
    .A2(net236));
 sg13g2_nor2_2 _11761_ (.A(net112),
    .B(_03621_),
    .Y(_03622_));
 sg13g2_a21o_1 _11762_ (.A2(_03616_),
    .A1(net118),
    .B1(_03622_),
    .X(_00085_));
 sg13g2_nand4_1 _11763_ (.B(crash_dump_o_90_),
    .C(net774),
    .A(crash_dump_o_89_),
    .Y(_03623_),
    .D(_03611_));
 sg13g2_xor2_1 _11764_ (.B(_03623_),
    .A(crash_dump_o_91_),
    .X(_03624_));
 sg13g2_nand2b_1 _11765_ (.Y(_03625_),
    .B(net1395),
    .A_N(boot_addr_i_27_));
 sg13g2_o21ai_1 _11766_ (.B1(net1456),
    .Y(_03626_),
    .A1(csr_mtvec_27_),
    .A2(_03482_));
 sg13g2_nand2_1 _11767_ (.Y(_03627_),
    .A(data_addr_o_27_),
    .B(net1554));
 sg13g2_a22oi_1 _11768_ (.Y(_03628_),
    .B1(net1487),
    .B2(crash_dump_o_27_),
    .A2(net1548),
    .A1(csr_depc_27_));
 sg13g2_nand4_1 _11769_ (.B(_03626_),
    .C(_03627_),
    .A(net239),
    .Y(_03629_),
    .D(_03628_));
 sg13g2_nand3_1 _11770_ (.B(_03625_),
    .C(_03629_),
    .A(net108),
    .Y(_03630_));
 sg13g2_o21ai_1 _11771_ (.B1(_03630_),
    .Y(_00086_),
    .A1(net105),
    .A2(_03624_));
 sg13g2_and4_1 _11772_ (.A(crash_dump_o_89_),
    .B(crash_dump_o_90_),
    .C(crash_dump_o_91_),
    .D(_03611_),
    .X(_03631_));
 sg13g2_nand2_2 _11773_ (.Y(_03632_),
    .A(net776),
    .B(_03631_));
 sg13g2_xor2_1 _11774_ (.B(_03632_),
    .A(crash_dump_o_92_),
    .X(_03633_));
 sg13g2_o21ai_1 _11775_ (.B1(_03322_),
    .Y(_03634_),
    .A1(csr_mtvec_28_),
    .A2(_03482_));
 sg13g2_nand2_1 _11776_ (.Y(_03635_),
    .A(data_addr_o_28_),
    .B(net1552));
 sg13g2_a22oi_1 _11777_ (.Y(_03636_),
    .B1(net1485),
    .B2(crash_dump_o_28_),
    .A2(net1546),
    .A1(csr_depc_28_));
 sg13g2_nand4_1 _11778_ (.B(_03634_),
    .C(_03635_),
    .A(net239),
    .Y(_03637_),
    .D(_03636_));
 sg13g2_o21ai_1 _11779_ (.B1(_03637_),
    .Y(_03638_),
    .A1(boot_addr_i_28_),
    .A2(net236));
 sg13g2_nand2b_2 _11780_ (.Y(_03639_),
    .B(net108),
    .A_N(_03638_));
 sg13g2_o21ai_1 _11781_ (.B1(_03639_),
    .Y(_00087_),
    .A1(net106),
    .A2(_03633_));
 sg13g2_nand2_1 _11782_ (.Y(_03640_),
    .A(crash_dump_o_92_),
    .B(_03631_));
 sg13g2_nand2b_1 _11783_ (.Y(_03641_),
    .B(net1395),
    .A_N(boot_addr_i_29_));
 sg13g2_nand2_1 _11784_ (.Y(_03642_),
    .A(csr_mtvec_29_),
    .B(net1392));
 sg13g2_nand2_1 _11785_ (.Y(_03643_),
    .A(data_addr_o_29_),
    .B(net1553));
 sg13g2_a22oi_1 _11786_ (.Y(_03644_),
    .B1(net1485),
    .B2(crash_dump_o_29_),
    .A2(net1546),
    .A1(csr_depc_29_));
 sg13g2_nand4_1 _11787_ (.B(_03642_),
    .C(_03643_),
    .A(net239),
    .Y(_03645_),
    .D(_03644_));
 sg13g2_nand3_1 _11788_ (.B(_03641_),
    .C(_03645_),
    .A(net108),
    .Y(_03646_));
 sg13g2_nand2_1 _11789_ (.Y(_03647_),
    .A(_03640_),
    .B(net2470));
 sg13g2_a21oi_1 _11790_ (.A1(net2488),
    .A2(_03647_),
    .Y(_03648_),
    .B1(crash_dump_o_93_));
 sg13g2_and4_1 _11791_ (.A(crash_dump_o_92_),
    .B(crash_dump_o_93_),
    .C(net776),
    .D(_03631_),
    .X(_03649_));
 sg13g2_o21ai_1 _11792_ (.B1(net2470),
    .Y(_03650_),
    .A1(net106),
    .A2(_03649_));
 sg13g2_nor2b_1 _11793_ (.A(_03648_),
    .B_N(_03650_),
    .Y(_00088_));
 sg13g2_xnor2_1 _11794_ (.Y(_03651_),
    .A(crash_dump_o_94_),
    .B(_03649_));
 sg13g2_nand2b_1 _11795_ (.Y(_03652_),
    .B(net1395),
    .A_N(boot_addr_i_30_));
 sg13g2_nand2_1 _11796_ (.Y(_03653_),
    .A(csr_mtvec_30_),
    .B(net1394));
 sg13g2_nand2_1 _11797_ (.Y(_03654_),
    .A(data_addr_o_30_),
    .B(net1553));
 sg13g2_a22oi_1 _11798_ (.Y(_03655_),
    .B1(net1486),
    .B2(crash_dump_o_30_),
    .A2(net1547),
    .A1(csr_depc_30_));
 sg13g2_nand4_1 _11799_ (.B(_03653_),
    .C(_03654_),
    .A(net239),
    .Y(_03656_),
    .D(_03655_));
 sg13g2_nand3_1 _11800_ (.B(_03652_),
    .C(_03656_),
    .A(net108),
    .Y(_03657_));
 sg13g2_o21ai_1 _11801_ (.B1(_03657_),
    .Y(_00089_),
    .A1(net106),
    .A2(_03651_));
 sg13g2_nand2_2 _11802_ (.Y(_03658_),
    .A(crash_dump_o_94_),
    .B(_03649_));
 sg13g2_xor2_1 _11803_ (.B(_03658_),
    .A(crash_dump_o_95_),
    .X(_03659_));
 sg13g2_nand2b_1 _11804_ (.Y(_03660_),
    .B(net1395),
    .A_N(boot_addr_i_31_));
 sg13g2_nand2_1 _11805_ (.Y(_03661_),
    .A(csr_mtvec_31_),
    .B(net1392));
 sg13g2_nand2_1 _11806_ (.Y(_03662_),
    .A(net36),
    .B(net1552));
 sg13g2_a22oi_1 _11807_ (.Y(_03663_),
    .B1(net1486),
    .B2(crash_dump_o_31_),
    .A2(net1547),
    .A1(csr_depc_31_));
 sg13g2_nand4_1 _11808_ (.B(_03661_),
    .C(_03662_),
    .A(net238),
    .Y(_03664_),
    .D(_03663_));
 sg13g2_nand3_1 _11809_ (.B(_03660_),
    .C(_03664_),
    .A(net108),
    .Y(_03665_));
 sg13g2_o21ai_1 _11810_ (.B1(net2491),
    .Y(_00090_),
    .A1(net105),
    .A2(_03659_));
 sg13g2_buf_2 fanout1052 (.A(\cs_registers_i/_0883_ ),
    .X(net1052));
 sg13g2_nor2b_1 _11812_ (.A(net775),
    .B_N(crash_dump_o_96_),
    .Y(_00091_));
 sg13g2_mux2_1 _11813_ (.A0(crash_dump_o_97_),
    .A1(net561),
    .S(net768),
    .X(_00092_));
 sg13g2_mux2_1 _11814_ (.A0(crash_dump_o_98_),
    .A1(crash_dump_o_66_),
    .S(net773),
    .X(_00093_));
 sg13g2_mux2_1 _11815_ (.A0(crash_dump_o_99_),
    .A1(crash_dump_o_67_),
    .S(net771),
    .X(_00094_));
 sg13g2_buf_4 fanout1051 (.X(net1051),
    .A(\cs_registers_i/_0883_ ));
 sg13g2_inv_1 _11817_ (.Y(csr_access),
    .A(net1402));
 sg13g2_buf_8 fanout1050 (.A(\cs_registers_i/_0903_ ),
    .X(net1050));
 sg13g2_buf_8 fanout1049 (.A(\cs_registers_i/_0961_ ),
    .X(net1049));
 sg13g2_nor2_1 _11820_ (.A(net1403),
    .B(net1461),
    .Y(csr_addr_0_));
 sg13g2_nor2_2 _11821_ (.A(net1403),
    .B(_02134_),
    .Y(csr_addr_10_));
 sg13g2_nor2_1 _11822_ (.A(net1402),
    .B(_02998_),
    .Y(csr_addr_11_));
 sg13g2_nor2_2 _11823_ (.A(net1403),
    .B(_03061_),
    .Y(csr_addr_1_));
 sg13g2_nor2_2 _11824_ (.A(net1402),
    .B(_02412_),
    .Y(csr_addr_2_));
 sg13g2_nor2_1 _11825_ (.A(net1402),
    .B(_03244_),
    .Y(csr_addr_3_));
 sg13g2_nor2_2 _11826_ (.A(net1402),
    .B(_02261_),
    .Y(csr_addr_4_));
 sg13g2_nor2_1 _11827_ (.A(net1402),
    .B(_02367_),
    .Y(csr_addr_5_));
 sg13g2_nor2_1 _11828_ (.A(net1402),
    .B(_02387_),
    .Y(csr_addr_6_));
 sg13g2_nor2_2 _11829_ (.A(net1403),
    .B(_02164_),
    .Y(csr_addr_7_));
 sg13g2_nor2_2 _11830_ (.A(net1403),
    .B(_02159_),
    .Y(csr_addr_8_));
 sg13g2_nor2_2 _11831_ (.A(net1402),
    .B(_02148_),
    .Y(csr_addr_9_));
 sg13g2_buf_2 fanout1048 (.A(\cs_registers_i/_0983_ ),
    .X(net1048));
 sg13g2_buf_8 fanout1047 (.A(\cs_registers_i/_0983_ ),
    .X(net1047));
 sg13g2_buf_4 fanout1046 (.X(net1046),
    .A(\cs_registers_i/_1031_ ));
 sg13g2_buf_2 fanout1045 (.A(\cs_registers_i/_1052_ ),
    .X(net1045));
 sg13g2_buf_8 fanout1044 (.A(\cs_registers_i/_1052_ ),
    .X(net1044));
 sg13g2_buf_4 fanout1043 (.X(net1043),
    .A(\cs_registers_i/_1079_ ));
 sg13g2_nor2b_1 _11838_ (.A(net440),
    .B_N(\id_stage_i.controller_i.instr_i_0_ ),
    .Y(_03676_));
 sg13g2_a21oi_1 _11839_ (.A1(net440),
    .A2(\id_stage_i.controller_i.instr_compressed_i_0_ ),
    .Y(_03677_),
    .B1(_03676_));
 sg13g2_nor3_1 _11840_ (.A(_03329_),
    .B(net1898),
    .C(_03677_),
    .Y(_03678_));
 sg13g2_a221oi_1 _11841_ (.B2(crash_dump_o_32_),
    .C1(_03678_),
    .B1(net324),
    .A1(crash_dump_o_96_),
    .Y(_03679_),
    .A2(net1898));
 sg13g2_nor2_1 _11842_ (.A(net1645),
    .B(_03679_),
    .Y(csr_mtval_0_));
 sg13g2_buf_4 fanout1042 (.X(net1042),
    .A(\cs_registers_i/_1152_ ));
 sg13g2_nand2_1 _11844_ (.Y(_03681_),
    .A(crash_dump_o_42_),
    .B(net328));
 sg13g2_nor2_2 _11845_ (.A(_03329_),
    .B(net1898),
    .Y(_03682_));
 sg13g2_nand2_1 _11846_ (.Y(_03683_),
    .A(net440),
    .B(\id_stage_i.controller_i.instr_compressed_i_10_ ));
 sg13g2_o21ai_1 _11847_ (.B1(_03683_),
    .Y(_03684_),
    .A1(net439),
    .A2(_02284_));
 sg13g2_and2_1 _11848_ (.A(crash_dump_o_97_),
    .B(crash_dump_o_98_),
    .X(_03685_));
 sg13g2_and4_1 _11849_ (.A(crash_dump_o_100_),
    .B(crash_dump_o_99_),
    .C(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .D(_03685_),
    .X(_03686_));
 sg13g2_and2_1 _11850_ (.A(crash_dump_o_101_),
    .B(_03686_),
    .X(_03687_));
 sg13g2_nand3_1 _11851_ (.B(crash_dump_o_103_),
    .C(_03687_),
    .A(crash_dump_o_102_),
    .Y(_03688_));
 sg13g2_nor2_1 _11852_ (.A(_03200_),
    .B(_03688_),
    .Y(_03689_));
 sg13g2_nand2_1 _11853_ (.Y(_03690_),
    .A(crash_dump_o_105_),
    .B(_03689_));
 sg13g2_xnor2_1 _11854_ (.Y(_03691_),
    .A(crash_dump_o_106_),
    .B(_03690_));
 sg13g2_a22oi_1 _11855_ (.Y(_03692_),
    .B1(_03691_),
    .B2(net1902),
    .A2(_03684_),
    .A1(_03682_));
 sg13g2_o21ai_1 _11856_ (.B1(_03310_),
    .Y(_03693_),
    .A1(_03331_),
    .A2(net328));
 sg13g2_a21oi_1 _11857_ (.A1(_03681_),
    .A2(_03692_),
    .Y(csr_mtval_10_),
    .B1(net1544));
 sg13g2_nand2_1 _11858_ (.Y(_03694_),
    .A(crash_dump_o_43_),
    .B(net328));
 sg13g2_mux2_1 _11859_ (.A0(net553),
    .A1(\id_stage_i.controller_i.instr_compressed_i_11_ ),
    .S(net439),
    .X(_03695_));
 sg13g2_nand3_1 _11860_ (.B(crash_dump_o_106_),
    .C(_03689_),
    .A(crash_dump_o_105_),
    .Y(_03696_));
 sg13g2_xnor2_1 _11861_ (.Y(_03697_),
    .A(crash_dump_o_107_),
    .B(_03696_));
 sg13g2_a22oi_1 _11862_ (.Y(_03698_),
    .B1(_03697_),
    .B2(net1902),
    .A2(_03695_),
    .A1(_03682_));
 sg13g2_buf_2 fanout1041 (.A(\cs_registers_i/_1181_ ),
    .X(net1041));
 sg13g2_a21oi_1 _11864_ (.A1(_03694_),
    .A2(_03698_),
    .Y(csr_mtval_11_),
    .B1(net1642));
 sg13g2_nor2_1 _11865_ (.A(_01212_),
    .B(_03696_),
    .Y(_03700_));
 sg13g2_xnor2_1 _11866_ (.Y(_03701_),
    .A(crash_dump_o_108_),
    .B(_03700_));
 sg13g2_buf_8 fanout1040 (.A(\cs_registers_i/_1181_ ),
    .X(net1040));
 sg13g2_buf_4 fanout1039 (.X(net1039),
    .A(\cs_registers_i/_1203_ ));
 sg13g2_mux2_1 _11869_ (.A0(net2098),
    .A1(\id_stage_i.controller_i.instr_compressed_i_12_ ),
    .S(net440),
    .X(_03704_));
 sg13g2_a21oi_1 _11870_ (.A1(net2100),
    .A2(_03704_),
    .Y(_03705_),
    .B1(net1897));
 sg13g2_a21oi_1 _11871_ (.A1(net1900),
    .A2(_03701_),
    .Y(_03706_),
    .B1(_03705_));
 sg13g2_a21oi_1 _11872_ (.A1(crash_dump_o_44_),
    .A2(net325),
    .Y(_03707_),
    .B1(_03706_));
 sg13g2_nor2_1 _11873_ (.A(net1643),
    .B(_03707_),
    .Y(csr_mtval_12_));
 sg13g2_nand2_1 _11874_ (.Y(_03708_),
    .A(crash_dump_o_108_),
    .B(_03700_));
 sg13g2_xor2_1 _11875_ (.B(_03708_),
    .A(crash_dump_o_109_),
    .X(_03709_));
 sg13g2_nand2_1 _11876_ (.Y(_03710_),
    .A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .B(\id_stage_i.controller_i.instr_compressed_i_13_ ));
 sg13g2_o21ai_1 _11877_ (.B1(_03710_),
    .Y(_03711_),
    .A1(net440),
    .A2(_01361_));
 sg13g2_a21oi_1 _11878_ (.A1(net2100),
    .A2(_03711_),
    .Y(_03712_),
    .B1(net1897));
 sg13g2_a21oi_1 _11879_ (.A1(net1900),
    .A2(_03709_),
    .Y(_03713_),
    .B1(_03712_));
 sg13g2_a21oi_1 _11880_ (.A1(crash_dump_o_45_),
    .A2(net325),
    .Y(_03714_),
    .B1(_03713_));
 sg13g2_nor2_1 _11881_ (.A(net1643),
    .B(_03714_),
    .Y(csr_mtval_13_));
 sg13g2_buf_4 fanout1038 (.X(net1038),
    .A(net1039));
 sg13g2_nand3_1 _11883_ (.B(crash_dump_o_109_),
    .C(_03700_),
    .A(crash_dump_o_108_),
    .Y(_03716_));
 sg13g2_xnor2_1 _11884_ (.Y(_03717_),
    .A(crash_dump_o_110_),
    .B(_03716_));
 sg13g2_nand2_1 _11885_ (.Y(_03718_),
    .A(net1900),
    .B(_03717_));
 sg13g2_mux2_1 _11886_ (.A0(net2089),
    .A1(\id_stage_i.controller_i.instr_compressed_i_14_ ),
    .S(net439),
    .X(_03719_));
 sg13g2_a22oi_1 _11887_ (.Y(_03720_),
    .B1(_03682_),
    .B2(_03719_),
    .A2(net326),
    .A1(crash_dump_o_46_));
 sg13g2_a21oi_1 _11888_ (.A1(_03718_),
    .A2(_03720_),
    .Y(csr_mtval_14_),
    .B1(net1544));
 sg13g2_nor2_1 _11889_ (.A(_03207_),
    .B(_03716_),
    .Y(_03721_));
 sg13g2_xnor2_1 _11890_ (.Y(_03722_),
    .A(crash_dump_o_111_),
    .B(_03721_));
 sg13g2_mux2_1 _11891_ (.A0(net2081),
    .A1(\id_stage_i.controller_i.instr_compressed_i_15_ ),
    .S(net440),
    .X(_03723_));
 sg13g2_a21oi_1 _11892_ (.A1(net2101),
    .A2(_03723_),
    .Y(_03724_),
    .B1(net1897));
 sg13g2_a21oi_1 _11893_ (.A1(net1900),
    .A2(_03722_),
    .Y(_03725_),
    .B1(_03724_));
 sg13g2_a21oi_1 _11894_ (.A1(crash_dump_o_47_),
    .A2(net325),
    .Y(_03726_),
    .B1(_03725_));
 sg13g2_nor2_1 _11895_ (.A(net1643),
    .B(_03726_),
    .Y(csr_mtval_15_));
 sg13g2_nor3_2 _11896_ (.A(_03207_),
    .B(_01226_),
    .C(_03716_),
    .Y(_03727_));
 sg13g2_xor2_1 _11897_ (.B(_03727_),
    .A(crash_dump_o_112_),
    .X(_03728_));
 sg13g2_nand2_1 _11898_ (.Y(_03729_),
    .A(net1901),
    .B(_03728_));
 sg13g2_nor2_1 _11899_ (.A(net438),
    .B(_03385_),
    .Y(_03730_));
 sg13g2_buf_4 fanout1037 (.X(net1037),
    .A(\cs_registers_i/_1224_ ));
 sg13g2_a22oi_1 _11901_ (.Y(_03732_),
    .B1(net1641),
    .B2(net536),
    .A2(net326),
    .A1(crash_dump_o_48_));
 sg13g2_a21oi_2 _11902_ (.B1(net1544),
    .Y(csr_mtval_16_),
    .A2(_03732_),
    .A1(_03729_));
 sg13g2_nand2_1 _11903_ (.Y(_03733_),
    .A(net530),
    .B(net2100));
 sg13g2_o21ai_1 _11904_ (.B1(net1880),
    .Y(_03734_),
    .A1(net438),
    .A2(_03733_));
 sg13g2_nand2_1 _11905_ (.Y(_03735_),
    .A(crash_dump_o_112_),
    .B(_03727_));
 sg13g2_xor2_1 _11906_ (.B(_03735_),
    .A(crash_dump_o_113_),
    .X(_03736_));
 sg13g2_nand2_1 _11907_ (.Y(_03737_),
    .A(net1900),
    .B(_03736_));
 sg13g2_a22oi_1 _11908_ (.Y(_03738_),
    .B1(_03734_),
    .B2(_03737_),
    .A2(net326),
    .A1(crash_dump_o_49_));
 sg13g2_nor2_1 _11909_ (.A(net1643),
    .B(_03738_),
    .Y(csr_mtval_17_));
 sg13g2_nand3_1 _11910_ (.B(crash_dump_o_113_),
    .C(_03727_),
    .A(crash_dump_o_112_),
    .Y(_03739_));
 sg13g2_xnor2_1 _11911_ (.Y(_03740_),
    .A(crash_dump_o_114_),
    .B(_03739_));
 sg13g2_nand2_1 _11912_ (.Y(_03741_),
    .A(net1901),
    .B(_03740_));
 sg13g2_a22oi_1 _11913_ (.Y(_03742_),
    .B1(net1641),
    .B2(\id_stage_i.controller_i.instr_i_18_ ),
    .A2(net326),
    .A1(crash_dump_o_50_));
 sg13g2_a21oi_1 _11914_ (.A1(_03741_),
    .A2(_03742_),
    .Y(csr_mtval_18_),
    .B1(net1544));
 sg13g2_nor2_1 _11915_ (.A(_01240_),
    .B(_03739_),
    .Y(_03743_));
 sg13g2_xor2_1 _11916_ (.B(_03743_),
    .A(crash_dump_o_115_),
    .X(_03744_));
 sg13g2_nand2_1 _11917_ (.Y(_03745_),
    .A(net1900),
    .B(_03744_));
 sg13g2_a22oi_1 _11918_ (.Y(_03746_),
    .B1(net1641),
    .B2(\id_stage_i.controller_i.instr_i_19_ ),
    .A2(net325),
    .A1(crash_dump_o_51_));
 sg13g2_a21oi_1 _11919_ (.A1(_03745_),
    .A2(_03746_),
    .Y(csr_mtval_19_),
    .B1(net1643));
 sg13g2_nor2b_1 _11920_ (.A(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .B_N(crash_dump_o_97_),
    .Y(_03747_));
 sg13g2_a21oi_1 _11921_ (.A1(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .A2(\csr_mtval_1__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_MUX__Y_B ),
    .Y(_03748_),
    .B1(_03747_));
 sg13g2_mux2_1 _11922_ (.A0(\id_stage_i.controller_i.instr_i_1_ ),
    .A1(\id_stage_i.controller_i.instr_compressed_i_1_ ),
    .S(net438),
    .X(_03749_));
 sg13g2_a21oi_1 _11923_ (.A1(\id_stage_i.controller_i.illegal_insn_q ),
    .A2(_03749_),
    .Y(_03750_),
    .B1(net1897));
 sg13g2_a21oi_1 _11924_ (.A1(net1898),
    .A2(_03748_),
    .Y(_03751_),
    .B1(_03750_));
 sg13g2_a21oi_1 _11925_ (.A1(crash_dump_o_33_),
    .A2(net325),
    .Y(_03752_),
    .B1(_03751_));
 sg13g2_nor2_1 _11926_ (.A(net1645),
    .B(_03752_),
    .Y(csr_mtval_1_));
 sg13g2_nand2_1 _11927_ (.Y(_03753_),
    .A(crash_dump_o_115_),
    .B(_03743_));
 sg13g2_xnor2_1 _11928_ (.Y(_03754_),
    .A(crash_dump_o_116_),
    .B(_03753_));
 sg13g2_nand2_1 _11929_ (.Y(_03755_),
    .A(net1900),
    .B(_03754_));
 sg13g2_buf_4 fanout1036 (.X(net1036),
    .A(\cs_registers_i/_1244_ ));
 sg13g2_a22oi_1 _11931_ (.Y(_03757_),
    .B1(net1641),
    .B2(net513),
    .A2(net327),
    .A1(crash_dump_o_52_));
 sg13g2_a21oi_1 _11932_ (.A1(_03755_),
    .A2(_03757_),
    .Y(csr_mtval_20_),
    .B1(net1544));
 sg13g2_nand3_1 _11933_ (.B(crash_dump_o_116_),
    .C(_03743_),
    .A(crash_dump_o_115_),
    .Y(_03758_));
 sg13g2_xnor2_1 _11934_ (.Y(_03759_),
    .A(crash_dump_o_117_),
    .B(_03758_));
 sg13g2_nand2_1 _11935_ (.Y(_03760_),
    .A(net1899),
    .B(_03759_));
 sg13g2_a22oi_1 _11936_ (.Y(_03761_),
    .B1(net1640),
    .B2(net453),
    .A2(net327),
    .A1(crash_dump_o_53_));
 sg13g2_a21oi_1 _11937_ (.A1(_03760_),
    .A2(_03761_),
    .Y(csr_mtval_21_),
    .B1(net1643));
 sg13g2_nor2_1 _11938_ (.A(_01255_),
    .B(_03758_),
    .Y(_03762_));
 sg13g2_xor2_1 _11939_ (.B(_03762_),
    .A(crash_dump_o_118_),
    .X(_03763_));
 sg13g2_nand2_1 _11940_ (.Y(_03764_),
    .A(net1901),
    .B(_03763_));
 sg13g2_a22oi_1 _11941_ (.Y(_03765_),
    .B1(net1641),
    .B2(net447),
    .A2(net327),
    .A1(crash_dump_o_54_));
 sg13g2_a21oi_1 _11942_ (.A1(_03764_),
    .A2(_03765_),
    .Y(csr_mtval_22_),
    .B1(net1544));
 sg13g2_nand2_1 _11943_ (.Y(_03766_),
    .A(crash_dump_o_118_),
    .B(_03762_));
 sg13g2_xnor2_1 _11944_ (.Y(_03767_),
    .A(crash_dump_o_119_),
    .B(_03766_));
 sg13g2_nand2_1 _11945_ (.Y(_03768_),
    .A(net1899),
    .B(_03767_));
 sg13g2_a22oi_1 _11946_ (.Y(_03769_),
    .B1(net1640),
    .B2(net2008),
    .A2(net327),
    .A1(crash_dump_o_55_));
 sg13g2_a21oi_1 _11947_ (.A1(_03768_),
    .A2(_03769_),
    .Y(csr_mtval_23_),
    .B1(net1642));
 sg13g2_and3_1 _11948_ (.X(_03770_),
    .A(crash_dump_o_118_),
    .B(crash_dump_o_119_),
    .C(_03762_));
 sg13g2_xor2_1 _11949_ (.B(_03770_),
    .A(crash_dump_o_120_),
    .X(_03771_));
 sg13g2_nand2_1 _11950_ (.Y(_03772_),
    .A(net1901),
    .B(_03771_));
 sg13g2_a22oi_1 _11951_ (.Y(_03773_),
    .B1(net1640),
    .B2(\id_stage_i.controller_i.instr_i_24_ ),
    .A2(net327),
    .A1(crash_dump_o_56_));
 sg13g2_a21oi_1 _11952_ (.A1(_03772_),
    .A2(_03773_),
    .Y(csr_mtval_24_),
    .B1(net1643));
 sg13g2_nand2_1 _11953_ (.Y(_03774_),
    .A(crash_dump_o_120_),
    .B(_03770_));
 sg13g2_xnor2_1 _11954_ (.Y(_03775_),
    .A(crash_dump_o_121_),
    .B(_03774_));
 sg13g2_nand2_1 _11955_ (.Y(_03776_),
    .A(net1899),
    .B(_03775_));
 sg13g2_a22oi_1 _11956_ (.Y(_03777_),
    .B1(net1640),
    .B2(net2006),
    .A2(net327),
    .A1(crash_dump_o_57_));
 sg13g2_a21oi_1 _11957_ (.A1(_03776_),
    .A2(_03777_),
    .Y(csr_mtval_25_),
    .B1(net1642));
 sg13g2_and3_1 _11958_ (.X(_03778_),
    .A(crash_dump_o_120_),
    .B(crash_dump_o_121_),
    .C(_03770_));
 sg13g2_xor2_1 _11959_ (.B(_03778_),
    .A(crash_dump_o_122_),
    .X(_03779_));
 sg13g2_nand2_1 _11960_ (.Y(_03780_),
    .A(net1899),
    .B(_03779_));
 sg13g2_a22oi_1 _11961_ (.Y(_03781_),
    .B1(net1640),
    .B2(\id_stage_i.controller_i.instr_i_26_ ),
    .A2(net326),
    .A1(crash_dump_o_58_));
 sg13g2_a21oi_1 _11962_ (.A1(_03780_),
    .A2(_03781_),
    .Y(csr_mtval_26_),
    .B1(_03693_));
 sg13g2_nand2_1 _11963_ (.Y(_03782_),
    .A(crash_dump_o_122_),
    .B(_03778_));
 sg13g2_xnor2_1 _11964_ (.Y(_03783_),
    .A(crash_dump_o_123_),
    .B(_03782_));
 sg13g2_nand2_1 _11965_ (.Y(_03784_),
    .A(net1899),
    .B(_03783_));
 sg13g2_a22oi_1 _11966_ (.Y(_03785_),
    .B1(net1640),
    .B2(\id_stage_i.controller_i.instr_i_27_ ),
    .A2(net326),
    .A1(crash_dump_o_59_));
 sg13g2_a21oi_2 _11967_ (.B1(net1642),
    .Y(csr_mtval_27_),
    .A2(_03785_),
    .A1(_03784_));
 sg13g2_nand3_1 _11968_ (.B(crash_dump_o_123_),
    .C(_03778_),
    .A(crash_dump_o_122_),
    .Y(_03786_));
 sg13g2_xnor2_1 _11969_ (.Y(_03787_),
    .A(crash_dump_o_124_),
    .B(_03786_));
 sg13g2_nand2_1 _11970_ (.Y(_03788_),
    .A(net1900),
    .B(_03787_));
 sg13g2_a22oi_1 _11971_ (.Y(_03789_),
    .B1(net1641),
    .B2(\id_stage_i.controller_i.instr_i_28_ ),
    .A2(net326),
    .A1(crash_dump_o_60_));
 sg13g2_a21oi_1 _11972_ (.A1(_03788_),
    .A2(_03789_),
    .Y(csr_mtval_28_),
    .B1(net1642));
 sg13g2_nor2_1 _11973_ (.A(_01284_),
    .B(_03786_),
    .Y(_03790_));
 sg13g2_xor2_1 _11974_ (.B(_03790_),
    .A(crash_dump_o_125_),
    .X(_03791_));
 sg13g2_nand2_1 _11975_ (.Y(_03792_),
    .A(net1899),
    .B(_03791_));
 sg13g2_a22oi_1 _11976_ (.Y(_03793_),
    .B1(net1640),
    .B2(\id_stage_i.controller_i.instr_i_29_ ),
    .A2(net326),
    .A1(crash_dump_o_61_));
 sg13g2_a21oi_1 _11977_ (.A1(_03792_),
    .A2(_03793_),
    .Y(csr_mtval_29_),
    .B1(net1642));
 sg13g2_nand2_1 _11978_ (.Y(_03794_),
    .A(crash_dump_o_97_),
    .B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ));
 sg13g2_xor2_1 _11979_ (.B(_03794_),
    .A(crash_dump_o_98_),
    .X(_03795_));
 sg13g2_mux2_1 _11980_ (.A0(\id_stage_i.controller_i.instr_i_2_ ),
    .A1(\id_stage_i.controller_i.instr_compressed_i_2_ ),
    .S(net438),
    .X(_03796_));
 sg13g2_a21oi_1 _11981_ (.A1(net2101),
    .A2(_03796_),
    .Y(_03797_),
    .B1(net1897));
 sg13g2_a21oi_1 _11982_ (.A1(net1903),
    .A2(_03795_),
    .Y(_03798_),
    .B1(_03797_));
 sg13g2_a21oi_1 _11983_ (.A1(crash_dump_o_34_),
    .A2(net324),
    .Y(_03799_),
    .B1(_03798_));
 sg13g2_nor2_1 _11984_ (.A(net1644),
    .B(_03799_),
    .Y(csr_mtval_2_));
 sg13g2_nand2_1 _11985_ (.Y(_03800_),
    .A(crash_dump_o_125_),
    .B(_03790_));
 sg13g2_xnor2_1 _11986_ (.Y(_03801_),
    .A(crash_dump_o_126_),
    .B(_03800_));
 sg13g2_nand2_1 _11987_ (.Y(_03802_),
    .A(net1899),
    .B(_03801_));
 sg13g2_a22oi_1 _11988_ (.Y(_03803_),
    .B1(net1640),
    .B2(net441),
    .A2(net325),
    .A1(crash_dump_o_62_));
 sg13g2_a21oi_1 _11989_ (.A1(_03802_),
    .A2(_03803_),
    .Y(csr_mtval_30_),
    .B1(net1642));
 sg13g2_nand3_1 _11990_ (.B(crash_dump_o_126_),
    .C(_03790_),
    .A(crash_dump_o_125_),
    .Y(_03804_));
 sg13g2_xnor2_1 _11991_ (.Y(_03805_),
    .A(crash_dump_o_127_),
    .B(_03804_));
 sg13g2_nand2_1 _11992_ (.Y(_03806_),
    .A(net1899),
    .B(_03805_));
 sg13g2_a22oi_1 _11993_ (.Y(_03807_),
    .B1(net1641),
    .B2(net2002),
    .A2(net325),
    .A1(crash_dump_o_63_));
 sg13g2_a21oi_1 _11994_ (.A1(_03806_),
    .A2(_03807_),
    .Y(csr_mtval_31_),
    .B1(net1642));
 sg13g2_nand2_1 _11995_ (.Y(_03808_),
    .A(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .B(_03685_));
 sg13g2_xor2_1 _11996_ (.B(_03808_),
    .A(crash_dump_o_99_),
    .X(_03809_));
 sg13g2_mux2_1 _11997_ (.A0(net1998),
    .A1(\id_stage_i.controller_i.instr_compressed_i_3_ ),
    .S(net439),
    .X(_03810_));
 sg13g2_nand3_1 _11998_ (.B(net1879),
    .C(_03810_),
    .A(net2101),
    .Y(_03811_));
 sg13g2_o21ai_1 _11999_ (.B1(_03811_),
    .Y(_03812_),
    .A1(net1880),
    .A2(_03809_));
 sg13g2_a21oi_1 _12000_ (.A1(crash_dump_o_35_),
    .A2(net324),
    .Y(_03813_),
    .B1(_03812_));
 sg13g2_nor2_1 _12001_ (.A(net1644),
    .B(_03813_),
    .Y(csr_mtval_3_));
 sg13g2_nand3_1 _12002_ (.B(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .C(_03685_),
    .A(crash_dump_o_99_),
    .Y(_03814_));
 sg13g2_xor2_1 _12003_ (.B(_03814_),
    .A(crash_dump_o_100_),
    .X(_03815_));
 sg13g2_mux2_1 _12004_ (.A0(net1997),
    .A1(\id_stage_i.controller_i.instr_compressed_i_4_ ),
    .S(net439),
    .X(_03816_));
 sg13g2_nand3_1 _12005_ (.B(net1879),
    .C(_03816_),
    .A(net2101),
    .Y(_03817_));
 sg13g2_o21ai_1 _12006_ (.B1(_03817_),
    .Y(_03818_),
    .A1(net1879),
    .A2(_03815_));
 sg13g2_a21oi_1 _12007_ (.A1(crash_dump_o_36_),
    .A2(net324),
    .Y(_03819_),
    .B1(_03818_));
 sg13g2_nor2_1 _12008_ (.A(net1644),
    .B(_03819_),
    .Y(csr_mtval_4_));
 sg13g2_xnor2_1 _12009_ (.Y(_03820_),
    .A(crash_dump_o_101_),
    .B(_03686_));
 sg13g2_mux2_1 _12010_ (.A0(net1996),
    .A1(\id_stage_i.controller_i.instr_compressed_i_5_ ),
    .S(net439),
    .X(_03821_));
 sg13g2_nand3_1 _12011_ (.B(net1879),
    .C(_03821_),
    .A(net2100),
    .Y(_03822_));
 sg13g2_o21ai_1 _12012_ (.B1(_03822_),
    .Y(_03823_),
    .A1(net1879),
    .A2(_03820_));
 sg13g2_a21oi_1 _12013_ (.A1(crash_dump_o_37_),
    .A2(net324),
    .Y(_03824_),
    .B1(_03823_));
 sg13g2_nor2_1 _12014_ (.A(net1544),
    .B(_03824_),
    .Y(csr_mtval_5_));
 sg13g2_xnor2_1 _12015_ (.Y(_03825_),
    .A(crash_dump_o_102_),
    .B(_03687_));
 sg13g2_mux2_1 _12016_ (.A0(net1995),
    .A1(\id_stage_i.controller_i.instr_compressed_i_6_ ),
    .S(net438),
    .X(_03826_));
 sg13g2_a21oi_1 _12017_ (.A1(net2100),
    .A2(_03826_),
    .Y(_03827_),
    .B1(net1897));
 sg13g2_a21oi_1 _12018_ (.A1(net1902),
    .A2(_03825_),
    .Y(_03828_),
    .B1(_03827_));
 sg13g2_a21oi_1 _12019_ (.A1(crash_dump_o_38_),
    .A2(net324),
    .Y(_03829_),
    .B1(_03828_));
 sg13g2_nor2_1 _12020_ (.A(net1644),
    .B(_03829_),
    .Y(csr_mtval_6_));
 sg13g2_nand2_1 _12021_ (.Y(_03830_),
    .A(crash_dump_o_39_),
    .B(net328));
 sg13g2_nand2_1 _12022_ (.Y(_03831_),
    .A(crash_dump_o_102_),
    .B(_03687_));
 sg13g2_xnor2_1 _12023_ (.Y(_03832_),
    .A(crash_dump_o_103_),
    .B(_03831_));
 sg13g2_mux2_1 _12024_ (.A0(net1993),
    .A1(\id_stage_i.controller_i.instr_compressed_i_7_ ),
    .S(net438),
    .X(_03833_));
 sg13g2_a22oi_1 _12025_ (.Y(_03834_),
    .B1(_03833_),
    .B2(_03682_),
    .A2(_03832_),
    .A1(net1903));
 sg13g2_a21oi_1 _12026_ (.A1(_03830_),
    .A2(_03834_),
    .Y(csr_mtval_7_),
    .B1(net1644));
 sg13g2_xnor2_1 _12027_ (.Y(_03835_),
    .A(_03200_),
    .B(_03688_));
 sg13g2_nand2_1 _12028_ (.Y(_03836_),
    .A(net440),
    .B(\id_stage_i.controller_i.instr_compressed_i_8_ ));
 sg13g2_o21ai_1 _12029_ (.B1(_03836_),
    .Y(_03837_),
    .A1(net439),
    .A2(_02333_));
 sg13g2_a21oi_1 _12030_ (.A1(net2100),
    .A2(_03837_),
    .Y(_03838_),
    .B1(net1897));
 sg13g2_a21oi_1 _12031_ (.A1(net1902),
    .A2(_03835_),
    .Y(_03839_),
    .B1(_03838_));
 sg13g2_a21oi_1 _12032_ (.A1(crash_dump_o_40_),
    .A2(net324),
    .Y(_03840_),
    .B1(_03839_));
 sg13g2_nor2_2 _12033_ (.A(net1544),
    .B(_03840_),
    .Y(csr_mtval_8_));
 sg13g2_xnor2_1 _12034_ (.Y(_03841_),
    .A(crash_dump_o_105_),
    .B(_03689_));
 sg13g2_mux2_1 _12035_ (.A0(net1992),
    .A1(\id_stage_i.controller_i.instr_compressed_i_9_ ),
    .S(net439),
    .X(_03842_));
 sg13g2_nand3_1 _12036_ (.B(net1879),
    .C(_03842_),
    .A(net2100),
    .Y(_03843_));
 sg13g2_o21ai_1 _12037_ (.B1(_03843_),
    .Y(_03844_),
    .A1(net1879),
    .A2(_03841_));
 sg13g2_a21oi_1 _12038_ (.A1(crash_dump_o_41_),
    .A2(net324),
    .Y(_03845_),
    .B1(_03844_));
 sg13g2_nor2_1 _12039_ (.A(net1644),
    .B(_03845_),
    .Y(csr_mtval_9_));
 sg13g2_nor4_1 _12040_ (.A(_01464_),
    .B(net1904),
    .C(_01468_),
    .D(_03298_),
    .Y(csr_mtvec_init));
 sg13g2_inv_2 _12041_ (.Y(csr_op_0_),
    .A(_01605_));
 sg13g2_inv_4 _12042_ (.A(_01602_),
    .Y(csr_op_1_));
 sg13g2_a21oi_2 _12043_ (.B1(_02857_),
    .Y(_03846_),
    .A2(_03184_),
    .A1(_03189_));
 sg13g2_nor2_2 _12044_ (.A(_01751_),
    .B(_03846_),
    .Y(_03847_));
 sg13g2_inv_4 _12045_ (.A(_03184_),
    .Y(_03848_));
 sg13g2_and2_2 _12046_ (.A(_01751_),
    .B(_03848_),
    .X(_03849_));
 sg13g2_nor2_2 _12047_ (.A(_03847_),
    .B(_03849_),
    .Y(_03850_));
 sg13g2_o21ai_1 _12048_ (.B1(_01635_),
    .Y(_03851_),
    .A1(_02863_),
    .A2(_03850_));
 sg13g2_inv_2 _12049_ (.Y(csr_op_en),
    .A(_03851_));
 sg13g2_nor2_2 _12050_ (.A(_03304_),
    .B(_03305_),
    .Y(csr_restore_dret_id));
 sg13g2_inv_1 _12051_ (.Y(_03852_),
    .A(_01484_));
 sg13g2_nor2_1 _12052_ (.A(_01445_),
    .B(_01447_),
    .Y(_03853_));
 sg13g2_or3_1 _12053_ (.A(_01573_),
    .B(net2103),
    .C(_03853_),
    .X(_03854_));
 sg13g2_nor2_1 _12054_ (.A(_03852_),
    .B(_03854_),
    .Y(csr_save_id));
 sg13g2_nor4_2 _12055_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_0_ ),
    .C(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .Y(_03855_),
    .D(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_B ));
 sg13g2_inv_2 _12056_ (.Y(_03856_),
    .A(_03855_));
 sg13g2_nand2_1 _12057_ (.Y(csr_save_if),
    .A(_03339_),
    .B(_03856_));
 sg13g2_and2_1 _12058_ (.A(_01456_),
    .B(_03310_),
    .X(_03857_));
 sg13g2_or3_1 _12059_ (.A(csr_save_id),
    .B(net1483),
    .C(_03857_),
    .X(csr_save_cause));
 sg13g2_nor2_2 _12060_ (.A(net549),
    .B(net2098),
    .Y(_03858_));
 sg13g2_and3_1 _12061_ (.X(_03859_),
    .A(_01161_),
    .B(net1905),
    .C(_01159_));
 sg13g2_o21ai_1 _12062_ (.B1(_03859_),
    .Y(_03860_),
    .A1(_01664_),
    .A2(_03858_));
 sg13g2_nor3_1 _12063_ (.A(\load_store_unit_i.handle_misaligned_q ),
    .B(_01373_),
    .C(_03858_),
    .Y(_03861_));
 sg13g2_a21oi_1 _12064_ (.A1(_03858_),
    .A2(net1128),
    .Y(_03862_),
    .B1(_03861_));
 sg13g2_nor2_1 _12065_ (.A(_01162_),
    .B(_03862_),
    .Y(_03863_));
 sg13g2_buf_8 fanout1035 (.A(\cs_registers_i/_1244_ ),
    .X(net1035));
 sg13g2_buf_2 fanout1034 (.A(\cs_registers_i/_1272_ ),
    .X(net1034));
 sg13g2_a22oi_1 _12068_ (.Y(_03866_),
    .B1(_03863_),
    .B2(net1113),
    .A2(_03860_),
    .A1(\data_be_o_$_MUX__Y_A ));
 sg13g2_inv_16 _12069_ (.A(_03866_),
    .Y(data_be_o_3_));
 sg13g2_buf_4 fanout1033 (.X(net1033),
    .A(\cs_registers_i/_1272_ ));
 sg13g2_o21ai_1 _12071_ (.B1(_03239_),
    .Y(_03868_),
    .A1(_01664_),
    .A2(_03858_));
 sg13g2_o21ai_1 _12072_ (.B1(_03859_),
    .Y(_03869_),
    .A1(_03858_),
    .A2(net1147));
 sg13g2_a22oi_1 _12073_ (.Y(_03870_),
    .B1(_03869_),
    .B2(_03239_),
    .A2(_03868_),
    .A1(net1147));
 sg13g2_nand2_1 _12074_ (.Y(_03871_),
    .A(\load_store_unit_i.handle_misaligned_q ),
    .B(_03860_));
 sg13g2_and2_2 _12075_ (.A(_03859_),
    .B(_03858_),
    .X(_03872_));
 sg13g2_nand2_1 _12076_ (.Y(_03873_),
    .A(net1147),
    .B(_03872_));
 sg13g2_o21ai_1 _12077_ (.B1(_03873_),
    .Y(_03874_),
    .A1(net1147),
    .A2(_03871_));
 sg13g2_nand2_1 _12078_ (.Y(_03875_),
    .A(net1113),
    .B(_03874_));
 sg13g2_o21ai_1 _12079_ (.B1(_03875_),
    .Y(data_be_o_2_),
    .A1(\load_store_unit_i.handle_misaligned_q ),
    .A2(_03870_));
 sg13g2_inv_1 _12080_ (.Y(_03876_),
    .A(\load_store_unit_i.handle_misaligned_q ));
 sg13g2_nor2_1 _12081_ (.A(_03876_),
    .B(_03872_),
    .Y(_03877_));
 sg13g2_a21oi_1 _12082_ (.A1(net1147),
    .A2(_03872_),
    .Y(_03878_),
    .B1(_03877_));
 sg13g2_nand2_1 _12083_ (.Y(_03879_),
    .A(_03239_),
    .B(_03878_));
 sg13g2_o21ai_1 _12084_ (.B1(_03879_),
    .Y(data_be_o_1_),
    .A1(_03239_),
    .A2(_03871_));
 sg13g2_mux2_2 _12085_ (.A0(_03877_),
    .A1(_03871_),
    .S(_03078_),
    .X(data_be_o_0_));
 sg13g2_nand2b_2 _12086_ (.Y(data_req_o),
    .B(_03222_),
    .A_N(_03218_));
 sg13g2_buf_4 fanout1032 (.X(net1032),
    .A(\cs_registers_i/_1286_ ));
 sg13g2_mux2_1 _12088_ (.A0(net289),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_15_ ),
    .S(net1107),
    .X(_03881_));
 sg13g2_inv_1 _12089_ (.Y(_03882_),
    .A(net1493));
 sg13g2_buf_4 fanout1031 (.X(net1031),
    .A(\cs_registers_i/_1348_ ));
 sg13g2_nand2_1 _12091_ (.Y(_03884_),
    .A(net283),
    .B(net1103));
 sg13g2_o21ai_1 _12092_ (.B1(_03884_),
    .Y(_03885_),
    .A1(_03882_),
    .A2(net1103));
 sg13g2_buf_4 fanout1030 (.X(net1030),
    .A(\cs_registers_i/_1396_ ));
 sg13g2_mux2_2 _12094_ (.A0(_03881_),
    .A1(_03885_),
    .S(net1126),
    .X(data_wdata_o_31_));
 sg13g2_nand2_1 _12095_ (.Y(_03887_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .B(net1102));
 sg13g2_o21ai_1 _12096_ (.B1(_03887_),
    .Y(_03888_),
    .A1(_01856_),
    .A2(net1102));
 sg13g2_mux2_1 _12097_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_22_ ),
    .A1(net1513),
    .S(net1108),
    .X(_03889_));
 sg13g2_mux2_2 _12098_ (.A0(_03888_),
    .A1(_03889_),
    .S(net1124),
    .X(data_wdata_o_30_));
 sg13g2_nand2_1 _12099_ (.Y(_03890_),
    .A(net1509),
    .B(net1106));
 sg13g2_o21ai_1 _12100_ (.B1(_03890_),
    .Y(_03891_),
    .A1(_02636_),
    .A2(net1106));
 sg13g2_buf_2 fanout1029 (.A(\cs_registers_i/_0738_ ),
    .X(net1029));
 sg13g2_nand2_1 _12102_ (.Y(_03893_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .B(net1105));
 sg13g2_o21ai_1 _12103_ (.B1(_03893_),
    .Y(_03894_),
    .A1(_02097_),
    .A2(net1102));
 sg13g2_mux2_2 _12104_ (.A0(_03891_),
    .A1(_03894_),
    .S(net1124),
    .X(data_wdata_o_21_));
 sg13g2_mux2_1 _12105_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ),
    .S(net1109),
    .X(_03895_));
 sg13g2_mux2_1 _12106_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .S(net1109),
    .X(_03896_));
 sg13g2_mux2_2 _12107_ (.A0(_03895_),
    .A1(_03896_),
    .S(net1127),
    .X(data_wdata_o_20_));
 sg13g2_inv_1 _12108_ (.Y(_03897_),
    .A(net1519));
 sg13g2_nand2_1 _12109_ (.Y(_03898_),
    .A(net1505),
    .B(net1104));
 sg13g2_o21ai_1 _12110_ (.B1(_03898_),
    .Y(_03899_),
    .A1(_03897_),
    .A2(net1104));
 sg13g2_nand2_1 _12111_ (.Y(_03900_),
    .A(net1499),
    .B(net1109));
 sg13g2_o21ai_1 _12112_ (.B1(_03900_),
    .Y(_03901_),
    .A1(_02478_),
    .A2(net1109));
 sg13g2_mux2_2 _12113_ (.A0(_03899_),
    .A1(_03901_),
    .S(net1125),
    .X(data_wdata_o_19_));
 sg13g2_mux2_1 _12114_ (.A0(net1514),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ),
    .S(net1108),
    .X(_03902_));
 sg13g2_nand2_1 _12115_ (.Y(_03903_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_26_ ),
    .B(net1110));
 sg13g2_o21ai_1 _12116_ (.B1(_03903_),
    .Y(_03904_),
    .A1(_02190_),
    .A2(net1110));
 sg13g2_mux2_2 _12117_ (.A0(_03902_),
    .A1(_03904_),
    .S(net1127),
    .X(data_wdata_o_18_));
 sg13g2_inv_1 _12118_ (.Y(_03905_),
    .A(net284));
 sg13g2_nand2_1 _12119_ (.Y(_03906_),
    .A(net1502),
    .B(net1107));
 sg13g2_o21ai_1 _12120_ (.B1(_03906_),
    .Y(_03907_),
    .A1(net234),
    .A2(net1107));
 sg13g2_inv_1 _12121_ (.Y(_03908_),
    .A(net1465));
 sg13g2_nand2_1 _12122_ (.Y(_03909_),
    .A(net1496),
    .B(net1104));
 sg13g2_o21ai_1 _12123_ (.B1(_03909_),
    .Y(_03910_),
    .A1(_03908_),
    .A2(net1104));
 sg13g2_mux2_2 _12124_ (.A0(_03907_),
    .A1(_03910_),
    .S(net1125),
    .X(data_wdata_o_17_));
 sg13g2_inv_2 _12125_ (.Y(_03911_),
    .A(net1470));
 sg13g2_nand2_1 _12126_ (.Y(_03912_),
    .A(net280),
    .B(net1106));
 sg13g2_o21ai_1 _12127_ (.B1(_03912_),
    .Y(_03913_),
    .A1(_03911_),
    .A2(net1106));
 sg13g2_inv_1 _12128_ (.Y(_03914_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ));
 sg13g2_nand2_1 _12129_ (.Y(_03915_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .B(net1103));
 sg13g2_o21ai_1 _12130_ (.B1(_03915_),
    .Y(_03916_),
    .A1(_03914_),
    .A2(net1103));
 sg13g2_mux2_2 _12131_ (.A0(_03913_),
    .A1(_03916_),
    .S(net1124),
    .X(data_wdata_o_16_));
 sg13g2_mux2_1 _12132_ (.A0(net1469),
    .A1(net289),
    .S(net1107),
    .X(_03917_));
 sg13g2_mux2_2 _12133_ (.A0(net283),
    .A1(net1493),
    .S(net1103),
    .X(_03918_));
 sg13g2_mux2_2 _12134_ (.A0(_03917_),
    .A1(_03918_),
    .S(net1124),
    .X(data_wdata_o_15_));
 sg13g2_inv_1 _12135_ (.Y(_03919_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ));
 sg13g2_nand2_1 _12136_ (.Y(_03920_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ),
    .B(net1102));
 sg13g2_o21ai_1 _12137_ (.B1(_03920_),
    .Y(_03921_),
    .A1(_03919_),
    .A2(net1102));
 sg13g2_mux2_1 _12138_ (.A0(net1512),
    .A1(net1491),
    .S(net1108),
    .X(_03922_));
 sg13g2_mux2_2 _12139_ (.A0(_03921_),
    .A1(_03922_),
    .S(net1124),
    .X(data_wdata_o_14_));
 sg13g2_mux2_1 _12140_ (.A0(net1509),
    .A1(net1521),
    .S(net1106),
    .X(_03923_));
 sg13g2_buf_4 fanout1028 (.X(net1028),
    .A(\cs_registers_i/_0738_ ));
 sg13g2_mux2_2 _12142_ (.A0(_03894_),
    .A1(_03923_),
    .S(net1125),
    .X(data_wdata_o_13_));
 sg13g2_mux2_1 _12143_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ),
    .S(net1109),
    .X(_03925_));
 sg13g2_mux2_2 _12144_ (.A0(_03896_),
    .A1(_03925_),
    .S(net1127),
    .X(data_wdata_o_12_));
 sg13g2_nand2_1 _12145_ (.Y(_03926_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .B(net1105));
 sg13g2_o21ai_1 _12146_ (.B1(_03926_),
    .Y(_03927_),
    .A1(_01959_),
    .A2(net1105));
 sg13g2_mux2_2 _12147_ (.A0(_03891_),
    .A1(_03927_),
    .S(net1146),
    .X(data_wdata_o_29_));
 sg13g2_nand2_1 _12148_ (.Y(_03928_),
    .A(net1519),
    .B(net1106));
 sg13g2_o21ai_1 _12149_ (.B1(_03928_),
    .Y(_03929_),
    .A1(_02283_),
    .A2(net1106));
 sg13g2_mux2_2 _12150_ (.A0(_03901_),
    .A1(_03929_),
    .S(net1125),
    .X(data_wdata_o_11_));
 sg13g2_nand2_1 _12151_ (.Y(_03930_),
    .A(net1514),
    .B(net1108));
 sg13g2_o21ai_1 _12152_ (.B1(_03930_),
    .Y(_03931_),
    .A1(_02320_),
    .A2(net1108));
 sg13g2_mux2_2 _12153_ (.A0(_03904_),
    .A1(_03931_),
    .S(net1127),
    .X(data_wdata_o_10_));
 sg13g2_inv_1 _12154_ (.Y(_03932_),
    .A(net1503));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(\cs_registers_i/_1009_ ));
 sg13g2_nand2_1 _12156_ (.Y(_03934_),
    .A(net286),
    .B(net1107));
 sg13g2_o21ai_1 _12157_ (.B1(_03934_),
    .Y(_03935_),
    .A1(net1380),
    .A2(net1107));
 sg13g2_mux2_2 _12158_ (.A0(_03910_),
    .A1(_03935_),
    .S(net1126),
    .X(data_wdata_o_9_));
 sg13g2_mux2_1 _12159_ (.A0(net280),
    .A1(net1470),
    .S(net1106),
    .X(_03936_));
 sg13g2_mux2_2 _12160_ (.A0(_03916_),
    .A1(_03936_),
    .S(net1124),
    .X(data_wdata_o_8_));
 sg13g2_mux2_2 _12161_ (.A0(_03881_),
    .A1(_03918_),
    .S(net1146),
    .X(data_wdata_o_7_));
 sg13g2_mux2_2 _12162_ (.A0(_03888_),
    .A1(_03922_),
    .S(net1146),
    .X(data_wdata_o_6_));
 sg13g2_mux2_2 _12163_ (.A0(_03923_),
    .A1(_03927_),
    .S(net1125),
    .X(data_wdata_o_5_));
 sg13g2_mux2_1 _12164_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .S(net1109),
    .X(_03937_));
 sg13g2_mux2_2 _12165_ (.A0(_03925_),
    .A1(_03937_),
    .S(net1127),
    .X(data_wdata_o_4_));
 sg13g2_mux2_1 _12166_ (.A0(net1499),
    .A1(net1468),
    .S(net1107),
    .X(_03938_));
 sg13g2_mux2_2 _12167_ (.A0(_03929_),
    .A1(_03938_),
    .S(net1126),
    .X(data_wdata_o_3_));
 sg13g2_nand2_1 _12168_ (.Y(_03939_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_10_ ),
    .B(net1112));
 sg13g2_o21ai_1 _12169_ (.B1(_03939_),
    .Y(_03940_),
    .A1(_02002_),
    .A2(net1112));
 sg13g2_mux2_2 _12170_ (.A0(_03931_),
    .A1(_03940_),
    .S(net1127),
    .X(data_wdata_o_2_));
 sg13g2_mux2_2 _12171_ (.A0(_03895_),
    .A1(_03937_),
    .S(net1146),
    .X(data_wdata_o_28_));
 sg13g2_nand2_1 _12172_ (.Y(_03941_),
    .A(net1464),
    .B(net1103));
 sg13g2_o21ai_1 _12173_ (.B1(_03941_),
    .Y(_03942_),
    .A1(_01990_),
    .A2(net1102));
 sg13g2_mux2_2 _12174_ (.A0(_03935_),
    .A1(_03942_),
    .S(net1125),
    .X(data_wdata_o_1_));
 sg13g2_nand2_1 _12175_ (.Y(_03943_),
    .A(net1463),
    .B(net1102));
 sg13g2_o21ai_1 _12176_ (.B1(_03943_),
    .Y(_03944_),
    .A1(_02058_),
    .A2(net1102));
 sg13g2_mux2_2 _12177_ (.A0(_03936_),
    .A1(_03944_),
    .S(net1124),
    .X(data_wdata_o_0_));
 sg13g2_mux2_2 _12178_ (.A0(_03899_),
    .A1(_03938_),
    .S(net1146),
    .X(data_wdata_o_27_));
 sg13g2_mux2_2 _12179_ (.A0(_03902_),
    .A1(_03940_),
    .S(net1145),
    .X(data_wdata_o_26_));
 sg13g2_mux2_2 _12180_ (.A0(_03907_),
    .A1(_03942_),
    .S(net1145),
    .X(data_wdata_o_25_));
 sg13g2_mux2_2 _12181_ (.A0(_03913_),
    .A1(_03944_),
    .S(net1145),
    .X(data_wdata_o_24_));
 sg13g2_mux2_2 _12182_ (.A0(_03885_),
    .A1(_03917_),
    .S(net1125),
    .X(data_wdata_o_23_));
 sg13g2_mux2_2 _12183_ (.A0(_03889_),
    .A1(_03921_),
    .S(net1124),
    .X(data_wdata_o_22_));
 sg13g2_nor3_2 _12184_ (.A(_01372_),
    .B(_01774_),
    .C(net1490),
    .Y(data_we_o));
 sg13g2_inv_1 _12185_ (.Y(_03945_),
    .A(debug_req_i));
 sg13g2_o21ai_1 _12186_ (.B1(_03855_),
    .Y(debug_cause_0_),
    .A1(_03945_),
    .A2(net8));
 sg13g2_o21ai_1 _12187_ (.B1(_03855_),
    .Y(_03946_),
    .A1(debug_req_i),
    .A2(net9));
 sg13g2_inv_1 _12188_ (.Y(debug_cause_1_),
    .A(_03946_));
 sg13g2_nor3_1 _12189_ (.A(debug_req_i),
    .B(net10),
    .C(_03856_),
    .Y(debug_cause_2_));
 sg13g2_a21oi_2 _12190_ (.B1(_03852_),
    .Y(debug_csr_save),
    .A2(_03854_),
    .A1(net2104));
 sg13g2_a21oi_1 _12191_ (.A1(_01463_),
    .A2(_01485_),
    .Y(_03947_),
    .B1(debug_mode));
 sg13g2_nor2_1 _12192_ (.A(csr_restore_dret_id),
    .B(_03947_),
    .Y(_00095_));
 sg13g2_nand2b_1 _12193_ (.Y(_03948_),
    .B(_01333_),
    .A_N(net2098));
 sg13g2_nand2_2 _12194_ (.Y(_03949_),
    .A(_01357_),
    .B(_03948_));
 sg13g2_nor2b_2 _12195_ (.A(_01530_),
    .B_N(_03949_),
    .Y(_03950_));
 sg13g2_and2_2 _12196_ (.A(net288),
    .B(_03950_),
    .X(_03951_));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(\cs_registers_i/_1128_ ));
 sg13g2_buf_4 fanout1025 (.X(net1025),
    .A(\cs_registers_i/_1369_ ));
 sg13g2_nand2_1 _12199_ (.Y(_03954_),
    .A(net1145),
    .B(net1454));
 sg13g2_o21ai_1 _12200_ (.B1(_03954_),
    .Y(_03955_),
    .A1(net280),
    .A2(net1454));
 sg13g2_nand3_1 _12201_ (.B(net410),
    .C(_01541_),
    .A(_01524_),
    .Y(_03956_));
 sg13g2_nor2_2 _12202_ (.A(_01568_),
    .B(net341),
    .Y(_03957_));
 sg13g2_nor3_1 _12203_ (.A(net2105),
    .B(net2111),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(_03958_));
 sg13g2_nand3_1 _12204_ (.B(_03957_),
    .C(_03958_),
    .A(net358),
    .Y(_03959_));
 sg13g2_buf_2 fanout1024 (.A(rf_wdata_wb_3_),
    .X(net1024));
 sg13g2_buf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sg13g2_buf_2 fanout1022 (.A(net1024),
    .X(net1022));
 sg13g2_nand2_1 _12208_ (.Y(_03963_),
    .A(\ex_block_i.alu_i.imd_val_q_i_0_ ),
    .B(net1228));
 sg13g2_o21ai_1 _12209_ (.B1(_03963_),
    .Y(_00096_),
    .A1(_03955_),
    .A2(net1228));
 sg13g2_nand2_1 _12210_ (.Y(_03964_),
    .A(_02895_),
    .B(net1451));
 sg13g2_o21ai_1 _12211_ (.B1(_03964_),
    .Y(_03965_),
    .A1(net258),
    .A2(net1451));
 sg13g2_nand2_1 _12212_ (.Y(_03966_),
    .A(\ex_block_i.alu_i.imd_val_q_i_10_ ),
    .B(net1225));
 sg13g2_o21ai_1 _12213_ (.B1(_03966_),
    .Y(_00097_),
    .A1(net1225),
    .A2(_03965_));
 sg13g2_nand2_2 _12214_ (.Y(_03967_),
    .A(net289),
    .B(_03950_));
 sg13g2_buf_1 fanout1021 (.A(net1022),
    .X(net1021));
 sg13g2_buf_2 fanout1020 (.A(net1022),
    .X(net1020));
 sg13g2_nand2_1 _12217_ (.Y(_03970_),
    .A(_02478_),
    .B(net1450));
 sg13g2_o21ai_1 _12218_ (.B1(_03970_),
    .Y(_03971_),
    .A1(data_addr_o_11_),
    .A2(net1450));
 sg13g2_nand2_1 _12219_ (.Y(_03972_),
    .A(\ex_block_i.alu_i.imd_val_q_i_11_ ),
    .B(net1229));
 sg13g2_o21ai_1 _12220_ (.B1(_03972_),
    .Y(_00098_),
    .A1(net1229),
    .A2(_03971_));
 sg13g2_buf_2 fanout1019 (.A(rf_wdata_wb_4_),
    .X(net1019));
 sg13g2_mux2_1 _12222_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .A1(data_addr_o_12_),
    .S(net1451),
    .X(_03974_));
 sg13g2_buf_2 fanout1018 (.A(net1019),
    .X(net1018));
 sg13g2_mux2_1 _12224_ (.A0(_03974_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_12_ ),
    .S(net1223),
    .X(_00099_));
 sg13g2_nand2_1 _12225_ (.Y(_03976_),
    .A(_02097_),
    .B(net1449));
 sg13g2_o21ai_1 _12226_ (.B1(_03976_),
    .Y(_03977_),
    .A1(data_addr_o_13_),
    .A2(net1449));
 sg13g2_nand2_1 _12227_ (.Y(_03978_),
    .A(\ex_block_i.alu_i.imd_val_q_i_13_ ),
    .B(net1227));
 sg13g2_o21ai_1 _12228_ (.B1(_03978_),
    .Y(_00100_),
    .A1(net1227),
    .A2(_03977_));
 sg13g2_nand2_1 _12229_ (.Y(_03979_),
    .A(_03265_),
    .B(net1453));
 sg13g2_o21ai_1 _12230_ (.B1(_03979_),
    .Y(_03980_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .A2(net1453));
 sg13g2_buf_2 fanout1017 (.A(net1019),
    .X(net1017));
 sg13g2_nand2_1 _12232_ (.Y(_03982_),
    .A(\ex_block_i.alu_i.imd_val_q_i_14_ ),
    .B(net1227));
 sg13g2_o21ai_1 _12233_ (.B1(_03982_),
    .Y(_00101_),
    .A1(net1227),
    .A2(_03980_));
 sg13g2_nand2b_1 _12234_ (.Y(_03983_),
    .B(net1447),
    .A_N(net1469));
 sg13g2_o21ai_1 _12235_ (.B1(_03983_),
    .Y(_03984_),
    .A1(data_addr_o_15_),
    .A2(net1447));
 sg13g2_nand2_1 _12236_ (.Y(_03985_),
    .A(\ex_block_i.alu_i.imd_val_q_i_15_ ),
    .B(net1223));
 sg13g2_o21ai_1 _12237_ (.B1(_03985_),
    .Y(_00102_),
    .A1(net1223),
    .A2(_03984_));
 sg13g2_nand2_1 _12238_ (.Y(_03986_),
    .A(_03911_),
    .B(net1450));
 sg13g2_o21ai_1 _12239_ (.B1(_03986_),
    .Y(_03987_),
    .A1(data_addr_o_16_),
    .A2(net1450));
 sg13g2_nand2_1 _12240_ (.Y(_03988_),
    .A(\ex_block_i.alu_i.imd_val_q_i_16_ ),
    .B(net1230));
 sg13g2_o21ai_1 _12241_ (.B1(_03988_),
    .Y(_00103_),
    .A1(net1230),
    .A2(_03987_));
 sg13g2_nand2_1 _12242_ (.Y(_03989_),
    .A(data_addr_o_17_),
    .B(net1455));
 sg13g2_o21ai_1 _12243_ (.B1(_03989_),
    .Y(_03990_),
    .A1(net234),
    .A2(net1455));
 sg13g2_mux2_1 _12244_ (.A0(_03990_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_17_ ),
    .S(net1230),
    .X(_00104_));
 sg13g2_mux2_1 _12245_ (.A0(net1516),
    .A1(data_addr_o_18_),
    .S(net1455),
    .X(_03991_));
 sg13g2_mux2_1 _12246_ (.A0(_03991_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_18_ ),
    .S(net1230),
    .X(_00105_));
 sg13g2_nand2_1 _12247_ (.Y(_03992_),
    .A(data_addr_o_19_),
    .B(net1455));
 sg13g2_o21ai_1 _12248_ (.B1(_03992_),
    .Y(_03993_),
    .A1(_03897_),
    .A2(net1455));
 sg13g2_mux2_1 _12249_ (.A0(_03993_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_19_ ),
    .S(net1230),
    .X(_00106_));
 sg13g2_nand2_1 _12250_ (.Y(_03994_),
    .A(net1109),
    .B(net1455));
 sg13g2_o21ai_1 _12251_ (.B1(_03994_),
    .Y(_03995_),
    .A1(net1381),
    .A2(net1455));
 sg13g2_mux2_1 _12252_ (.A0(_03995_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_1_ ),
    .S(net1230),
    .X(_00107_));
 sg13g2_nand2_1 _12253_ (.Y(_03996_),
    .A(net287),
    .B(net1449));
 sg13g2_o21ai_1 _12254_ (.B1(_03996_),
    .Y(_03997_),
    .A1(_03274_),
    .A2(net1449));
 sg13g2_mux2_1 _12255_ (.A0(_03997_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_20_ ),
    .S(net1228),
    .X(_00108_));
 sg13g2_nand2_1 _12256_ (.Y(_03998_),
    .A(data_addr_o_21_),
    .B(net1454));
 sg13g2_o21ai_1 _12257_ (.B1(_03998_),
    .Y(_03999_),
    .A1(_02636_),
    .A2(net1454));
 sg13g2_mux2_1 _12258_ (.A0(_03999_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_21_ ),
    .S(net1229),
    .X(_00109_));
 sg13g2_nand2_1 _12259_ (.Y(_04000_),
    .A(net1491),
    .B(net1450));
 sg13g2_o21ai_1 _12260_ (.B1(_04000_),
    .Y(_04001_),
    .A1(_03174_),
    .A2(net1450));
 sg13g2_mux2_1 _12261_ (.A0(_04001_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_22_ ),
    .S(net1229),
    .X(_00110_));
 sg13g2_nand2_1 _12262_ (.Y(_04002_),
    .A(_03278_),
    .B(net1452));
 sg13g2_o21ai_1 _12263_ (.B1(_04002_),
    .Y(_04003_),
    .A1(net1494),
    .A2(net1452));
 sg13g2_nand2_1 _12264_ (.Y(_04004_),
    .A(\ex_block_i.alu_i.imd_val_q_i_23_ ),
    .B(net1226));
 sg13g2_o21ai_1 _12265_ (.B1(_04004_),
    .Y(_00111_),
    .A1(net1226),
    .A2(_04003_));
 sg13g2_nand2_1 _12266_ (.Y(_04005_),
    .A(_02058_),
    .B(net1447));
 sg13g2_o21ai_1 _12267_ (.B1(_04005_),
    .Y(_04006_),
    .A1(data_addr_o_24_),
    .A2(net1447));
 sg13g2_nand2_1 _12268_ (.Y(_04007_),
    .A(\ex_block_i.alu_i.imd_val_q_i_24_ ),
    .B(net1223));
 sg13g2_o21ai_1 _12269_ (.B1(_04007_),
    .Y(_00112_),
    .A1(net1223),
    .A2(_04006_));
 sg13g2_nand2_1 _12270_ (.Y(_04008_),
    .A(_01990_),
    .B(net1448));
 sg13g2_o21ai_1 _12271_ (.B1(_04008_),
    .Y(_04009_),
    .A1(data_addr_o_25_),
    .A2(net1448));
 sg13g2_nand2_1 _12272_ (.Y(_04010_),
    .A(\ex_block_i.alu_i.imd_val_q_i_25_ ),
    .B(net1226));
 sg13g2_o21ai_1 _12273_ (.B1(_04010_),
    .Y(_00113_),
    .A1(net1226),
    .A2(_04009_));
 sg13g2_nand2_1 _12274_ (.Y(_04011_),
    .A(_03182_),
    .B(net1452));
 sg13g2_o21ai_1 _12275_ (.B1(_04011_),
    .Y(_04012_),
    .A1(net1497),
    .A2(net1452));
 sg13g2_nand2_1 _12276_ (.Y(_04013_),
    .A(\ex_block_i.alu_i.imd_val_q_i_26_ ),
    .B(net1226));
 sg13g2_o21ai_1 _12277_ (.B1(_04013_),
    .Y(_00114_),
    .A1(net1226),
    .A2(_04012_));
 sg13g2_nand2b_1 _12278_ (.Y(_04014_),
    .B(net1447),
    .A_N(net1499));
 sg13g2_o21ai_1 _12279_ (.B1(_04014_),
    .Y(_04015_),
    .A1(net2487),
    .A2(net1447));
 sg13g2_nand2_1 _12280_ (.Y(_04016_),
    .A(\ex_block_i.alu_i.imd_val_q_i_27_ ),
    .B(net1224));
 sg13g2_o21ai_1 _12281_ (.B1(_04016_),
    .Y(_00115_),
    .A1(net1224),
    .A2(_04015_));
 sg13g2_mux2_1 _12282_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .A1(data_addr_o_28_),
    .S(net1451),
    .X(_04017_));
 sg13g2_mux2_1 _12283_ (.A0(_04017_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_28_ ),
    .S(net1223),
    .X(_00116_));
 sg13g2_nand2_1 _12284_ (.Y(_04018_),
    .A(_01959_),
    .B(net1447));
 sg13g2_o21ai_1 _12285_ (.B1(_04018_),
    .Y(_04019_),
    .A1(data_addr_o_29_),
    .A2(net1447));
 sg13g2_nand2_1 _12286_ (.Y(_04020_),
    .A(\ex_block_i.alu_i.imd_val_q_i_29_ ),
    .B(net1224));
 sg13g2_o21ai_1 _12287_ (.B1(_04020_),
    .Y(_00117_),
    .A1(net1224),
    .A2(_04019_));
 sg13g2_nand2_1 _12288_ (.Y(_04021_),
    .A(data_addr_o_2_),
    .B(net1454));
 sg13g2_o21ai_1 _12289_ (.B1(_04021_),
    .Y(_04022_),
    .A1(_02320_),
    .A2(net1454));
 sg13g2_mux2_1 _12290_ (.A0(_04022_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_2_ ),
    .S(net1229),
    .X(_00118_));
 sg13g2_nand2_1 _12291_ (.Y(_04023_),
    .A(_01856_),
    .B(net1449));
 sg13g2_o21ai_1 _12292_ (.B1(_04023_),
    .Y(_04024_),
    .A1(net2494),
    .A2(net1449));
 sg13g2_nand2_1 _12293_ (.Y(_04025_),
    .A(\ex_block_i.alu_i.imd_val_q_i_30_ ),
    .B(net1229));
 sg13g2_o21ai_1 _12294_ (.B1(_04025_),
    .Y(_00119_),
    .A1(net1228),
    .A2(_04024_));
 sg13g2_inv_1 _12295_ (.Y(_04026_),
    .A(_03950_));
 sg13g2_o21ai_1 _12296_ (.B1(net288),
    .Y(_04027_),
    .A1(net36),
    .A2(_04026_));
 sg13g2_nand2_1 _12297_ (.Y(_04028_),
    .A(\ex_block_i.alu_i.imd_val_q_i_31_ ),
    .B(net1228));
 sg13g2_o21ai_1 _12298_ (.B1(_04028_),
    .Y(_00120_),
    .A1(net1228),
    .A2(_04027_));
 sg13g2_nand2_2 _12299_ (.Y(_04029_),
    .A(net410),
    .B(_01541_));
 sg13g2_nor2_2 _12300_ (.A(net2088),
    .B(_04029_),
    .Y(_04030_));
 sg13g2_buf_2 fanout1016 (.A(net1019),
    .X(net1016));
 sg13g2_nand2_2 _12302_ (.Y(_04032_),
    .A(_01569_),
    .B(net1578));
 sg13g2_or2_2 _12303_ (.X(_04033_),
    .B(_04029_),
    .A(net2093));
 sg13g2_nor2_1 _12304_ (.A(_01568_),
    .B(_04033_),
    .Y(_04034_));
 sg13g2_inv_2 _12305_ (.Y(_04035_),
    .A(_04034_));
 sg13g2_a21oi_2 _12306_ (.B1(net368),
    .Y(_04036_),
    .A2(_04035_),
    .A1(net142));
 sg13g2_buf_2 fanout1015 (.A(net1019),
    .X(net1015));
 sg13g2_buf_1 fanout1014 (.A(_04069_),
    .X(net1014));
 sg13g2_nor2_2 _12309_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ),
    .Y(_04039_));
 sg13g2_nor2_1 _12310_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ),
    .Y(_04040_));
 sg13g2_or3_1 _12311_ (.A(_01531_),
    .B(_04039_),
    .C(_04040_),
    .X(_04041_));
 sg13g2_buf_2 fanout1013 (.A(net1014),
    .X(net1013));
 sg13g2_buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sg13g2_nand2_1 _12314_ (.Y(_04044_),
    .A(net341),
    .B(net1540));
 sg13g2_a21oi_1 _12315_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .Y(_04045_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ));
 sg13g2_mux2_2 _12316_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .S(net423),
    .X(_04046_));
 sg13g2_buf_2 fanout1011 (.A(net1014),
    .X(net1011));
 sg13g2_buf_2 fanout1010 (.A(net1014),
    .X(net1010));
 sg13g2_buf_2 fanout1009 (.A(_04069_),
    .X(net1009));
 sg13g2_a21oi_2 _12320_ (.B1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .Y(_04050_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ));
 sg13g2_mux2_2 _12321_ (.A0(net280),
    .A1(net1471),
    .S(net1876),
    .X(_04051_));
 sg13g2_buf_1 fanout1008 (.A(net1009),
    .X(net1008));
 sg13g2_nand2_2 _12323_ (.Y(_04053_),
    .A(net232),
    .B(net1379));
 sg13g2_nor2_2 _12324_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ),
    .Y(_04054_));
 sg13g2_inv_1 _12325_ (.Y(_04055_),
    .A(_04054_));
 sg13g2_a21o_1 _12326_ (.A2(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .X(_04056_));
 sg13g2_buf_2 fanout1007 (.A(net1009),
    .X(net1007));
 sg13g2_buf_2 fanout1006 (.A(_04081_),
    .X(net1006));
 sg13g2_buf_4 fanout1005 (.X(net1005),
    .A(_04081_));
 sg13g2_buf_2 fanout1004 (.A(rf_wdata_wb_1_),
    .X(net1004));
 sg13g2_o21ai_1 _12331_ (.B1(net1871),
    .Y(_04061_),
    .A1(_01531_),
    .A2(_04055_));
 sg13g2_nor3_1 _12332_ (.A(_01527_),
    .B(_01530_),
    .C(_04055_),
    .Y(_04062_));
 sg13g2_a22oi_1 _12333_ (.Y(_04063_),
    .B1(net321),
    .B2(\ex_block_i.alu_i.imd_val_q_i_32_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_48_ ));
 sg13g2_xor2_1 _12334_ (.B(_04063_),
    .A(_04053_),
    .X(_04064_));
 sg13g2_nor2_1 _12335_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ),
    .B(net2110),
    .Y(_04065_));
 sg13g2_nand2b_2 _12336_ (.Y(_04066_),
    .B(_04065_),
    .A_N(net2111));
 sg13g2_o21ai_1 _12337_ (.B1(net36),
    .Y(_04067_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_31_ ),
    .A2(_01846_));
 sg13g2_nand2_1 _12338_ (.Y(_04068_),
    .A(\ex_block_i.alu_i.imd_val_q_i_31_ ),
    .B(_01846_));
 sg13g2_and2_1 _12339_ (.A(_04067_),
    .B(_04068_),
    .X(_04069_));
 sg13g2_buf_2 fanout1003 (.A(net1004),
    .X(net1003));
 sg13g2_buf_2 fanout1002 (.A(net1003),
    .X(net1002));
 sg13g2_nor2_1 _12342_ (.A(\ex_block_i.alu_i.imd_val_q_i_32_ ),
    .B(net1010),
    .Y(_04072_));
 sg13g2_a21oi_1 _12343_ (.A1(net1145),
    .A2(net1010),
    .Y(_04073_),
    .B1(_04072_));
 sg13g2_nand2_1 _12344_ (.Y(_04074_),
    .A(_01524_),
    .B(_01130_));
 sg13g2_nor2_1 _12345_ (.A(_01368_),
    .B(net549),
    .Y(_04075_));
 sg13g2_o21ai_1 _12346_ (.B1(_04075_),
    .Y(_04076_),
    .A1(net2092),
    .A2(net2095));
 sg13g2_nor3_2 _12347_ (.A(_01530_),
    .B(_04074_),
    .C(_04076_),
    .Y(_04077_));
 sg13g2_buf_2 fanout1001 (.A(net1004),
    .X(net1001));
 sg13g2_buf_2 fanout1000 (.A(net1001),
    .X(net1000));
 sg13g2_buf_8 fanout999 (.A(rf_wdata_wb_5_),
    .X(net999));
 sg13g2_nand2_2 _12351_ (.Y(_04081_),
    .A(_04067_),
    .B(_04068_));
 sg13g2_buf_16 fanout998 (.X(net998),
    .A(net999));
 sg13g2_nor3_2 _12353_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_3_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .C(net1006),
    .Y(_04083_));
 sg13g2_nor2_1 _12354_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ),
    .Y(_04084_));
 sg13g2_and2_2 _12355_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .B(_04084_),
    .X(_04085_));
 sg13g2_buf_16 fanout997 (.X(net997),
    .A(net999));
 sg13g2_a21oi_1 _12357_ (.A1(_04083_),
    .A2(_04085_),
    .Y(_04087_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_0_ ));
 sg13g2_buf_16 fanout996 (.X(net996),
    .A(net999));
 sg13g2_buf_16 fanout995 (.X(net995),
    .A(net999));
 sg13g2_nand2_1 _12360_ (.Y(_04090_),
    .A(_04087_),
    .B(net306));
 sg13g2_o21ai_1 _12361_ (.B1(_04090_),
    .Y(_04091_),
    .A1(_04073_),
    .A2(net306));
 sg13g2_buf_2 fanout994 (.A(rf_wdata_wb_7_),
    .X(net994));
 sg13g2_buf_2 fanout993 (.A(net994),
    .X(net993));
 sg13g2_buf_2 fanout992 (.A(rf_wdata_wb_7_),
    .X(net992));
 sg13g2_buf_2 fanout991 (.A(rf_wdata_wb_7_),
    .X(net991));
 sg13g2_mux4_1 _12366_ (.S0(net555),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_1_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_2_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_3_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_0_ ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .X(_04096_));
 sg13g2_mux4_1 _12367_ (.S0(net555),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_5_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_6_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_7_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_4_ ),
    .S1(net2113),
    .X(_04097_));
 sg13g2_mux4_1 _12368_ (.S0(net2113),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_9_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_11_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_10_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_8_ ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0_ ),
    .X(_04098_));
 sg13g2_mux4_1 _12369_ (.S0(net555),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_13_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_14_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_15_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_12_ ),
    .S1(net2113),
    .X(_04099_));
 sg13g2_a21oi_1 _12370_ (.A1(net554),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .Y(_04100_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ));
 sg13g2_xnor2_1 _12371_ (.Y(_04101_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .B(_04100_));
 sg13g2_nor2b_1 _12372_ (.A(_04100_),
    .B_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .Y(_04102_));
 sg13g2_nor2_1 _12373_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ),
    .B(_04102_),
    .Y(_04103_));
 sg13g2_xnor2_1 _12374_ (.Y(_04104_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_A ),
    .B(_04103_));
 sg13g2_mux4_1 _12375_ (.S0(_04101_),
    .A0(_04096_),
    .A1(_04097_),
    .A2(_04098_),
    .A3(_04099_),
    .S1(_04104_),
    .X(_04105_));
 sg13g2_mux4_1 _12376_ (.S0(net554),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_17_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_18_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_19_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_16_ ),
    .S1(net2113),
    .X(_04106_));
 sg13g2_mux4_1 _12377_ (.S0(net554),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_21_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_22_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_23_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_20_ ),
    .S1(net2113),
    .X(_04107_));
 sg13g2_mux4_1 _12378_ (.S0(net554),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_25_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_26_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_27_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_24_ ),
    .S1(net2113),
    .X(_04108_));
 sg13g2_mux4_1 _12379_ (.S0(net2113),
    .A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_29_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31_ ),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_30_ ),
    .A3(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_28_ ),
    .S1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0_ ),
    .X(_04109_));
 sg13g2_mux4_1 _12380_ (.S0(_04101_),
    .A0(_04106_),
    .A1(_04107_),
    .A2(_04108_),
    .A3(_04109_),
    .S1(_04104_),
    .X(_04110_));
 sg13g2_inv_1 _12381_ (.Y(_04111_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_A ));
 sg13g2_inv_2 _12382_ (.Y(_04112_),
    .A(net2112));
 sg13g2_o21ai_1 _12383_ (.B1(_04112_),
    .Y(_04113_),
    .A1(_04111_),
    .A2(_04103_));
 sg13g2_xor2_1 _12384_ (.B(_04113_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_A ),
    .X(_04114_));
 sg13g2_mux2_1 _12385_ (.A0(_04105_),
    .A1(_04110_),
    .S(_04114_),
    .X(_04115_));
 sg13g2_nor3_2 _12386_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ),
    .C(net2110),
    .Y(_04116_));
 sg13g2_buf_4 fanout990 (.X(net990),
    .A(\register_file_i/_2801_ ));
 sg13g2_nor2b_2 _12388_ (.A(_01530_),
    .B_N(_01658_),
    .Y(_04118_));
 sg13g2_nand2_1 _12389_ (.Y(_04119_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .B(_04118_));
 sg13g2_nand2_1 _12390_ (.Y(_04120_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_change_sign_$_AND__Y_B ),
    .B(net1448));
 sg13g2_and2_1 _12391_ (.A(net304),
    .B(_04120_),
    .X(_04121_));
 sg13g2_nand4_1 _12392_ (.B(net1453),
    .C(net304),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_change_sign_$_AND__Y_B ),
    .Y(_04122_),
    .D(net1445));
 sg13g2_o21ai_1 _12393_ (.B1(_04122_),
    .Y(_04123_),
    .A1(net1445),
    .A2(_04121_));
 sg13g2_buf_4 fanout989 (.X(net989),
    .A(net990));
 sg13g2_buf_2 fanout988 (.A(net989),
    .X(net988));
 sg13g2_nor2_1 _12396_ (.A(\ex_block_i.alu_i.imd_val_q_i_32_ ),
    .B(net1261),
    .Y(_04126_));
 sg13g2_a21oi_1 _12397_ (.A1(net1145),
    .A2(net1261),
    .Y(_04127_),
    .B1(_04126_));
 sg13g2_a21o_1 _12398_ (.A2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .A1(net2111),
    .B1(net2105),
    .X(_04128_));
 sg13g2_inv_1 _12399_ (.Y(_04129_),
    .A(net2110));
 sg13g2_nor2_1 _12400_ (.A(net2105),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Y(_04130_));
 sg13g2_nor2_1 _12401_ (.A(_04129_),
    .B(_04130_),
    .Y(_04131_));
 sg13g2_a221oi_1 _12402_ (.B2(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ),
    .C1(_04131_),
    .B1(_04128_),
    .A1(net2111),
    .Y(_04132_),
    .A2(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ));
 sg13g2_buf_4 fanout987 (.X(net987),
    .A(net989));
 sg13g2_inv_1 _12404_ (.Y(_04134_),
    .A(net1575));
 sg13g2_nor2_2 _12405_ (.A(net337),
    .B(net1478),
    .Y(_04135_));
 sg13g2_nand3_1 _12406_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31_ ),
    .C(_01535_),
    .A(net1881),
    .Y(_04136_));
 sg13g2_nor3_2 _12407_ (.A(net2107),
    .B(net2111),
    .C(net2110),
    .Y(_04137_));
 sg13g2_o21ai_1 _12408_ (.B1(net1636),
    .Y(_04138_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .A2(net305));
 sg13g2_nand3_1 _12409_ (.B(_04136_),
    .C(_04138_),
    .A(_04135_),
    .Y(_04139_));
 sg13g2_a221oi_1 _12410_ (.B2(_04127_),
    .C1(_04139_),
    .B1(net420),
    .A1(net1884),
    .Y(_04140_),
    .A2(_04115_));
 sg13g2_o21ai_1 _12411_ (.B1(_04140_),
    .Y(_04141_),
    .A1(net1708),
    .A2(_04091_));
 sg13g2_o21ai_1 _12412_ (.B1(_04141_),
    .Y(_04142_),
    .A1(_04044_),
    .A2(_04064_));
 sg13g2_nor3_1 _12413_ (.A(_01531_),
    .B(_04039_),
    .C(_04040_),
    .Y(_04143_));
 sg13g2_nor2_2 _12414_ (.A(net1578),
    .B(net298),
    .Y(_04144_));
 sg13g2_buf_8 fanout986 (.A(net990),
    .X(net986));
 sg13g2_o21ai_1 _12416_ (.B1(net1186),
    .Y(_04146_),
    .A1(_04135_),
    .A2(_04144_));
 sg13g2_a22oi_1 _12417_ (.Y(_00121_),
    .B1(_04146_),
    .B2(_02304_),
    .A2(_04142_),
    .A1(net1186));
 sg13g2_inv_2 _12418_ (.Y(_04147_),
    .A(\ex_block_i.alu_i.imd_val_q_i_33_ ));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(net986));
 sg13g2_buf_4 fanout984 (.X(net984),
    .A(\register_file_i/_2890_ ));
 sg13g2_buf_2 fanout983 (.A(net984),
    .X(net983));
 sg13g2_and2_2 _12422_ (.A(net554),
    .B(_04084_),
    .X(_04151_));
 sg13g2_buf_4 fanout982 (.X(net982),
    .A(net984));
 sg13g2_a21oi_1 _12424_ (.A1(_04083_),
    .A2(_04151_),
    .Y(_04153_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_1_ ));
 sg13g2_nand2_1 _12425_ (.Y(_04154_),
    .A(net1111),
    .B(net1011));
 sg13g2_o21ai_1 _12426_ (.B1(_04154_),
    .Y(_04155_),
    .A1(_04147_),
    .A2(net1011));
 sg13g2_nor2_1 _12427_ (.A(net308),
    .B(_04155_),
    .Y(_04156_));
 sg13g2_a21oi_1 _12428_ (.A1(net315),
    .A2(_04153_),
    .Y(_04157_),
    .B1(_04156_));
 sg13g2_nand2_1 _12429_ (.Y(_04158_),
    .A(net1890),
    .B(_04157_));
 sg13g2_buf_4 fanout981 (.X(net981),
    .A(net984));
 sg13g2_nand2_1 _12431_ (.Y(_04160_),
    .A(net1111),
    .B(net1262));
 sg13g2_o21ai_1 _12432_ (.B1(_04160_),
    .Y(_04161_),
    .A1(_04147_),
    .A2(net1262));
 sg13g2_buf_2 fanout980 (.A(net981),
    .X(net980));
 sg13g2_o21ai_1 _12434_ (.B1(net1636),
    .Y(_04163_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ),
    .A2(net305));
 sg13g2_nand3_1 _12435_ (.B(_04135_),
    .C(_04163_),
    .A(net1185),
    .Y(_04164_));
 sg13g2_a221oi_1 _12436_ (.B2(_04161_),
    .C1(_04164_),
    .B1(net420),
    .A1(net1885),
    .Y(_04165_),
    .A2(_04073_));
 sg13g2_o21ai_1 _12437_ (.B1(net358),
    .Y(_04166_),
    .A1(_03957_),
    .A2(_04034_));
 sg13g2_buf_4 fanout979 (.X(net979),
    .A(net981));
 sg13g2_buf_4 fanout978 (.X(net978),
    .A(\register_file_i/_2917_ ));
 sg13g2_nor2_1 _12440_ (.A(_04053_),
    .B(_04063_),
    .Y(_04169_));
 sg13g2_mux2_1 _12441_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ),
    .S(net423),
    .X(_04170_));
 sg13g2_buf_4 fanout977 (.X(net977),
    .A(net978));
 sg13g2_buf_4 fanout976 (.X(net976),
    .A(\register_file_i/_2917_ ));
 sg13g2_nand2_1 _12444_ (.Y(_04173_),
    .A(net1379),
    .B(net278));
 sg13g2_mux2_1 _12445_ (.A0(net285),
    .A1(net1501),
    .S(net1869),
    .X(_04174_));
 sg13g2_buf_4 fanout975 (.X(net975),
    .A(net976));
 sg13g2_nand2_1 _12447_ (.Y(_04176_),
    .A(net232),
    .B(net1440));
 sg13g2_xnor2_1 _12448_ (.Y(_04177_),
    .A(_04173_),
    .B(_04176_));
 sg13g2_buf_4 fanout974 (.X(net974),
    .A(net976));
 sg13g2_buf_4 fanout973 (.X(net973),
    .A(\register_file_i/_2921_ ));
 sg13g2_buf_4 fanout972 (.X(net972),
    .A(net973));
 sg13g2_buf_4 fanout971 (.X(net971),
    .A(net973));
 sg13g2_mux2_1 _12453_ (.A0(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .A1(\ex_block_i.alu_i.imd_val_q_i_33_ ),
    .S(_01531_),
    .X(_04182_));
 sg13g2_a22oi_1 _12454_ (.Y(_04183_),
    .B1(_04054_),
    .B2(_04182_),
    .A2(net1873),
    .A1(\ex_block_i.alu_i.imd_val_q_i_49_ ));
 sg13g2_xor2_1 _12455_ (.B(_04183_),
    .A(_04177_),
    .X(_04184_));
 sg13g2_xnor2_1 _12456_ (.Y(_04185_),
    .A(_04169_),
    .B(_04184_));
 sg13g2_buf_4 fanout970 (.X(net970),
    .A(net973));
 sg13g2_buf_4 fanout969 (.X(net969),
    .A(net970));
 sg13g2_a21oi_1 _12459_ (.A1(_04144_),
    .A2(_04185_),
    .Y(_04188_),
    .B1(net376));
 sg13g2_nor2_1 _12460_ (.A(net93),
    .B(_04188_),
    .Y(_04189_));
 sg13g2_a221oi_1 _12461_ (.B2(_04165_),
    .C1(_04189_),
    .B1(_04158_),
    .A1(_04147_),
    .Y(_00122_),
    .A2(_04146_));
 sg13g2_inv_2 _12462_ (.Y(_04190_),
    .A(\ex_block_i.alu_i.imd_val_q_i_34_ ));
 sg13g2_buf_4 fanout968 (.X(net968),
    .A(net970));
 sg13g2_nand2_1 _12464_ (.Y(_04192_),
    .A(data_addr_o_2_),
    .B(net1011));
 sg13g2_o21ai_1 _12465_ (.B1(_04192_),
    .Y(_04193_),
    .A1(_04190_),
    .A2(net1011));
 sg13g2_inv_2 _12466_ (.Y(_04194_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ));
 sg13g2_nor3_2 _12467_ (.A(net2112),
    .B(_04194_),
    .C(net1005),
    .Y(_04195_));
 sg13g2_a21oi_1 _12468_ (.A1(_04085_),
    .A2(_04195_),
    .Y(_04196_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_2_ ));
 sg13g2_nand2_1 _12469_ (.Y(_04197_),
    .A(net315),
    .B(_04196_));
 sg13g2_o21ai_1 _12470_ (.B1(_04197_),
    .Y(_04198_),
    .A1(net305),
    .A2(_04193_));
 sg13g2_nand2_1 _12471_ (.Y(_04199_),
    .A(data_addr_o_2_),
    .B(net1262));
 sg13g2_o21ai_1 _12472_ (.B1(_04199_),
    .Y(_04200_),
    .A1(_04190_),
    .A2(net1261));
 sg13g2_buf_2 fanout967 (.A(\register_file_i/_2941_ ),
    .X(net967));
 sg13g2_buf_4 fanout966 (.X(net966),
    .A(net967));
 sg13g2_o21ai_1 _12475_ (.B1(net1636),
    .Y(_04203_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ),
    .A2(net308));
 sg13g2_nand2_1 _12476_ (.Y(_04204_),
    .A(net1575),
    .B(_04203_));
 sg13g2_a221oi_1 _12477_ (.B2(net420),
    .C1(_04204_),
    .B1(_04200_),
    .A1(net1885),
    .Y(_04205_),
    .A2(_04155_));
 sg13g2_o21ai_1 _12478_ (.B1(_04205_),
    .Y(_04206_),
    .A1(net1708),
    .A2(_04198_));
 sg13g2_buf_4 fanout965 (.X(net965),
    .A(\register_file_i/_2941_ ));
 sg13g2_buf_4 fanout964 (.X(net964),
    .A(net965));
 sg13g2_nand2_1 _12481_ (.Y(_04209_),
    .A(_04177_),
    .B(_04183_));
 sg13g2_nor2_1 _12482_ (.A(_04177_),
    .B(_04183_),
    .Y(_04210_));
 sg13g2_a21o_1 _12483_ (.A2(_04209_),
    .A1(_04169_),
    .B1(_04210_),
    .X(_04211_));
 sg13g2_nor2_1 _12484_ (.A(net1380),
    .B(net1504),
    .Y(_04212_));
 sg13g2_nor2_1 _12485_ (.A(net1502),
    .B(_02320_),
    .Y(_04213_));
 sg13g2_a21oi_1 _12486_ (.A1(net276),
    .A2(_04212_),
    .Y(_04214_),
    .B1(_04213_));
 sg13g2_inv_1 _12487_ (.Y(_04215_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_inv_2 _12488_ (.Y(_04216_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ));
 sg13g2_mux2_2 _12489_ (.A0(_04215_),
    .A1(_04216_),
    .S(net423),
    .X(_04217_));
 sg13g2_mux2_2 _12490_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ),
    .S(net423),
    .X(_04218_));
 sg13g2_buf_4 fanout963 (.X(net963),
    .A(net965));
 sg13g2_and3_1 _12492_ (.X(_04220_),
    .A(net279),
    .B(net273),
    .C(_04212_));
 sg13g2_a21oi_1 _12493_ (.A1(_04217_),
    .A2(_04213_),
    .Y(_04221_),
    .B1(_04220_));
 sg13g2_o21ai_1 _12494_ (.B1(_04221_),
    .Y(_04222_),
    .A1(net279),
    .A2(_04214_));
 sg13g2_nor2_1 _12495_ (.A(net1877),
    .B(_04222_),
    .Y(_04223_));
 sg13g2_nand2_1 _12496_ (.Y(_04224_),
    .A(net234),
    .B(net1515));
 sg13g2_nor2_1 _12497_ (.A(net234),
    .B(net1514),
    .Y(_04225_));
 sg13g2_nand2_1 _12498_ (.Y(_04226_),
    .A(net276),
    .B(_04225_));
 sg13g2_a21oi_1 _12499_ (.A1(_04224_),
    .A2(_04226_),
    .Y(_04227_),
    .B1(net1470));
 sg13g2_nand3_1 _12500_ (.B(net273),
    .C(_04225_),
    .A(net1470),
    .Y(_04228_));
 sg13g2_o21ai_1 _12501_ (.B1(_04228_),
    .Y(_04229_),
    .A1(net273),
    .A2(_04224_));
 sg13g2_nor3_1 _12502_ (.A(net1870),
    .B(_04227_),
    .C(_04229_),
    .Y(_04230_));
 sg13g2_nor2b_2 _12503_ (.A(net1470),
    .B_N(net284),
    .Y(_04231_));
 sg13g2_nand3_1 _12504_ (.B(net1877),
    .C(_04231_),
    .A(net1514),
    .Y(_04232_));
 sg13g2_nor2_1 _12505_ (.A(net279),
    .B(net1380),
    .Y(_04233_));
 sg13g2_nand3_1 _12506_ (.B(net1870),
    .C(_04233_),
    .A(net1504),
    .Y(_04234_));
 sg13g2_a21oi_1 _12507_ (.A1(_04232_),
    .A2(_04234_),
    .Y(_04235_),
    .B1(net276));
 sg13g2_and2_1 _12508_ (.A(net279),
    .B(net1869),
    .X(_04236_));
 sg13g2_nor2_1 _12509_ (.A(_03911_),
    .B(net1870),
    .Y(_04237_));
 sg13g2_nor2_2 _12510_ (.A(net1477),
    .B(net1378),
    .Y(_04238_));
 sg13g2_inv_1 _12511_ (.Y(_04239_),
    .A(net1440));
 sg13g2_xor2_1 _12512_ (.B(net1514),
    .A(net284),
    .X(_04240_));
 sg13g2_xor2_1 _12513_ (.B(net1504),
    .A(net1501),
    .X(_04241_));
 sg13g2_mux2_1 _12514_ (.A0(_04240_),
    .A1(_04241_),
    .S(net1869),
    .X(_04242_));
 sg13g2_buf_2 fanout962 (.A(\register_file_i/_2947_ ),
    .X(net962));
 sg13g2_buf_4 fanout961 (.X(net961),
    .A(net962));
 sg13g2_nor4_1 _12517_ (.A(_04238_),
    .B(_04239_),
    .C(net274),
    .D(net228),
    .Y(_04245_));
 sg13g2_nor2_1 _12518_ (.A(_04235_),
    .B(_04245_),
    .Y(_04246_));
 sg13g2_o21ai_1 _12519_ (.B1(_04246_),
    .Y(_04247_),
    .A1(_04223_),
    .A2(_04230_));
 sg13g2_nand2_1 _12520_ (.Y(_04248_),
    .A(net1379),
    .B(net273));
 sg13g2_buf_4 fanout960 (.X(net960),
    .A(\register_file_i/_2947_ ));
 sg13g2_buf_4 fanout959 (.X(net959),
    .A(net960));
 sg13g2_buf_4 fanout958 (.X(net958),
    .A(net960));
 sg13g2_nor2b_1 _12524_ (.A(net427),
    .B_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .Y(_04252_));
 sg13g2_a21oi_2 _12525_ (.B1(_04252_),
    .Y(_04253_),
    .A2(net427),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ));
 sg13g2_nand2_1 _12526_ (.Y(_04254_),
    .A(net276),
    .B(net1440));
 sg13g2_inv_1 _12527_ (.Y(_04255_),
    .A(net229));
 sg13g2_a22oi_1 _12528_ (.Y(_04256_),
    .B1(_04255_),
    .B2(_04239_),
    .A2(_04254_),
    .A1(net1376));
 sg13g2_nand4_1 _12529_ (.B(net278),
    .C(net1440),
    .A(net1376),
    .Y(_04257_),
    .D(_04248_));
 sg13g2_o21ai_1 _12530_ (.B1(_04257_),
    .Y(_04258_),
    .A1(_04248_),
    .A2(_04256_));
 sg13g2_a21oi_2 _12531_ (.B1(_04258_),
    .Y(_04259_),
    .A2(_04247_),
    .A1(net232));
 sg13g2_nand2_1 _12532_ (.Y(_04260_),
    .A(\ex_block_i.alu_i.imd_val_q_i_34_ ),
    .B(_01531_));
 sg13g2_o21ai_1 _12533_ (.B1(_04260_),
    .Y(_04261_),
    .A1(_02572_),
    .A2(_01531_));
 sg13g2_a22oi_1 _12534_ (.Y(_04262_),
    .B1(_04054_),
    .B2(_04261_),
    .A2(net1873),
    .A1(\ex_block_i.alu_i.imd_val_q_i_50_ ));
 sg13g2_xor2_1 _12535_ (.B(_04262_),
    .A(_04259_),
    .X(_04263_));
 sg13g2_xnor2_1 _12536_ (.Y(_04264_),
    .A(_04211_),
    .B(_04263_));
 sg13g2_nand3_1 _12537_ (.B(net1542),
    .C(_04264_),
    .A(net342),
    .Y(_04265_));
 sg13g2_o21ai_1 _12538_ (.B1(_04265_),
    .Y(_04266_),
    .A1(net338),
    .A2(_04206_));
 sg13g2_a22oi_1 _12539_ (.Y(_00123_),
    .B1(_04266_),
    .B2(net1186),
    .A2(_04146_),
    .A1(_04190_));
 sg13g2_a21oi_1 _12540_ (.A1(_04151_),
    .A2(_04195_),
    .Y(_04267_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_3_ ));
 sg13g2_buf_2 fanout957 (.A(\register_file_i/_2952_ ),
    .X(net957));
 sg13g2_buf_4 fanout956 (.X(net956),
    .A(net957));
 sg13g2_buf_2 fanout955 (.A(\register_file_i/_2952_ ),
    .X(net955));
 sg13g2_nand2_1 _12544_ (.Y(_04271_),
    .A(data_addr_o_3_),
    .B(net1011));
 sg13g2_o21ai_1 _12545_ (.B1(_04271_),
    .Y(_04272_),
    .A1(_02280_),
    .A2(net1011));
 sg13g2_nor2_1 _12546_ (.A(net309),
    .B(_04272_),
    .Y(_04273_));
 sg13g2_a21oi_1 _12547_ (.A1(net314),
    .A2(_04267_),
    .Y(_04274_),
    .B1(_04273_));
 sg13g2_o21ai_1 _12548_ (.B1(net1638),
    .Y(_04275_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .A2(net309));
 sg13g2_buf_4 fanout954 (.X(net954),
    .A(net955));
 sg13g2_buf_2 fanout953 (.A(net955),
    .X(net953));
 sg13g2_buf_4 fanout952 (.X(net952),
    .A(net955));
 sg13g2_nand2_1 _12552_ (.Y(_04279_),
    .A(net2490),
    .B(net1262));
 sg13g2_o21ai_1 _12553_ (.B1(_04279_),
    .Y(_04280_),
    .A1(_02280_),
    .A2(net1262));
 sg13g2_nand2_1 _12554_ (.Y(_04281_),
    .A(net422),
    .B(_04280_));
 sg13g2_nand3_1 _12555_ (.B(_04275_),
    .C(_04281_),
    .A(_04135_),
    .Y(_04282_));
 sg13g2_a221oi_1 _12556_ (.B2(net1890),
    .C1(_04282_),
    .B1(_04274_),
    .A1(net1885),
    .Y(_04283_),
    .A2(_04193_));
 sg13g2_nor2_1 _12557_ (.A(_04259_),
    .B(_04262_),
    .Y(_04284_));
 sg13g2_nand2_1 _12558_ (.Y(_04285_),
    .A(_04259_),
    .B(_04262_));
 sg13g2_o21ai_1 _12559_ (.B1(_04285_),
    .Y(_04286_),
    .A1(_04211_),
    .A2(_04284_));
 sg13g2_nand2_1 _12560_ (.Y(_04287_),
    .A(net231),
    .B(net226));
 sg13g2_nand2_1 _12561_ (.Y(_04288_),
    .A(net1518),
    .B(net1877));
 sg13g2_o21ai_1 _12562_ (.B1(_04288_),
    .Y(_04289_),
    .A1(_02283_),
    .A2(net1876));
 sg13g2_buf_2 fanout951 (.A(\register_file_i/_2981_ ),
    .X(net951));
 sg13g2_buf_4 fanout950 (.X(net950),
    .A(net951));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(\register_file_i/_2981_ ));
 sg13g2_xnor2_1 _12566_ (.Y(_04293_),
    .A(net1380),
    .B(_04217_));
 sg13g2_xnor2_1 _12567_ (.Y(_04294_),
    .A(net234),
    .B(_04217_));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(net949));
 sg13g2_inv_2 _12569_ (.Y(_04296_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ));
 sg13g2_mux2_2 _12570_ (.A0(_02293_),
    .A1(_04296_),
    .S(net424),
    .X(_04297_));
 sg13g2_a21oi_1 _12571_ (.A1(_04297_),
    .A2(net1440),
    .Y(_04298_),
    .B1(net1379));
 sg13g2_a221oi_1 _12572_ (.B2(net1378),
    .C1(_04298_),
    .B1(_04294_),
    .A1(net1477),
    .Y(_04299_),
    .A2(_04293_));
 sg13g2_xnor2_1 _12573_ (.Y(_04300_),
    .A(net168),
    .B(_04299_));
 sg13g2_nor2_1 _12574_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ),
    .Y(_04301_));
 sg13g2_nor3_1 _12575_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ),
    .C(net426),
    .Y(_04302_));
 sg13g2_a21o_2 _12576_ (.A2(_04301_),
    .A1(net426),
    .B1(_04302_),
    .X(_04303_));
 sg13g2_nand3_1 _12577_ (.B(_04248_),
    .C(_04303_),
    .A(net1440),
    .Y(_04304_));
 sg13g2_o21ai_1 _12578_ (.B1(_04304_),
    .Y(_04305_),
    .A1(_04287_),
    .A2(_04300_));
 sg13g2_mux2_2 _12579_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ),
    .S(net423),
    .X(_04306_));
 sg13g2_xnor2_1 _12580_ (.Y(_04307_),
    .A(net1500),
    .B(net270));
 sg13g2_xnor2_1 _12581_ (.Y(_04308_),
    .A(net285),
    .B(net271));
 sg13g2_a21oi_1 _12582_ (.A1(net1439),
    .A2(_04217_),
    .Y(_04309_),
    .B1(net1379));
 sg13g2_a221oi_1 _12583_ (.B2(net1377),
    .C1(_04309_),
    .B1(_04308_),
    .A1(net1476),
    .Y(_04310_),
    .A2(_04307_));
 sg13g2_nand2b_1 _12584_ (.Y(_04311_),
    .B(net1518),
    .A_N(net1514));
 sg13g2_nand3b_1 _12585_ (.B(net1514),
    .C(net284),
    .Y(_04312_),
    .A_N(net1518));
 sg13g2_o21ai_1 _12586_ (.B1(_04312_),
    .Y(_04313_),
    .A1(net284),
    .A2(_04311_));
 sg13g2_nand2b_1 _12587_ (.Y(_04314_),
    .B(net1506),
    .A_N(net1504));
 sg13g2_nand3b_1 _12588_ (.B(net1504),
    .C(net1502),
    .Y(_04315_),
    .A_N(net1505));
 sg13g2_o21ai_1 _12589_ (.B1(_04315_),
    .Y(_04316_),
    .A1(net1502),
    .A2(_04314_));
 sg13g2_mux2_2 _12590_ (.A0(_04313_),
    .A1(_04316_),
    .S(net1869),
    .X(_04317_));
 sg13g2_buf_4 fanout947 (.X(net947),
    .A(net949));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(\register_file_i/_2992_ ));
 sg13g2_and2_1 _12593_ (.A(net275),
    .B(net226),
    .X(_04320_));
 sg13g2_a21o_1 _12594_ (.A2(_04317_),
    .A1(net231),
    .B1(_04320_),
    .X(_04321_));
 sg13g2_xnor2_1 _12595_ (.Y(_04322_),
    .A(_04310_),
    .B(_04321_));
 sg13g2_xor2_1 _12596_ (.B(_04322_),
    .A(_04305_),
    .X(_04323_));
 sg13g2_a22oi_1 _12597_ (.Y(_04324_),
    .B1(net321),
    .B2(\ex_block_i.alu_i.imd_val_q_i_35_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_51_ ));
 sg13g2_xor2_1 _12598_ (.B(_04324_),
    .A(_04323_),
    .X(_04325_));
 sg13g2_xnor2_1 _12599_ (.Y(_04326_),
    .A(_04286_),
    .B(_04325_));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(net946));
 sg13g2_o21ai_1 _12601_ (.B1(net1615),
    .Y(_04328_),
    .A1(_04044_),
    .A2(_04326_));
 sg13g2_or2_1 _12602_ (.X(_04329_),
    .B(_04328_),
    .A(_04283_));
 sg13g2_a22oi_1 _12603_ (.Y(_00124_),
    .B1(_04329_),
    .B2(net1186),
    .A2(_04146_),
    .A1(_02280_));
 sg13g2_inv_2 _12604_ (.Y(_04330_),
    .A(\ex_block_i.alu_i.imd_val_q_i_36_ ));
 sg13g2_nand2_1 _12605_ (.Y(_04331_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ));
 sg13g2_nor2_2 _12606_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ),
    .B(_04331_),
    .Y(_04332_));
 sg13g2_a21oi_1 _12607_ (.A1(_04083_),
    .A2(_04332_),
    .Y(_04333_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_4_ ));
 sg13g2_nand2_1 _12608_ (.Y(_04334_),
    .A(data_addr_o_4_),
    .B(net1010));
 sg13g2_o21ai_1 _12609_ (.B1(_04334_),
    .Y(_04335_),
    .A1(_04330_),
    .A2(net1010));
 sg13g2_nor2_1 _12610_ (.A(net305),
    .B(_04335_),
    .Y(_04336_));
 sg13g2_a21oi_1 _12611_ (.A1(net315),
    .A2(_04333_),
    .Y(_04337_),
    .B1(_04336_));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(net946));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(net946));
 sg13g2_nand2_1 _12614_ (.Y(_04340_),
    .A(data_addr_o_4_),
    .B(net1261));
 sg13g2_o21ai_1 _12615_ (.B1(_04340_),
    .Y(_04341_),
    .A1(_04330_),
    .A2(net1261));
 sg13g2_nand2_1 _12616_ (.Y(_04342_),
    .A(_04116_),
    .B(_04341_));
 sg13g2_o21ai_1 _12617_ (.B1(net1636),
    .Y(_04343_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ),
    .A2(net305));
 sg13g2_nand3_1 _12618_ (.B(_04342_),
    .C(_04343_),
    .A(net1569),
    .Y(_04344_));
 sg13g2_a221oi_1 _12619_ (.B2(net1890),
    .C1(_04344_),
    .B1(_04337_),
    .A1(net1884),
    .Y(_04345_),
    .A2(_04272_));
 sg13g2_buf_2 fanout942 (.A(net943),
    .X(net942));
 sg13g2_o21ai_1 _12621_ (.B1(net1579),
    .Y(_04347_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .A2(net1571));
 sg13g2_buf_4 fanout941 (.X(net941),
    .A(net943));
 sg13g2_o21ai_1 _12623_ (.B1(_04209_),
    .Y(_04349_),
    .A1(_04169_),
    .A2(_04210_));
 sg13g2_inv_1 _12624_ (.Y(_04350_),
    .A(_04349_));
 sg13g2_o21ai_1 _12625_ (.B1(_04285_),
    .Y(_04351_),
    .A1(_04284_),
    .A2(_04350_));
 sg13g2_a21o_1 _12626_ (.A2(_04351_),
    .A1(_04323_),
    .B1(_04324_),
    .X(_04352_));
 sg13g2_o21ai_1 _12627_ (.B1(_04352_),
    .Y(_04353_),
    .A1(_04323_),
    .A2(_04351_));
 sg13g2_inv_4 _12628_ (.A(net166),
    .Y(_04354_));
 sg13g2_nand4_1 _12629_ (.B(net228),
    .C(_04354_),
    .A(net232),
    .Y(_04355_),
    .D(_04299_));
 sg13g2_and2_1 _12630_ (.A(_04304_),
    .B(_04355_),
    .X(_04356_));
 sg13g2_o21ai_1 _12631_ (.B1(net168),
    .Y(_04357_),
    .A1(_04287_),
    .A2(_04299_));
 sg13g2_nand2b_1 _12632_ (.Y(_04358_),
    .B(_04322_),
    .A_N(_04357_));
 sg13g2_o21ai_1 _12633_ (.B1(_04358_),
    .Y(_04359_),
    .A1(_04322_),
    .A2(_04356_));
 sg13g2_nand2_1 _12634_ (.Y(_04360_),
    .A(net1509),
    .B(net1866));
 sg13g2_o21ai_1 _12635_ (.B1(_04360_),
    .Y(_04361_),
    .A1(_02636_),
    .A2(net1866));
 sg13g2_buf_4 fanout940 (.X(net940),
    .A(\register_file_i/_2999_ ));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(\register_file_i/_2999_ ));
 sg13g2_mux2_1 _12638_ (.A0(net167),
    .A1(_04321_),
    .S(_04310_),
    .X(_04364_));
 sg13g2_a22oi_1 _12639_ (.Y(_04365_),
    .B1(net164),
    .B2(net277),
    .A2(net227),
    .A1(net272));
 sg13g2_xnor2_1 _12640_ (.Y(_04366_),
    .A(_04364_),
    .B(_04365_));
 sg13g2_nor2b_1 _12641_ (.A(net426),
    .B_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .Y(_04367_));
 sg13g2_a21oi_2 _12642_ (.B1(_04367_),
    .Y(_04368_),
    .A2(net426),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ));
 sg13g2_mux2_2 _12643_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ),
    .S(net423),
    .X(_04369_));
 sg13g2_buf_4 fanout938 (.X(net938),
    .A(\register_file_i/_2999_ ));
 sg13g2_xnor2_1 _12645_ (.Y(_04371_),
    .A(net234),
    .B(net268));
 sg13g2_a221oi_1 _12646_ (.B2(net1470),
    .C1(net1870),
    .B1(_04371_),
    .A1(_04231_),
    .Y(_04372_),
    .A2(_04368_));
 sg13g2_xnor2_1 _12647_ (.Y(_04373_),
    .A(net1380),
    .B(net268));
 sg13g2_a221oi_1 _12648_ (.B2(net279),
    .C1(net1877),
    .B1(_04373_),
    .A1(_04233_),
    .Y(_04374_),
    .A2(_04368_));
 sg13g2_nor2_2 _12649_ (.A(_04372_),
    .B(_04374_),
    .Y(_04375_));
 sg13g2_xor2_1 _12650_ (.B(net287),
    .A(net1517),
    .X(_04376_));
 sg13g2_xor2_1 _12651_ (.B(net1507),
    .A(net1505),
    .X(_04377_));
 sg13g2_mux2_1 _12652_ (.A0(_04376_),
    .A1(_04377_),
    .S(net1867),
    .X(_04378_));
 sg13g2_buf_2 fanout937 (.A(net938),
    .X(net937));
 sg13g2_nand2_1 _12654_ (.Y(_04380_),
    .A(net231),
    .B(net222));
 sg13g2_xnor2_1 _12655_ (.Y(_04381_),
    .A(net224),
    .B(_04380_));
 sg13g2_xnor2_1 _12656_ (.Y(_04382_),
    .A(_04375_),
    .B(_04381_));
 sg13g2_xnor2_1 _12657_ (.Y(_04383_),
    .A(_04366_),
    .B(_04382_));
 sg13g2_and2_1 _12658_ (.A(net223),
    .B(_04383_),
    .X(_04384_));
 sg13g2_nor2_1 _12659_ (.A(net223),
    .B(_04383_),
    .Y(_04385_));
 sg13g2_nor2_1 _12660_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 sg13g2_xnor2_1 _12661_ (.Y(_04387_),
    .A(_04359_),
    .B(_04386_));
 sg13g2_nand2_1 _12662_ (.Y(_04388_),
    .A(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .B(net319));
 sg13g2_nand2_1 _12663_ (.Y(_04389_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .B(net303));
 sg13g2_nand3_1 _12664_ (.B(_04388_),
    .C(_04389_),
    .A(_04387_),
    .Y(_04390_));
 sg13g2_a21o_1 _12665_ (.A2(_04389_),
    .A1(_04388_),
    .B1(_04387_),
    .X(_04391_));
 sg13g2_nand2_1 _12666_ (.Y(_04392_),
    .A(_04390_),
    .B(_04391_));
 sg13g2_xnor2_1 _12667_ (.Y(_04393_),
    .A(_04353_),
    .B(_04392_));
 sg13g2_nand2_1 _12668_ (.Y(_04394_),
    .A(net1541),
    .B(_04393_));
 sg13g2_o21ai_1 _12669_ (.B1(_04394_),
    .Y(_04395_),
    .A1(_04330_),
    .A2(net1541));
 sg13g2_nand2_2 _12670_ (.Y(_04396_),
    .A(net342),
    .B(_04395_));
 sg13g2_o21ai_1 _12671_ (.B1(_04396_),
    .Y(_04397_),
    .A1(_04345_),
    .A2(_04347_));
 sg13g2_nand3_1 _12672_ (.B(net1185),
    .C(_04397_),
    .A(net1615),
    .Y(_04398_));
 sg13g2_o21ai_1 _12673_ (.B1(_04398_),
    .Y(_00125_),
    .A1(_04330_),
    .A2(net1185));
 sg13g2_inv_1 _12674_ (.Y(_04399_),
    .A(\ex_block_i.alu_i.imd_val_q_i_37_ ));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(net938));
 sg13g2_nor2_2 _12676_ (.A(net367),
    .B(net1576),
    .Y(_04401_));
 sg13g2_buf_2 fanout935 (.A(\register_file_i/_3003_ ),
    .X(net935));
 sg13g2_buf_2 fanout934 (.A(net935),
    .X(net934));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(net935));
 sg13g2_buf_4 fanout932 (.X(net932),
    .A(net935));
 sg13g2_buf_2 fanout931 (.A(net932),
    .X(net931));
 sg13g2_inv_1 _12682_ (.Y(_04407_),
    .A(_04324_));
 sg13g2_a21oi_1 _12683_ (.A1(_04211_),
    .A2(_04285_),
    .Y(_04408_),
    .B1(_04284_));
 sg13g2_nor2_1 _12684_ (.A(_04323_),
    .B(_04408_),
    .Y(_04409_));
 sg13g2_nand2_1 _12685_ (.Y(_04410_),
    .A(_04323_),
    .B(_04408_));
 sg13g2_o21ai_1 _12686_ (.B1(_04410_),
    .Y(_04411_),
    .A1(_04407_),
    .A2(_04409_));
 sg13g2_inv_1 _12687_ (.Y(_04412_),
    .A(_04390_));
 sg13g2_a21oi_1 _12688_ (.A1(_04391_),
    .A2(_04411_),
    .Y(_04413_),
    .B1(_04412_));
 sg13g2_a22oi_1 _12689_ (.Y(_04414_),
    .B1(net321),
    .B2(\ex_block_i.alu_i.imd_val_q_i_37_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_53_ ));
 sg13g2_inv_2 _12690_ (.Y(_04415_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ));
 sg13g2_inv_1 _12691_ (.Y(_04416_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ));
 sg13g2_mux2_2 _12692_ (.A0(_04415_),
    .A1(_04416_),
    .S(net424),
    .X(_04417_));
 sg13g2_xnor2_1 _12693_ (.Y(_04418_),
    .A(net1500),
    .B(_04417_));
 sg13g2_xnor2_1 _12694_ (.Y(_04419_),
    .A(net286),
    .B(_04417_));
 sg13g2_nand2b_1 _12695_ (.Y(_04420_),
    .B(net1501),
    .A_N(net279));
 sg13g2_nor2_1 _12696_ (.A(net1876),
    .B(_04420_),
    .Y(_04421_));
 sg13g2_a21oi_2 _12697_ (.B1(_04421_),
    .Y(_04422_),
    .A2(_04231_),
    .A1(net1877));
 sg13g2_nor2_1 _12698_ (.A(net267),
    .B(_04422_),
    .Y(_04423_));
 sg13g2_a221oi_1 _12699_ (.B2(net1377),
    .C1(_04423_),
    .B1(_04419_),
    .A1(net1477),
    .Y(_04424_),
    .A2(_04418_));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(net932));
 sg13g2_and2_1 _12701_ (.A(net226),
    .B(net270),
    .X(_04426_));
 sg13g2_a21o_1 _12702_ (.A2(net165),
    .A1(_04218_),
    .B1(_04426_),
    .X(_04427_));
 sg13g2_xnor2_1 _12703_ (.Y(_04428_),
    .A(net1505),
    .B(net1509));
 sg13g2_xor2_1 _12704_ (.B(net1521),
    .A(net1518),
    .X(_04429_));
 sg13g2_nor2_1 _12705_ (.A(net1867),
    .B(_04429_),
    .Y(_04430_));
 sg13g2_a21oi_2 _12706_ (.B1(_04430_),
    .Y(_04431_),
    .A2(_04428_),
    .A1(net1867));
 sg13g2_nand2b_1 _12707_ (.Y(_04432_),
    .B(net1520),
    .A_N(net287));
 sg13g2_nand3b_1 _12708_ (.B(net287),
    .C(net1517),
    .Y(_04433_),
    .A_N(net1520));
 sg13g2_o21ai_1 _12709_ (.B1(_04433_),
    .Y(_04434_),
    .A1(net1517),
    .A2(_04432_));
 sg13g2_nand2b_1 _12710_ (.Y(_04435_),
    .B(net1509),
    .A_N(net1507));
 sg13g2_nand3b_1 _12711_ (.B(net1507),
    .C(net1505),
    .Y(_04436_),
    .A_N(net1508));
 sg13g2_o21ai_1 _12712_ (.B1(_04436_),
    .Y(_04437_),
    .A1(net1505),
    .A2(_04435_));
 sg13g2_mux2_2 _12713_ (.A0(_04434_),
    .A1(_04437_),
    .S(net1867),
    .X(_04438_));
 sg13g2_buf_4 fanout929 (.X(net929),
    .A(\register_file_i/_3007_ ));
 sg13g2_and2_1 _12715_ (.A(net275),
    .B(net222),
    .X(_04440_));
 sg13g2_a21o_1 _12716_ (.A2(_04438_),
    .A1(net230),
    .B1(_04440_),
    .X(_04441_));
 sg13g2_xnor2_1 _12717_ (.Y(_04442_),
    .A(net1341),
    .B(_04441_));
 sg13g2_xnor2_1 _12718_ (.Y(_04443_),
    .A(_04427_),
    .B(_04442_));
 sg13g2_xnor2_1 _12719_ (.Y(_04444_),
    .A(_04424_),
    .B(_04443_));
 sg13g2_xor2_1 _12720_ (.B(_04380_),
    .A(net223),
    .X(_04445_));
 sg13g2_nand2b_1 _12721_ (.Y(_04446_),
    .B(_04365_),
    .A_N(_04310_));
 sg13g2_o21ai_1 _12722_ (.B1(net226),
    .Y(_04447_),
    .A1(net275),
    .A2(net273));
 sg13g2_nand2b_1 _12723_ (.Y(_04448_),
    .B(net164),
    .A_N(_04303_));
 sg13g2_a21oi_1 _12724_ (.A1(_04447_),
    .A2(_04448_),
    .Y(_04449_),
    .B1(net166));
 sg13g2_or2_1 _12725_ (.X(_04450_),
    .B(_04365_),
    .A(_04310_));
 sg13g2_nand3_1 _12726_ (.B(net273),
    .C(net226),
    .A(net277),
    .Y(_04451_));
 sg13g2_nand3_1 _12727_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ),
    .C(net425),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .Y(_04452_));
 sg13g2_nand3b_1 _12728_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .Y(_04453_),
    .A_N(net424));
 sg13g2_nand3_1 _12729_ (.B(_04452_),
    .C(_04453_),
    .A(_04297_),
    .Y(_04454_));
 sg13g2_a21o_1 _12730_ (.A2(net277),
    .A1(net230),
    .B1(net227),
    .X(_04455_));
 sg13g2_nand3_1 _12731_ (.B(_04454_),
    .C(_04455_),
    .A(net164),
    .Y(_04456_));
 sg13g2_and3_1 _12732_ (.X(_04457_),
    .A(net166),
    .B(_04451_),
    .C(_04456_));
 sg13g2_a22oi_1 _12733_ (.Y(_04458_),
    .B1(_04450_),
    .B2(_04457_),
    .A2(_04449_),
    .A1(_04446_));
 sg13g2_or2_1 _12734_ (.X(_04459_),
    .B(_04374_),
    .A(_04372_));
 sg13g2_o21ai_1 _12735_ (.B1(_04459_),
    .Y(_04460_),
    .A1(_04445_),
    .A2(_04458_));
 sg13g2_nand2_1 _12736_ (.Y(_04461_),
    .A(_04445_),
    .B(_04458_));
 sg13g2_a21oi_1 _12737_ (.A1(net230),
    .A2(net164),
    .Y(_04462_),
    .B1(_04320_));
 sg13g2_nor3_1 _12738_ (.A(net166),
    .B(_04462_),
    .C(_04365_),
    .Y(_04463_));
 sg13g2_and3_1 _12739_ (.X(_04464_),
    .A(net166),
    .B(_04462_),
    .C(_04365_));
 sg13g2_o21ai_1 _12740_ (.B1(_04310_),
    .Y(_04465_),
    .A1(_04463_),
    .A2(_04464_));
 sg13g2_inv_1 _12741_ (.Y(_04466_),
    .A(_04465_));
 sg13g2_a21oi_1 _12742_ (.A1(_04460_),
    .A2(_04461_),
    .Y(_04467_),
    .B1(_04466_));
 sg13g2_or3_1 _12743_ (.A(_04459_),
    .B(_04445_),
    .C(_04465_),
    .X(_04468_));
 sg13g2_inv_1 _12744_ (.Y(_04469_),
    .A(_04468_));
 sg13g2_or3_1 _12745_ (.A(_04444_),
    .B(_04467_),
    .C(_04469_),
    .X(_04470_));
 sg13g2_o21ai_1 _12746_ (.B1(_04444_),
    .Y(_04471_),
    .A1(_04467_),
    .A2(_04469_));
 sg13g2_and2_1 _12747_ (.A(_04470_),
    .B(_04471_),
    .X(_04472_));
 sg13g2_nor3_1 _12748_ (.A(_04304_),
    .B(_04322_),
    .C(_04355_),
    .Y(_04473_));
 sg13g2_inv_1 _12749_ (.Y(_04474_),
    .A(_04473_));
 sg13g2_nor2_1 _12750_ (.A(_04359_),
    .B(_04384_),
    .Y(_04475_));
 sg13g2_a21oi_1 _12751_ (.A1(_04385_),
    .A2(_04474_),
    .Y(_04476_),
    .B1(_04475_));
 sg13g2_xnor2_1 _12752_ (.Y(_04477_),
    .A(_04472_),
    .B(_04476_));
 sg13g2_xor2_1 _12753_ (.B(_04477_),
    .A(_04414_),
    .X(_04478_));
 sg13g2_xnor2_1 _12754_ (.Y(_04479_),
    .A(_04413_),
    .B(_04478_));
 sg13g2_nor2_1 _12755_ (.A(net298),
    .B(_04479_),
    .Y(_04480_));
 sg13g2_a21oi_1 _12756_ (.A1(_04399_),
    .A2(net300),
    .Y(_04481_),
    .B1(_04480_));
 sg13g2_nand2_1 _12757_ (.Y(_04482_),
    .A(net1184),
    .B(_04481_));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(net929));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(\register_file_i/_3007_ ));
 sg13g2_buf_2 fanout926 (.A(net927),
    .X(net926));
 sg13g2_inv_1 _12761_ (.Y(_04486_),
    .A(net554));
 sg13g2_inv_1 _12762_ (.Y(_04487_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ));
 sg13g2_nor3_2 _12763_ (.A(_04486_),
    .B(_04487_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ),
    .Y(_04488_));
 sg13g2_nand2_1 _12764_ (.Y(_04489_),
    .A(net1009),
    .B(_04488_));
 sg13g2_nor3_1 _12765_ (.A(net2112),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .C(_04489_),
    .Y(_04490_));
 sg13g2_nor2_1 _12766_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_5_ ),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_nand2_1 _12767_ (.Y(_04492_),
    .A(data_addr_o_5_),
    .B(net1013));
 sg13g2_o21ai_1 _12768_ (.B1(_04492_),
    .Y(_04493_),
    .A1(_04399_),
    .A2(net1013));
 sg13g2_nor2_1 _12769_ (.A(net307),
    .B(_04493_),
    .Y(_04494_));
 sg13g2_a21oi_1 _12770_ (.A1(net314),
    .A2(_04491_),
    .Y(_04495_),
    .B1(_04494_));
 sg13g2_buf_4 fanout925 (.X(net925),
    .A(net927));
 sg13g2_nand2_1 _12772_ (.Y(_04497_),
    .A(data_addr_o_5_),
    .B(net1263));
 sg13g2_o21ai_1 _12773_ (.B1(_04497_),
    .Y(_04498_),
    .A1(_04399_),
    .A2(net1263));
 sg13g2_nand2_1 _12774_ (.Y(_04499_),
    .A(net421),
    .B(_04498_));
 sg13g2_buf_4 fanout924 (.X(net924),
    .A(\register_file_i/_3012_ ));
 sg13g2_o21ai_1 _12776_ (.B1(net1635),
    .Y(_04501_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ),
    .A2(net311));
 sg13g2_nand3_1 _12777_ (.B(_04499_),
    .C(_04501_),
    .A(net1570),
    .Y(_04502_));
 sg13g2_a221oi_1 _12778_ (.B2(net1889),
    .C1(_04502_),
    .B1(_04495_),
    .A1(net1886),
    .Y(_04503_),
    .A2(_04335_));
 sg13g2_buf_2 fanout923 (.A(net924),
    .X(net923));
 sg13g2_o21ai_1 _12780_ (.B1(net1189),
    .Y(_04505_),
    .A1(net339),
    .A2(_04503_));
 sg13g2_o21ai_1 _12781_ (.B1(_04505_),
    .Y(_04506_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_37_ ),
    .A2(net1573));
 sg13g2_a22oi_1 _12782_ (.Y(_00126_),
    .B1(_04482_),
    .B2(_04506_),
    .A2(net97),
    .A1(_04399_));
 sg13g2_inv_2 _12783_ (.Y(_04507_),
    .A(\ex_block_i.alu_i.imd_val_q_i_38_ ));
 sg13g2_nor2b_1 _12784_ (.A(_04477_),
    .B_N(_04414_),
    .Y(_04508_));
 sg13g2_a21oi_1 _12785_ (.A1(_04323_),
    .A2(_04408_),
    .Y(_04509_),
    .B1(_04324_));
 sg13g2_o21ai_1 _12786_ (.B1(_04390_),
    .Y(_04510_),
    .A1(_04409_),
    .A2(_04509_));
 sg13g2_and2_1 _12787_ (.A(_04391_),
    .B(_04510_),
    .X(_04511_));
 sg13g2_nand2b_1 _12788_ (.Y(_04512_),
    .B(_04477_),
    .A_N(_04414_));
 sg13g2_o21ai_1 _12789_ (.B1(_04512_),
    .Y(_04513_),
    .A1(_04508_),
    .A2(_04511_));
 sg13g2_buf_4 fanout922 (.X(net922),
    .A(net924));
 sg13g2_a22oi_1 _12791_ (.Y(_04515_),
    .B1(net321),
    .B2(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .A2(net302),
    .A1(\ex_block_i.alu_i.imd_val_q_i_54_ ));
 sg13g2_a21oi_1 _12792_ (.A1(_04445_),
    .A2(_04458_),
    .Y(_04516_),
    .B1(_04459_));
 sg13g2_o21ai_1 _12793_ (.B1(_04465_),
    .Y(_04517_),
    .A1(_04445_),
    .A2(_04458_));
 sg13g2_o21ai_1 _12794_ (.B1(_04444_),
    .Y(_04518_),
    .A1(_04516_),
    .A2(_04517_));
 sg13g2_and2_2 _12795_ (.A(_04468_),
    .B(_04518_),
    .X(_04519_));
 sg13g2_buf_8 fanout921 (.A(\register_file_i/_3012_ ),
    .X(net921));
 sg13g2_xor2_1 _12797_ (.B(net1491),
    .A(net1520),
    .X(_04521_));
 sg13g2_xor2_1 _12798_ (.B(net1512),
    .A(net1508),
    .X(_04522_));
 sg13g2_mux2_1 _12799_ (.A0(_04521_),
    .A1(_04522_),
    .S(net1871),
    .X(_04523_));
 sg13g2_buf_4 fanout920 (.X(net920),
    .A(net921));
 sg13g2_buf_4 fanout919 (.X(net919),
    .A(\register_file_i/_3017_ ));
 sg13g2_and2_1 _12802_ (.A(net233),
    .B(net219),
    .X(_04526_));
 sg13g2_mux2_2 _12803_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ),
    .S(net423),
    .X(_04527_));
 sg13g2_buf_2 fanout918 (.A(net919),
    .X(net918));
 sg13g2_xnor2_1 _12805_ (.Y(_04529_),
    .A(net1500),
    .B(net1475));
 sg13g2_xnor2_1 _12806_ (.Y(_04530_),
    .A(net286),
    .B(net1475));
 sg13g2_a21oi_1 _12807_ (.A1(net1439),
    .A2(_04417_),
    .Y(_04531_),
    .B1(_04051_));
 sg13g2_a221oi_1 _12808_ (.B2(net1377),
    .C1(_04531_),
    .B1(_04530_),
    .A1(net1476),
    .Y(_04532_),
    .A2(_04529_));
 sg13g2_inv_1 _12809_ (.Y(_04533_),
    .A(_04532_));
 sg13g2_and2_1 _12810_ (.A(net226),
    .B(net267),
    .X(_04534_));
 sg13g2_a21o_1 _12811_ (.A2(net165),
    .A1(net271),
    .B1(_04534_),
    .X(_04535_));
 sg13g2_buf_4 fanout917 (.X(net917),
    .A(net919));
 sg13g2_and2_1 _12813_ (.A(net272),
    .B(net222),
    .X(_04537_));
 sg13g2_a21o_1 _12814_ (.A2(net163),
    .A1(net277),
    .B1(_04537_),
    .X(_04538_));
 sg13g2_xor2_1 _12815_ (.B(_04538_),
    .A(net1341),
    .X(_04539_));
 sg13g2_xnor2_1 _12816_ (.Y(_04540_),
    .A(_04535_),
    .B(_04539_));
 sg13g2_xnor2_1 _12817_ (.Y(_04541_),
    .A(_04533_),
    .B(_04540_));
 sg13g2_xnor2_1 _12818_ (.Y(_04542_),
    .A(net223),
    .B(_04441_));
 sg13g2_xnor2_1 _12819_ (.Y(_04543_),
    .A(net167),
    .B(_04427_));
 sg13g2_o21ai_1 _12820_ (.B1(_04543_),
    .Y(_04544_),
    .A1(_04424_),
    .A2(_04542_));
 sg13g2_nand2_1 _12821_ (.Y(_04545_),
    .A(_04424_),
    .B(_04542_));
 sg13g2_and2_2 _12822_ (.A(_04544_),
    .B(_04545_),
    .X(_04546_));
 sg13g2_xnor2_1 _12823_ (.Y(_04547_),
    .A(net52),
    .B(_04546_));
 sg13g2_xnor2_1 _12824_ (.Y(_04548_),
    .A(net1222),
    .B(_04547_));
 sg13g2_xnor2_1 _12825_ (.Y(_04549_),
    .A(_04519_),
    .B(_04548_));
 sg13g2_inv_1 _12826_ (.Y(_04550_),
    .A(_04472_));
 sg13g2_nand2_1 _12827_ (.Y(_04551_),
    .A(net225),
    .B(_04383_));
 sg13g2_nor2_1 _12828_ (.A(_04551_),
    .B(_04474_),
    .Y(_04552_));
 sg13g2_o21ai_1 _12829_ (.B1(_04476_),
    .Y(_04553_),
    .A1(_04550_),
    .A2(_04552_));
 sg13g2_xnor2_1 _12830_ (.Y(_04554_),
    .A(_04549_),
    .B(_04553_));
 sg13g2_nor2_1 _12831_ (.A(_04515_),
    .B(_04554_),
    .Y(_04555_));
 sg13g2_nand2_1 _12832_ (.Y(_04556_),
    .A(_04515_),
    .B(_04554_));
 sg13g2_nand2b_1 _12833_ (.Y(_04557_),
    .B(_04556_),
    .A_N(_04555_));
 sg13g2_xnor2_1 _12834_ (.Y(_04558_),
    .A(_04513_),
    .B(_04557_));
 sg13g2_nand2_1 _12835_ (.Y(_04559_),
    .A(net1542),
    .B(_04558_));
 sg13g2_o21ai_1 _12836_ (.B1(_04559_),
    .Y(_04560_),
    .A1(_04507_),
    .A2(net1542));
 sg13g2_nand2_1 _12837_ (.Y(_04561_),
    .A(net1184),
    .B(_04560_));
 sg13g2_a21oi_1 _12838_ (.A1(_04195_),
    .A2(_04332_),
    .Y(_04562_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_6_ ));
 sg13g2_nand2_1 _12839_ (.Y(_04563_),
    .A(data_addr_o_6_),
    .B(net1013));
 sg13g2_o21ai_1 _12840_ (.B1(_04563_),
    .Y(_04564_),
    .A1(_04507_),
    .A2(net1013));
 sg13g2_nor2_1 _12841_ (.A(net307),
    .B(_04564_),
    .Y(_04565_));
 sg13g2_a21oi_1 _12842_ (.A1(net314),
    .A2(_04562_),
    .Y(_04566_),
    .B1(_04565_));
 sg13g2_nand2_1 _12843_ (.Y(_04567_),
    .A(data_addr_o_6_),
    .B(net1263));
 sg13g2_o21ai_1 _12844_ (.B1(_04567_),
    .Y(_04568_),
    .A1(_04507_),
    .A2(net1263));
 sg13g2_nand2_1 _12845_ (.Y(_04569_),
    .A(net421),
    .B(_04568_));
 sg13g2_o21ai_1 _12846_ (.B1(net1637),
    .Y(_04570_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ),
    .A2(net311));
 sg13g2_nand3_1 _12847_ (.B(_04569_),
    .C(_04570_),
    .A(net1570),
    .Y(_04571_));
 sg13g2_a221oi_1 _12848_ (.B2(net1889),
    .C1(_04571_),
    .B1(_04566_),
    .A1(net1886),
    .Y(_04572_),
    .A2(_04493_));
 sg13g2_o21ai_1 _12849_ (.B1(net1187),
    .Y(_04573_),
    .A1(net339),
    .A2(_04572_));
 sg13g2_o21ai_1 _12850_ (.B1(_04573_),
    .Y(_04574_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .A2(net1573));
 sg13g2_a22oi_1 _12851_ (.Y(_00127_),
    .B1(_04561_),
    .B2(_04574_),
    .A2(net97),
    .A1(_04507_));
 sg13g2_a21oi_1 _12852_ (.A1(_04512_),
    .A2(_04511_),
    .Y(_04575_),
    .B1(_04508_));
 sg13g2_o21ai_1 _12853_ (.B1(_04556_),
    .Y(_04576_),
    .A1(_04555_),
    .A2(_04575_));
 sg13g2_nor2b_1 _12854_ (.A(_04472_),
    .B_N(_04476_),
    .Y(_04577_));
 sg13g2_inv_1 _12855_ (.Y(_04578_),
    .A(_04549_));
 sg13g2_o21ai_1 _12856_ (.B1(_04578_),
    .Y(_04579_),
    .A1(_04577_),
    .A2(_04552_));
 sg13g2_nand2_1 _12857_ (.Y(_04580_),
    .A(_04468_),
    .B(_04518_));
 sg13g2_buf_4 fanout916 (.X(net916),
    .A(\register_file_i/_3017_ ));
 sg13g2_buf_4 fanout915 (.X(net915),
    .A(net916));
 sg13g2_nand2b_1 _12860_ (.Y(_04583_),
    .B(net281),
    .A_N(net1512));
 sg13g2_nand3b_1 _12861_ (.B(net1512),
    .C(net1508),
    .Y(_04584_),
    .A_N(net281));
 sg13g2_o21ai_1 _12862_ (.B1(_04584_),
    .Y(_04585_),
    .A1(net1508),
    .A2(_04583_));
 sg13g2_nand2b_1 _12863_ (.Y(_04586_),
    .B(net1492),
    .A_N(net1491));
 sg13g2_nand3b_1 _12864_ (.B(net1491),
    .C(net1520),
    .Y(_04587_),
    .A_N(net1492));
 sg13g2_o21ai_1 _12865_ (.B1(_04587_),
    .Y(_04588_),
    .A1(net1520),
    .A2(_04586_));
 sg13g2_mux2_2 _12866_ (.A0(_04585_),
    .A1(_04588_),
    .S(net1872),
    .X(_04589_));
 sg13g2_buf_4 fanout914 (.X(net914),
    .A(net915));
 sg13g2_buf_4 fanout913 (.X(net913),
    .A(\register_file_i/_3021_ ));
 sg13g2_nand2_1 _12869_ (.Y(_04592_),
    .A(net283),
    .B(net1866));
 sg13g2_o21ai_1 _12870_ (.B1(_04592_),
    .Y(_04593_),
    .A1(_03882_),
    .A2(net1866));
 sg13g2_buf_2 fanout912 (.A(net913),
    .X(net912));
 sg13g2_nand2_1 _12872_ (.Y(_04595_),
    .A(net217),
    .B(net156));
 sg13g2_nor3_1 _12873_ (.A(net276),
    .B(net161),
    .C(_04595_),
    .Y(_04596_));
 sg13g2_a21oi_1 _12874_ (.A1(net161),
    .A2(_04595_),
    .Y(_04597_),
    .B1(_04596_));
 sg13g2_nand2_2 _12875_ (.Y(_04598_),
    .A(net275),
    .B(net219));
 sg13g2_a21o_1 _12876_ (.A2(net159),
    .A1(net231),
    .B1(_04598_),
    .X(_04599_));
 sg13g2_o21ai_1 _12877_ (.B1(_04599_),
    .Y(_04600_),
    .A1(_04253_),
    .A2(_04597_));
 sg13g2_buf_4 fanout911 (.X(net911),
    .A(net913));
 sg13g2_xnor2_1 _12879_ (.Y(_04602_),
    .A(net223),
    .B(_04538_));
 sg13g2_xnor2_1 _12880_ (.Y(_04603_),
    .A(net167),
    .B(_04535_));
 sg13g2_o21ai_1 _12881_ (.B1(_04533_),
    .Y(_04604_),
    .A1(_04602_),
    .A2(_04603_));
 sg13g2_nand2_1 _12882_ (.Y(_04605_),
    .A(_04602_),
    .B(_04603_));
 sg13g2_and2_1 _12883_ (.A(_04604_),
    .B(_04605_),
    .X(_04606_));
 sg13g2_nand2_1 _12884_ (.Y(_04607_),
    .A(net280),
    .B(net1870));
 sg13g2_mux2_2 _12885_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ),
    .S(net424),
    .X(_04608_));
 sg13g2_buf_8 fanout910 (.A(\register_file_i/_3021_ ),
    .X(net910));
 sg13g2_xnor2_1 _12887_ (.Y(_04610_),
    .A(net1381),
    .B(net266));
 sg13g2_xnor2_1 _12888_ (.Y(_04611_),
    .A(net285),
    .B(net266));
 sg13g2_nand2b_1 _12889_ (.Y(_04612_),
    .B(net1440),
    .A_N(net1475));
 sg13g2_a22oi_1 _12890_ (.Y(_04613_),
    .B1(_04612_),
    .B2(_04238_),
    .A2(_04611_),
    .A1(net1378));
 sg13g2_o21ai_1 _12891_ (.B1(_04613_),
    .Y(_04614_),
    .A1(_04607_),
    .A2(_04610_));
 sg13g2_buf_4 fanout909 (.X(net909),
    .A(net910));
 sg13g2_a22oi_1 _12893_ (.Y(_04616_),
    .B1(net162),
    .B2(_04218_),
    .A2(net220),
    .A1(net270));
 sg13g2_nand2_1 _12894_ (.Y(_04617_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ),
    .B(net424));
 sg13g2_o21ai_1 _12895_ (.B1(_04617_),
    .Y(_04618_),
    .A1(_04415_),
    .A2(net424));
 sg13g2_a22oi_1 _12896_ (.Y(_04619_),
    .B1(net253),
    .B2(net227),
    .A2(net268),
    .A1(net164));
 sg13g2_xor2_1 _12897_ (.B(_04619_),
    .A(net1341),
    .X(_04620_));
 sg13g2_xnor2_1 _12898_ (.Y(_04621_),
    .A(_04616_),
    .B(_04620_));
 sg13g2_xnor2_1 _12899_ (.Y(_04622_),
    .A(_04614_),
    .B(_04621_));
 sg13g2_xnor2_1 _12900_ (.Y(_04623_),
    .A(_04606_),
    .B(_04622_));
 sg13g2_xnor2_1 _12901_ (.Y(_04624_),
    .A(_04600_),
    .B(_04623_));
 sg13g2_nand3_1 _12902_ (.B(net52),
    .C(net1123),
    .A(net1222),
    .Y(_04625_));
 sg13g2_nand2_2 _12903_ (.Y(_04626_),
    .A(_04544_),
    .B(_04545_));
 sg13g2_nor2_2 _12904_ (.A(net51),
    .B(_04626_),
    .Y(_04627_));
 sg13g2_xor2_1 _12905_ (.B(_04623_),
    .A(_04600_),
    .X(_04628_));
 sg13g2_nand3_1 _12906_ (.B(_04627_),
    .C(_04628_),
    .A(net1222),
    .Y(_04629_));
 sg13g2_nand3_1 _12907_ (.B(_04625_),
    .C(_04629_),
    .A(_04580_),
    .Y(_04630_));
 sg13g2_nand2_2 _12908_ (.Y(_04631_),
    .A(net231),
    .B(net217));
 sg13g2_a21oi_2 _12909_ (.B1(_04424_),
    .Y(_04632_),
    .A2(_04542_),
    .A1(_04543_));
 sg13g2_inv_1 _12910_ (.Y(_04633_),
    .A(_04632_));
 sg13g2_or2_1 _12911_ (.X(_04634_),
    .B(_04542_),
    .A(_04543_));
 sg13g2_a221oi_1 _12912_ (.B2(_04634_),
    .C1(_04628_),
    .B1(_04633_),
    .A1(_04631_),
    .Y(_04635_),
    .A2(net52));
 sg13g2_xnor2_1 _12913_ (.Y(_04636_),
    .A(_04532_),
    .B(_04540_));
 sg13g2_nand3_1 _12914_ (.B(_04636_),
    .C(net1123),
    .A(_04526_),
    .Y(_04637_));
 sg13g2_nand3b_1 _12915_ (.B(_04637_),
    .C(_04519_),
    .Y(_04638_),
    .A_N(_04635_));
 sg13g2_nor2_1 _12916_ (.A(_04543_),
    .B(_04542_),
    .Y(_04639_));
 sg13g2_nor2_2 _12917_ (.A(_04632_),
    .B(_04639_),
    .Y(_04640_));
 sg13g2_nor2_1 _12918_ (.A(net52),
    .B(_04640_),
    .Y(_04641_));
 sg13g2_o21ai_1 _12919_ (.B1(_04519_),
    .Y(_04642_),
    .A1(net1123),
    .A2(_04641_));
 sg13g2_and2_1 _12920_ (.A(net51),
    .B(_04640_),
    .X(_04643_));
 sg13g2_nor3_1 _12921_ (.A(_04519_),
    .B(net1123),
    .C(_04643_),
    .Y(_04644_));
 sg13g2_a221oi_1 _12922_ (.B2(_04643_),
    .C1(_04644_),
    .B1(net1123),
    .A1(net232),
    .Y(_04645_),
    .A2(net219));
 sg13g2_nand3_1 _12923_ (.B(_04580_),
    .C(net1123),
    .A(net1222),
    .Y(_04646_));
 sg13g2_nand3_1 _12924_ (.B(net51),
    .C(_04628_),
    .A(_04519_),
    .Y(_04647_));
 sg13g2_a21oi_1 _12925_ (.A1(_04646_),
    .A2(_04647_),
    .Y(_04648_),
    .B1(_04546_));
 sg13g2_a221oi_1 _12926_ (.B2(_04645_),
    .C1(_04648_),
    .B1(_04642_),
    .A1(_04630_),
    .Y(_04649_),
    .A2(_04638_));
 sg13g2_xor2_1 _12927_ (.B(_04649_),
    .A(_04579_),
    .X(_04650_));
 sg13g2_buf_4 fanout908 (.X(net908),
    .A(\register_file_i/_3026_ ));
 sg13g2_a22oi_1 _12929_ (.Y(_04652_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .A2(net302),
    .A1(\ex_block_i.alu_i.imd_val_q_i_55_ ));
 sg13g2_nor2b_1 _12930_ (.A(_04650_),
    .B_N(_04652_),
    .Y(_04653_));
 sg13g2_nand2b_1 _12931_ (.Y(_04654_),
    .B(_04650_),
    .A_N(_04652_));
 sg13g2_nor2b_1 _12932_ (.A(_04653_),
    .B_N(_04654_),
    .Y(_04655_));
 sg13g2_xor2_1 _12933_ (.B(_04655_),
    .A(_04576_),
    .X(_04656_));
 sg13g2_nor2_1 _12934_ (.A(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .B(net1542),
    .Y(_04657_));
 sg13g2_a21oi_1 _12935_ (.A1(net1543),
    .A2(_04656_),
    .Y(_04658_),
    .B1(_04657_));
 sg13g2_nand2_1 _12936_ (.Y(_04659_),
    .A(net1184),
    .B(_04658_));
 sg13g2_buf_4 fanout907 (.X(net907),
    .A(net908));
 sg13g2_a21oi_1 _12938_ (.A1(_04195_),
    .A2(_04488_),
    .Y(_04661_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_7_ ));
 sg13g2_buf_4 fanout906 (.X(net906),
    .A(net907));
 sg13g2_nand2_1 _12940_ (.Y(_04663_),
    .A(data_addr_o_7_),
    .B(net1013));
 sg13g2_o21ai_1 _12941_ (.B1(_04663_),
    .Y(_04664_),
    .A1(_02204_),
    .A2(net1012));
 sg13g2_nor2_1 _12942_ (.A(net307),
    .B(_04664_),
    .Y(_04665_));
 sg13g2_a21oi_1 _12943_ (.A1(net316),
    .A2(_04661_),
    .Y(_04666_),
    .B1(_04665_));
 sg13g2_buf_8 fanout905 (.A(\register_file_i/_3026_ ),
    .X(net905));
 sg13g2_nand2_1 _12945_ (.Y(_04668_),
    .A(data_addr_o_7_),
    .B(net1264));
 sg13g2_o21ai_1 _12946_ (.B1(_04668_),
    .Y(_04669_),
    .A1(_02204_),
    .A2(net1263));
 sg13g2_nand2_1 _12947_ (.Y(_04670_),
    .A(net421),
    .B(_04669_));
 sg13g2_o21ai_1 _12948_ (.B1(net1637),
    .Y(_04671_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ),
    .A2(net310));
 sg13g2_nand3_1 _12949_ (.B(_04670_),
    .C(_04671_),
    .A(net1574),
    .Y(_04672_));
 sg13g2_a221oi_1 _12950_ (.B2(net1889),
    .C1(_04672_),
    .B1(_04666_),
    .A1(net1886),
    .Y(_04673_),
    .A2(_04564_));
 sg13g2_o21ai_1 _12951_ (.B1(net1189),
    .Y(_04674_),
    .A1(net339),
    .A2(_04673_));
 sg13g2_o21ai_1 _12952_ (.B1(_04674_),
    .Y(_04675_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .A2(net1572));
 sg13g2_a22oi_1 _12953_ (.Y(_00128_),
    .B1(_04659_),
    .B2(_04675_),
    .A2(net97),
    .A1(_02204_));
 sg13g2_nand2_1 _12954_ (.Y(_04676_),
    .A(net2490),
    .B(net1454));
 sg13g2_o21ai_1 _12955_ (.B1(_04676_),
    .Y(_04677_),
    .A1(_02283_),
    .A2(net1454));
 sg13g2_mux2_1 _12956_ (.A0(_04677_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_3_ ),
    .S(net1229),
    .X(_00129_));
 sg13g2_inv_1 _12957_ (.Y(_04678_),
    .A(\ex_block_i.alu_i.imd_val_q_i_40_ ));
 sg13g2_a21oi_2 _12958_ (.B1(_04653_),
    .Y(_04679_),
    .A2(_04654_),
    .A1(_04576_));
 sg13g2_xnor2_1 _12959_ (.Y(_04680_),
    .A(_04526_),
    .B(_04546_));
 sg13g2_nand2_1 _12960_ (.Y(_04681_),
    .A(_04631_),
    .B(_04626_));
 sg13g2_mux2_1 _12961_ (.A0(_04680_),
    .A1(_04681_),
    .S(_04636_),
    .X(_04682_));
 sg13g2_nor2_1 _12962_ (.A(_04624_),
    .B(_04682_),
    .Y(_04683_));
 sg13g2_nor4_1 _12963_ (.A(_04631_),
    .B(net51),
    .C(_04626_),
    .D(_04628_),
    .Y(_04684_));
 sg13g2_xnor2_1 _12964_ (.Y(_04685_),
    .A(net168),
    .B(_04365_));
 sg13g2_nand3_1 _12965_ (.B(_04381_),
    .C(_04685_),
    .A(_04375_),
    .Y(_04686_));
 sg13g2_nand3_1 _12966_ (.B(_04445_),
    .C(_04685_),
    .A(_04459_),
    .Y(_04687_));
 sg13g2_o21ai_1 _12967_ (.B1(_04687_),
    .Y(_04688_),
    .A1(_04382_),
    .A2(_04685_));
 sg13g2_nand2_1 _12968_ (.Y(_04689_),
    .A(_04444_),
    .B(_04688_));
 sg13g2_o21ai_1 _12969_ (.B1(_04689_),
    .Y(_04690_),
    .A1(_04444_),
    .A2(_04686_));
 sg13g2_xnor2_1 _12970_ (.Y(_04691_),
    .A(net168),
    .B(_04462_));
 sg13g2_and3_1 _12971_ (.X(_04692_),
    .A(_04310_),
    .B(_04690_),
    .C(_04691_));
 sg13g2_o21ai_1 _12972_ (.B1(_04692_),
    .Y(_04693_),
    .A1(_04683_),
    .A2(_04684_));
 sg13g2_o21ai_1 _12973_ (.B1(_04693_),
    .Y(_04694_),
    .A1(_04579_),
    .A2(_04649_));
 sg13g2_o21ai_1 _12974_ (.B1(_04375_),
    .Y(_04695_),
    .A1(_04381_),
    .A2(_04685_));
 sg13g2_nand2_1 _12975_ (.Y(_04696_),
    .A(_04381_),
    .B(_04685_));
 sg13g2_nand2_1 _12976_ (.Y(_04697_),
    .A(_04695_),
    .B(_04696_));
 sg13g2_and2_1 _12977_ (.A(_04444_),
    .B(_04697_),
    .X(_04698_));
 sg13g2_a21oi_1 _12978_ (.A1(_04444_),
    .A2(_04697_),
    .Y(_04699_),
    .B1(_04636_));
 sg13g2_a21oi_1 _12979_ (.A1(_04640_),
    .A2(_04699_),
    .Y(_04700_),
    .B1(_04641_));
 sg13g2_a22oi_1 _12980_ (.Y(_04701_),
    .B1(_04700_),
    .B2(net1222),
    .A2(_04698_),
    .A1(_04547_));
 sg13g2_nand4_1 _12981_ (.B(_04627_),
    .C(net1123),
    .A(net1222),
    .Y(_04702_),
    .D(_04698_));
 sg13g2_o21ai_1 _12982_ (.B1(_04702_),
    .Y(_04703_),
    .A1(net1123),
    .A2(_04701_));
 sg13g2_mux2_2 _12983_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ),
    .S(net424),
    .X(_04704_));
 sg13g2_xnor2_1 _12984_ (.Y(_04705_),
    .A(net1381),
    .B(net251));
 sg13g2_xnor2_1 _12985_ (.Y(_04706_),
    .A(net285),
    .B(net251));
 sg13g2_nand2b_1 _12986_ (.Y(_04707_),
    .B(net1439),
    .A_N(net264));
 sg13g2_a22oi_1 _12987_ (.Y(_04708_),
    .B1(_04707_),
    .B2(_04238_),
    .A2(_04706_),
    .A1(net1378));
 sg13g2_o21ai_1 _12988_ (.B1(_04708_),
    .Y(_04709_),
    .A1(_04607_),
    .A2(_04705_));
 sg13g2_a22oi_1 _12989_ (.Y(_04710_),
    .B1(net1475),
    .B2(net227),
    .A2(net254),
    .A1(net164));
 sg13g2_a22oi_1 _12990_ (.Y(_04711_),
    .B1(net162),
    .B2(net271),
    .A2(net220),
    .A1(net267));
 sg13g2_xor2_1 _12991_ (.B(_04711_),
    .A(net1341),
    .X(_04712_));
 sg13g2_xnor2_1 _12992_ (.Y(_04713_),
    .A(_04710_),
    .B(_04712_));
 sg13g2_xnor2_1 _12993_ (.Y(_04714_),
    .A(_04709_),
    .B(_04713_));
 sg13g2_xnor2_1 _12994_ (.Y(_04715_),
    .A(net224),
    .B(_04616_));
 sg13g2_xnor2_1 _12995_ (.Y(_04716_),
    .A(net167),
    .B(_04619_));
 sg13g2_nor2_1 _12996_ (.A(_04715_),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_nand2_1 _12997_ (.Y(_04718_),
    .A(_04715_),
    .B(_04716_));
 sg13g2_o21ai_1 _12998_ (.B1(_04718_),
    .Y(_04719_),
    .A1(_04614_),
    .A2(_04717_));
 sg13g2_xor2_1 _12999_ (.B(_04719_),
    .A(_04714_),
    .X(_04720_));
 sg13g2_and2_1 _13000_ (.A(net272),
    .B(net217),
    .X(_04721_));
 sg13g2_a21o_2 _13001_ (.A2(_04589_),
    .A1(net277),
    .B1(_04721_),
    .X(_04722_));
 sg13g2_xor2_1 _13002_ (.B(net1463),
    .A(net281),
    .X(_04723_));
 sg13g2_xor2_1 _13003_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .A(net1492),
    .X(_04724_));
 sg13g2_mux2_2 _13004_ (.A0(_04723_),
    .A1(_04724_),
    .S(net1875),
    .X(_04725_));
 sg13g2_inv_4 _13005_ (.A(net1339),
    .Y(_04726_));
 sg13g2_nor2_2 _13006_ (.A(net1376),
    .B(_04726_),
    .Y(_04727_));
 sg13g2_a21oi_1 _13007_ (.A1(net1376),
    .A2(_04598_),
    .Y(_04728_),
    .B1(_04727_));
 sg13g2_buf_4 fanout904 (.X(net904),
    .A(net905));
 sg13g2_nor3_1 _13009_ (.A(net1520),
    .B(net1491),
    .C(net1493),
    .Y(_04730_));
 sg13g2_nand3_1 _13010_ (.B(net1491),
    .C(net1492),
    .A(net1520),
    .Y(_04731_));
 sg13g2_nand2b_1 _13011_ (.Y(_04732_),
    .B(_04731_),
    .A_N(_04730_));
 sg13g2_or3_1 _13012_ (.A(net1508),
    .B(net1512),
    .C(net281),
    .X(_04733_));
 sg13g2_nand3_1 _13013_ (.B(net1512),
    .C(net282),
    .A(net1508),
    .Y(_04734_));
 sg13g2_nand3_1 _13014_ (.B(_04733_),
    .C(_04734_),
    .A(net1866),
    .Y(_04735_));
 sg13g2_o21ai_1 _13015_ (.B1(_04735_),
    .Y(_04736_),
    .A1(net1866),
    .A2(_04732_));
 sg13g2_nand2_1 _13016_ (.Y(_04737_),
    .A(net157),
    .B(_04736_));
 sg13g2_mux2_1 _13017_ (.A0(_04728_),
    .A1(_04727_),
    .S(_04737_),
    .X(_04738_));
 sg13g2_xnor2_1 _13018_ (.Y(_04739_),
    .A(_04722_),
    .B(_04738_));
 sg13g2_xnor2_1 _13019_ (.Y(_04740_),
    .A(_04720_),
    .B(_04739_));
 sg13g2_a21o_1 _13020_ (.A2(_04603_),
    .A1(_04533_),
    .B1(_04602_),
    .X(_04741_));
 sg13g2_o21ai_1 _13021_ (.B1(_04741_),
    .Y(_04742_),
    .A1(_04533_),
    .A2(_04603_));
 sg13g2_a22oi_1 _13022_ (.Y(_04743_),
    .B1(_04600_),
    .B2(_04742_),
    .A2(_04546_),
    .A1(_04636_));
 sg13g2_nor2_1 _13023_ (.A(_04600_),
    .B(_04742_),
    .Y(_04744_));
 sg13g2_o21ai_1 _13024_ (.B1(_04622_),
    .Y(_04745_),
    .A1(_04743_),
    .A2(_04744_));
 sg13g2_nand2_2 _13025_ (.Y(_04746_),
    .A(_04604_),
    .B(_04605_));
 sg13g2_nor2_1 _13026_ (.A(_04746_),
    .B(_04622_),
    .Y(_04747_));
 sg13g2_nand3_1 _13027_ (.B(_04600_),
    .C(_04747_),
    .A(_04627_),
    .Y(_04748_));
 sg13g2_or3_1 _13028_ (.A(_04627_),
    .B(_04600_),
    .C(_04606_),
    .X(_04749_));
 sg13g2_nand3_1 _13029_ (.B(_04748_),
    .C(_04749_),
    .A(_04745_),
    .Y(_04750_));
 sg13g2_xor2_1 _13030_ (.B(_04750_),
    .A(_04740_),
    .X(_04751_));
 sg13g2_xor2_1 _13031_ (.B(_04751_),
    .A(_04703_),
    .X(_04752_));
 sg13g2_xnor2_1 _13032_ (.Y(_04753_),
    .A(_04694_),
    .B(_04752_));
 sg13g2_a22oi_1 _13033_ (.Y(_04754_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .A2(net302),
    .A1(net556));
 sg13g2_xor2_1 _13034_ (.B(_04754_),
    .A(_04753_),
    .X(_04755_));
 sg13g2_xor2_1 _13035_ (.B(_04755_),
    .A(_04679_),
    .X(_04756_));
 sg13g2_nor2_1 _13036_ (.A(net298),
    .B(_04756_),
    .Y(_04757_));
 sg13g2_a21oi_1 _13037_ (.A1(_04678_),
    .A2(net300),
    .Y(_04758_),
    .B1(_04757_));
 sg13g2_nand2_1 _13038_ (.Y(_04759_),
    .A(net1184),
    .B(_04758_));
 sg13g2_nand2_2 _13039_ (.Y(_04760_),
    .A(net2112),
    .B(_04194_));
 sg13g2_nor2_2 _13040_ (.A(net1006),
    .B(_04760_),
    .Y(_04761_));
 sg13g2_a21oi_1 _13041_ (.A1(_04085_),
    .A2(_04761_),
    .Y(_04762_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_8_ ));
 sg13g2_mux2_1 _13042_ (.A0(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .A1(data_addr_o_8_),
    .S(net1013),
    .X(_04763_));
 sg13g2_nor2_1 _13043_ (.A(net307),
    .B(_04763_),
    .Y(_04764_));
 sg13g2_a21oi_1 _13044_ (.A1(net316),
    .A2(_04762_),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nor2_1 _13045_ (.A(net1445),
    .B(_04121_),
    .Y(_04766_));
 sg13g2_nor2b_1 _13046_ (.A(_04766_),
    .B_N(_04122_),
    .Y(_04767_));
 sg13g2_buf_4 fanout903 (.X(net903),
    .A(\register_file_i/_3030_ ));
 sg13g2_buf_4 fanout902 (.X(net902),
    .A(net903));
 sg13g2_nor2_1 _13049_ (.A(data_addr_o_8_),
    .B(net1221),
    .Y(_04770_));
 sg13g2_a21oi_1 _13050_ (.A1(_04678_),
    .A2(net1220),
    .Y(_04771_),
    .B1(_04770_));
 sg13g2_nand2_1 _13051_ (.Y(_04772_),
    .A(net421),
    .B(_04771_));
 sg13g2_buf_8 fanout901 (.A(\register_file_i/_3030_ ),
    .X(net901));
 sg13g2_o21ai_1 _13053_ (.B1(net1639),
    .Y(_04774_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ),
    .A2(net310));
 sg13g2_nand3_1 _13054_ (.B(_04772_),
    .C(_04774_),
    .A(net1573),
    .Y(_04775_));
 sg13g2_a221oi_1 _13055_ (.B2(net1890),
    .C1(_04775_),
    .B1(_04765_),
    .A1(net1887),
    .Y(_04776_),
    .A2(_04664_));
 sg13g2_o21ai_1 _13056_ (.B1(net1189),
    .Y(_04777_),
    .A1(net339),
    .A2(_04776_));
 sg13g2_o21ai_1 _13057_ (.B1(_04777_),
    .Y(_04778_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .A2(net1572));
 sg13g2_a22oi_1 _13058_ (.Y(_00130_),
    .B1(_04759_),
    .B2(_04778_),
    .A2(net96),
    .A1(_04678_));
 sg13g2_inv_1 _13059_ (.Y(_04779_),
    .A(\ex_block_i.alu_i.imd_val_q_i_41_ ));
 sg13g2_nor2_1 _13060_ (.A(_04753_),
    .B(_04754_),
    .Y(_04780_));
 sg13g2_nor2_1 _13061_ (.A(_04679_),
    .B(_04780_),
    .Y(_04781_));
 sg13g2_a21oi_2 _13062_ (.B1(_04781_),
    .Y(_04782_),
    .A2(_04754_),
    .A1(_04753_));
 sg13g2_a22oi_1 _13063_ (.Y(_04783_),
    .B1(net322),
    .B2(net2115),
    .A2(net302),
    .A1(\ex_block_i.alu_i.imd_val_q_i_57_ ));
 sg13g2_a21oi_2 _13064_ (.B1(_04717_),
    .Y(_04784_),
    .A2(_04718_),
    .A1(_04614_));
 sg13g2_nand2b_1 _13065_ (.Y(_04785_),
    .B(_04784_),
    .A_N(_04714_));
 sg13g2_mux2_2 _13066_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ),
    .S(net423),
    .X(_04786_));
 sg13g2_buf_2 fanout900 (.A(net901),
    .X(net900));
 sg13g2_xnor2_1 _13068_ (.Y(_04788_),
    .A(net1500),
    .B(net1438));
 sg13g2_xnor2_1 _13069_ (.Y(_04789_),
    .A(net285),
    .B(net1438));
 sg13g2_nor2_1 _13070_ (.A(_02175_),
    .B(net427),
    .Y(_04790_));
 sg13g2_a21oi_2 _13071_ (.B1(_04790_),
    .Y(_04791_),
    .A2(net426),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ));
 sg13g2_a21oi_1 _13072_ (.A1(net1439),
    .A2(_04791_),
    .Y(_04792_),
    .B1(_04051_));
 sg13g2_a221oi_1 _13073_ (.B2(net1378),
    .C1(_04792_),
    .B1(_04789_),
    .A1(net1477),
    .Y(_04793_),
    .A2(_04788_));
 sg13g2_buf_4 fanout899 (.X(net899),
    .A(net901));
 sg13g2_a22oi_1 _13075_ (.Y(_04795_),
    .B1(net162),
    .B2(net269),
    .A2(net254),
    .A1(net222));
 sg13g2_a22oi_1 _13076_ (.Y(_04796_),
    .B1(net264),
    .B2(net227),
    .A2(net1475),
    .A1(net164));
 sg13g2_xnor2_1 _13077_ (.Y(_04797_),
    .A(net1342),
    .B(_04796_));
 sg13g2_xnor2_1 _13078_ (.Y(_04798_),
    .A(_04795_),
    .B(_04797_));
 sg13g2_xnor2_1 _13079_ (.Y(_04799_),
    .A(_04793_),
    .B(_04798_));
 sg13g2_xnor2_1 _13080_ (.Y(_04800_),
    .A(net167),
    .B(_04710_));
 sg13g2_xnor2_1 _13081_ (.Y(_04801_),
    .A(net224),
    .B(_04711_));
 sg13g2_nor2_1 _13082_ (.A(_04800_),
    .B(_04801_),
    .Y(_04802_));
 sg13g2_nand2_1 _13083_ (.Y(_04803_),
    .A(_04800_),
    .B(_04801_));
 sg13g2_o21ai_1 _13084_ (.B1(_04803_),
    .Y(_04804_),
    .A1(_04709_),
    .A2(_04802_));
 sg13g2_xor2_1 _13085_ (.B(_04804_),
    .A(_04799_),
    .X(_04805_));
 sg13g2_nand2_1 _13086_ (.Y(_04806_),
    .A(net1496),
    .B(net1874));
 sg13g2_o21ai_1 _13087_ (.B1(_04806_),
    .Y(_04807_),
    .A1(_03908_),
    .A2(net1874));
 sg13g2_buf_4 fanout898 (.X(net898),
    .A(\register_file_i/_3034_ ));
 sg13g2_xnor2_1 _13089_ (.Y(_04809_),
    .A(_04722_),
    .B(net1338));
 sg13g2_nor2_1 _13090_ (.A(net157),
    .B(_04727_),
    .Y(_04810_));
 sg13g2_a21oi_1 _13091_ (.A1(_04727_),
    .A2(_04809_),
    .Y(_04811_),
    .B1(_04810_));
 sg13g2_and2_1 _13092_ (.A(net270),
    .B(net217),
    .X(_04812_));
 sg13g2_a21o_1 _13093_ (.A2(net161),
    .A1(net274),
    .B1(_04812_),
    .X(_04813_));
 sg13g2_nand2b_1 _13094_ (.Y(_04814_),
    .B(net1465),
    .A_N(net1463));
 sg13g2_nand3b_1 _13095_ (.B(net1463),
    .C(net282),
    .Y(_04815_),
    .A_N(net1465));
 sg13g2_o21ai_1 _13096_ (.B1(_04815_),
    .Y(_04816_),
    .A1(net281),
    .A2(_04814_));
 sg13g2_nand2b_1 _13097_ (.Y(_04817_),
    .B(net1495),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ));
 sg13g2_nand3b_1 _13098_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .C(net1492),
    .Y(_04818_),
    .A_N(net1495));
 sg13g2_o21ai_1 _13099_ (.B1(_04818_),
    .Y(_04819_),
    .A1(net1492),
    .A2(_04817_));
 sg13g2_mux2_1 _13100_ (.A0(_04816_),
    .A1(_04819_),
    .S(net1873),
    .X(_04820_));
 sg13g2_nand2_1 _13101_ (.Y(_04821_),
    .A(net230),
    .B(net139));
 sg13g2_o21ai_1 _13102_ (.B1(_04821_),
    .Y(_04822_),
    .A1(_04297_),
    .A2(_04726_));
 sg13g2_xor2_1 _13103_ (.B(_04822_),
    .A(_04813_),
    .X(_04823_));
 sg13g2_xnor2_1 _13104_ (.Y(_04824_),
    .A(_04811_),
    .B(_04823_));
 sg13g2_inv_1 _13105_ (.Y(_04825_),
    .A(_04824_));
 sg13g2_xnor2_1 _13106_ (.Y(_04826_),
    .A(_04805_),
    .B(_04825_));
 sg13g2_xnor2_1 _13107_ (.Y(_04827_),
    .A(_04785_),
    .B(_04826_));
 sg13g2_buf_4 fanout897 (.X(net897),
    .A(net898));
 sg13g2_a21oi_2 _13109_ (.B1(_04721_),
    .Y(_04829_),
    .A2(net161),
    .A1(net275));
 sg13g2_nand2_1 _13110_ (.Y(_04830_),
    .A(net1376),
    .B(_04598_));
 sg13g2_o21ai_1 _13111_ (.B1(_04830_),
    .Y(_04831_),
    .A1(_04727_),
    .A2(_04736_));
 sg13g2_and2_1 _13112_ (.A(_04724_),
    .B(_04732_),
    .X(_04832_));
 sg13g2_nand4_1 _13113_ (.B(net1512),
    .C(net282),
    .A(net1508),
    .Y(_04833_),
    .D(_03914_));
 sg13g2_or4_1 _13114_ (.A(net1508),
    .B(net1512),
    .C(net283),
    .D(_03914_),
    .X(_04834_));
 sg13g2_a21oi_1 _13115_ (.A1(_04833_),
    .A2(_04834_),
    .Y(_04835_),
    .B1(net1873));
 sg13g2_a21oi_1 _13116_ (.A1(net1875),
    .A2(_04832_),
    .Y(_04836_),
    .B1(_04835_));
 sg13g2_nor3_1 _13117_ (.A(net1376),
    .B(_04829_),
    .C(_04836_),
    .Y(_04837_));
 sg13g2_a21o_1 _13118_ (.A2(_04831_),
    .A1(_04829_),
    .B1(_04837_),
    .X(_04838_));
 sg13g2_nand2_1 _13119_ (.Y(_04839_),
    .A(net159),
    .B(_04838_));
 sg13g2_nor3_2 _13120_ (.A(_04746_),
    .B(_04622_),
    .C(_04839_),
    .Y(_04840_));
 sg13g2_nor2_1 _13121_ (.A(_04720_),
    .B(_04840_),
    .Y(_04841_));
 sg13g2_nand3_1 _13122_ (.B(_04726_),
    .C(_04736_),
    .A(net158),
    .Y(_04842_));
 sg13g2_o21ai_1 _13123_ (.B1(_04842_),
    .Y(_04843_),
    .A1(net157),
    .A2(_04726_));
 sg13g2_nor3_1 _13124_ (.A(_04722_),
    .B(_04726_),
    .C(_04737_),
    .Y(_04844_));
 sg13g2_a21oi_1 _13125_ (.A1(_04722_),
    .A2(_04843_),
    .Y(_04845_),
    .B1(_04844_));
 sg13g2_nor4_1 _13126_ (.A(net233),
    .B(_04598_),
    .C(_04829_),
    .D(_04737_),
    .Y(_04846_));
 sg13g2_a21oi_1 _13127_ (.A1(_04829_),
    .A2(_04810_),
    .Y(_04847_),
    .B1(_04846_));
 sg13g2_o21ai_1 _13128_ (.B1(_04847_),
    .Y(_04848_),
    .A1(net1376),
    .A2(_04845_));
 sg13g2_inv_1 _13129_ (.Y(_04849_),
    .A(_04848_));
 sg13g2_inv_1 _13130_ (.Y(_04850_),
    .A(_04838_));
 sg13g2_o21ai_1 _13131_ (.B1(_04850_),
    .Y(_04851_),
    .A1(_04746_),
    .A2(_04622_));
 sg13g2_and3_1 _13132_ (.X(_04852_),
    .A(_04720_),
    .B(_04849_),
    .C(_04851_));
 sg13g2_o21ai_1 _13133_ (.B1(_04848_),
    .Y(_04853_),
    .A1(_04746_),
    .A2(_04622_));
 sg13g2_o21ai_1 _13134_ (.B1(_04853_),
    .Y(_04854_),
    .A1(_04841_),
    .A2(_04852_));
 sg13g2_xnor2_1 _13135_ (.Y(_04855_),
    .A(_04827_),
    .B(_04854_));
 sg13g2_o21ai_1 _13136_ (.B1(_04623_),
    .Y(_04856_),
    .A1(_04627_),
    .A2(_04600_));
 sg13g2_nand3_1 _13137_ (.B(_04600_),
    .C(_04622_),
    .A(_04627_),
    .Y(_04857_));
 sg13g2_and2_1 _13138_ (.A(_04856_),
    .B(_04857_),
    .X(_04858_));
 sg13g2_mux2_2 _13139_ (.A0(_04858_),
    .A1(_04748_),
    .S(_04740_),
    .X(_04859_));
 sg13g2_nor2b_1 _13140_ (.A(_04855_),
    .B_N(_04859_),
    .Y(_04860_));
 sg13g2_nand2b_1 _13141_ (.Y(_04861_),
    .B(_04855_),
    .A_N(_04859_));
 sg13g2_nor2b_1 _13142_ (.A(_04860_),
    .B_N(_04861_),
    .Y(_04862_));
 sg13g2_inv_1 _13143_ (.Y(_04863_),
    .A(_04862_));
 sg13g2_inv_1 _13144_ (.Y(_04864_),
    .A(_04703_));
 sg13g2_inv_1 _13145_ (.Y(_04865_),
    .A(_04751_));
 sg13g2_or2_1 _13146_ (.X(_04866_),
    .B(_04355_),
    .A(_04322_));
 sg13g2_nand2_1 _13147_ (.Y(_04867_),
    .A(_04358_),
    .B(_04866_));
 sg13g2_nor2_1 _13148_ (.A(_04384_),
    .B(_04867_),
    .Y(_04868_));
 sg13g2_or4_1 _13149_ (.A(_04385_),
    .B(_04472_),
    .C(_04549_),
    .D(_04868_),
    .X(_04869_));
 sg13g2_and2_1 _13150_ (.A(_04693_),
    .B(_04869_),
    .X(_04870_));
 sg13g2_a221oi_1 _13151_ (.B2(_04649_),
    .C1(_04870_),
    .B1(_04693_),
    .A1(_04864_),
    .Y(_04871_),
    .A2(_04865_));
 sg13g2_a22oi_1 _13152_ (.Y(_04872_),
    .B1(_04640_),
    .B2(_04519_),
    .A2(_04626_),
    .A1(_04631_));
 sg13g2_or2_1 _13153_ (.X(_04873_),
    .B(_04640_),
    .A(net51));
 sg13g2_nand2_1 _13154_ (.Y(_04874_),
    .A(_04526_),
    .B(_04873_));
 sg13g2_a22oi_1 _13155_ (.Y(_04875_),
    .B1(_04874_),
    .B2(_04519_),
    .A2(_04627_),
    .A1(_04631_));
 sg13g2_o21ai_1 _13156_ (.B1(_04875_),
    .Y(_04876_),
    .A1(_04636_),
    .A2(_04872_));
 sg13g2_a221oi_1 _13157_ (.B2(_04358_),
    .C1(_04385_),
    .B1(_04866_),
    .A1(_04470_),
    .Y(_04877_),
    .A2(_04471_));
 sg13g2_and3_1 _13158_ (.X(_04878_),
    .A(_04551_),
    .B(_04470_),
    .C(_04471_));
 sg13g2_nor2_1 _13159_ (.A(_04304_),
    .B(_04322_),
    .Y(_04879_));
 sg13g2_o21ai_1 _13160_ (.B1(_04879_),
    .Y(_04880_),
    .A1(_04386_),
    .A2(_04867_));
 sg13g2_nor4_1 _13161_ (.A(_04549_),
    .B(_04877_),
    .C(_04878_),
    .D(_04880_),
    .Y(_04881_));
 sg13g2_a21o_1 _13162_ (.A2(_04881_),
    .A1(_04876_),
    .B1(_04751_),
    .X(_04882_));
 sg13g2_nand3_1 _13163_ (.B(_04518_),
    .C(_04627_),
    .A(_04468_),
    .Y(_04883_));
 sg13g2_nand2_1 _13164_ (.Y(_04884_),
    .A(net1222),
    .B(net51));
 sg13g2_a21oi_1 _13165_ (.A1(_04883_),
    .A2(_04884_),
    .Y(_04885_),
    .B1(_04640_));
 sg13g2_nor2_1 _13166_ (.A(net51),
    .B(_04546_),
    .Y(_04886_));
 sg13g2_a21oi_1 _13167_ (.A1(net51),
    .A2(_04681_),
    .Y(_04887_),
    .B1(_04886_));
 sg13g2_nor2_1 _13168_ (.A(net1222),
    .B(_04626_),
    .Y(_04888_));
 sg13g2_nor4_1 _13169_ (.A(_04631_),
    .B(_04546_),
    .C(_04632_),
    .D(_04639_),
    .Y(_04889_));
 sg13g2_o21ai_1 _13170_ (.B1(_04636_),
    .Y(_04890_),
    .A1(_04888_),
    .A2(_04889_));
 sg13g2_o21ai_1 _13171_ (.B1(_04890_),
    .Y(_04891_),
    .A1(_04519_),
    .A2(_04887_));
 sg13g2_or3_1 _13172_ (.A(_04628_),
    .B(_04885_),
    .C(_04891_),
    .X(_04892_));
 sg13g2_o21ai_1 _13173_ (.B1(_04628_),
    .Y(_04893_),
    .A1(_04885_),
    .A2(_04891_));
 sg13g2_and4_1 _13174_ (.A(_04751_),
    .B(_04881_),
    .C(_04892_),
    .D(_04893_),
    .X(_04894_));
 sg13g2_a21oi_2 _13175_ (.B1(_04894_),
    .Y(_04895_),
    .A2(_04882_),
    .A1(_04703_));
 sg13g2_nor2b_2 _13176_ (.A(_04871_),
    .B_N(_04895_),
    .Y(_04896_));
 sg13g2_xnor2_1 _13177_ (.Y(_04897_),
    .A(_04863_),
    .B(_04896_));
 sg13g2_nor2_1 _13178_ (.A(_04783_),
    .B(_04897_),
    .Y(_04898_));
 sg13g2_nand2_1 _13179_ (.Y(_04899_),
    .A(_04783_),
    .B(_04897_));
 sg13g2_nand2b_1 _13180_ (.Y(_04900_),
    .B(_04899_),
    .A_N(_04898_));
 sg13g2_xnor2_1 _13181_ (.Y(_04901_),
    .A(_04782_),
    .B(_04900_));
 sg13g2_nor2_1 _13182_ (.A(net298),
    .B(_04901_),
    .Y(_04902_));
 sg13g2_a21oi_1 _13183_ (.A1(_04779_),
    .A2(net300),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_nand2_1 _13184_ (.Y(_04904_),
    .A(net1184),
    .B(_04903_));
 sg13g2_a21oi_1 _13185_ (.A1(_04151_),
    .A2(_04761_),
    .Y(_04905_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_9_ ));
 sg13g2_nand2_1 _13186_ (.Y(_04906_),
    .A(data_addr_o_9_),
    .B(net1014));
 sg13g2_o21ai_1 _13187_ (.B1(_04906_),
    .Y(_04907_),
    .A1(_04779_),
    .A2(net1012));
 sg13g2_nor2_1 _13188_ (.A(net307),
    .B(_04907_),
    .Y(_04908_));
 sg13g2_a21oi_1 _13189_ (.A1(net316),
    .A2(_04905_),
    .Y(_04909_),
    .B1(_04908_));
 sg13g2_nand2_1 _13190_ (.Y(_04910_),
    .A(data_addr_o_9_),
    .B(net1264));
 sg13g2_o21ai_1 _13191_ (.B1(_04910_),
    .Y(_04911_),
    .A1(_04779_),
    .A2(net1264));
 sg13g2_nand2_1 _13192_ (.Y(_04912_),
    .A(net421),
    .B(_04911_));
 sg13g2_o21ai_1 _13193_ (.B1(net1638),
    .Y(_04913_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ),
    .A2(net310));
 sg13g2_nand3_1 _13194_ (.B(_04912_),
    .C(_04913_),
    .A(net1574),
    .Y(_04914_));
 sg13g2_a221oi_1 _13195_ (.B2(net1891),
    .C1(_04914_),
    .B1(_04909_),
    .A1(net1887),
    .Y(_04915_),
    .A2(_04763_));
 sg13g2_o21ai_1 _13196_ (.B1(net1187),
    .Y(_04916_),
    .A1(net338),
    .A2(_04915_));
 sg13g2_o21ai_1 _13197_ (.B1(_04916_),
    .Y(_04917_),
    .A1(net2115),
    .A2(net1574));
 sg13g2_a22oi_1 _13198_ (.Y(_00131_),
    .B1(_04904_),
    .B2(_04917_),
    .A2(net96),
    .A1(_04779_));
 sg13g2_inv_1 _13199_ (.Y(_04918_),
    .A(\ex_block_i.alu_i.imd_val_q_i_42_ ));
 sg13g2_xnor2_1 _13200_ (.Y(_04919_),
    .A(_04714_),
    .B(_04719_));
 sg13g2_and2_1 _13201_ (.A(_04849_),
    .B(_04851_),
    .X(_04920_));
 sg13g2_o21ai_1 _13202_ (.B1(_04853_),
    .Y(_04921_),
    .A1(_04919_),
    .A2(_04920_));
 sg13g2_inv_1 _13203_ (.Y(_04922_),
    .A(_04859_));
 sg13g2_nand2_1 _13204_ (.Y(_04923_),
    .A(_04827_),
    .B(_04922_));
 sg13g2_nor2b_2 _13205_ (.A(_04714_),
    .B_N(_04784_),
    .Y(_04924_));
 sg13g2_nor2_1 _13206_ (.A(_04924_),
    .B(_04840_),
    .Y(_04925_));
 sg13g2_nand2b_1 _13207_ (.Y(_04926_),
    .B(_04714_),
    .A_N(_04784_));
 sg13g2_nor2b_1 _13208_ (.A(_04925_),
    .B_N(_04926_),
    .Y(_04927_));
 sg13g2_nand2_1 _13209_ (.Y(_04928_),
    .A(_04924_),
    .B(_04826_));
 sg13g2_o21ai_1 _13210_ (.B1(_04928_),
    .Y(_04929_),
    .A1(_04826_),
    .A2(_04927_));
 sg13g2_nand2_1 _13211_ (.Y(_04930_),
    .A(_04919_),
    .B(_04840_));
 sg13g2_nor3_1 _13212_ (.A(_04921_),
    .B(_04923_),
    .C(_04930_),
    .Y(_04931_));
 sg13g2_a221oi_1 _13213_ (.B2(_04859_),
    .C1(_04931_),
    .B1(_04929_),
    .A1(_04921_),
    .Y(_04932_),
    .A2(_04923_));
 sg13g2_a22oi_1 _13214_ (.Y(_04933_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_58_ ));
 sg13g2_inv_1 _13215_ (.Y(_04934_),
    .A(_04933_));
 sg13g2_nand2_1 _13216_ (.Y(_04935_),
    .A(_04805_),
    .B(_04824_));
 sg13g2_o21ai_1 _13217_ (.B1(_04785_),
    .Y(_04936_),
    .A1(_04805_),
    .A2(_04824_));
 sg13g2_nand2_1 _13218_ (.Y(_04937_),
    .A(_04935_),
    .B(_04936_));
 sg13g2_nor3_1 _13219_ (.A(net1376),
    .B(_04726_),
    .C(net1338),
    .Y(_04938_));
 sg13g2_mux2_1 _13220_ (.A0(_04938_),
    .A1(net1338),
    .S(_04823_),
    .X(_04939_));
 sg13g2_nor2b_1 _13221_ (.A(_04727_),
    .B_N(net1338),
    .Y(_04940_));
 sg13g2_a22oi_1 _13222_ (.Y(_04941_),
    .B1(_04940_),
    .B2(_04823_),
    .A2(_04939_),
    .A1(_04829_));
 sg13g2_inv_1 _13223_ (.Y(_04942_),
    .A(_04823_));
 sg13g2_mux2_1 _13224_ (.A0(net1338),
    .A1(_04938_),
    .S(_04823_),
    .X(_04943_));
 sg13g2_a221oi_1 _13225_ (.B2(_04722_),
    .C1(net157),
    .B1(_04943_),
    .A1(_04942_),
    .Y(_04944_),
    .A2(_04940_));
 sg13g2_a21oi_2 _13226_ (.B1(_04944_),
    .Y(_04945_),
    .A2(_04941_),
    .A1(net159));
 sg13g2_mux2_2 _13227_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ),
    .S(net425),
    .X(_04946_));
 sg13g2_buf_2 fanout896 (.A(net897),
    .X(net896));
 sg13g2_xnor2_1 _13229_ (.Y(_04948_),
    .A(net1500),
    .B(net250));
 sg13g2_xnor2_1 _13230_ (.Y(_04949_),
    .A(net285),
    .B(net249));
 sg13g2_inv_1 _13231_ (.Y(_04950_),
    .A(net1438));
 sg13g2_a21oi_1 _13232_ (.A1(net1439),
    .A2(_04950_),
    .Y(_04951_),
    .B1(_04051_));
 sg13g2_a221oi_1 _13233_ (.B2(net1378),
    .C1(_04951_),
    .B1(_04949_),
    .A1(net1476),
    .Y(_04952_),
    .A2(_04948_));
 sg13g2_and2_1 _13234_ (.A(net226),
    .B(net252),
    .X(_04953_));
 sg13g2_a21o_1 _13235_ (.A2(net266),
    .A1(_04317_),
    .B1(_04953_),
    .X(_04954_));
 sg13g2_a22oi_1 _13236_ (.Y(_04955_),
    .B1(net1475),
    .B2(net220),
    .A2(net163),
    .A1(net253));
 sg13g2_xor2_1 _13237_ (.B(_04955_),
    .A(net1342),
    .X(_04956_));
 sg13g2_xnor2_1 _13238_ (.Y(_04957_),
    .A(_04954_),
    .B(_04956_));
 sg13g2_xnor2_1 _13239_ (.Y(_04958_),
    .A(_04952_),
    .B(_04957_));
 sg13g2_xnor2_1 _13240_ (.Y(_04959_),
    .A(net224),
    .B(_04795_));
 sg13g2_xnor2_1 _13241_ (.Y(_04960_),
    .A(net166),
    .B(_04796_));
 sg13g2_a21oi_1 _13242_ (.A1(_04959_),
    .A2(_04960_),
    .Y(_04961_),
    .B1(_04793_));
 sg13g2_nor2_1 _13243_ (.A(_04959_),
    .B(_04960_),
    .Y(_04962_));
 sg13g2_nor2_2 _13244_ (.A(_04961_),
    .B(_04962_),
    .Y(_04963_));
 sg13g2_xnor2_1 _13245_ (.Y(_04964_),
    .A(_04958_),
    .B(_04963_));
 sg13g2_inv_1 _13246_ (.Y(_04965_),
    .A(_04964_));
 sg13g2_xnor2_1 _13247_ (.Y(_04966_),
    .A(_04945_),
    .B(_04965_));
 sg13g2_a21oi_2 _13248_ (.B1(_04802_),
    .Y(_04967_),
    .A2(_04803_),
    .A1(_04709_));
 sg13g2_nand2b_2 _13249_ (.Y(_04968_),
    .B(_04967_),
    .A_N(_04799_));
 sg13g2_xor2_1 _13250_ (.B(_04822_),
    .A(net1336),
    .X(_04969_));
 sg13g2_xor2_1 _13251_ (.B(_04813_),
    .A(net156),
    .X(_04970_));
 sg13g2_nand2_1 _13252_ (.Y(_04971_),
    .A(_04969_),
    .B(_04970_));
 sg13g2_buf_4 fanout895 (.X(net895),
    .A(net897));
 sg13g2_buf_8 fanout894 (.A(net898),
    .X(net894));
 sg13g2_and2_1 _13255_ (.A(net272),
    .B(net1340),
    .X(_04974_));
 sg13g2_a21o_1 _13256_ (.A2(net141),
    .A1(net277),
    .B1(_04974_),
    .X(_04975_));
 sg13g2_and2_1 _13257_ (.A(net267),
    .B(net217),
    .X(_04976_));
 sg13g2_a21o_1 _13258_ (.A2(net161),
    .A1(net271),
    .B1(_04976_),
    .X(_04977_));
 sg13g2_nor3_1 _13259_ (.A(net1493),
    .B(_01990_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_26_ ),
    .Y(_04978_));
 sg13g2_nand3_1 _13260_ (.B(_01990_),
    .C(net1497),
    .A(net1493),
    .Y(_04979_));
 sg13g2_nor2b_1 _13261_ (.A(_04978_),
    .B_N(_04979_),
    .Y(_04980_));
 sg13g2_nor3_1 _13262_ (.A(net258),
    .B(net282),
    .C(_03908_),
    .Y(_04981_));
 sg13g2_and3_1 _13263_ (.X(_04982_),
    .A(net258),
    .B(net282),
    .C(_03908_));
 sg13g2_nor3_1 _13264_ (.A(net1874),
    .B(_04981_),
    .C(_04982_),
    .Y(_04983_));
 sg13g2_a21oi_1 _13265_ (.A1(net1875),
    .A2(_04980_),
    .Y(_04984_),
    .B1(_04983_));
 sg13g2_xnor2_1 _13266_ (.Y(_04985_),
    .A(net1493),
    .B(net1497));
 sg13g2_xor2_1 _13267_ (.B(net1464),
    .A(net258),
    .X(_04986_));
 sg13g2_nor2_1 _13268_ (.A(net1874),
    .B(_04986_),
    .Y(_04987_));
 sg13g2_a21oi_1 _13269_ (.A1(net1874),
    .A2(_04985_),
    .Y(_04988_),
    .B1(_04987_));
 sg13g2_nand2_1 _13270_ (.Y(_04989_),
    .A(net230),
    .B(_04988_));
 sg13g2_xor2_1 _13271_ (.B(net1464),
    .A(net281),
    .X(_04990_));
 sg13g2_xnor2_1 _13272_ (.Y(_04991_),
    .A(net1492),
    .B(net1495));
 sg13g2_nand2_1 _13273_ (.Y(_04992_),
    .A(net1875),
    .B(_04991_));
 sg13g2_o21ai_1 _13274_ (.B1(_04992_),
    .Y(_04993_),
    .A1(net1875),
    .A2(_04990_));
 sg13g2_a22oi_1 _13275_ (.Y(_04994_),
    .B1(_04989_),
    .B2(_04993_),
    .A2(_04984_),
    .A1(net233));
 sg13g2_xor2_1 _13276_ (.B(_04994_),
    .A(_04977_),
    .X(_04995_));
 sg13g2_xnor2_1 _13277_ (.Y(_04996_),
    .A(_04975_),
    .B(_04995_));
 sg13g2_xor2_1 _13278_ (.B(_04996_),
    .A(_04971_),
    .X(_04997_));
 sg13g2_nand2b_1 _13279_ (.Y(_04998_),
    .B(_04997_),
    .A_N(_04968_));
 sg13g2_nand2b_1 _13280_ (.Y(_04999_),
    .B(_04968_),
    .A_N(_04997_));
 sg13g2_and2_1 _13281_ (.A(_04998_),
    .B(_04999_),
    .X(_05000_));
 sg13g2_xnor2_1 _13282_ (.Y(_05001_),
    .A(_04966_),
    .B(_05000_));
 sg13g2_xor2_1 _13283_ (.B(_05001_),
    .A(_04937_),
    .X(_05002_));
 sg13g2_xnor2_1 _13284_ (.Y(_05003_),
    .A(_04934_),
    .B(_05002_));
 sg13g2_xnor2_1 _13285_ (.Y(_05004_),
    .A(_04932_),
    .B(_05003_));
 sg13g2_inv_1 _13286_ (.Y(_05005_),
    .A(_04783_));
 sg13g2_nand2_1 _13287_ (.Y(_05006_),
    .A(_05005_),
    .B(_04862_));
 sg13g2_nor2_1 _13288_ (.A(_05005_),
    .B(_04862_),
    .Y(_05007_));
 sg13g2_a21oi_1 _13289_ (.A1(_04896_),
    .A2(_05006_),
    .Y(_05008_),
    .B1(_05007_));
 sg13g2_nor2_1 _13290_ (.A(_04896_),
    .B(_05006_),
    .Y(_05009_));
 sg13g2_a22oi_1 _13291_ (.Y(_05010_),
    .B1(_05009_),
    .B2(_04782_),
    .A2(_05007_),
    .A1(_04896_));
 sg13g2_o21ai_1 _13292_ (.B1(_05010_),
    .Y(_05011_),
    .A1(_04782_),
    .A2(_05008_));
 sg13g2_xor2_1 _13293_ (.B(_05011_),
    .A(_05004_),
    .X(_05012_));
 sg13g2_nor2_1 _13294_ (.A(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .B(net1541),
    .Y(_05013_));
 sg13g2_a21oi_1 _13295_ (.A1(net1541),
    .A2(_05012_),
    .Y(_05014_),
    .B1(_05013_));
 sg13g2_nand2_1 _13296_ (.Y(_05015_),
    .A(net1183),
    .B(_05014_));
 sg13g2_nor3_2 _13297_ (.A(_04112_),
    .B(_04194_),
    .C(net1005),
    .Y(_05016_));
 sg13g2_a21oi_1 _13298_ (.A1(_04085_),
    .A2(_05016_),
    .Y(_05017_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_10_ ));
 sg13g2_buf_4 fanout893 (.X(net893),
    .A(net894));
 sg13g2_nor2_1 _13300_ (.A(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .B(net1012),
    .Y(_05019_));
 sg13g2_a21oi_1 _13301_ (.A1(_02895_),
    .A2(net1012),
    .Y(_05020_),
    .B1(_05019_));
 sg13g2_nor2_1 _13302_ (.A(net312),
    .B(_05020_),
    .Y(_05021_));
 sg13g2_a21oi_1 _13303_ (.A1(net316),
    .A2(_05017_),
    .Y(_05022_),
    .B1(_05021_));
 sg13g2_nor2_1 _13304_ (.A(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .B(net1263),
    .Y(_05023_));
 sg13g2_a21oi_1 _13305_ (.A1(_02895_),
    .A2(net1263),
    .Y(_05024_),
    .B1(_05023_));
 sg13g2_nand2_1 _13306_ (.Y(_05025_),
    .A(net421),
    .B(_05024_));
 sg13g2_o21ai_1 _13307_ (.B1(net1637),
    .Y(_05026_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ),
    .A2(net310));
 sg13g2_nand3_1 _13308_ (.B(_05025_),
    .C(_05026_),
    .A(net1570),
    .Y(_05027_));
 sg13g2_a221oi_1 _13309_ (.B2(net1889),
    .C1(_05027_),
    .B1(_05022_),
    .A1(net1886),
    .Y(_05028_),
    .A2(_04907_));
 sg13g2_o21ai_1 _13310_ (.B1(net1189),
    .Y(_05029_),
    .A1(net338),
    .A2(_05028_));
 sg13g2_o21ai_1 _13311_ (.B1(_05029_),
    .Y(_05030_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .A2(net1572));
 sg13g2_a22oi_1 _13312_ (.Y(_00132_),
    .B1(_05015_),
    .B2(_05030_),
    .A2(net96),
    .A1(_04918_));
 sg13g2_inv_1 _13313_ (.Y(_05031_),
    .A(\ex_block_i.alu_i.imd_val_q_i_43_ ));
 sg13g2_o21ai_1 _13314_ (.B1(_04899_),
    .Y(_05032_),
    .A1(_04782_),
    .A2(_04898_));
 sg13g2_a21oi_1 _13315_ (.A1(_04861_),
    .A2(_04896_),
    .Y(_05033_),
    .B1(_04860_));
 sg13g2_nor2_1 _13316_ (.A(_04921_),
    .B(_04929_),
    .Y(_05034_));
 sg13g2_xnor2_1 _13317_ (.Y(_05035_),
    .A(_05002_),
    .B(_05034_));
 sg13g2_xnor2_1 _13318_ (.Y(_05036_),
    .A(_05033_),
    .B(_05035_));
 sg13g2_nand2_1 _13319_ (.Y(_05037_),
    .A(_04934_),
    .B(_05036_));
 sg13g2_nor2_1 _13320_ (.A(_04934_),
    .B(_05036_),
    .Y(_05038_));
 sg13g2_a21oi_1 _13321_ (.A1(_05032_),
    .A2(_05037_),
    .Y(_05039_),
    .B1(_05038_));
 sg13g2_a22oi_1 _13322_ (.Y(_05040_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_59_ ));
 sg13g2_mux2_2 _13323_ (.A0(net1467),
    .A1(net1498),
    .S(net1874),
    .X(_05041_));
 sg13g2_buf_4 fanout892 (.X(net892),
    .A(\register_file_i/_3038_ ));
 sg13g2_inv_4 _13325_ (.A(net1375),
    .Y(_05043_));
 sg13g2_mux2_2 _13326_ (.A0(_04971_),
    .A1(_05043_),
    .S(_04996_),
    .X(_05044_));
 sg13g2_xor2_1 _13327_ (.B(_04977_),
    .A(net157),
    .X(_05045_));
 sg13g2_xor2_1 _13328_ (.B(net1497),
    .A(net1495),
    .X(_05046_));
 sg13g2_mux2_2 _13329_ (.A0(_04986_),
    .A1(_05046_),
    .S(net1874),
    .X(_05047_));
 sg13g2_nand2_1 _13330_ (.Y(_05048_),
    .A(net231),
    .B(net1335));
 sg13g2_xnor2_1 _13331_ (.Y(_05049_),
    .A(net1375),
    .B(_05048_));
 sg13g2_xor2_1 _13332_ (.B(_04975_),
    .A(net1336),
    .X(_05050_));
 sg13g2_a21oi_1 _13333_ (.A1(_05045_),
    .A2(_05049_),
    .Y(_05051_),
    .B1(_05050_));
 sg13g2_nor2_1 _13334_ (.A(_05045_),
    .B(_05049_),
    .Y(_05052_));
 sg13g2_nor2_1 _13335_ (.A(_05051_),
    .B(_05052_),
    .Y(_05053_));
 sg13g2_xnor2_1 _13336_ (.Y(_05054_),
    .A(_04993_),
    .B(net1374));
 sg13g2_buf_4 fanout891 (.X(net891),
    .A(net892));
 sg13g2_a22oi_1 _13338_ (.Y(_05056_),
    .B1(net160),
    .B2(net268),
    .A2(net218),
    .A1(net253));
 sg13g2_xnor2_1 _13339_ (.Y(_05057_),
    .A(_05054_),
    .B(_05056_));
 sg13g2_nand2b_1 _13340_ (.Y(_05058_),
    .B(net1498),
    .A_N(net1497));
 sg13g2_nand3b_1 _13341_ (.B(net1497),
    .C(net1495),
    .Y(_05059_),
    .A_N(net1498));
 sg13g2_o21ai_1 _13342_ (.B1(_05059_),
    .Y(_05060_),
    .A1(net1495),
    .A2(_05058_));
 sg13g2_nand2b_1 _13343_ (.Y(_05061_),
    .B(net1467),
    .A_N(net1464));
 sg13g2_nand3b_1 _13344_ (.B(net1464),
    .C(net258),
    .Y(_05062_),
    .A_N(net1467));
 sg13g2_o21ai_1 _13345_ (.B1(_05062_),
    .Y(_05063_),
    .A1(net258),
    .A2(_05061_));
 sg13g2_mux2_2 _13346_ (.A0(_05060_),
    .A1(_05063_),
    .S(net1865),
    .X(_05064_));
 sg13g2_and2_1 _13347_ (.A(net275),
    .B(net1335),
    .X(_05065_));
 sg13g2_a21o_1 _13348_ (.A2(net138),
    .A1(net230),
    .B1(_05065_),
    .X(_05066_));
 sg13g2_and2_1 _13349_ (.A(net270),
    .B(net1339),
    .X(_05067_));
 sg13g2_a21o_1 _13350_ (.A2(net141),
    .A1(net274),
    .B1(_05067_),
    .X(_05068_));
 sg13g2_xnor2_1 _13351_ (.Y(_05069_),
    .A(_05066_),
    .B(_05068_));
 sg13g2_xnor2_1 _13352_ (.Y(_05070_),
    .A(_05057_),
    .B(_05069_));
 sg13g2_xnor2_1 _13353_ (.Y(_05071_),
    .A(_05053_),
    .B(_05070_));
 sg13g2_xnor2_1 _13354_ (.Y(_05072_),
    .A(_05044_),
    .B(_05071_));
 sg13g2_nand2b_2 _13355_ (.Y(_05073_),
    .B(_04963_),
    .A_N(_04958_));
 sg13g2_xnor2_1 _13356_ (.Y(_05074_),
    .A(net224),
    .B(_04955_));
 sg13g2_xnor2_1 _13357_ (.Y(_05075_),
    .A(_04354_),
    .B(_04954_));
 sg13g2_o21ai_1 _13358_ (.B1(_04952_),
    .Y(_05076_),
    .A1(_05074_),
    .A2(_05075_));
 sg13g2_nand2_1 _13359_ (.Y(_05077_),
    .A(_05074_),
    .B(_05075_));
 sg13g2_nand2_1 _13360_ (.Y(_05078_),
    .A(_05076_),
    .B(_05077_));
 sg13g2_mux2_2 _13361_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ),
    .S(net425),
    .X(_05079_));
 sg13g2_xnor2_1 _13362_ (.Y(_05080_),
    .A(net1381),
    .B(net246));
 sg13g2_buf_4 fanout890 (.X(net890),
    .A(net891));
 sg13g2_xnor2_1 _13364_ (.Y(_05082_),
    .A(_03905_),
    .B(net247));
 sg13g2_nor2_1 _13365_ (.A(_04422_),
    .B(net248),
    .Y(_05083_));
 sg13g2_a221oi_1 _13366_ (.B2(net1377),
    .C1(_05083_),
    .B1(_05082_),
    .A1(net1476),
    .Y(_05084_),
    .A2(_05080_));
 sg13g2_buf_8 fanout889 (.A(net892),
    .X(net889));
 sg13g2_a22oi_1 _13368_ (.Y(_05086_),
    .B1(net1438),
    .B2(net228),
    .A2(_04704_),
    .A1(net165));
 sg13g2_buf_4 fanout888 (.X(net888),
    .A(net889));
 sg13g2_buf_2 fanout887 (.A(rf_wdata_wb_2_),
    .X(net887));
 sg13g2_buf_2 fanout886 (.A(net887),
    .X(net886));
 sg13g2_a22oi_1 _13372_ (.Y(_05090_),
    .B1(net264),
    .B2(net221),
    .A2(net1474),
    .A1(net163));
 sg13g2_xnor2_1 _13373_ (.Y(_05091_),
    .A(net1342),
    .B(_05090_));
 sg13g2_xnor2_1 _13374_ (.Y(_05092_),
    .A(_05086_),
    .B(_05091_));
 sg13g2_xnor2_1 _13375_ (.Y(_05093_),
    .A(_05084_),
    .B(_05092_));
 sg13g2_xnor2_1 _13376_ (.Y(_05094_),
    .A(_05078_),
    .B(_05093_));
 sg13g2_xnor2_1 _13377_ (.Y(_05095_),
    .A(_05073_),
    .B(_05094_));
 sg13g2_xnor2_1 _13378_ (.Y(_05096_),
    .A(_05072_),
    .B(_05095_));
 sg13g2_inv_1 _13379_ (.Y(_05097_),
    .A(_04968_));
 sg13g2_a21o_1 _13380_ (.A2(_05097_),
    .A1(_04945_),
    .B1(_04964_),
    .X(_05098_));
 sg13g2_nand2b_1 _13381_ (.Y(_05099_),
    .B(_04968_),
    .A_N(_04945_));
 sg13g2_a21oi_1 _13382_ (.A1(_05098_),
    .A2(_05099_),
    .Y(_05100_),
    .B1(_04997_));
 sg13g2_nand2_1 _13383_ (.Y(_05101_),
    .A(_04937_),
    .B(_05100_));
 sg13g2_nand3_1 _13384_ (.B(_04936_),
    .C(_04999_),
    .A(_04935_),
    .Y(_05102_));
 sg13g2_a21oi_1 _13385_ (.A1(_04998_),
    .A2(_05102_),
    .Y(_05103_),
    .B1(_04965_));
 sg13g2_nor2_1 _13386_ (.A(_04937_),
    .B(_04998_),
    .Y(_05104_));
 sg13g2_o21ai_1 _13387_ (.B1(_04945_),
    .Y(_05105_),
    .A1(_05103_),
    .A2(_05104_));
 sg13g2_o21ai_1 _13388_ (.B1(_04997_),
    .Y(_05106_),
    .A1(_04924_),
    .A2(_04825_));
 sg13g2_nand2b_1 _13389_ (.Y(_05107_),
    .B(_04799_),
    .A_N(_04967_));
 sg13g2_a21oi_1 _13390_ (.A1(_04924_),
    .A2(_04825_),
    .Y(_05108_),
    .B1(_05107_));
 sg13g2_a21o_1 _13391_ (.A2(_05106_),
    .A1(_04968_),
    .B1(_05108_),
    .X(_05109_));
 sg13g2_nor2_1 _13392_ (.A(_04945_),
    .B(_04964_),
    .Y(_05110_));
 sg13g2_a22oi_1 _13393_ (.Y(_05111_),
    .B1(_05109_),
    .B2(_05110_),
    .A2(_05104_),
    .A1(_04964_));
 sg13g2_nand3_1 _13394_ (.B(_05105_),
    .C(_05111_),
    .A(_05101_),
    .Y(_05112_));
 sg13g2_xor2_1 _13395_ (.B(_05112_),
    .A(_05096_),
    .X(_05113_));
 sg13g2_o21ai_1 _13396_ (.B1(_05002_),
    .Y(_05114_),
    .A1(_04827_),
    .A2(_04922_));
 sg13g2_nand2b_1 _13397_ (.Y(_05115_),
    .B(_04827_),
    .A_N(_04930_));
 sg13g2_a21oi_1 _13398_ (.A1(_04859_),
    .A2(_05115_),
    .Y(_05116_),
    .B1(_04929_));
 sg13g2_nor2_1 _13399_ (.A(_05002_),
    .B(_05116_),
    .Y(_05117_));
 sg13g2_a21o_1 _13400_ (.A2(_05114_),
    .A1(_04921_),
    .B1(_05117_),
    .X(_05118_));
 sg13g2_a21oi_1 _13401_ (.A1(_04840_),
    .A2(_04926_),
    .Y(_05119_),
    .B1(_04924_));
 sg13g2_nand2b_1 _13402_ (.Y(_05120_),
    .B(_05119_),
    .A_N(_04826_));
 sg13g2_a21oi_1 _13403_ (.A1(_04928_),
    .A2(_05120_),
    .Y(_05121_),
    .B1(_04921_));
 sg13g2_a21o_1 _13404_ (.A2(_04854_),
    .A1(_04827_),
    .B1(_05121_),
    .X(_05122_));
 sg13g2_a22oi_1 _13405_ (.Y(_05123_),
    .B1(_05122_),
    .B2(_04922_),
    .A2(_05034_),
    .A1(_05002_));
 sg13g2_nand3b_1 _13406_ (.B(_05123_),
    .C(_04895_),
    .Y(_05124_),
    .A_N(_04871_));
 sg13g2_nor2b_2 _13407_ (.A(_05118_),
    .B_N(_05124_),
    .Y(_05125_));
 sg13g2_xnor2_1 _13408_ (.Y(_05126_),
    .A(_05113_),
    .B(_05125_));
 sg13g2_xnor2_1 _13409_ (.Y(_05127_),
    .A(_05040_),
    .B(_05126_));
 sg13g2_xnor2_1 _13410_ (.Y(_05128_),
    .A(_05039_),
    .B(_05127_));
 sg13g2_nor2_1 _13411_ (.A(net298),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_a21oi_1 _13412_ (.A1(_05031_),
    .A2(net300),
    .Y(_05130_),
    .B1(_05129_));
 sg13g2_nand2_1 _13413_ (.Y(_05131_),
    .A(net1184),
    .B(_05130_));
 sg13g2_a21oi_1 _13414_ (.A1(_04151_),
    .A2(_05016_),
    .Y(_05132_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_11_ ));
 sg13g2_mux2_1 _13415_ (.A0(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .A1(data_addr_o_11_),
    .S(net1013),
    .X(_05133_));
 sg13g2_nor2_1 _13416_ (.A(net312),
    .B(_05133_),
    .Y(_05134_));
 sg13g2_a21oi_1 _13417_ (.A1(net316),
    .A2(_05132_),
    .Y(_05135_),
    .B1(_05134_));
 sg13g2_nor2_1 _13418_ (.A(data_addr_o_11_),
    .B(net1220),
    .Y(_05136_));
 sg13g2_a21oi_1 _13419_ (.A1(_05031_),
    .A2(net1220),
    .Y(_05137_),
    .B1(_05136_));
 sg13g2_nand2_1 _13420_ (.Y(_05138_),
    .A(net421),
    .B(_05137_));
 sg13g2_o21ai_1 _13421_ (.B1(net1638),
    .Y(_05139_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ),
    .A2(net310));
 sg13g2_nand3_1 _13422_ (.B(_05138_),
    .C(_05139_),
    .A(net1573),
    .Y(_05140_));
 sg13g2_a221oi_1 _13423_ (.B2(net1889),
    .C1(_05140_),
    .B1(_05135_),
    .A1(net1886),
    .Y(_05141_),
    .A2(_05020_));
 sg13g2_o21ai_1 _13424_ (.B1(net1189),
    .Y(_05142_),
    .A1(net338),
    .A2(_05141_));
 sg13g2_o21ai_1 _13425_ (.B1(_05142_),
    .Y(_05143_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .A2(net1572));
 sg13g2_a22oi_1 _13426_ (.Y(_00133_),
    .B1(_05131_),
    .B2(_05143_),
    .A2(net96),
    .A1(_05031_));
 sg13g2_a21oi_1 _13427_ (.A1(_04332_),
    .A2(_04761_),
    .Y(_05144_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_12_ ));
 sg13g2_mux2_1 _13428_ (.A0(net2114),
    .A1(data_addr_o_12_),
    .S(net1010),
    .X(_05145_));
 sg13g2_nor2_1 _13429_ (.A(net308),
    .B(_05145_),
    .Y(_05146_));
 sg13g2_a21oi_1 _13430_ (.A1(net315),
    .A2(_05144_),
    .Y(_05147_),
    .B1(_05146_));
 sg13g2_mux2_1 _13431_ (.A0(net2114),
    .A1(data_addr_o_12_),
    .S(net1263),
    .X(_05148_));
 sg13g2_nand2_1 _13432_ (.Y(_05149_),
    .A(net420),
    .B(_05148_));
 sg13g2_o21ai_1 _13433_ (.B1(net1636),
    .Y(_05150_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ),
    .A2(net305));
 sg13g2_nand3_1 _13434_ (.B(_05149_),
    .C(_05150_),
    .A(net1569),
    .Y(_05151_));
 sg13g2_a221oi_1 _13435_ (.B2(net1889),
    .C1(_05151_),
    .B1(_05147_),
    .A1(net1886),
    .Y(_05152_),
    .A2(_05133_));
 sg13g2_nor2_2 _13436_ (.A(net93),
    .B(net1478),
    .Y(_05153_));
 sg13g2_buf_2 fanout885 (.A(net887),
    .X(net885));
 sg13g2_o21ai_1 _13438_ (.B1(net1579),
    .Y(_05155_),
    .A1(net2114),
    .A2(net1181));
 sg13g2_buf_2 fanout884 (.A(rf_wdata_wb_2_),
    .X(net884));
 sg13g2_nand3_1 _13440_ (.B(_04863_),
    .C(_04896_),
    .A(_05005_),
    .Y(_05157_));
 sg13g2_o21ai_1 _13441_ (.B1(_05157_),
    .Y(_05158_),
    .A1(_05005_),
    .A2(_04897_));
 sg13g2_mux2_1 _13442_ (.A0(_05009_),
    .A1(_05158_),
    .S(_05004_),
    .X(_05159_));
 sg13g2_and2_1 _13443_ (.A(_04679_),
    .B(_04755_),
    .X(_05160_));
 sg13g2_o21ai_1 _13444_ (.B1(_04783_),
    .Y(_05161_),
    .A1(_04753_),
    .A2(_04754_));
 sg13g2_nand2b_1 _13445_ (.Y(_05162_),
    .B(_05161_),
    .A_N(_04897_));
 sg13g2_nand2_1 _13446_ (.Y(_05163_),
    .A(_04780_),
    .B(_05005_));
 sg13g2_o21ai_1 _13447_ (.B1(_04861_),
    .Y(_05164_),
    .A1(_04860_),
    .A2(_04896_));
 sg13g2_xor2_1 _13448_ (.B(_05164_),
    .A(_05035_),
    .X(_05165_));
 sg13g2_a22oi_1 _13449_ (.Y(_05166_),
    .B1(_05165_),
    .B2(_04933_),
    .A2(_05163_),
    .A1(_05162_));
 sg13g2_a221oi_1 _13450_ (.B2(_05160_),
    .C1(_05166_),
    .B1(_05159_),
    .A1(_04934_),
    .Y(_05167_),
    .A2(_05036_));
 sg13g2_a21o_1 _13451_ (.A2(_05126_),
    .A1(_05040_),
    .B1(_05167_),
    .X(_05168_));
 sg13g2_o21ai_1 _13452_ (.B1(_05168_),
    .Y(_05169_),
    .A1(_05040_),
    .A2(_05126_));
 sg13g2_and2_1 _13453_ (.A(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .B(net303),
    .X(_05170_));
 sg13g2_a21o_2 _13454_ (.A2(net323),
    .A1(\ex_block_i.alu_i.imd_val_q_i_44_ ),
    .B1(_05170_),
    .X(_05171_));
 sg13g2_nand2_1 _13455_ (.Y(_05172_),
    .A(_04945_),
    .B(_04997_));
 sg13g2_a21oi_1 _13456_ (.A1(_05096_),
    .A2(_05172_),
    .Y(_05173_),
    .B1(_04968_));
 sg13g2_nor2_1 _13457_ (.A(_04945_),
    .B(_04997_),
    .Y(_05174_));
 sg13g2_nor2_1 _13458_ (.A(_05096_),
    .B(_05174_),
    .Y(_05175_));
 sg13g2_o21ai_1 _13459_ (.B1(_04964_),
    .Y(_05176_),
    .A1(_05173_),
    .A2(_05175_));
 sg13g2_o21ai_1 _13460_ (.B1(_05172_),
    .Y(_05177_),
    .A1(_04968_),
    .A2(_05174_));
 sg13g2_nand2b_1 _13461_ (.Y(_05178_),
    .B(_05177_),
    .A_N(_05096_));
 sg13g2_nand2_1 _13462_ (.Y(_05179_),
    .A(_05094_),
    .B(_05071_));
 sg13g2_inv_1 _13463_ (.Y(_05180_),
    .A(_05179_));
 sg13g2_o21ai_1 _13464_ (.B1(_05044_),
    .Y(_05181_),
    .A1(_05094_),
    .A2(_05071_));
 sg13g2_nand2_1 _13465_ (.Y(_05182_),
    .A(_05181_),
    .B(_05179_));
 sg13g2_or2_1 _13466_ (.X(_05183_),
    .B(_05071_),
    .A(_05094_));
 sg13g2_nor3_1 _13467_ (.A(_05073_),
    .B(_05044_),
    .C(_05183_),
    .Y(_05184_));
 sg13g2_a221oi_1 _13468_ (.B2(_05073_),
    .C1(_05184_),
    .B1(_05182_),
    .A1(_05044_),
    .Y(_05185_),
    .A2(_05180_));
 sg13g2_and2_1 _13469_ (.A(_05053_),
    .B(_05070_),
    .X(_05186_));
 sg13g2_o21ai_1 _13470_ (.B1(_05074_),
    .Y(_05187_),
    .A1(_04952_),
    .A2(_05075_));
 sg13g2_nand2_1 _13471_ (.Y(_05188_),
    .A(_04952_),
    .B(_05075_));
 sg13g2_nand2_1 _13472_ (.Y(_05189_),
    .A(_05187_),
    .B(_05188_));
 sg13g2_nand2_2 _13473_ (.Y(_05190_),
    .A(_05093_),
    .B(_05189_));
 sg13g2_xor2_1 _13474_ (.B(_05190_),
    .A(_05186_),
    .X(_05191_));
 sg13g2_mux2_2 _13475_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_28_ ),
    .S(net425),
    .X(_05192_));
 sg13g2_buf_2 fanout883 (.A(rf_wdata_wb_6_),
    .X(net883));
 sg13g2_xnor2_1 _13477_ (.Y(_05194_),
    .A(net1501),
    .B(net1436));
 sg13g2_xnor2_1 _13478_ (.Y(_05195_),
    .A(net286),
    .B(net1436));
 sg13g2_nor2b_1 _13479_ (.A(net426),
    .B_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ),
    .Y(_05196_));
 sg13g2_a21oi_2 _13480_ (.B1(_05196_),
    .Y(_05197_),
    .A2(net426),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_a21oi_1 _13481_ (.A1(_04174_),
    .A2(_05197_),
    .Y(_05198_),
    .B1(net1379));
 sg13g2_a221oi_1 _13482_ (.B2(net1377),
    .C1(_05198_),
    .B1(_05195_),
    .A1(net1476),
    .Y(_05199_),
    .A2(_05194_));
 sg13g2_a22oi_1 _13483_ (.Y(_05200_),
    .B1(net248),
    .B2(net228),
    .A2(net1438),
    .A1(net165));
 sg13g2_and2_1 _13484_ (.A(net222),
    .B(net252),
    .X(_05201_));
 sg13g2_a21o_1 _13485_ (.A2(net266),
    .A1(_04438_),
    .B1(_05201_),
    .X(_05202_));
 sg13g2_xor2_1 _13486_ (.B(_05202_),
    .A(net1342),
    .X(_05203_));
 sg13g2_xnor2_1 _13487_ (.Y(_05204_),
    .A(_05200_),
    .B(_05203_));
 sg13g2_xnor2_1 _13488_ (.Y(_05205_),
    .A(_05199_),
    .B(_05204_));
 sg13g2_inv_4 _13489_ (.A(net223),
    .Y(_05206_));
 sg13g2_xnor2_1 _13490_ (.Y(_05207_),
    .A(_05206_),
    .B(_05090_));
 sg13g2_xnor2_1 _13491_ (.Y(_05208_),
    .A(_04354_),
    .B(_05086_));
 sg13g2_o21ai_1 _13492_ (.B1(_05208_),
    .Y(_05209_),
    .A1(_05084_),
    .A2(_05207_));
 sg13g2_nand2_1 _13493_ (.Y(_05210_),
    .A(_05084_),
    .B(_05207_));
 sg13g2_nand2_1 _13494_ (.Y(_05211_),
    .A(_05209_),
    .B(_05210_));
 sg13g2_xor2_1 _13495_ (.B(_05211_),
    .A(_05205_),
    .X(_05212_));
 sg13g2_xnor2_1 _13496_ (.Y(_05213_),
    .A(net1336),
    .B(_05068_));
 sg13g2_xor2_1 _13497_ (.B(_05056_),
    .A(net156),
    .X(_05214_));
 sg13g2_xnor2_1 _13498_ (.Y(_05215_),
    .A(net1375),
    .B(_05066_));
 sg13g2_o21ai_1 _13499_ (.B1(_05215_),
    .Y(_05216_),
    .A1(_05213_),
    .A2(_05214_));
 sg13g2_nand2_1 _13500_ (.Y(_05217_),
    .A(_05213_),
    .B(_05214_));
 sg13g2_nand2_1 _13501_ (.Y(_05218_),
    .A(_05216_),
    .B(_05217_));
 sg13g2_xnor2_1 _13502_ (.Y(_05219_),
    .A(net1467),
    .B(net282));
 sg13g2_xor2_1 _13503_ (.B(net1498),
    .A(net1492),
    .X(_05220_));
 sg13g2_nor2_1 _13504_ (.A(net1866),
    .B(_05220_),
    .Y(_05221_));
 sg13g2_a21oi_1 _13505_ (.A1(net1866),
    .A2(_05219_),
    .Y(_05222_),
    .B1(_05221_));
 sg13g2_xnor2_1 _13506_ (.Y(_05223_),
    .A(net1338),
    .B(_05222_));
 sg13g2_a22oi_1 _13507_ (.Y(_05224_),
    .B1(net160),
    .B2(net254),
    .A2(net1474),
    .A1(net217));
 sg13g2_xor2_1 _13508_ (.B(_05224_),
    .A(_05223_),
    .X(_05225_));
 sg13g2_and2_1 _13509_ (.A(net267),
    .B(net1340),
    .X(_05226_));
 sg13g2_a21o_1 _13510_ (.A2(net141),
    .A1(net271),
    .B1(_05226_),
    .X(_05227_));
 sg13g2_and2_1 _13511_ (.A(net272),
    .B(net1335),
    .X(_05228_));
 sg13g2_a21o_1 _13512_ (.A2(net138),
    .A1(net277),
    .B1(_05228_),
    .X(_05229_));
 sg13g2_xnor2_1 _13513_ (.Y(_05230_),
    .A(_05227_),
    .B(_05229_));
 sg13g2_xnor2_1 _13514_ (.Y(_05231_),
    .A(_05225_),
    .B(_05230_));
 sg13g2_xor2_1 _13515_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .A(net1467),
    .X(_05232_));
 sg13g2_xor2_1 _13516_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .A(net1498),
    .X(_05233_));
 sg13g2_mux2_2 _13517_ (.A0(_05232_),
    .A1(_05233_),
    .S(net1872),
    .X(_05234_));
 sg13g2_buf_2 fanout882 (.A(net883),
    .X(net882));
 sg13g2_and2_1 _13519_ (.A(net233),
    .B(net1333),
    .X(_05236_));
 sg13g2_xnor2_1 _13520_ (.Y(_05237_),
    .A(_05231_),
    .B(_05236_));
 sg13g2_xor2_1 _13521_ (.B(_05237_),
    .A(_05218_),
    .X(_05238_));
 sg13g2_xnor2_1 _13522_ (.Y(_05239_),
    .A(_05212_),
    .B(_05238_));
 sg13g2_xnor2_1 _13523_ (.Y(_05240_),
    .A(_05191_),
    .B(_05239_));
 sg13g2_inv_1 _13524_ (.Y(_05241_),
    .A(_05240_));
 sg13g2_xnor2_1 _13525_ (.Y(_05242_),
    .A(_05185_),
    .B(_05241_));
 sg13g2_a21oi_2 _13526_ (.B1(_05242_),
    .Y(_05243_),
    .A2(_05178_),
    .A1(_05176_));
 sg13g2_and3_1 _13527_ (.X(_05244_),
    .A(_05176_),
    .B(_05178_),
    .C(_05242_));
 sg13g2_nor2_2 _13528_ (.A(_05243_),
    .B(_05244_),
    .Y(_05245_));
 sg13g2_nand3b_1 _13529_ (.B(_05124_),
    .C(_05113_),
    .Y(_05246_),
    .A_N(_05118_));
 sg13g2_nand2b_1 _13530_ (.Y(_05247_),
    .B(_04825_),
    .A_N(_04805_));
 sg13g2_nand2_1 _13531_ (.Y(_05248_),
    .A(_04924_),
    .B(_04935_));
 sg13g2_and2_1 _13532_ (.A(_04945_),
    .B(_04964_),
    .X(_05249_));
 sg13g2_mux2_1 _13533_ (.A0(_05110_),
    .A1(_05249_),
    .S(_05096_),
    .X(_05250_));
 sg13g2_nor2_1 _13534_ (.A(_04997_),
    .B(_05097_),
    .Y(_05251_));
 sg13g2_inv_1 _13535_ (.Y(_05252_),
    .A(_04998_));
 sg13g2_mux2_1 _13536_ (.A0(_05251_),
    .A1(_05252_),
    .S(_05096_),
    .X(_05253_));
 sg13g2_a22oi_1 _13537_ (.Y(_05254_),
    .B1(_05253_),
    .B2(_04966_),
    .A2(_05250_),
    .A1(_05000_));
 sg13g2_a21o_1 _13538_ (.A2(_05248_),
    .A1(_05247_),
    .B1(_05254_),
    .X(_05255_));
 sg13g2_nand2_1 _13539_ (.Y(_05256_),
    .A(_05246_),
    .B(_05255_));
 sg13g2_xor2_1 _13540_ (.B(_05256_),
    .A(_05245_),
    .X(_05257_));
 sg13g2_and2_1 _13541_ (.A(_05171_),
    .B(_05257_),
    .X(_05258_));
 sg13g2_a21oi_2 _13542_ (.B1(_05170_),
    .Y(_05259_),
    .A2(net323),
    .A1(net2114));
 sg13g2_nand2b_1 _13543_ (.Y(_05260_),
    .B(_05259_),
    .A_N(_05257_));
 sg13g2_nor2b_1 _13544_ (.A(_05258_),
    .B_N(_05260_),
    .Y(_05261_));
 sg13g2_xnor2_1 _13545_ (.Y(_05262_),
    .A(_05169_),
    .B(_05261_));
 sg13g2_nor3_1 _13546_ (.A(net93),
    .B(net300),
    .C(_05262_),
    .Y(_05263_));
 sg13g2_a21o_1 _13547_ (.A2(_04143_),
    .A1(net2114),
    .B1(_05263_),
    .X(_05264_));
 sg13g2_a22oi_1 _13548_ (.Y(_05265_),
    .B1(net1182),
    .B2(_05264_),
    .A2(net97),
    .A1(net2114));
 sg13g2_o21ai_1 _13549_ (.B1(_05265_),
    .Y(_00134_),
    .A1(_05152_),
    .A2(_05155_));
 sg13g2_o21ai_1 _13550_ (.B1(_05260_),
    .Y(_05266_),
    .A1(_05169_),
    .A2(_05258_));
 sg13g2_and2_1 _13551_ (.A(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .B(net319),
    .X(_05267_));
 sg13g2_a21o_2 _13552_ (.A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .B1(_05267_),
    .X(_05268_));
 sg13g2_nand3_1 _13553_ (.B(_05178_),
    .C(_05242_),
    .A(_05176_),
    .Y(_05269_));
 sg13g2_inv_1 _13554_ (.Y(_05270_),
    .A(_05243_));
 sg13g2_nand3_1 _13555_ (.B(_05270_),
    .C(_05255_),
    .A(_05246_),
    .Y(_05271_));
 sg13g2_nand2_1 _13556_ (.Y(_05272_),
    .A(_05269_),
    .B(_05271_));
 sg13g2_nor2_2 _13557_ (.A(_05205_),
    .B(_05211_),
    .Y(_05273_));
 sg13g2_xnor2_1 _13558_ (.Y(_05274_),
    .A(net1375),
    .B(_05229_));
 sg13g2_xor2_1 _13559_ (.B(_05224_),
    .A(net156),
    .X(_05275_));
 sg13g2_xnor2_1 _13560_ (.Y(_05276_),
    .A(_05043_),
    .B(_05229_));
 sg13g2_xnor2_1 _13561_ (.Y(_05277_),
    .A(net158),
    .B(_05224_));
 sg13g2_xor2_1 _13562_ (.B(_05227_),
    .A(net1336),
    .X(_05278_));
 sg13g2_o21ai_1 _13563_ (.B1(_05278_),
    .Y(_05279_),
    .A1(_05276_),
    .A2(_05277_));
 sg13g2_o21ai_1 _13564_ (.B1(_05279_),
    .Y(_05280_),
    .A1(_05274_),
    .A2(_05275_));
 sg13g2_a22oi_1 _13565_ (.Y(_05281_),
    .B1(net264),
    .B2(net218),
    .A2(net161),
    .A1(net1473));
 sg13g2_xor2_1 _13566_ (.B(_05281_),
    .A(_05223_),
    .X(_05282_));
 sg13g2_and2_1 _13567_ (.A(net270),
    .B(net1335),
    .X(_05283_));
 sg13g2_a21o_1 _13568_ (.A2(net138),
    .A1(net274),
    .B1(_05283_),
    .X(_05284_));
 sg13g2_a22oi_1 _13569_ (.Y(_05285_),
    .B1(net139),
    .B2(net268),
    .A2(net1340),
    .A1(net253));
 sg13g2_xor2_1 _13570_ (.B(_05285_),
    .A(_05284_),
    .X(_05286_));
 sg13g2_xnor2_1 _13571_ (.Y(_05287_),
    .A(_05282_),
    .B(_05286_));
 sg13g2_nand2_1 _13572_ (.Y(_05288_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .B(net1865));
 sg13g2_o21ai_1 _13573_ (.B1(_05288_),
    .Y(_05289_),
    .A1(_01959_),
    .A2(net1865));
 sg13g2_nand2b_1 _13574_ (.Y(_05290_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ));
 sg13g2_nand3b_1 _13575_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ),
    .C(net1467),
    .Y(_05291_),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ));
 sg13g2_o21ai_1 _13576_ (.B1(_05291_),
    .Y(_05292_),
    .A1(net1467),
    .A2(_05290_));
 sg13g2_nand2b_1 _13577_ (.Y(_05293_),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ));
 sg13g2_nand3b_1 _13578_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ),
    .C(net1498),
    .Y(_05294_),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ));
 sg13g2_o21ai_1 _13579_ (.B1(_05294_),
    .Y(_05295_),
    .A1(net1498),
    .A2(_05293_));
 sg13g2_mux2_1 _13580_ (.A0(_05292_),
    .A1(_05295_),
    .S(net1872),
    .X(_05296_));
 sg13g2_a22oi_1 _13581_ (.Y(_05297_),
    .B1(net134),
    .B2(net231),
    .A2(net1333),
    .A1(net275));
 sg13g2_xnor2_1 _13582_ (.Y(_05298_),
    .A(net1329),
    .B(_05297_));
 sg13g2_xnor2_1 _13583_ (.Y(_05299_),
    .A(_05287_),
    .B(_05298_));
 sg13g2_xnor2_1 _13584_ (.Y(_05300_),
    .A(_05280_),
    .B(_05299_));
 sg13g2_xnor2_1 _13585_ (.Y(_05301_),
    .A(_05273_),
    .B(_05300_));
 sg13g2_mux2_2 _13586_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ),
    .S(net425),
    .X(_05302_));
 sg13g2_buf_2 fanout881 (.A(rf_wdata_wb_6_),
    .X(net881));
 sg13g2_xnor2_1 _13588_ (.Y(_05304_),
    .A(net1500),
    .B(net1434));
 sg13g2_xnor2_1 _13589_ (.Y(_05305_),
    .A(net285),
    .B(net1434));
 sg13g2_inv_1 _13590_ (.Y(_05306_),
    .A(net1436));
 sg13g2_a21oi_1 _13591_ (.A1(net1439),
    .A2(_05306_),
    .Y(_05307_),
    .B1(net1379));
 sg13g2_a221oi_1 _13592_ (.B2(net1377),
    .C1(_05307_),
    .B1(_05305_),
    .A1(net1476),
    .Y(_05308_),
    .A2(_05304_));
 sg13g2_buf_2 fanout880 (.A(rf_wdata_wb_6_),
    .X(net880));
 sg13g2_a22oi_1 _13594_ (.Y(_05310_),
    .B1(_04786_),
    .B2(net221),
    .A2(net251),
    .A1(net163));
 sg13g2_and2_1 _13595_ (.A(net226),
    .B(net246),
    .X(_05311_));
 sg13g2_a21o_1 _13596_ (.A2(net249),
    .A1(_04317_),
    .B1(_05311_),
    .X(_05312_));
 sg13g2_xor2_1 _13597_ (.B(_05312_),
    .A(net1341),
    .X(_05313_));
 sg13g2_xnor2_1 _13598_ (.Y(_05314_),
    .A(_05310_),
    .B(_05313_));
 sg13g2_xnor2_1 _13599_ (.Y(_05315_),
    .A(_05308_),
    .B(_05314_));
 sg13g2_xnor2_1 _13600_ (.Y(_05316_),
    .A(net168),
    .B(_05200_));
 sg13g2_xnor2_1 _13601_ (.Y(_05317_),
    .A(_05206_),
    .B(_05202_));
 sg13g2_a21oi_1 _13602_ (.A1(_05316_),
    .A2(_05317_),
    .Y(_05318_),
    .B1(_05199_));
 sg13g2_nor2_1 _13603_ (.A(_05316_),
    .B(_05317_),
    .Y(_05319_));
 sg13g2_nor2_1 _13604_ (.A(_05318_),
    .B(_05319_),
    .Y(_05320_));
 sg13g2_xnor2_1 _13605_ (.Y(_05321_),
    .A(_05315_),
    .B(_05320_));
 sg13g2_nand2_1 _13606_ (.Y(_05322_),
    .A(net232),
    .B(net1333));
 sg13g2_buf_1 fanout879 (.A(rf_wdata_wb_8_),
    .X(net879));
 sg13g2_or2_1 _13608_ (.X(_05324_),
    .B(_05214_),
    .A(_05213_));
 sg13g2_a21o_1 _13609_ (.A2(_05214_),
    .A1(_05213_),
    .B1(_05215_),
    .X(_05325_));
 sg13g2_nand2_1 _13610_ (.Y(_05326_),
    .A(_05324_),
    .B(_05325_));
 sg13g2_nand4_1 _13611_ (.B(_05217_),
    .C(_05231_),
    .A(_05216_),
    .Y(_05327_),
    .D(net1330));
 sg13g2_o21ai_1 _13612_ (.B1(_05327_),
    .Y(_05328_),
    .A1(net1330),
    .A2(_05326_));
 sg13g2_nor2_1 _13613_ (.A(_05236_),
    .B(net1329),
    .Y(_05329_));
 sg13g2_inv_1 _13614_ (.Y(_05330_),
    .A(_05329_));
 sg13g2_nand3_1 _13615_ (.B(_05236_),
    .C(_05325_),
    .A(_05324_),
    .Y(_05331_));
 sg13g2_a21oi_1 _13616_ (.A1(_05330_),
    .A2(_05331_),
    .Y(_05332_),
    .B1(_05231_));
 sg13g2_a21oi_1 _13617_ (.A1(_05322_),
    .A2(_05328_),
    .Y(_05333_),
    .B1(_05332_));
 sg13g2_xnor2_1 _13618_ (.Y(_05334_),
    .A(_05321_),
    .B(_05333_));
 sg13g2_xnor2_1 _13619_ (.Y(_05335_),
    .A(_05301_),
    .B(_05334_));
 sg13g2_inv_1 _13620_ (.Y(_05336_),
    .A(_05186_));
 sg13g2_nand2_1 _13621_ (.Y(_05337_),
    .A(_05212_),
    .B(_05238_));
 sg13g2_nor3_1 _13622_ (.A(_05336_),
    .B(_05190_),
    .C(_05337_),
    .Y(_05338_));
 sg13g2_nor2_1 _13623_ (.A(_05212_),
    .B(_05238_),
    .Y(_05339_));
 sg13g2_a21oi_1 _13624_ (.A1(_05190_),
    .A2(_05337_),
    .Y(_05340_),
    .B1(_05339_));
 sg13g2_nand2_1 _13625_ (.Y(_05341_),
    .A(_05190_),
    .B(_05339_));
 sg13g2_o21ai_1 _13626_ (.B1(_05341_),
    .Y(_05342_),
    .A1(_05186_),
    .A2(_05340_));
 sg13g2_nor2_1 _13627_ (.A(_05338_),
    .B(_05342_),
    .Y(_05343_));
 sg13g2_xnor2_1 _13628_ (.Y(_05344_),
    .A(_05335_),
    .B(_05343_));
 sg13g2_a21oi_1 _13629_ (.A1(_05183_),
    .A2(_05240_),
    .Y(_05345_),
    .B1(_05044_));
 sg13g2_a21oi_1 _13630_ (.A1(_05179_),
    .A2(_05241_),
    .Y(_05346_),
    .B1(_05345_));
 sg13g2_nand2b_1 _13631_ (.Y(_05347_),
    .B(_05179_),
    .A_N(_05044_));
 sg13g2_a21o_1 _13632_ (.A2(_05347_),
    .A1(_05183_),
    .B1(_05240_),
    .X(_05348_));
 sg13g2_o21ai_1 _13633_ (.B1(_05348_),
    .Y(_05349_),
    .A1(_05073_),
    .A2(_05346_));
 sg13g2_nor2_2 _13634_ (.A(_05344_),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_nand2_1 _13635_ (.Y(_05351_),
    .A(_05344_),
    .B(_05349_));
 sg13g2_inv_1 _13636_ (.Y(_05352_),
    .A(_05351_));
 sg13g2_nor2_1 _13637_ (.A(_05350_),
    .B(_05352_),
    .Y(_05353_));
 sg13g2_xnor2_1 _13638_ (.Y(_05354_),
    .A(_05272_),
    .B(_05353_));
 sg13g2_xnor2_1 _13639_ (.Y(_05355_),
    .A(_05268_),
    .B(_05354_));
 sg13g2_xnor2_1 _13640_ (.Y(_05356_),
    .A(_05266_),
    .B(_05355_));
 sg13g2_nand2_1 _13641_ (.Y(_05357_),
    .A(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .B(net298));
 sg13g2_o21ai_1 _13642_ (.B1(_05357_),
    .Y(_05358_),
    .A1(net297),
    .A2(_05356_));
 sg13g2_nand2_1 _13643_ (.Y(_05359_),
    .A(net1183),
    .B(_05358_));
 sg13g2_nor2_1 _13644_ (.A(_04489_),
    .B(_04760_),
    .Y(_05360_));
 sg13g2_nor2_1 _13645_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_13_ ),
    .B(_05360_),
    .Y(_05361_));
 sg13g2_mux2_1 _13646_ (.A0(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .A1(data_addr_o_13_),
    .S(net1010),
    .X(_05362_));
 sg13g2_nor2_1 _13647_ (.A(net312),
    .B(_05362_),
    .Y(_05363_));
 sg13g2_a21oi_1 _13648_ (.A1(net316),
    .A2(_05361_),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_nor2_1 _13649_ (.A(data_addr_o_13_),
    .B(net1220),
    .Y(_05365_));
 sg13g2_a21oi_1 _13650_ (.A1(_02115_),
    .A2(net1220),
    .Y(_05366_),
    .B1(_05365_));
 sg13g2_nand2_1 _13651_ (.Y(_05367_),
    .A(_04116_),
    .B(_05366_));
 sg13g2_o21ai_1 _13652_ (.B1(net1637),
    .Y(_05368_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ),
    .A2(net310));
 sg13g2_nand3_1 _13653_ (.B(_05367_),
    .C(_05368_),
    .A(net1570),
    .Y(_05369_));
 sg13g2_a221oi_1 _13654_ (.B2(net1890),
    .C1(_05369_),
    .B1(_05364_),
    .A1(net1884),
    .Y(_05370_),
    .A2(_05145_));
 sg13g2_o21ai_1 _13655_ (.B1(net1187),
    .Y(_05371_),
    .A1(net338),
    .A2(_05370_));
 sg13g2_o21ai_1 _13656_ (.B1(_05371_),
    .Y(_05372_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .A2(net1575));
 sg13g2_a22oi_1 _13657_ (.Y(_00135_),
    .B1(_05359_),
    .B2(_05372_),
    .A2(net96),
    .A1(_02115_));
 sg13g2_nor2_1 _13658_ (.A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(net1010),
    .Y(_05373_));
 sg13g2_a21oi_1 _13659_ (.A1(_03265_),
    .A2(net1010),
    .Y(_05374_),
    .B1(_05373_));
 sg13g2_a21oi_1 _13660_ (.A1(_04332_),
    .A2(_05016_),
    .Y(_05375_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_14_ ));
 sg13g2_nand2_1 _13661_ (.Y(_05376_),
    .A(net314),
    .B(_05375_));
 sg13g2_o21ai_1 _13662_ (.B1(_05376_),
    .Y(_05377_),
    .A1(net306),
    .A2(_05374_));
 sg13g2_nor2_1 _13663_ (.A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(net1261),
    .Y(_05378_));
 sg13g2_a21oi_1 _13664_ (.A1(_03265_),
    .A2(net1261),
    .Y(_05379_),
    .B1(_05378_));
 sg13g2_o21ai_1 _13665_ (.B1(net1636),
    .Y(_05380_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ),
    .A2(net304));
 sg13g2_nand2_1 _13666_ (.Y(_05381_),
    .A(net1571),
    .B(_05380_));
 sg13g2_a221oi_1 _13667_ (.B2(net419),
    .C1(_05381_),
    .B1(_05379_),
    .A1(net1884),
    .Y(_05382_),
    .A2(_05362_));
 sg13g2_o21ai_1 _13668_ (.B1(_05382_),
    .Y(_05383_),
    .A1(net1708),
    .A2(_05377_));
 sg13g2_a21oi_1 _13669_ (.A1(net1578),
    .A2(_05383_),
    .Y(_05384_),
    .B1(net93));
 sg13g2_and2_1 _13670_ (.A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(net319),
    .X(_05385_));
 sg13g2_a21o_2 _13671_ (.A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .B1(_05385_),
    .X(_05386_));
 sg13g2_nand2b_1 _13672_ (.Y(_05387_),
    .B(_05335_),
    .A_N(_05338_));
 sg13g2_nor2b_1 _13673_ (.A(_05342_),
    .B_N(_05387_),
    .Y(_05388_));
 sg13g2_nand2b_2 _13674_ (.Y(_05389_),
    .B(_05322_),
    .A_N(_05327_));
 sg13g2_a21o_1 _13675_ (.A2(_05331_),
    .A1(_05330_),
    .B1(_05231_),
    .X(_05390_));
 sg13g2_and2_1 _13676_ (.A(_05324_),
    .B(_05325_),
    .X(_05391_));
 sg13g2_nand2_1 _13677_ (.Y(_05392_),
    .A(_05329_),
    .B(_05391_));
 sg13g2_nand3_1 _13678_ (.B(_05390_),
    .C(_05392_),
    .A(_05300_),
    .Y(_05393_));
 sg13g2_inv_1 _13679_ (.Y(_05394_),
    .A(_05321_));
 sg13g2_a21oi_1 _13680_ (.A1(_05389_),
    .A2(_05393_),
    .Y(_05395_),
    .B1(_05394_));
 sg13g2_xor2_1 _13681_ (.B(_05299_),
    .A(_05280_),
    .X(_05396_));
 sg13g2_nor2_1 _13682_ (.A(_05396_),
    .B(_05389_),
    .Y(_05397_));
 sg13g2_o21ai_1 _13683_ (.B1(_05273_),
    .Y(_05398_),
    .A1(_05395_),
    .A2(_05397_));
 sg13g2_a221oi_1 _13684_ (.B2(_05396_),
    .C1(_05332_),
    .B1(_05389_),
    .A1(_05329_),
    .Y(_05399_),
    .A2(_05391_));
 sg13g2_a21o_1 _13685_ (.A2(_05392_),
    .A1(_05390_),
    .B1(_05300_),
    .X(_05400_));
 sg13g2_o21ai_1 _13686_ (.B1(_05400_),
    .Y(_05401_),
    .A1(_05321_),
    .A2(_05399_));
 sg13g2_inv_1 _13687_ (.Y(_05402_),
    .A(_05273_));
 sg13g2_nor2_1 _13688_ (.A(_05321_),
    .B(_05400_),
    .Y(_05403_));
 sg13g2_a221oi_1 _13689_ (.B2(_05402_),
    .C1(_05403_),
    .B1(_05401_),
    .A1(_05321_),
    .Y(_05404_),
    .A2(_05397_));
 sg13g2_nor2b_2 _13690_ (.A(_05315_),
    .B_N(_05320_),
    .Y(_05405_));
 sg13g2_o21ai_1 _13691_ (.B1(_05287_),
    .Y(_05406_),
    .A1(_05298_),
    .A2(_05280_));
 sg13g2_nand2_1 _13692_ (.Y(_05407_),
    .A(_05298_),
    .B(_05280_));
 sg13g2_nand2_1 _13693_ (.Y(_05408_),
    .A(_05406_),
    .B(_05407_));
 sg13g2_xnor2_1 _13694_ (.Y(_05409_),
    .A(_05405_),
    .B(_05408_));
 sg13g2_nor2_1 _13695_ (.A(_02072_),
    .B(net425),
    .Y(_05410_));
 sg13g2_a21oi_2 _13696_ (.B1(_05410_),
    .Y(_05411_),
    .A2(net425),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ));
 sg13g2_xnor2_1 _13697_ (.Y(_05412_),
    .A(net1500),
    .B(_05411_));
 sg13g2_xnor2_1 _13698_ (.Y(_05413_),
    .A(net286),
    .B(_05411_));
 sg13g2_nor2_1 _13699_ (.A(_04422_),
    .B(net1434),
    .Y(_05414_));
 sg13g2_a221oi_1 _13700_ (.B2(net1377),
    .C1(_05414_),
    .B1(_05413_),
    .A1(net1476),
    .Y(_05415_),
    .A2(_05412_));
 sg13g2_a22oi_1 _13701_ (.Y(_05416_),
    .B1(_05192_),
    .B2(net228),
    .A2(net247),
    .A1(net165));
 sg13g2_a22oi_1 _13702_ (.Y(_05417_),
    .B1(net248),
    .B2(net221),
    .A2(net1438),
    .A1(net162));
 sg13g2_xnor2_1 _13703_ (.Y(_05418_),
    .A(net1341),
    .B(_05417_));
 sg13g2_xnor2_1 _13704_ (.Y(_05419_),
    .A(_05416_),
    .B(_05418_));
 sg13g2_xnor2_1 _13705_ (.Y(_05420_),
    .A(_05415_),
    .B(_05419_));
 sg13g2_xnor2_1 _13706_ (.Y(_05421_),
    .A(_05206_),
    .B(_05310_));
 sg13g2_xnor2_1 _13707_ (.Y(_05422_),
    .A(_04354_),
    .B(_05312_));
 sg13g2_nand2_1 _13708_ (.Y(_05423_),
    .A(_05308_),
    .B(_05422_));
 sg13g2_nor2_1 _13709_ (.A(_05308_),
    .B(_05422_),
    .Y(_05424_));
 sg13g2_a21oi_1 _13710_ (.A1(_05421_),
    .A2(_05423_),
    .Y(_05425_),
    .B1(_05424_));
 sg13g2_xnor2_1 _13711_ (.Y(_05426_),
    .A(_05420_),
    .B(_05425_));
 sg13g2_xnor2_1 _13712_ (.Y(_05427_),
    .A(net158),
    .B(_05281_));
 sg13g2_xnor2_1 _13713_ (.Y(_05428_),
    .A(_05043_),
    .B(_05284_));
 sg13g2_xnor2_1 _13714_ (.Y(_05429_),
    .A(net1336),
    .B(_05285_));
 sg13g2_a21oi_1 _13715_ (.A1(_05427_),
    .A2(_05428_),
    .Y(_05430_),
    .B1(_05429_));
 sg13g2_nor2_1 _13716_ (.A(_05427_),
    .B(_05428_),
    .Y(_05431_));
 sg13g2_nor2_1 _13717_ (.A(_05430_),
    .B(_05431_),
    .Y(_05432_));
 sg13g2_nand2_1 _13718_ (.Y(_05433_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .B(net1871));
 sg13g2_nand2_1 _13719_ (.Y(_05434_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ),
    .B(net1872));
 sg13g2_nand3_1 _13720_ (.B(_05433_),
    .C(_05434_),
    .A(net230),
    .Y(_05435_));
 sg13g2_o21ai_1 _13721_ (.B1(_05435_),
    .Y(_05436_),
    .A1(net233),
    .A2(net1330));
 sg13g2_and2_1 _13722_ (.A(net272),
    .B(net1333),
    .X(_05437_));
 sg13g2_a21o_1 _13723_ (.A2(net136),
    .A1(net277),
    .B1(_05437_),
    .X(_05438_));
 sg13g2_xnor2_1 _13724_ (.Y(_05439_),
    .A(_05436_),
    .B(_05438_));
 sg13g2_xnor2_1 _13725_ (.Y(_05440_),
    .A(_04993_),
    .B(_05043_));
 sg13g2_and2_1 _13726_ (.A(net217),
    .B(net252),
    .X(_05441_));
 sg13g2_a21o_1 _13727_ (.A2(net266),
    .A1(net161),
    .B1(_05441_),
    .X(_05442_));
 sg13g2_xnor2_1 _13728_ (.Y(_05443_),
    .A(_05440_),
    .B(_05442_));
 sg13g2_a22oi_1 _13729_ (.Y(_05444_),
    .B1(net139),
    .B2(net254),
    .A2(net1340),
    .A1(net1473));
 sg13g2_and2_1 _13730_ (.A(net267),
    .B(net1335),
    .X(_05445_));
 sg13g2_a21o_1 _13731_ (.A2(net138),
    .A1(net271),
    .B1(_05445_),
    .X(_05446_));
 sg13g2_xor2_1 _13732_ (.B(_05446_),
    .A(_05444_),
    .X(_05447_));
 sg13g2_xnor2_1 _13733_ (.Y(_05448_),
    .A(_05443_),
    .B(_05447_));
 sg13g2_xnor2_1 _13734_ (.Y(_05449_),
    .A(_05439_),
    .B(_05448_));
 sg13g2_xor2_1 _13735_ (.B(_05449_),
    .A(_05432_),
    .X(_05450_));
 sg13g2_nor2_1 _13736_ (.A(_05426_),
    .B(_05450_),
    .Y(_05451_));
 sg13g2_and2_1 _13737_ (.A(_05426_),
    .B(_05450_),
    .X(_05452_));
 sg13g2_nor2_1 _13738_ (.A(_05451_),
    .B(_05452_),
    .Y(_05453_));
 sg13g2_xnor2_1 _13739_ (.Y(_05454_),
    .A(_05409_),
    .B(_05453_));
 sg13g2_a21oi_1 _13740_ (.A1(_05398_),
    .A2(_05404_),
    .Y(_05455_),
    .B1(_05454_));
 sg13g2_and3_1 _13741_ (.X(_05456_),
    .A(_05398_),
    .B(_05404_),
    .C(_05454_));
 sg13g2_nor2_1 _13742_ (.A(_05455_),
    .B(_05456_),
    .Y(_05457_));
 sg13g2_xnor2_1 _13743_ (.Y(_05458_),
    .A(_05388_),
    .B(_05457_));
 sg13g2_o21ai_1 _13744_ (.B1(_05351_),
    .Y(_05459_),
    .A1(_05272_),
    .A2(_05350_));
 sg13g2_xnor2_1 _13745_ (.Y(_05460_),
    .A(_05458_),
    .B(_05459_));
 sg13g2_nand2_1 _13746_ (.Y(_05461_),
    .A(_05386_),
    .B(_05460_));
 sg13g2_a21oi_1 _13747_ (.A1(_05269_),
    .A2(_05271_),
    .Y(_05462_),
    .B1(_05352_));
 sg13g2_or3_1 _13748_ (.A(_05350_),
    .B(_05458_),
    .C(_05462_),
    .X(_05463_));
 sg13g2_o21ai_1 _13749_ (.B1(_05458_),
    .Y(_05464_),
    .A1(_05350_),
    .A2(_05462_));
 sg13g2_a21o_1 _13750_ (.A2(_05464_),
    .A1(_05463_),
    .B1(_05386_),
    .X(_05465_));
 sg13g2_nand2_1 _13751_ (.Y(_05466_),
    .A(_05461_),
    .B(_05465_));
 sg13g2_nor2_1 _13752_ (.A(_05268_),
    .B(_05354_),
    .Y(_05467_));
 sg13g2_nand2_1 _13753_ (.Y(_05468_),
    .A(_05268_),
    .B(_05354_));
 sg13g2_o21ai_1 _13754_ (.B1(_05468_),
    .Y(_05469_),
    .A1(_05266_),
    .A2(_05467_));
 sg13g2_xnor2_1 _13755_ (.Y(_05470_),
    .A(_05466_),
    .B(_05469_));
 sg13g2_o21ai_1 _13756_ (.B1(net1182),
    .Y(_05471_),
    .A1(net297),
    .A2(_05470_));
 sg13g2_nand3_1 _13757_ (.B(net1182),
    .C(_05470_),
    .A(net1541),
    .Y(_05472_));
 sg13g2_a221oi_1 _13758_ (.B2(net299),
    .C1(net93),
    .B1(_05384_),
    .A1(net1478),
    .Y(_05473_),
    .A2(_05472_));
 sg13g2_nor2_1 _13759_ (.A(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .B(_05473_),
    .Y(_05474_));
 sg13g2_a21oi_1 _13760_ (.A1(_05384_),
    .A2(_05471_),
    .Y(_00136_),
    .B1(_05474_));
 sg13g2_inv_1 _13761_ (.Y(_05475_),
    .A(\ex_block_i.alu_i.imd_val_q_i_47_ ));
 sg13g2_nor2_1 _13762_ (.A(_05040_),
    .B(_05259_),
    .Y(_05476_));
 sg13g2_inv_1 _13763_ (.Y(_05477_),
    .A(_05040_));
 sg13g2_nor3_1 _13764_ (.A(_05477_),
    .B(_05113_),
    .C(_05125_),
    .Y(_05478_));
 sg13g2_a21oi_1 _13765_ (.A1(_05247_),
    .A2(_05248_),
    .Y(_05479_),
    .B1(_05254_));
 sg13g2_o21ai_1 _13766_ (.B1(_05479_),
    .Y(_05480_),
    .A1(_05259_),
    .A2(_05478_));
 sg13g2_o21ai_1 _13767_ (.B1(_05480_),
    .Y(_05481_),
    .A1(_05246_),
    .A2(_05476_));
 sg13g2_inv_1 _13768_ (.Y(_05482_),
    .A(_05113_));
 sg13g2_or3_1 _13769_ (.A(_05482_),
    .B(_05259_),
    .C(_05245_),
    .X(_05483_));
 sg13g2_o21ai_1 _13770_ (.B1(_05483_),
    .Y(_05484_),
    .A1(_05040_),
    .A2(_05113_));
 sg13g2_nor3_1 _13771_ (.A(_05243_),
    .B(_05244_),
    .C(_05479_),
    .Y(_05485_));
 sg13g2_nand2_1 _13772_ (.Y(_05486_),
    .A(_05482_),
    .B(_05485_));
 sg13g2_o21ai_1 _13773_ (.B1(_05486_),
    .Y(_05487_),
    .A1(_05245_),
    .A2(_05255_));
 sg13g2_a22oi_1 _13774_ (.Y(_05488_),
    .B1(_05171_),
    .B2(_05485_),
    .A2(_05113_),
    .A1(_05477_));
 sg13g2_nor2_1 _13775_ (.A(_05125_),
    .B(_05488_),
    .Y(_05489_));
 sg13g2_a221oi_1 _13776_ (.B2(_05171_),
    .C1(_05489_),
    .B1(_05487_),
    .A1(_05125_),
    .Y(_05490_),
    .A2(_05484_));
 sg13g2_o21ai_1 _13777_ (.B1(_05255_),
    .Y(_05491_),
    .A1(_05243_),
    .A2(_05244_));
 sg13g2_nor2_1 _13778_ (.A(_05171_),
    .B(_05491_),
    .Y(_05492_));
 sg13g2_o21ai_1 _13779_ (.B1(_05171_),
    .Y(_05493_),
    .A1(_05113_),
    .A2(_05491_));
 sg13g2_nand3_1 _13780_ (.B(_05482_),
    .C(_05493_),
    .A(_05040_),
    .Y(_05494_));
 sg13g2_nor2b_1 _13781_ (.A(_05492_),
    .B_N(_05494_),
    .Y(_05495_));
 sg13g2_and4_1 _13782_ (.A(_05040_),
    .B(_05113_),
    .C(_05125_),
    .D(_05259_),
    .X(_05496_));
 sg13g2_a21oi_1 _13783_ (.A1(_05482_),
    .A2(_05492_),
    .Y(_05497_),
    .B1(_05496_));
 sg13g2_o21ai_1 _13784_ (.B1(_05497_),
    .Y(_05498_),
    .A1(_05125_),
    .A2(_05495_));
 sg13g2_a221oi_1 _13785_ (.B2(_05167_),
    .C1(_05498_),
    .B1(_05490_),
    .A1(_05245_),
    .Y(_05499_),
    .A2(_05481_));
 sg13g2_o21ai_1 _13786_ (.B1(_05354_),
    .Y(_05500_),
    .A1(_05268_),
    .A2(_05499_));
 sg13g2_nand2_1 _13787_ (.Y(_05501_),
    .A(_05268_),
    .B(_05499_));
 sg13g2_nand2_1 _13788_ (.Y(_05502_),
    .A(_05500_),
    .B(_05501_));
 sg13g2_inv_1 _13789_ (.Y(_05503_),
    .A(_05461_));
 sg13g2_a21oi_1 _13790_ (.A1(_05465_),
    .A2(_05502_),
    .Y(_05504_),
    .B1(_05503_));
 sg13g2_buf_2 fanout878 (.A(net879),
    .X(net878));
 sg13g2_a22oi_1 _13792_ (.Y(_05506_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .A2(net301),
    .A1(\ex_block_i.alu_i.imd_val_q_i_63_ ));
 sg13g2_inv_1 _13793_ (.Y(_05507_),
    .A(_05506_));
 sg13g2_o21ai_1 _13794_ (.B1(_05423_),
    .Y(_05508_),
    .A1(_05421_),
    .A2(_05424_));
 sg13g2_nand2_2 _13795_ (.Y(_05509_),
    .A(_05420_),
    .B(_05508_));
 sg13g2_xor2_1 _13796_ (.B(_05444_),
    .A(net1336),
    .X(_05510_));
 sg13g2_xnor2_1 _13797_ (.Y(_05511_),
    .A(_05043_),
    .B(_05446_));
 sg13g2_xor2_1 _13798_ (.B(_05442_),
    .A(net156),
    .X(_05512_));
 sg13g2_nor2_1 _13799_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sg13g2_nand2_1 _13800_ (.Y(_05514_),
    .A(_05511_),
    .B(_05512_));
 sg13g2_o21ai_1 _13801_ (.B1(_05514_),
    .Y(_05515_),
    .A1(_05510_),
    .A2(_05513_));
 sg13g2_nor3_1 _13802_ (.A(_01959_),
    .B(_01856_),
    .C(net288),
    .Y(_05516_));
 sg13g2_nand3_1 _13803_ (.B(_01856_),
    .C(net288),
    .A(_01959_),
    .Y(_05517_));
 sg13g2_nor2b_1 _13804_ (.A(_05516_),
    .B_N(_05517_),
    .Y(_05518_));
 sg13g2_nor3_1 _13805_ (.A(_02097_),
    .B(_03919_),
    .C(net1469),
    .Y(_05519_));
 sg13g2_and3_1 _13806_ (.X(_05520_),
    .A(_02097_),
    .B(_03919_),
    .C(net1469));
 sg13g2_nor3_1 _13807_ (.A(net1872),
    .B(_05519_),
    .C(_05520_),
    .Y(_05521_));
 sg13g2_a21oi_2 _13808_ (.B1(_05521_),
    .Y(_05522_),
    .A2(_05518_),
    .A1(net1872));
 sg13g2_xnor2_1 _13809_ (.Y(_05523_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ));
 sg13g2_xor2_1 _13810_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .X(_05524_));
 sg13g2_nor2_1 _13811_ (.A(net1872),
    .B(_05524_),
    .Y(_05525_));
 sg13g2_a21oi_2 _13812_ (.B1(_05525_),
    .Y(_05526_),
    .A2(_05523_),
    .A1(net1872));
 sg13g2_and2_1 _13813_ (.A(net275),
    .B(net1258),
    .X(_05527_));
 sg13g2_a21o_1 _13814_ (.A2(net92),
    .A1(net230),
    .B1(_05527_),
    .X(_05528_));
 sg13g2_xnor2_1 _13815_ (.Y(_05529_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ),
    .B(net1469));
 sg13g2_xor2_1 _13816_ (.B(net288),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ),
    .X(_05530_));
 sg13g2_nor2_1 _13817_ (.A(net1865),
    .B(_05530_),
    .Y(_05531_));
 sg13g2_a21oi_2 _13818_ (.B1(_05531_),
    .Y(_05532_),
    .A2(_05529_),
    .A1(net1865));
 sg13g2_and2_1 _13819_ (.A(net270),
    .B(net1333),
    .X(_05533_));
 sg13g2_a21o_1 _13820_ (.A2(net136),
    .A1(net274),
    .B1(_05533_),
    .X(_05534_));
 sg13g2_xor2_1 _13821_ (.B(_05534_),
    .A(_05532_),
    .X(_05535_));
 sg13g2_xnor2_1 _13822_ (.Y(_05536_),
    .A(_05528_),
    .B(_05535_));
 sg13g2_a22oi_1 _13823_ (.Y(_05537_),
    .B1(net137),
    .B2(net268),
    .A2(_05047_),
    .A1(net253));
 sg13g2_xnor2_1 _13824_ (.Y(_05538_),
    .A(_05054_),
    .B(_05537_));
 sg13g2_a22oi_1 _13825_ (.Y(_05539_),
    .B1(net1437),
    .B2(net218),
    .A2(net251),
    .A1(net160));
 sg13g2_a22oi_1 _13826_ (.Y(_05540_),
    .B1(net139),
    .B2(net1474),
    .A2(net1340),
    .A1(net264));
 sg13g2_xnor2_1 _13827_ (.Y(_05541_),
    .A(_05539_),
    .B(_05540_));
 sg13g2_xnor2_1 _13828_ (.Y(_05542_),
    .A(_05538_),
    .B(_05541_));
 sg13g2_xnor2_1 _13829_ (.Y(_05543_),
    .A(_05536_),
    .B(_05542_));
 sg13g2_xnor2_1 _13830_ (.Y(_05544_),
    .A(_05515_),
    .B(_05543_));
 sg13g2_xnor2_1 _13831_ (.Y(_05545_),
    .A(_05509_),
    .B(_05544_));
 sg13g2_xnor2_1 _13832_ (.Y(_05546_),
    .A(net168),
    .B(_05416_));
 sg13g2_xnor2_1 _13833_ (.Y(_05547_),
    .A(net224),
    .B(_05417_));
 sg13g2_nand2_1 _13834_ (.Y(_05548_),
    .A(_05546_),
    .B(_05547_));
 sg13g2_nor2_1 _13835_ (.A(_05546_),
    .B(_05547_),
    .Y(_05549_));
 sg13g2_a21o_2 _13836_ (.A2(_05548_),
    .A1(_05415_),
    .B1(_05549_),
    .X(_05550_));
 sg13g2_a22oi_1 _13837_ (.Y(_05551_),
    .B1(net246),
    .B2(net221),
    .A2(net249),
    .A1(net163));
 sg13g2_xnor2_1 _13838_ (.Y(_05552_),
    .A(net223),
    .B(_05551_));
 sg13g2_inv_1 _13839_ (.Y(_05553_),
    .A(_05552_));
 sg13g2_a22oi_1 _13840_ (.Y(_05554_),
    .B1(net1433),
    .B2(net227),
    .A2(net1436),
    .A1(net165));
 sg13g2_xnor2_1 _13841_ (.Y(_05555_),
    .A(net166),
    .B(_05554_));
 sg13g2_mux2_2 _13842_ (.A0(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .S(net424),
    .X(_05556_));
 sg13g2_buf_2 fanout877 (.A(net879),
    .X(net877));
 sg13g2_xnor2_1 _13844_ (.Y(_05558_),
    .A(net1500),
    .B(net244));
 sg13g2_xnor2_1 _13845_ (.Y(_05559_),
    .A(net285),
    .B(net244));
 sg13g2_a21oi_1 _13846_ (.A1(net1439),
    .A2(_05411_),
    .Y(_05560_),
    .B1(net1379));
 sg13g2_a221oi_1 _13847_ (.B2(net1377),
    .C1(_05560_),
    .B1(_05559_),
    .A1(net1476),
    .Y(_05561_),
    .A2(_05558_));
 sg13g2_xor2_1 _13848_ (.B(_05561_),
    .A(_05555_),
    .X(_05562_));
 sg13g2_xnor2_1 _13849_ (.Y(_05563_),
    .A(_05553_),
    .B(_05562_));
 sg13g2_xnor2_1 _13850_ (.Y(_05564_),
    .A(_05550_),
    .B(_05563_));
 sg13g2_xnor2_1 _13851_ (.Y(_05565_),
    .A(net1329),
    .B(_05438_));
 sg13g2_nand2_1 _13852_ (.Y(_05566_),
    .A(net1469),
    .B(net1869));
 sg13g2_nand2_1 _13853_ (.Y(_05567_),
    .A(net289),
    .B(net1876));
 sg13g2_and2_1 _13854_ (.A(_05566_),
    .B(_05567_),
    .X(_05568_));
 sg13g2_buf_2 fanout876 (.A(rf_wdata_wb_8_),
    .X(net876));
 sg13g2_nand2_1 _13856_ (.Y(_05570_),
    .A(net231),
    .B(net1258));
 sg13g2_mux2_2 _13857_ (.A0(_05565_),
    .A1(net1327),
    .S(_05570_),
    .X(_05571_));
 sg13g2_or2_1 _13858_ (.X(_05572_),
    .B(_05448_),
    .A(_05439_));
 sg13g2_xor2_1 _13859_ (.B(_05281_),
    .A(net156),
    .X(_05573_));
 sg13g2_nor2_1 _13860_ (.A(_05429_),
    .B(_05428_),
    .Y(_05574_));
 sg13g2_nand2_1 _13861_ (.Y(_05575_),
    .A(_05429_),
    .B(_05428_));
 sg13g2_o21ai_1 _13862_ (.B1(_05575_),
    .Y(_05576_),
    .A1(_05573_),
    .A2(_05574_));
 sg13g2_and2_1 _13863_ (.A(_05439_),
    .B(_05448_),
    .X(_05577_));
 sg13g2_a21oi_2 _13864_ (.B1(_05577_),
    .Y(_05578_),
    .A2(_05576_),
    .A1(_05572_));
 sg13g2_xnor2_1 _13865_ (.Y(_05579_),
    .A(_05571_),
    .B(_05578_));
 sg13g2_xnor2_1 _13866_ (.Y(_05580_),
    .A(_05564_),
    .B(_05579_));
 sg13g2_xnor2_1 _13867_ (.Y(_05581_),
    .A(_05545_),
    .B(_05580_));
 sg13g2_a21oi_1 _13868_ (.A1(_05276_),
    .A2(_05277_),
    .Y(_05582_),
    .B1(_05278_));
 sg13g2_a21o_1 _13869_ (.A2(_05275_),
    .A1(_05274_),
    .B1(_05582_),
    .X(_05583_));
 sg13g2_nand2b_1 _13870_ (.Y(_05584_),
    .B(_05583_),
    .A_N(_05298_));
 sg13g2_nor2b_1 _13871_ (.A(_05583_),
    .B_N(_05298_),
    .Y(_05585_));
 sg13g2_a21o_1 _13872_ (.A2(_05584_),
    .A1(_05287_),
    .B1(_05585_),
    .X(_05586_));
 sg13g2_nand3_1 _13873_ (.B(_05451_),
    .C(_05586_),
    .A(_05405_),
    .Y(_05587_));
 sg13g2_inv_1 _13874_ (.Y(_05588_),
    .A(_05405_));
 sg13g2_inv_1 _13875_ (.Y(_05589_),
    .A(_05452_));
 sg13g2_o21ai_1 _13876_ (.B1(_05589_),
    .Y(_05590_),
    .A1(_05405_),
    .A2(_05451_));
 sg13g2_o21ai_1 _13877_ (.B1(_05584_),
    .Y(_05591_),
    .A1(_05287_),
    .A2(_05585_));
 sg13g2_a22oi_1 _13878_ (.Y(_05592_),
    .B1(_05590_),
    .B2(_05591_),
    .A2(_05452_),
    .A1(_05588_));
 sg13g2_nand2_1 _13879_ (.Y(_05593_),
    .A(_05587_),
    .B(_05592_));
 sg13g2_xor2_1 _13880_ (.B(_05593_),
    .A(_05581_),
    .X(_05594_));
 sg13g2_nand2_1 _13881_ (.Y(_05595_),
    .A(_05394_),
    .B(_05396_));
 sg13g2_and2_1 _13882_ (.A(_05390_),
    .B(_05392_),
    .X(_05596_));
 sg13g2_o21ai_1 _13883_ (.B1(_05454_),
    .Y(_05597_),
    .A1(_05273_),
    .A2(_05596_));
 sg13g2_o21ai_1 _13884_ (.B1(_05597_),
    .Y(_05598_),
    .A1(_05402_),
    .A2(_05389_));
 sg13g2_nor2_1 _13885_ (.A(_05394_),
    .B(_05396_),
    .Y(_05599_));
 sg13g2_nand2_1 _13886_ (.Y(_05600_),
    .A(_05273_),
    .B(_05596_));
 sg13g2_nor2_1 _13887_ (.A(_05454_),
    .B(_05599_),
    .Y(_05601_));
 sg13g2_a21oi_1 _13888_ (.A1(_05389_),
    .A2(_05600_),
    .Y(_05602_),
    .B1(_05601_));
 sg13g2_a221oi_1 _13889_ (.B2(_05454_),
    .C1(_05602_),
    .B1(_05599_),
    .A1(_05595_),
    .Y(_05603_),
    .A2(_05598_));
 sg13g2_and2_1 _13890_ (.A(_05594_),
    .B(_05603_),
    .X(_05604_));
 sg13g2_or2_1 _13891_ (.X(_05605_),
    .B(_05603_),
    .A(_05594_));
 sg13g2_nand2b_1 _13892_ (.Y(_05606_),
    .B(_05605_),
    .A_N(_05604_));
 sg13g2_nor4_1 _13893_ (.A(_05244_),
    .B(_05350_),
    .C(_05352_),
    .D(_05458_),
    .Y(_05607_));
 sg13g2_nand2b_1 _13894_ (.Y(_05608_),
    .B(_05338_),
    .A_N(_05335_));
 sg13g2_o21ai_1 _13895_ (.B1(_05608_),
    .Y(_05609_),
    .A1(_05455_),
    .A2(_05456_));
 sg13g2_a22oi_1 _13896_ (.Y(_05610_),
    .B1(_05609_),
    .B2(_05349_),
    .A2(_05457_),
    .A1(_05387_));
 sg13g2_nand3b_1 _13897_ (.B(_05349_),
    .C(_05457_),
    .Y(_05611_),
    .A_N(_05335_));
 sg13g2_o21ai_1 _13898_ (.B1(_05611_),
    .Y(_05612_),
    .A1(_05342_),
    .A2(_05610_));
 sg13g2_a21oi_1 _13899_ (.A1(_05271_),
    .A2(_05607_),
    .Y(_05613_),
    .B1(_05612_));
 sg13g2_xor2_1 _13900_ (.B(net35),
    .A(_05606_),
    .X(_05614_));
 sg13g2_xnor2_1 _13901_ (.Y(_05615_),
    .A(_05507_),
    .B(_05614_));
 sg13g2_xnor2_1 _13902_ (.Y(_05616_),
    .A(_05504_),
    .B(_05615_));
 sg13g2_nand2_1 _13903_ (.Y(_05617_),
    .A(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .B(net298));
 sg13g2_o21ai_1 _13904_ (.B1(_05617_),
    .Y(_05618_),
    .A1(net298),
    .A2(_05616_));
 sg13g2_mux2_1 _13905_ (.A0(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .A1(data_addr_o_15_),
    .S(net1008),
    .X(_05619_));
 sg13g2_nand4_1 _13906_ (.B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .C(net1009),
    .A(net2112),
    .Y(_05620_),
    .D(_04488_));
 sg13g2_nand3b_1 _13907_ (.B(net313),
    .C(_05620_),
    .Y(_05621_),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_15_ ));
 sg13g2_o21ai_1 _13908_ (.B1(_05621_),
    .Y(_05622_),
    .A1(net308),
    .A2(_05619_));
 sg13g2_nor2_1 _13909_ (.A(data_addr_o_15_),
    .B(net1218),
    .Y(_05623_));
 sg13g2_a21oi_1 _13910_ (.A1(_05475_),
    .A2(net1218),
    .Y(_05624_),
    .B1(_05623_));
 sg13g2_o21ai_1 _13911_ (.B1(net1635),
    .Y(_05625_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ),
    .A2(net309));
 sg13g2_nand2_1 _13912_ (.Y(_05626_),
    .A(net1181),
    .B(_05625_));
 sg13g2_a221oi_1 _13913_ (.B2(net420),
    .C1(_05626_),
    .B1(_05624_),
    .A1(net1884),
    .Y(_05627_),
    .A2(_05374_));
 sg13g2_o21ai_1 _13914_ (.B1(_05627_),
    .Y(_05628_),
    .A1(net1708),
    .A2(_05622_));
 sg13g2_a22oi_1 _13915_ (.Y(_05629_),
    .B1(net1478),
    .B2(_05475_),
    .A2(net1185),
    .A1(net337));
 sg13g2_a22oi_1 _13916_ (.Y(_05630_),
    .B1(_05628_),
    .B2(_05629_),
    .A2(_05618_),
    .A1(_04401_));
 sg13g2_a21oi_1 _13917_ (.A1(_05475_),
    .A2(net95),
    .Y(_00137_),
    .B1(_05630_));
 sg13g2_mux2_1 _13918_ (.A0(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .A1(data_addr_o_16_),
    .S(net1011),
    .X(_05631_));
 sg13g2_and3_2 _13919_ (.X(_05632_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .B(_04487_),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ));
 sg13g2_buf_2 fanout875 (.A(rf_wdata_wb_8_),
    .X(net875));
 sg13g2_a21oi_1 _13921_ (.A1(_04083_),
    .A2(_05632_),
    .Y(_05634_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_16_ ));
 sg13g2_nand2_1 _13922_ (.Y(_05635_),
    .A(net313),
    .B(_05634_));
 sg13g2_o21ai_1 _13923_ (.B1(_05635_),
    .Y(_05636_),
    .A1(net309),
    .A2(_05631_));
 sg13g2_inv_1 _13924_ (.Y(_05637_),
    .A(\ex_block_i.alu_i.imd_val_q_i_48_ ));
 sg13g2_nor2_1 _13925_ (.A(data_addr_o_16_),
    .B(net1220),
    .Y(_05638_));
 sg13g2_a21oi_1 _13926_ (.A1(_05637_),
    .A2(net1220),
    .Y(_05639_),
    .B1(_05638_));
 sg13g2_o21ai_1 _13927_ (.B1(net1636),
    .Y(_05640_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ),
    .A2(net306));
 sg13g2_nand2_1 _13928_ (.Y(_05641_),
    .A(net1574),
    .B(_05640_));
 sg13g2_a221oi_1 _13929_ (.B2(net422),
    .C1(_05641_),
    .B1(_05639_),
    .A1(net1884),
    .Y(_05642_),
    .A2(_05619_));
 sg13g2_o21ai_1 _13930_ (.B1(_05642_),
    .Y(_05643_),
    .A1(_04066_),
    .A2(_05636_));
 sg13g2_a21oi_1 _13931_ (.A1(_05637_),
    .A2(net1478),
    .Y(_05644_),
    .B1(net337));
 sg13g2_a22oi_1 _13932_ (.Y(_05645_),
    .B1(net322),
    .B2(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .A2(_04039_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ));
 sg13g2_inv_1 _13933_ (.Y(_05646_),
    .A(_05587_));
 sg13g2_o21ai_1 _13934_ (.B1(_05592_),
    .Y(_05647_),
    .A1(_05581_),
    .A2(_05646_));
 sg13g2_and2_1 _13935_ (.A(net288),
    .B(net1873),
    .X(_05648_));
 sg13g2_and4_2 _13936_ (.A(net410),
    .B(_01529_),
    .C(_03949_),
    .D(_05648_),
    .X(_05649_));
 sg13g2_inv_1 _13937_ (.Y(_05650_),
    .A(_04231_));
 sg13g2_nand2_1 _13938_ (.Y(_05651_),
    .A(net1470),
    .B(net234));
 sg13g2_o21ai_1 _13939_ (.B1(_05651_),
    .Y(_05652_),
    .A1(_05650_),
    .A2(net242));
 sg13g2_nand2_1 _13940_ (.Y(_05653_),
    .A(net280),
    .B(net1380));
 sg13g2_o21ai_1 _13941_ (.B1(_05653_),
    .Y(_05654_),
    .A1(_04420_),
    .A2(net242));
 sg13g2_mux2_1 _13942_ (.A0(_05652_),
    .A1(_05654_),
    .S(net1870),
    .X(_05655_));
 sg13g2_a21oi_1 _13943_ (.A1(_04238_),
    .A2(net244),
    .Y(_05656_),
    .B1(_04239_));
 sg13g2_and2_1 _13944_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .B(net425),
    .X(_05657_));
 sg13g2_nand4_1 _13945_ (.B(_01529_),
    .C(_01658_),
    .A(net411),
    .Y(_05658_),
    .D(_05657_));
 sg13g2_mux2_2 _13946_ (.A0(_05655_),
    .A1(_05656_),
    .S(net1371),
    .X(_05659_));
 sg13g2_a21o_2 _13947_ (.A2(net426),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ),
    .B1(_05410_),
    .X(_05660_));
 sg13g2_a22oi_1 _13948_ (.Y(_05661_),
    .B1(net1322),
    .B2(net227),
    .A2(net1433),
    .A1(net165));
 sg13g2_a22oi_1 _13949_ (.Y(_05662_),
    .B1(net1435),
    .B2(net220),
    .A2(net247),
    .A1(net162));
 sg13g2_xnor2_1 _13950_ (.Y(_05663_),
    .A(net1341),
    .B(_05662_));
 sg13g2_xnor2_1 _13951_ (.Y(_05664_),
    .A(_05661_),
    .B(_05663_));
 sg13g2_xnor2_1 _13952_ (.Y(_05665_),
    .A(_05659_),
    .B(_05664_));
 sg13g2_xnor2_1 _13953_ (.Y(_05666_),
    .A(net1372),
    .B(_05665_));
 sg13g2_xor2_1 _13954_ (.B(_05534_),
    .A(net1329),
    .X(_05667_));
 sg13g2_xnor2_1 _13955_ (.Y(_05668_),
    .A(net1327),
    .B(_05528_));
 sg13g2_nand2_2 _13956_ (.Y(_05669_),
    .A(_05667_),
    .B(_05668_));
 sg13g2_xor2_1 _13957_ (.B(_05669_),
    .A(_05666_),
    .X(_05670_));
 sg13g2_o21ai_1 _13958_ (.B1(_05548_),
    .Y(_05671_),
    .A1(_05415_),
    .A2(_05549_));
 sg13g2_nand2_1 _13959_ (.Y(_05672_),
    .A(_05555_),
    .B(_05561_));
 sg13g2_nor2_1 _13960_ (.A(_05553_),
    .B(_05672_),
    .Y(_05673_));
 sg13g2_and2_1 _13961_ (.A(_05552_),
    .B(_05555_),
    .X(_05674_));
 sg13g2_or2_1 _13962_ (.X(_05675_),
    .B(_05555_),
    .A(_05552_));
 sg13g2_o21ai_1 _13963_ (.B1(_05675_),
    .Y(_05676_),
    .A1(_05561_),
    .A2(_05674_));
 sg13g2_nor2_1 _13964_ (.A(_05561_),
    .B(_05675_),
    .Y(_05677_));
 sg13g2_a221oi_1 _13965_ (.B2(_05550_),
    .C1(_05677_),
    .B1(_05676_),
    .A1(_05671_),
    .Y(_05678_),
    .A2(_05673_));
 sg13g2_xnor2_1 _13966_ (.Y(_05679_),
    .A(_05670_),
    .B(_05678_));
 sg13g2_nor2_1 _13967_ (.A(_05515_),
    .B(_05542_),
    .Y(_05680_));
 sg13g2_nand2_1 _13968_ (.Y(_05681_),
    .A(_05515_),
    .B(_05542_));
 sg13g2_o21ai_1 _13969_ (.B1(_05681_),
    .Y(_05682_),
    .A1(_05536_),
    .A2(_05680_));
 sg13g2_nand2_1 _13970_ (.Y(_05683_),
    .A(_05566_),
    .B(_05567_));
 sg13g2_nand4_1 _13971_ (.B(_01529_),
    .C(_03949_),
    .A(net411),
    .Y(_05684_),
    .D(_05648_));
 sg13g2_buf_2 fanout874 (.A(\register_file_i/_2817_ ),
    .X(net874));
 sg13g2_nand2_1 _13973_ (.Y(_05686_),
    .A(net1321),
    .B(net215));
 sg13g2_nor2_1 _13974_ (.A(net233),
    .B(net1257),
    .Y(_05687_));
 sg13g2_a22oi_1 _13975_ (.Y(_05688_),
    .B1(net90),
    .B2(net278),
    .A2(_05526_),
    .A1(net272));
 sg13g2_a22oi_1 _13976_ (.Y(_05689_),
    .B1(net134),
    .B2(net271),
    .A2(net1332),
    .A1(net267));
 sg13g2_xor2_1 _13977_ (.B(_05689_),
    .A(net1328),
    .X(_05690_));
 sg13g2_xnor2_1 _13978_ (.Y(_05691_),
    .A(_05688_),
    .B(_05690_));
 sg13g2_xnor2_1 _13979_ (.Y(_05692_),
    .A(_05687_),
    .B(_05691_));
 sg13g2_xor2_1 _13980_ (.B(_05539_),
    .A(net156),
    .X(_05693_));
 sg13g2_xnor2_1 _13981_ (.Y(_05694_),
    .A(net1336),
    .B(_05540_));
 sg13g2_xnor2_1 _13982_ (.Y(_05695_),
    .A(net1375),
    .B(_05537_));
 sg13g2_nand2_1 _13983_ (.Y(_05696_),
    .A(_05694_),
    .B(_05695_));
 sg13g2_nor2_1 _13984_ (.A(_05694_),
    .B(_05695_),
    .Y(_05697_));
 sg13g2_a21oi_1 _13985_ (.A1(_05693_),
    .A2(_05696_),
    .Y(_05698_),
    .B1(_05697_));
 sg13g2_a22oi_1 _13986_ (.Y(_05699_),
    .B1(net137),
    .B2(net254),
    .A2(_05047_),
    .A1(net1474));
 sg13g2_xnor2_1 _13987_ (.Y(_05700_),
    .A(_05054_),
    .B(_05699_));
 sg13g2_a22oi_1 _13988_ (.Y(_05701_),
    .B1(net248),
    .B2(net219),
    .A2(net1437),
    .A1(net161));
 sg13g2_buf_4 fanout873 (.X(net873),
    .A(net874));
 sg13g2_nand2_1 _13990_ (.Y(_05703_),
    .A(net265),
    .B(net139));
 sg13g2_o21ai_1 _13991_ (.B1(_05703_),
    .Y(_05704_),
    .A1(_04726_),
    .A2(_04791_));
 sg13g2_xor2_1 _13992_ (.B(_05704_),
    .A(_05701_),
    .X(_05705_));
 sg13g2_xnor2_1 _13993_ (.Y(_05706_),
    .A(_05700_),
    .B(_05705_));
 sg13g2_xor2_1 _13994_ (.B(_05706_),
    .A(_05698_),
    .X(_05707_));
 sg13g2_xnor2_1 _13995_ (.Y(_05708_),
    .A(_05692_),
    .B(_05707_));
 sg13g2_xnor2_1 _13996_ (.Y(_05709_),
    .A(_05682_),
    .B(_05708_));
 sg13g2_xnor2_1 _13997_ (.Y(_05710_),
    .A(_05679_),
    .B(_05709_));
 sg13g2_nor2_1 _13998_ (.A(_05571_),
    .B(_05578_),
    .Y(_05711_));
 sg13g2_a21oi_1 _13999_ (.A1(_05571_),
    .A2(_05578_),
    .Y(_05712_),
    .B1(_05509_));
 sg13g2_xor2_1 _14000_ (.B(_05543_),
    .A(_05515_),
    .X(_05713_));
 sg13g2_o21ai_1 _14001_ (.B1(_05713_),
    .Y(_05714_),
    .A1(_05711_),
    .A2(_05712_));
 sg13g2_nand2_1 _14002_ (.Y(_05715_),
    .A(_05439_),
    .B(_05448_));
 sg13g2_a21o_1 _14003_ (.A2(_05575_),
    .A1(_05573_),
    .B1(_05574_),
    .X(_05716_));
 sg13g2_nor2_1 _14004_ (.A(_05439_),
    .B(_05448_),
    .Y(_05717_));
 sg13g2_a21oi_2 _14005_ (.B1(_05717_),
    .Y(_05718_),
    .A2(_05716_),
    .A1(_05715_));
 sg13g2_nor2_1 _14006_ (.A(_05509_),
    .B(_05571_),
    .Y(_05719_));
 sg13g2_nand2_1 _14007_ (.Y(_05720_),
    .A(_05718_),
    .B(_05719_));
 sg13g2_nand2_1 _14008_ (.Y(_05721_),
    .A(_05714_),
    .B(_05720_));
 sg13g2_and2_1 _14009_ (.A(_05713_),
    .B(_05718_),
    .X(_05722_));
 sg13g2_inv_1 _14010_ (.Y(_05723_),
    .A(_05509_));
 sg13g2_nand2b_1 _14011_ (.Y(_05724_),
    .B(_05544_),
    .A_N(_05718_));
 sg13g2_o21ai_1 _14012_ (.B1(_05724_),
    .Y(_05725_),
    .A1(_05564_),
    .A2(_05722_));
 sg13g2_nor2_1 _14013_ (.A(_05564_),
    .B(_05713_),
    .Y(_05726_));
 sg13g2_a22oi_1 _14014_ (.Y(_05727_),
    .B1(_05726_),
    .B2(_05578_),
    .A2(_05725_),
    .A1(_05571_));
 sg13g2_inv_1 _14015_ (.Y(_05728_),
    .A(_05571_));
 sg13g2_or4_1 _14016_ (.A(_05564_),
    .B(_05728_),
    .C(_05713_),
    .D(_05718_),
    .X(_05729_));
 sg13g2_o21ai_1 _14017_ (.B1(_05729_),
    .Y(_05730_),
    .A1(_05723_),
    .A2(_05727_));
 sg13g2_a221oi_1 _14018_ (.B2(_05719_),
    .C1(_05730_),
    .B1(_05722_),
    .A1(_05564_),
    .Y(_05731_),
    .A2(_05721_));
 sg13g2_xnor2_1 _14019_ (.Y(_05732_),
    .A(_05710_),
    .B(_05731_));
 sg13g2_xnor2_1 _14020_ (.Y(_05733_),
    .A(_05647_),
    .B(_05732_));
 sg13g2_xor2_1 _14021_ (.B(_05733_),
    .A(_05645_),
    .X(_05734_));
 sg13g2_a21oi_1 _14022_ (.A1(_05266_),
    .A2(_05468_),
    .Y(_05735_),
    .B1(_05467_));
 sg13g2_o21ai_1 _14023_ (.B1(_05465_),
    .Y(_05736_),
    .A1(_05503_),
    .A2(_05735_));
 sg13g2_o21ai_1 _14024_ (.B1(_05605_),
    .Y(_05737_),
    .A1(_05506_),
    .A2(_05604_));
 sg13g2_nor2b_1 _14025_ (.A(net35),
    .B_N(_05737_),
    .Y(_05738_));
 sg13g2_nor2_1 _14026_ (.A(_05506_),
    .B(_05605_),
    .Y(_05739_));
 sg13g2_nor2_1 _14027_ (.A(_05738_),
    .B(_05739_),
    .Y(_05740_));
 sg13g2_and2_1 _14028_ (.A(_05506_),
    .B(_05604_),
    .X(_05741_));
 sg13g2_a21o_1 _14029_ (.A2(_05605_),
    .A1(_05506_),
    .B1(_05604_),
    .X(_05742_));
 sg13g2_a21oi_1 _14030_ (.A1(net35),
    .A2(_05742_),
    .Y(_05743_),
    .B1(_05741_));
 sg13g2_inv_1 _14031_ (.Y(_05744_),
    .A(_05743_));
 sg13g2_nor2b_1 _14032_ (.A(net35),
    .B_N(_05739_),
    .Y(_05745_));
 sg13g2_a221oi_1 _14033_ (.B2(_05736_),
    .C1(_05745_),
    .B1(_05744_),
    .A1(net35),
    .Y(_05746_),
    .A2(_05741_));
 sg13g2_o21ai_1 _14034_ (.B1(_05746_),
    .Y(_05747_),
    .A1(_05736_),
    .A2(_05740_));
 sg13g2_xnor2_1 _14035_ (.Y(_05748_),
    .A(_05734_),
    .B(_05747_));
 sg13g2_nor2_1 _14036_ (.A(net1542),
    .B(_04064_),
    .Y(_05749_));
 sg13g2_a21oi_1 _14037_ (.A1(net1542),
    .A2(_05748_),
    .Y(_05750_),
    .B1(_05749_));
 sg13g2_buf_2 fanout872 (.A(\register_file_i/_2817_ ),
    .X(net872));
 sg13g2_a22oi_1 _14039_ (.Y(_05752_),
    .B1(_05750_),
    .B2(net343),
    .A2(_05644_),
    .A1(_05643_));
 sg13g2_nor3_1 _14040_ (.A(net376),
    .B(net94),
    .C(_05752_),
    .Y(_05753_));
 sg13g2_a21o_1 _14041_ (.A2(net96),
    .A1(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .B1(_05753_),
    .X(_00138_));
 sg13g2_a21oi_1 _14042_ (.A1(_05605_),
    .A2(net35),
    .Y(_05754_),
    .B1(_05604_));
 sg13g2_xor2_1 _14043_ (.B(_05754_),
    .A(_05733_),
    .X(_05755_));
 sg13g2_nand2b_1 _14044_ (.Y(_05756_),
    .B(_05755_),
    .A_N(_05645_));
 sg13g2_nor2_1 _14045_ (.A(_05268_),
    .B(_05499_),
    .Y(_05757_));
 sg13g2_a21oi_1 _14046_ (.A1(_05268_),
    .A2(_05499_),
    .Y(_05758_),
    .B1(_05354_));
 sg13g2_a22oi_1 _14047_ (.Y(_05759_),
    .B1(_05507_),
    .B2(_05614_),
    .A2(_05460_),
    .A1(_05386_));
 sg13g2_o21ai_1 _14048_ (.B1(_05759_),
    .Y(_05760_),
    .A1(_05757_),
    .A2(_05758_));
 sg13g2_a21o_1 _14049_ (.A2(_05613_),
    .A1(_05603_),
    .B1(_05594_),
    .X(_05761_));
 sg13g2_o21ai_1 _14050_ (.B1(_05761_),
    .Y(_05762_),
    .A1(_05603_),
    .A2(net35));
 sg13g2_mux2_1 _14051_ (.A0(_05604_),
    .A1(_05762_),
    .S(_05734_),
    .X(_05763_));
 sg13g2_a21oi_1 _14052_ (.A1(_05463_),
    .A2(_05464_),
    .Y(_05764_),
    .B1(_05386_));
 sg13g2_nor2_1 _14053_ (.A(_05764_),
    .B(_05506_),
    .Y(_05765_));
 sg13g2_inv_1 _14054_ (.Y(_05766_),
    .A(_05603_));
 sg13g2_and2_1 _14055_ (.A(_05766_),
    .B(_05734_),
    .X(_05767_));
 sg13g2_nor2_1 _14056_ (.A(_05766_),
    .B(_05734_),
    .Y(_05768_));
 sg13g2_mux2_1 _14057_ (.A0(_05767_),
    .A1(_05768_),
    .S(net35),
    .X(_05769_));
 sg13g2_nand2b_1 _14058_ (.Y(_05770_),
    .B(_05769_),
    .A_N(_05594_));
 sg13g2_xnor2_1 _14059_ (.Y(_05771_),
    .A(_05766_),
    .B(_05613_));
 sg13g2_nand3b_1 _14060_ (.B(_05771_),
    .C(_05594_),
    .Y(_05772_),
    .A_N(_05734_));
 sg13g2_a22oi_1 _14061_ (.Y(_05773_),
    .B1(_05770_),
    .B2(_05772_),
    .A2(_05506_),
    .A1(_05764_));
 sg13g2_a21o_1 _14062_ (.A2(_05765_),
    .A1(_05763_),
    .B1(_05773_),
    .X(_05774_));
 sg13g2_nand2_1 _14063_ (.Y(_05775_),
    .A(_05760_),
    .B(_05774_));
 sg13g2_and2_1 _14064_ (.A(_05756_),
    .B(_05775_),
    .X(_05776_));
 sg13g2_nand2_2 _14065_ (.Y(_05777_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ),
    .B(_04039_));
 sg13g2_nand2_1 _14066_ (.Y(_05778_),
    .A(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .B(net320));
 sg13g2_a21oi_1 _14067_ (.A1(_05581_),
    .A2(_05612_),
    .Y(_05779_),
    .B1(_05732_));
 sg13g2_nand2_1 _14068_ (.Y(_05780_),
    .A(_05646_),
    .B(_05732_));
 sg13g2_o21ai_1 _14069_ (.B1(_05780_),
    .Y(_05781_),
    .A1(_05603_),
    .A2(_05779_));
 sg13g2_nor2b_1 _14070_ (.A(_05606_),
    .B_N(_05733_),
    .Y(_05782_));
 sg13g2_and2_1 _14071_ (.A(_05271_),
    .B(_05607_),
    .X(_05783_));
 sg13g2_a221oi_1 _14072_ (.B2(_05592_),
    .C1(_05766_),
    .B1(_05732_),
    .A1(_05581_),
    .Y(_05784_),
    .A2(_05612_));
 sg13g2_nor2_1 _14073_ (.A(_05646_),
    .B(_05732_),
    .Y(_05785_));
 sg13g2_nor2_1 _14074_ (.A(_05581_),
    .B(_05612_),
    .Y(_05786_));
 sg13g2_nor3_1 _14075_ (.A(_05784_),
    .B(_05785_),
    .C(_05786_),
    .Y(_05787_));
 sg13g2_a221oi_1 _14076_ (.B2(_05783_),
    .C1(_05787_),
    .B1(_05782_),
    .A1(_05592_),
    .Y(_05788_),
    .A2(_05781_));
 sg13g2_buf_4 fanout871 (.X(net871),
    .A(net872));
 sg13g2_nand2_1 _14078_ (.Y(_05790_),
    .A(_05544_),
    .B(_05578_));
 sg13g2_nor2_1 _14079_ (.A(_05544_),
    .B(_05578_),
    .Y(_05791_));
 sg13g2_a21oi_1 _14080_ (.A1(_05564_),
    .A2(_05790_),
    .Y(_05792_),
    .B1(_05791_));
 sg13g2_nand2_1 _14081_ (.Y(_05793_),
    .A(_05564_),
    .B(_05722_));
 sg13g2_o21ai_1 _14082_ (.B1(_05793_),
    .Y(_05794_),
    .A1(_05571_),
    .A2(_05792_));
 sg13g2_nor3_1 _14083_ (.A(_05571_),
    .B(_05544_),
    .C(_05578_),
    .Y(_05795_));
 sg13g2_a22oi_1 _14084_ (.Y(_05796_),
    .B1(_05795_),
    .B2(_05564_),
    .A2(_05794_),
    .A1(_05723_));
 sg13g2_o21ai_1 _14085_ (.B1(_05796_),
    .Y(_05797_),
    .A1(_05710_),
    .A2(_05730_));
 sg13g2_buf_2 fanout870 (.A(net872),
    .X(net870));
 sg13g2_o21ai_1 _14087_ (.B1(_05688_),
    .Y(_05799_),
    .A1(net233),
    .A2(net1373));
 sg13g2_nor3_1 _14088_ (.A(net233),
    .B(_05688_),
    .C(net1257),
    .Y(_05800_));
 sg13g2_a221oi_1 _14089_ (.B2(_05799_),
    .C1(_05800_),
    .B1(_05690_),
    .A1(net1327),
    .Y(_05801_),
    .A2(_05688_));
 sg13g2_nor2_1 _14090_ (.A(_03911_),
    .B(net286),
    .Y(_05802_));
 sg13g2_nor2b_1 _14091_ (.A(net1501),
    .B_N(net279),
    .Y(_05803_));
 sg13g2_and4_2 _14092_ (.A(net410),
    .B(_01529_),
    .C(_01658_),
    .D(_05657_),
    .X(_05804_));
 sg13g2_buf_4 fanout869 (.X(net869),
    .A(net872));
 sg13g2_mux4_1 _14094_ (.S0(net1869),
    .A0(net286),
    .A1(net1501),
    .A2(_05802_),
    .A3(_05803_),
    .S1(_05804_),
    .X(_05806_));
 sg13g2_buf_4 fanout868 (.X(net868),
    .A(\register_file_i/_2870_ ));
 sg13g2_a22oi_1 _14096_ (.Y(_05808_),
    .B1(net243),
    .B2(net227),
    .A2(net1322),
    .A1(net165));
 sg13g2_xnor2_1 _14097_ (.Y(_05809_),
    .A(_04354_),
    .B(_05808_));
 sg13g2_xnor2_1 _14098_ (.Y(_05810_),
    .A(_05806_),
    .B(_05809_));
 sg13g2_a22oi_1 _14099_ (.Y(_05811_),
    .B1(net1433),
    .B2(net220),
    .A2(net1435),
    .A1(net163));
 sg13g2_xnor2_1 _14100_ (.Y(_05812_),
    .A(_05206_),
    .B(_05811_));
 sg13g2_xnor2_1 _14101_ (.Y(_05813_),
    .A(net223),
    .B(_05662_));
 sg13g2_xnor2_1 _14102_ (.Y(_05814_),
    .A(net167),
    .B(_05661_));
 sg13g2_nor2_1 _14103_ (.A(_05813_),
    .B(_05814_),
    .Y(_05815_));
 sg13g2_a21oi_1 _14104_ (.A1(_05813_),
    .A2(_05814_),
    .Y(_05816_),
    .B1(_05659_));
 sg13g2_nor2_1 _14105_ (.A(_05815_),
    .B(_05816_),
    .Y(_05817_));
 sg13g2_xnor2_1 _14106_ (.Y(_05818_),
    .A(_05812_),
    .B(_05817_));
 sg13g2_xnor2_1 _14107_ (.Y(_05819_),
    .A(_05810_),
    .B(_05818_));
 sg13g2_xnor2_1 _14108_ (.Y(_05820_),
    .A(_05801_),
    .B(_05819_));
 sg13g2_or2_1 _14109_ (.X(_05821_),
    .B(_05665_),
    .A(net215));
 sg13g2_and2_1 _14110_ (.A(net215),
    .B(_05665_),
    .X(_05822_));
 sg13g2_a21oi_2 _14111_ (.B1(_05822_),
    .Y(_05823_),
    .A2(_05821_),
    .A1(_05676_));
 sg13g2_xnor2_1 _14112_ (.Y(_05824_),
    .A(_05820_),
    .B(_05823_));
 sg13g2_nor2_1 _14113_ (.A(net276),
    .B(net1257),
    .Y(_05825_));
 sg13g2_a22oi_1 _14114_ (.Y(_05826_),
    .B1(net90),
    .B2(net274),
    .A2(_05526_),
    .A1(net270));
 sg13g2_xnor2_1 _14115_ (.Y(_05827_),
    .A(_05825_),
    .B(_05826_));
 sg13g2_a22oi_1 _14116_ (.Y(_05828_),
    .B1(net134),
    .B2(net268),
    .A2(net1332),
    .A1(net253));
 sg13g2_xor2_1 _14117_ (.B(_05828_),
    .A(net1328),
    .X(_05829_));
 sg13g2_xnor2_1 _14118_ (.Y(_05830_),
    .A(_05827_),
    .B(_05829_));
 sg13g2_xnor2_1 _14119_ (.Y(_05831_),
    .A(net1468),
    .B(net1464));
 sg13g2_xor2_1 _14120_ (.B(net1498),
    .A(net1495),
    .X(_05832_));
 sg13g2_nor2_1 _14121_ (.A(net1865),
    .B(_05832_),
    .Y(_05833_));
 sg13g2_a21oi_2 _14122_ (.B1(_05833_),
    .Y(_05834_),
    .A2(_05831_),
    .A1(net1865));
 sg13g2_xnor2_1 _14123_ (.Y(_05835_),
    .A(net158),
    .B(_05834_));
 sg13g2_buf_2 fanout867 (.A(net868),
    .X(net867));
 sg13g2_buf_2 fanout866 (.A(net867),
    .X(net866));
 sg13g2_a22oi_1 _14126_ (.Y(_05838_),
    .B1(net138),
    .B2(net1474),
    .A2(_05047_),
    .A1(net264));
 sg13g2_xnor2_1 _14127_ (.Y(_05839_),
    .A(_05835_),
    .B(_05838_));
 sg13g2_a22oi_1 _14128_ (.Y(_05840_),
    .B1(net140),
    .B2(net251),
    .A2(_04786_),
    .A1(net1340));
 sg13g2_and2_1 _14129_ (.A(net217),
    .B(net246),
    .X(_05841_));
 sg13g2_a21o_1 _14130_ (.A2(net249),
    .A1(_04589_),
    .B1(_05841_),
    .X(_05842_));
 sg13g2_xor2_1 _14131_ (.B(_05842_),
    .A(_05840_),
    .X(_05843_));
 sg13g2_xnor2_1 _14132_ (.Y(_05844_),
    .A(_05839_),
    .B(_05843_));
 sg13g2_inv_1 _14133_ (.Y(_05845_),
    .A(_05844_));
 sg13g2_buf_4 fanout865 (.X(net865),
    .A(net867));
 sg13g2_xor2_1 _14135_ (.B(_05704_),
    .A(_04807_),
    .X(_05847_));
 sg13g2_buf_4 fanout864 (.X(net864),
    .A(net868));
 sg13g2_xnor2_1 _14137_ (.Y(_05849_),
    .A(_05041_),
    .B(_05699_));
 sg13g2_xnor2_1 _14138_ (.Y(_05850_),
    .A(net158),
    .B(_05701_));
 sg13g2_a21oi_1 _14139_ (.A1(_05847_),
    .A2(_05849_),
    .Y(_05851_),
    .B1(_05850_));
 sg13g2_nor2_1 _14140_ (.A(_05847_),
    .B(_05849_),
    .Y(_05852_));
 sg13g2_nor2_2 _14141_ (.A(_05851_),
    .B(_05852_),
    .Y(_05853_));
 sg13g2_xnor2_1 _14142_ (.Y(_05854_),
    .A(_05845_),
    .B(_05853_));
 sg13g2_xnor2_1 _14143_ (.Y(_05855_),
    .A(_05830_),
    .B(_05854_));
 sg13g2_o21ai_1 _14144_ (.B1(_05696_),
    .Y(_05856_),
    .A1(_05693_),
    .A2(_05697_));
 sg13g2_o21ai_1 _14145_ (.B1(_05692_),
    .Y(_05857_),
    .A1(_05706_),
    .A2(_05856_));
 sg13g2_inv_1 _14146_ (.Y(_05858_),
    .A(_05857_));
 sg13g2_a21oi_2 _14147_ (.B1(_05858_),
    .Y(_05859_),
    .A2(_05856_),
    .A1(_05706_));
 sg13g2_xnor2_1 _14148_ (.Y(_05860_),
    .A(_05855_),
    .B(_05859_));
 sg13g2_xnor2_1 _14149_ (.Y(_05861_),
    .A(_05824_),
    .B(_05860_));
 sg13g2_xnor2_1 _14150_ (.Y(_05862_),
    .A(net1081),
    .B(_05861_));
 sg13g2_nor3_1 _14151_ (.A(_05553_),
    .B(_05550_),
    .C(_05669_),
    .Y(_05863_));
 sg13g2_nand2_1 _14152_ (.Y(_05864_),
    .A(_05552_),
    .B(_05562_));
 sg13g2_o21ai_1 _14153_ (.B1(_05864_),
    .Y(_05865_),
    .A1(_05672_),
    .A2(_05863_));
 sg13g2_nand3_1 _14154_ (.B(_05555_),
    .C(_05561_),
    .A(_05552_),
    .Y(_05866_));
 sg13g2_a221oi_1 _14155_ (.B2(_05550_),
    .C1(_05677_),
    .B1(_05676_),
    .A1(_05669_),
    .Y(_05867_),
    .A2(_05866_));
 sg13g2_o21ai_1 _14156_ (.B1(_05669_),
    .Y(_05868_),
    .A1(_05550_),
    .A2(_05677_));
 sg13g2_o21ai_1 _14157_ (.B1(_05868_),
    .Y(_05869_),
    .A1(_05666_),
    .A2(_05867_));
 sg13g2_a21oi_1 _14158_ (.A1(_05666_),
    .A2(_05865_),
    .Y(_05870_),
    .B1(_05869_));
 sg13g2_inv_1 _14159_ (.Y(_05871_),
    .A(_05870_));
 sg13g2_inv_1 _14160_ (.Y(_05872_),
    .A(_05542_));
 sg13g2_a21o_1 _14161_ (.A2(_05514_),
    .A1(_05510_),
    .B1(_05513_),
    .X(_05873_));
 sg13g2_a21oi_1 _14162_ (.A1(_05872_),
    .A2(_05873_),
    .Y(_05874_),
    .B1(_05536_));
 sg13g2_nor2_1 _14163_ (.A(_05872_),
    .B(_05873_),
    .Y(_05875_));
 sg13g2_nor2_1 _14164_ (.A(_05874_),
    .B(_05875_),
    .Y(_05876_));
 sg13g2_inv_1 _14165_ (.Y(_05877_),
    .A(_05876_));
 sg13g2_nand2_1 _14166_ (.Y(_05878_),
    .A(_05679_),
    .B(_05877_));
 sg13g2_nor2_1 _14167_ (.A(_05679_),
    .B(_05877_),
    .Y(_05879_));
 sg13g2_a21o_1 _14168_ (.A2(_05878_),
    .A1(_05708_),
    .B1(_05879_),
    .X(_05880_));
 sg13g2_xnor2_1 _14169_ (.Y(_05881_),
    .A(_05871_),
    .B(_05880_));
 sg13g2_xnor2_1 _14170_ (.Y(_05882_),
    .A(_05862_),
    .B(_05881_));
 sg13g2_xnor2_1 _14171_ (.Y(_05883_),
    .A(_05788_),
    .B(_05882_));
 sg13g2_a21oi_1 _14172_ (.A1(_05777_),
    .A2(_05778_),
    .Y(_05884_),
    .B1(_05883_));
 sg13g2_and3_1 _14173_ (.X(_05885_),
    .A(_05777_),
    .B(_05778_),
    .C(_05883_));
 sg13g2_nor2_1 _14174_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sg13g2_xnor2_1 _14175_ (.Y(_05887_),
    .A(_05776_),
    .B(_05886_));
 sg13g2_nand2_1 _14176_ (.Y(_05888_),
    .A(net1542),
    .B(_05887_));
 sg13g2_o21ai_1 _14177_ (.B1(_05888_),
    .Y(_05889_),
    .A1(net1542),
    .A2(_04185_));
 sg13g2_nand2_1 _14178_ (.Y(_05890_),
    .A(net1184),
    .B(_05889_));
 sg13g2_nand2_1 _14179_ (.Y(_05891_),
    .A(net554),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ));
 sg13g2_nor2_2 _14180_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ),
    .B(_05891_),
    .Y(_05892_));
 sg13g2_a21oi_1 _14181_ (.A1(_04083_),
    .A2(_05892_),
    .Y(_05893_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_17_ ));
 sg13g2_nand2_1 _14182_ (.Y(_05894_),
    .A(data_addr_o_17_),
    .B(net1012));
 sg13g2_o21ai_1 _14183_ (.B1(_05894_),
    .Y(_05895_),
    .A1(_02576_),
    .A2(net1012));
 sg13g2_nor2_1 _14184_ (.A(net312),
    .B(_05895_),
    .Y(_05896_));
 sg13g2_a21oi_1 _14185_ (.A1(net316),
    .A2(_05893_),
    .Y(_05897_),
    .B1(_05896_));
 sg13g2_nand2_1 _14186_ (.Y(_05898_),
    .A(data_addr_o_17_),
    .B(net1264));
 sg13g2_o21ai_1 _14187_ (.B1(_05898_),
    .Y(_05899_),
    .A1(_02576_),
    .A2(net1264));
 sg13g2_nand2_1 _14188_ (.Y(_05900_),
    .A(net422),
    .B(_05899_));
 sg13g2_o21ai_1 _14189_ (.B1(net1638),
    .Y(_05901_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ),
    .A2(net305));
 sg13g2_nand3_1 _14190_ (.B(_05900_),
    .C(_05901_),
    .A(net1574),
    .Y(_05902_));
 sg13g2_a221oi_1 _14191_ (.B2(net1890),
    .C1(_05902_),
    .B1(_05897_),
    .A1(net1884),
    .Y(_05903_),
    .A2(_05631_));
 sg13g2_o21ai_1 _14192_ (.B1(net1188),
    .Y(_05904_),
    .A1(net338),
    .A2(_05903_));
 sg13g2_o21ai_1 _14193_ (.B1(_05904_),
    .Y(_05905_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .A2(net1572));
 sg13g2_a22oi_1 _14194_ (.Y(_00139_),
    .B1(_05890_),
    .B2(_05905_),
    .A2(net96),
    .A1(_02576_));
 sg13g2_mux2_1 _14195_ (.A0(net1507),
    .A1(data_addr_o_4_),
    .S(net1451),
    .X(_05906_));
 sg13g2_mux2_1 _14196_ (.A0(_05906_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_4_ ),
    .S(net1223),
    .X(_00140_));
 sg13g2_a21o_1 _14197_ (.A2(_05778_),
    .A1(_05777_),
    .B1(_05883_),
    .X(_05907_));
 sg13g2_a21oi_1 _14198_ (.A1(_05776_),
    .A2(_05907_),
    .Y(_05908_),
    .B1(_05885_));
 sg13g2_nor2_1 _14199_ (.A(_01658_),
    .B(_03949_),
    .Y(_05909_));
 sg13g2_or3_1 _14200_ (.A(_01530_),
    .B(_05777_),
    .C(_05909_),
    .X(_05910_));
 sg13g2_nand2_1 _14201_ (.Y(_05911_),
    .A(\ex_block_i.alu_i.imd_val_q_i_50_ ),
    .B(net320));
 sg13g2_nor2_1 _14202_ (.A(net1873),
    .B(_04054_),
    .Y(_05912_));
 sg13g2_a21oi_1 _14203_ (.A1(net1568),
    .A2(_05911_),
    .Y(_05913_),
    .B1(net1566));
 sg13g2_nand2_1 _14204_ (.Y(_05914_),
    .A(_05859_),
    .B(_05824_));
 sg13g2_nor2_1 _14205_ (.A(_05859_),
    .B(_05824_),
    .Y(_05915_));
 sg13g2_a21o_1 _14206_ (.A2(_05914_),
    .A1(_05855_),
    .B1(_05915_),
    .X(_05916_));
 sg13g2_inv_1 _14207_ (.Y(_05917_),
    .A(_05819_));
 sg13g2_o21ai_1 _14208_ (.B1(_05801_),
    .Y(_05918_),
    .A1(_05917_),
    .A2(_05823_));
 sg13g2_nand2_1 _14209_ (.Y(_05919_),
    .A(_05917_),
    .B(_05823_));
 sg13g2_nand2_1 _14210_ (.Y(_05920_),
    .A(_05918_),
    .B(_05919_));
 sg13g2_inv_1 _14211_ (.Y(_05921_),
    .A(_05815_));
 sg13g2_and2_1 _14212_ (.A(_05813_),
    .B(_05814_),
    .X(_05922_));
 sg13g2_a21oi_2 _14213_ (.B1(_05922_),
    .Y(_05923_),
    .A2(_05921_),
    .A1(_05659_));
 sg13g2_mux4_1 _14214_ (.S0(net1869),
    .A0(net234),
    .A1(net1380),
    .A2(_05651_),
    .A3(_05653_),
    .S1(_05804_),
    .X(_05924_));
 sg13g2_nand2_1 _14215_ (.Y(_05925_),
    .A(_05809_),
    .B(_05812_));
 sg13g2_nor2_1 _14216_ (.A(_05809_),
    .B(_05812_),
    .Y(_05926_));
 sg13g2_a21oi_1 _14217_ (.A1(net89),
    .A2(_05925_),
    .Y(_05927_),
    .B1(_05926_));
 sg13g2_nor2_1 _14218_ (.A(net89),
    .B(_05925_),
    .Y(_05928_));
 sg13g2_a22oi_1 _14219_ (.Y(_05929_),
    .B1(_05928_),
    .B2(_05923_),
    .A2(_05926_),
    .A1(net89));
 sg13g2_o21ai_1 _14220_ (.B1(_05929_),
    .Y(_05930_),
    .A1(_05923_),
    .A2(_05927_));
 sg13g2_o21ai_1 _14221_ (.B1(_05826_),
    .Y(_05931_),
    .A1(net276),
    .A2(net1372));
 sg13g2_nor3_1 _14222_ (.A(net276),
    .B(net1257),
    .C(_05826_),
    .Y(_05932_));
 sg13g2_a221oi_1 _14223_ (.B2(_05931_),
    .C1(_05932_),
    .B1(_05829_),
    .A1(net1327),
    .Y(_05933_),
    .A2(_05826_));
 sg13g2_buf_4 fanout863 (.X(net863),
    .A(net868));
 sg13g2_nand2_1 _14225_ (.Y(_05935_),
    .A(net164),
    .B(net243));
 sg13g2_o21ai_1 _14226_ (.B1(_05935_),
    .Y(_05936_),
    .A1(_04255_),
    .A2(net1371));
 sg13g2_a22oi_1 _14227_ (.Y(_05937_),
    .B1(net1323),
    .B2(net220),
    .A2(net1433),
    .A1(net163));
 sg13g2_xnor2_1 _14228_ (.Y(_05938_),
    .A(net1341),
    .B(_05937_));
 sg13g2_xnor2_1 _14229_ (.Y(_05939_),
    .A(_05936_),
    .B(_05938_));
 sg13g2_xnor2_1 _14230_ (.Y(_05940_),
    .A(_05933_),
    .B(_05939_));
 sg13g2_xnor2_1 _14231_ (.Y(_05941_),
    .A(_05930_),
    .B(_05940_));
 sg13g2_nor2_1 _14232_ (.A(net272),
    .B(net1257),
    .Y(_05942_));
 sg13g2_a22oi_1 _14233_ (.Y(_05943_),
    .B1(net90),
    .B2(net271),
    .A2(_05526_),
    .A1(net267));
 sg13g2_xnor2_1 _14234_ (.Y(_05944_),
    .A(_05942_),
    .B(_05943_));
 sg13g2_a22oi_1 _14235_ (.Y(_05945_),
    .B1(net134),
    .B2(net254),
    .A2(net1331),
    .A1(net1473));
 sg13g2_xnor2_1 _14236_ (.Y(_05946_),
    .A(net1328),
    .B(_05945_));
 sg13g2_xnor2_1 _14237_ (.Y(_05947_),
    .A(_05944_),
    .B(_05946_));
 sg13g2_xor2_1 _14238_ (.B(_05842_),
    .A(net156),
    .X(_05948_));
 sg13g2_xnor2_1 _14239_ (.Y(_05949_),
    .A(net1375),
    .B(_05838_));
 sg13g2_xnor2_1 _14240_ (.Y(_05950_),
    .A(net1336),
    .B(_05840_));
 sg13g2_o21ai_1 _14241_ (.B1(_05950_),
    .Y(_05951_),
    .A1(_05948_),
    .A2(_05949_));
 sg13g2_nand2_1 _14242_ (.Y(_05952_),
    .A(_05948_),
    .B(_05949_));
 sg13g2_nand2_1 _14243_ (.Y(_05953_),
    .A(_05951_),
    .B(_05952_));
 sg13g2_and2_1 _14244_ (.A(net252),
    .B(net1334),
    .X(_05954_));
 sg13g2_a21o_1 _14245_ (.A2(net138),
    .A1(_04608_),
    .B1(_05954_),
    .X(_05955_));
 sg13g2_xor2_1 _14246_ (.B(_05955_),
    .A(_05835_),
    .X(_05956_));
 sg13g2_buf_4 fanout862 (.X(net862),
    .A(\register_file_i/_2879_ ));
 sg13g2_a22oi_1 _14248_ (.Y(_05958_),
    .B1(net249),
    .B2(net1339),
    .A2(net141),
    .A1(net1437));
 sg13g2_buf_4 fanout861 (.X(net861),
    .A(net862));
 sg13g2_a22oi_1 _14250_ (.Y(_05960_),
    .B1(net1436),
    .B2(net218),
    .A2(net247),
    .A1(net160));
 sg13g2_xnor2_1 _14251_ (.Y(_05961_),
    .A(_05958_),
    .B(_05960_));
 sg13g2_xnor2_1 _14252_ (.Y(_05962_),
    .A(_05956_),
    .B(_05961_));
 sg13g2_xor2_1 _14253_ (.B(_05962_),
    .A(_05953_),
    .X(_05963_));
 sg13g2_xnor2_1 _14254_ (.Y(_05964_),
    .A(_05947_),
    .B(_05963_));
 sg13g2_o21ai_1 _14255_ (.B1(_05830_),
    .Y(_05965_),
    .A1(_05845_),
    .A2(_05853_));
 sg13g2_nand2_1 _14256_ (.Y(_05966_),
    .A(_05845_),
    .B(_05853_));
 sg13g2_and2_1 _14257_ (.A(_05965_),
    .B(_05966_),
    .X(_05967_));
 sg13g2_xnor2_1 _14258_ (.Y(_05968_),
    .A(_05964_),
    .B(_05967_));
 sg13g2_xnor2_1 _14259_ (.Y(_05969_),
    .A(_05941_),
    .B(_05968_));
 sg13g2_xnor2_1 _14260_ (.Y(_05970_),
    .A(_05920_),
    .B(_05969_));
 sg13g2_xor2_1 _14261_ (.B(_05970_),
    .A(_05916_),
    .X(_05971_));
 sg13g2_inv_1 _14262_ (.Y(_05972_),
    .A(_05708_));
 sg13g2_o21ai_1 _14263_ (.B1(_05972_),
    .Y(_05973_),
    .A1(_05679_),
    .A2(_05877_));
 sg13g2_and3_1 _14264_ (.X(_05974_),
    .A(_05871_),
    .B(_05878_),
    .C(_05973_));
 sg13g2_nand2b_1 _14265_ (.Y(_05975_),
    .B(_05974_),
    .A_N(_05861_));
 sg13g2_nor2_1 _14266_ (.A(net1081),
    .B(_05975_),
    .Y(_05976_));
 sg13g2_nor2_2 _14267_ (.A(_05871_),
    .B(_05880_),
    .Y(_05977_));
 sg13g2_nand2_1 _14268_ (.Y(_05978_),
    .A(_05861_),
    .B(_05977_));
 sg13g2_nand2b_1 _14269_ (.Y(_05979_),
    .B(_05861_),
    .A_N(_05974_));
 sg13g2_inv_1 _14270_ (.Y(_05980_),
    .A(_05979_));
 sg13g2_o21ai_1 _14271_ (.B1(net1081),
    .Y(_05981_),
    .A1(_05977_),
    .A2(_05980_));
 sg13g2_nand2_1 _14272_ (.Y(_05982_),
    .A(_05978_),
    .B(_05981_));
 sg13g2_nor2_1 _14273_ (.A(_05976_),
    .B(_05982_),
    .Y(_05983_));
 sg13g2_nor2b_1 _14274_ (.A(_05978_),
    .B_N(net1081),
    .Y(_05984_));
 sg13g2_nor2_1 _14275_ (.A(_05861_),
    .B(_05977_),
    .Y(_05985_));
 sg13g2_nor2_1 _14276_ (.A(_05974_),
    .B(_05985_),
    .Y(_05986_));
 sg13g2_o21ai_1 _14277_ (.B1(_05975_),
    .Y(_05987_),
    .A1(net1081),
    .A2(_05986_));
 sg13g2_nor2_1 _14278_ (.A(_05984_),
    .B(_05987_),
    .Y(_05988_));
 sg13g2_mux2_1 _14279_ (.A0(_05983_),
    .A1(_05988_),
    .S(_05788_),
    .X(_05989_));
 sg13g2_xnor2_1 _14280_ (.Y(_05990_),
    .A(_05971_),
    .B(_05989_));
 sg13g2_nand2b_1 _14281_ (.Y(_05991_),
    .B(_05990_),
    .A_N(_05913_));
 sg13g2_and2_1 _14282_ (.A(_05788_),
    .B(_05987_),
    .X(_05992_));
 sg13g2_nor2b_1 _14283_ (.A(_05788_),
    .B_N(_05982_),
    .Y(_05993_));
 sg13g2_nor4_1 _14284_ (.A(_05984_),
    .B(_05976_),
    .C(_05992_),
    .D(_05993_),
    .Y(_05994_));
 sg13g2_xor2_1 _14285_ (.B(_05994_),
    .A(_05971_),
    .X(_05995_));
 sg13g2_nand2_1 _14286_ (.Y(_05996_),
    .A(_05913_),
    .B(_05995_));
 sg13g2_nand2_1 _14287_ (.Y(_05997_),
    .A(_05991_),
    .B(_05996_));
 sg13g2_xnor2_1 _14288_ (.Y(_05998_),
    .A(_05908_),
    .B(_05997_));
 sg13g2_nor2_1 _14289_ (.A(net297),
    .B(_05998_),
    .Y(_05999_));
 sg13g2_a21oi_1 _14290_ (.A1(net299),
    .A2(_04264_),
    .Y(_06000_),
    .B1(_05999_));
 sg13g2_nand2_1 _14291_ (.Y(_06001_),
    .A(net1183),
    .B(_06000_));
 sg13g2_a21oi_1 _14292_ (.A1(_04195_),
    .A2(_05632_),
    .Y(_06002_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_18_ ));
 sg13g2_nand2_1 _14293_ (.Y(_06003_),
    .A(data_addr_o_18_),
    .B(net1012));
 sg13g2_o21ai_1 _14294_ (.B1(_06003_),
    .Y(_06004_),
    .A1(_02572_),
    .A2(net1012));
 sg13g2_nor2_1 _14295_ (.A(net311),
    .B(_06004_),
    .Y(_06005_));
 sg13g2_a21oi_1 _14296_ (.A1(net316),
    .A2(_06002_),
    .Y(_06006_),
    .B1(_06005_));
 sg13g2_nand2_1 _14297_ (.Y(_06007_),
    .A(data_addr_o_18_),
    .B(net1264));
 sg13g2_o21ai_1 _14298_ (.B1(_06007_),
    .Y(_06008_),
    .A1(_02572_),
    .A2(net1264));
 sg13g2_nand2_1 _14299_ (.Y(_06009_),
    .A(net422),
    .B(_06008_));
 sg13g2_o21ai_1 _14300_ (.B1(net1638),
    .Y(_06010_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ),
    .A2(net305));
 sg13g2_nand3_1 _14301_ (.B(_06009_),
    .C(_06010_),
    .A(net1574),
    .Y(_06011_));
 sg13g2_a221oi_1 _14302_ (.B2(net1889),
    .C1(_06011_),
    .B1(_06006_),
    .A1(net1886),
    .Y(_06012_),
    .A2(_05895_));
 sg13g2_o21ai_1 _14303_ (.B1(net1188),
    .Y(_06013_),
    .A1(net338),
    .A2(_06012_));
 sg13g2_o21ai_1 _14304_ (.B1(_06013_),
    .Y(_06014_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_50_ ),
    .A2(net1575));
 sg13g2_a22oi_1 _14305_ (.Y(_00141_),
    .B1(_06001_),
    .B2(_06014_),
    .A2(net96),
    .A1(_02572_));
 sg13g2_inv_1 _14306_ (.Y(_06015_),
    .A(\ex_block_i.alu_i.imd_val_q_i_51_ ));
 sg13g2_nor2_2 _14307_ (.A(net1576),
    .B(_04033_),
    .Y(_06016_));
 sg13g2_nand2b_1 _14308_ (.Y(_06017_),
    .B(_05996_),
    .A_N(_05908_));
 sg13g2_nand2_1 _14309_ (.Y(_06018_),
    .A(_05991_),
    .B(_06017_));
 sg13g2_nand2_1 _14310_ (.Y(_06019_),
    .A(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .B(net320));
 sg13g2_a21oi_2 _14311_ (.B1(net1566),
    .Y(_06020_),
    .A2(_06019_),
    .A1(net1568));
 sg13g2_inv_1 _14312_ (.Y(_06021_),
    .A(_05862_));
 sg13g2_mux2_1 _14313_ (.A0(_05977_),
    .A1(_05974_),
    .S(_05971_),
    .X(_06022_));
 sg13g2_nand2b_1 _14314_ (.Y(_06023_),
    .B(_05971_),
    .A_N(_05861_));
 sg13g2_nand3b_1 _14315_ (.B(net1081),
    .C(_05861_),
    .Y(_06024_),
    .A_N(_05971_));
 sg13g2_o21ai_1 _14316_ (.B1(_06024_),
    .Y(_06025_),
    .A1(net1081),
    .A2(_06023_));
 sg13g2_nor2_1 _14317_ (.A(_05977_),
    .B(_05974_),
    .Y(_06026_));
 sg13g2_a22oi_1 _14318_ (.Y(_06027_),
    .B1(_06025_),
    .B2(_06026_),
    .A2(_06022_),
    .A1(_06021_));
 sg13g2_nand2b_1 _14319_ (.Y(_06028_),
    .B(_05979_),
    .A_N(net1081));
 sg13g2_and2_1 _14320_ (.A(_05975_),
    .B(_06028_),
    .X(_06029_));
 sg13g2_o21ai_1 _14321_ (.B1(_05971_),
    .Y(_06030_),
    .A1(_05977_),
    .A2(_06029_));
 sg13g2_nor2b_1 _14322_ (.A(_05984_),
    .B_N(_06030_),
    .Y(_06031_));
 sg13g2_and2_1 _14323_ (.A(_06027_),
    .B(_06031_),
    .X(_06032_));
 sg13g2_nand2b_1 _14324_ (.Y(_06033_),
    .B(_05978_),
    .A_N(_05797_));
 sg13g2_a21oi_1 _14325_ (.A1(_05986_),
    .A2(_06033_),
    .Y(_06034_),
    .B1(_05971_));
 sg13g2_nor2_1 _14326_ (.A(_05976_),
    .B(_06034_),
    .Y(_06035_));
 sg13g2_and2_1 _14327_ (.A(_06035_),
    .B(_06027_),
    .X(_06036_));
 sg13g2_o21ai_1 _14328_ (.B1(_05946_),
    .Y(_06037_),
    .A1(net1326),
    .A2(_05943_));
 sg13g2_nand3_1 _14329_ (.B(net215),
    .C(_06037_),
    .A(_04217_),
    .Y(_06038_));
 sg13g2_buf_4 fanout860 (.X(net860),
    .A(net861));
 sg13g2_nor2_1 _14331_ (.A(_05943_),
    .B(_05946_),
    .Y(_06040_));
 sg13g2_a21oi_1 _14332_ (.A1(net1327),
    .A2(_05943_),
    .Y(_06041_),
    .B1(_06040_));
 sg13g2_nand2_1 _14333_ (.Y(_06042_),
    .A(_06038_),
    .B(_06041_));
 sg13g2_inv_1 _14334_ (.Y(_06043_),
    .A(_05939_));
 sg13g2_nor2_1 _14335_ (.A(net89),
    .B(_06043_),
    .Y(_06044_));
 sg13g2_nor3_1 _14336_ (.A(_05806_),
    .B(_05809_),
    .C(_05939_),
    .Y(_06045_));
 sg13g2_xnor2_1 _14337_ (.Y(_06046_),
    .A(net225),
    .B(_05811_));
 sg13g2_o21ai_1 _14338_ (.B1(_06046_),
    .Y(_06047_),
    .A1(_06044_),
    .A2(_06045_));
 sg13g2_nand2b_1 _14339_ (.Y(_06048_),
    .B(_06044_),
    .A_N(_05809_));
 sg13g2_nand3_1 _14340_ (.B(_06047_),
    .C(_06048_),
    .A(_06042_),
    .Y(_06049_));
 sg13g2_a21oi_1 _14341_ (.A1(_06047_),
    .A2(_06048_),
    .Y(_06050_),
    .B1(_06042_));
 sg13g2_inv_1 _14342_ (.Y(_06051_),
    .A(_06050_));
 sg13g2_nand2_1 _14343_ (.Y(_06052_),
    .A(_06049_),
    .B(_06051_));
 sg13g2_nand2_1 _14344_ (.Y(_06053_),
    .A(_05962_),
    .B(_05947_));
 sg13g2_nor2_1 _14345_ (.A(_05962_),
    .B(_05947_),
    .Y(_06054_));
 sg13g2_a21oi_2 _14346_ (.B1(_06054_),
    .Y(_06055_),
    .A2(_06053_),
    .A1(_05953_));
 sg13g2_a22oi_1 _14347_ (.Y(_06056_),
    .B1(net134),
    .B2(net1473),
    .A2(net1331),
    .A1(net264));
 sg13g2_xnor2_1 _14348_ (.Y(_06057_),
    .A(_05532_),
    .B(_06056_));
 sg13g2_and2_1 _14349_ (.A(net253),
    .B(net1258),
    .X(_06058_));
 sg13g2_a21o_1 _14350_ (.A2(net92),
    .A1(net268),
    .B1(_06058_),
    .X(_06059_));
 sg13g2_o21ai_1 _14351_ (.B1(net216),
    .Y(_06060_),
    .A1(_04368_),
    .A2(net1326));
 sg13g2_xnor2_1 _14352_ (.Y(_06061_),
    .A(_06059_),
    .B(_06060_));
 sg13g2_xnor2_1 _14353_ (.Y(_06062_),
    .A(_06057_),
    .B(_06061_));
 sg13g2_xor2_1 _14354_ (.B(_05960_),
    .A(net157),
    .X(_06063_));
 sg13g2_xnor2_1 _14355_ (.Y(_06064_),
    .A(net1375),
    .B(_05955_));
 sg13g2_xor2_1 _14356_ (.B(_05958_),
    .A(net1337),
    .X(_06065_));
 sg13g2_o21ai_1 _14357_ (.B1(_06065_),
    .Y(_06066_),
    .A1(_06063_),
    .A2(_06064_));
 sg13g2_nand2_1 _14358_ (.Y(_06067_),
    .A(_06063_),
    .B(_06064_));
 sg13g2_nand2_2 _14359_ (.Y(_06068_),
    .A(_06066_),
    .B(_06067_));
 sg13g2_nand2_1 _14360_ (.Y(_06069_),
    .A(net140),
    .B(net249));
 sg13g2_o21ai_1 _14361_ (.B1(_06069_),
    .Y(_06070_),
    .A1(_04726_),
    .A2(_05197_));
 sg13g2_xnor2_1 _14362_ (.Y(_06071_),
    .A(_05054_),
    .B(_06070_));
 sg13g2_a22oi_1 _14363_ (.Y(_06072_),
    .B1(net1433),
    .B2(net218),
    .A2(_05192_),
    .A1(net160));
 sg13g2_a22oi_1 _14364_ (.Y(_06073_),
    .B1(net138),
    .B2(net251),
    .A2(net1335),
    .A1(net1437));
 sg13g2_xnor2_1 _14365_ (.Y(_06074_),
    .A(_06072_),
    .B(_06073_));
 sg13g2_xnor2_1 _14366_ (.Y(_06075_),
    .A(_06071_),
    .B(_06074_));
 sg13g2_xor2_1 _14367_ (.B(_06075_),
    .A(_06068_),
    .X(_06076_));
 sg13g2_xnor2_1 _14368_ (.Y(_06077_),
    .A(_06062_),
    .B(_06076_));
 sg13g2_nor3_1 _14369_ (.A(net284),
    .B(net1515),
    .C(net1517),
    .Y(_06078_));
 sg13g2_and3_1 _14370_ (.X(_06079_),
    .A(net284),
    .B(net1515),
    .C(net1517));
 sg13g2_nor3_1 _14371_ (.A(net1869),
    .B(_06078_),
    .C(_06079_),
    .Y(_06080_));
 sg13g2_nor3_1 _14372_ (.A(net1502),
    .B(net1504),
    .C(net1505),
    .Y(_06081_));
 sg13g2_nor3_1 _14373_ (.A(net1380),
    .B(_02320_),
    .C(_02283_),
    .Y(_06082_));
 sg13g2_nor3_1 _14374_ (.A(net1876),
    .B(_06081_),
    .C(_06082_),
    .Y(_06083_));
 sg13g2_o21ai_1 _14375_ (.B1(net214),
    .Y(_06084_),
    .A1(_06080_),
    .A2(_06083_));
 sg13g2_xnor2_1 _14376_ (.Y(_06085_),
    .A(net167),
    .B(_06084_));
 sg13g2_a22oi_1 _14377_ (.Y(_06086_),
    .B1(net243),
    .B2(net220),
    .A2(net1323),
    .A1(net163));
 sg13g2_xnor2_1 _14378_ (.Y(_06087_),
    .A(_05206_),
    .B(_06086_));
 sg13g2_inv_1 _14379_ (.Y(_06088_),
    .A(_06087_));
 sg13g2_xnor2_1 _14380_ (.Y(_06089_),
    .A(_06085_),
    .B(_06088_));
 sg13g2_xnor2_1 _14381_ (.Y(_06090_),
    .A(net225),
    .B(_05937_));
 sg13g2_xnor2_1 _14382_ (.Y(_06091_),
    .A(_04354_),
    .B(_05936_));
 sg13g2_nor2_1 _14383_ (.A(_06090_),
    .B(_06091_),
    .Y(_06092_));
 sg13g2_and3_1 _14384_ (.X(_06093_),
    .A(net89),
    .B(_06090_),
    .C(_06091_));
 sg13g2_a21oi_1 _14385_ (.A1(_05806_),
    .A2(_06092_),
    .Y(_06094_),
    .B1(_06093_));
 sg13g2_xnor2_1 _14386_ (.Y(_06095_),
    .A(_06089_),
    .B(_06094_));
 sg13g2_xnor2_1 _14387_ (.Y(_06096_),
    .A(_06077_),
    .B(_06095_));
 sg13g2_xnor2_1 _14388_ (.Y(_06097_),
    .A(_06055_),
    .B(_06096_));
 sg13g2_xnor2_1 _14389_ (.Y(_06098_),
    .A(_06052_),
    .B(_06097_));
 sg13g2_nand3_1 _14390_ (.B(_05812_),
    .C(_05939_),
    .A(_05806_),
    .Y(_06099_));
 sg13g2_nand3_1 _14391_ (.B(_06046_),
    .C(_06043_),
    .A(net89),
    .Y(_06100_));
 sg13g2_a21oi_1 _14392_ (.A1(_06099_),
    .A2(_06100_),
    .Y(_06101_),
    .B1(_05809_));
 sg13g2_nand2_1 _14393_ (.Y(_06102_),
    .A(_05809_),
    .B(_05923_));
 sg13g2_nand2_1 _14394_ (.Y(_06103_),
    .A(net89),
    .B(_05939_));
 sg13g2_nand3_1 _14395_ (.B(_05812_),
    .C(_06043_),
    .A(_05806_),
    .Y(_06104_));
 sg13g2_a22oi_1 _14396_ (.Y(_06105_),
    .B1(_06103_),
    .B2(_06104_),
    .A2(_06102_),
    .A1(_05933_));
 sg13g2_xnor2_1 _14397_ (.Y(_06106_),
    .A(_05806_),
    .B(_05812_));
 sg13g2_nand2_1 _14398_ (.Y(_06107_),
    .A(_05933_),
    .B(_06043_));
 sg13g2_a22oi_1 _14399_ (.Y(_06108_),
    .B1(_06107_),
    .B2(_05809_),
    .A2(_05923_),
    .A1(_05939_));
 sg13g2_nor2_1 _14400_ (.A(_06106_),
    .B(_06108_),
    .Y(_06109_));
 sg13g2_a21oi_1 _14401_ (.A1(_06046_),
    .A2(_05939_),
    .Y(_06110_),
    .B1(_05923_));
 sg13g2_nor2_1 _14402_ (.A(_05933_),
    .B(_06110_),
    .Y(_06111_));
 sg13g2_nor4_2 _14403_ (.A(_06101_),
    .B(_06105_),
    .C(_06109_),
    .Y(_06112_),
    .D(_06111_));
 sg13g2_or2_1 _14404_ (.X(_06113_),
    .B(_05967_),
    .A(_05964_));
 sg13g2_and2_1 _14405_ (.A(_05964_),
    .B(_05967_),
    .X(_06114_));
 sg13g2_a21oi_1 _14406_ (.A1(_05941_),
    .A2(_06113_),
    .Y(_06115_),
    .B1(_06114_));
 sg13g2_xnor2_1 _14407_ (.Y(_06116_),
    .A(_06112_),
    .B(_06115_));
 sg13g2_xnor2_1 _14408_ (.Y(_06117_),
    .A(_06098_),
    .B(_06116_));
 sg13g2_inv_1 _14409_ (.Y(_06118_),
    .A(_05969_));
 sg13g2_a21oi_1 _14410_ (.A1(_05561_),
    .A2(_05675_),
    .Y(_06119_),
    .B1(_05674_));
 sg13g2_o21ai_1 _14411_ (.B1(_05821_),
    .Y(_06120_),
    .A1(_05822_),
    .A2(_06119_));
 sg13g2_inv_1 _14412_ (.Y(_06121_),
    .A(_06120_));
 sg13g2_o21ai_1 _14413_ (.B1(_05801_),
    .Y(_06122_),
    .A1(_05917_),
    .A2(_06120_));
 sg13g2_o21ai_1 _14414_ (.B1(_06122_),
    .Y(_06123_),
    .A1(_05819_),
    .A2(_06121_));
 sg13g2_a21oi_1 _14415_ (.A1(_05916_),
    .A2(_06118_),
    .Y(_06124_),
    .B1(_06123_));
 sg13g2_nor2_1 _14416_ (.A(_05916_),
    .B(_06118_),
    .Y(_06125_));
 sg13g2_nor2_1 _14417_ (.A(_06124_),
    .B(_06125_),
    .Y(_06126_));
 sg13g2_xor2_1 _14418_ (.B(_06126_),
    .A(_06117_),
    .X(_06127_));
 sg13g2_mux4_1 _14419_ (.S0(_05788_),
    .A0(_06032_),
    .A1(_06031_),
    .A2(_06035_),
    .A3(_06036_),
    .S1(_06127_),
    .X(_06128_));
 sg13g2_xnor2_1 _14420_ (.Y(_06129_),
    .A(_06020_),
    .B(_06128_));
 sg13g2_xnor2_1 _14421_ (.Y(_06130_),
    .A(_06018_),
    .B(_06129_));
 sg13g2_nand2_1 _14422_ (.Y(_06131_),
    .A(net299),
    .B(_04326_));
 sg13g2_o21ai_1 _14423_ (.B1(_06131_),
    .Y(_06132_),
    .A1(net297),
    .A2(_06130_));
 sg13g2_nand2_2 _14424_ (.Y(_06133_),
    .A(_06016_),
    .B(_06132_));
 sg13g2_a21oi_1 _14425_ (.A1(_04195_),
    .A2(_05892_),
    .Y(_06134_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_19_ ));
 sg13g2_nand2_1 _14426_ (.Y(_06135_),
    .A(data_addr_o_19_),
    .B(net1008));
 sg13g2_o21ai_1 _14427_ (.B1(_06135_),
    .Y(_06136_),
    .A1(_06015_),
    .A2(net1008));
 sg13g2_nor2_1 _14428_ (.A(net311),
    .B(_06136_),
    .Y(_06137_));
 sg13g2_a21oi_1 _14429_ (.A1(net315),
    .A2(_06134_),
    .Y(_06138_),
    .B1(_06137_));
 sg13g2_nand2_1 _14430_ (.Y(_06139_),
    .A(data_addr_o_19_),
    .B(net1260));
 sg13g2_o21ai_1 _14431_ (.B1(_06139_),
    .Y(_06140_),
    .A1(_06015_),
    .A2(net1266));
 sg13g2_nand2_1 _14432_ (.Y(_06141_),
    .A(net422),
    .B(_06140_));
 sg13g2_o21ai_1 _14433_ (.B1(_04137_),
    .Y(_06142_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ),
    .A2(net304));
 sg13g2_nand3_1 _14434_ (.B(_06141_),
    .C(_06142_),
    .A(net1569),
    .Y(_06143_));
 sg13g2_a221oi_1 _14435_ (.B2(net1891),
    .C1(_06143_),
    .B1(_06138_),
    .A1(net1883),
    .Y(_06144_),
    .A2(_06004_));
 sg13g2_o21ai_1 _14436_ (.B1(net1187),
    .Y(_06145_),
    .A1(net339),
    .A2(_06144_));
 sg13g2_o21ai_1 _14437_ (.B1(_06145_),
    .Y(_06146_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .A2(net1571));
 sg13g2_a22oi_1 _14438_ (.Y(_00142_),
    .B1(_06133_),
    .B2(_06146_),
    .A2(net95),
    .A1(_06015_));
 sg13g2_inv_1 _14439_ (.Y(_06147_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ));
 sg13g2_or2_1 _14440_ (.X(_06148_),
    .B(_06128_),
    .A(_06020_));
 sg13g2_and2_1 _14441_ (.A(_05991_),
    .B(_06148_),
    .X(_06149_));
 sg13g2_nor2b_1 _14442_ (.A(_05990_),
    .B_N(_05913_),
    .Y(_06150_));
 sg13g2_nor2_1 _14443_ (.A(_05884_),
    .B(_06150_),
    .Y(_06151_));
 sg13g2_o21ai_1 _14444_ (.B1(_06151_),
    .Y(_06152_),
    .A1(_05776_),
    .A2(_05885_));
 sg13g2_and2_1 _14445_ (.A(_06020_),
    .B(_06128_),
    .X(_06153_));
 sg13g2_a21oi_2 _14446_ (.B1(_06153_),
    .Y(_06154_),
    .A2(_06152_),
    .A1(_06149_));
 sg13g2_nand2_1 _14447_ (.Y(_06155_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .B(net320));
 sg13g2_a21oi_2 _14448_ (.B1(net1566),
    .Y(_06156_),
    .A2(_06155_),
    .A1(net1568));
 sg13g2_or2_1 _14449_ (.X(_06157_),
    .B(_06127_),
    .A(_06027_));
 sg13g2_nor2_1 _14450_ (.A(_05855_),
    .B(_05915_),
    .Y(_06158_));
 sg13g2_a21oi_2 _14451_ (.B1(_06158_),
    .Y(_06159_),
    .A2(_05824_),
    .A1(_05859_));
 sg13g2_nand2_1 _14452_ (.Y(_06160_),
    .A(_06123_),
    .B(_06159_));
 sg13g2_nor2_1 _14453_ (.A(_06123_),
    .B(_06159_),
    .Y(_06161_));
 sg13g2_a21o_1 _14454_ (.A2(_06160_),
    .A1(_05969_),
    .B1(_06161_),
    .X(_06162_));
 sg13g2_xor2_1 _14455_ (.B(_06159_),
    .A(_05970_),
    .X(_06163_));
 sg13g2_a221oi_1 _14456_ (.B2(_05977_),
    .C1(_05984_),
    .B1(_06163_),
    .A1(_05971_),
    .Y(_06164_),
    .A2(_06029_));
 sg13g2_o21ai_1 _14457_ (.B1(_06164_),
    .Y(_06165_),
    .A1(_06117_),
    .A2(_06162_));
 sg13g2_nand2_1 _14458_ (.Y(_06166_),
    .A(_06117_),
    .B(_06162_));
 sg13g2_nand2_1 _14459_ (.Y(_06167_),
    .A(_06165_),
    .B(_06166_));
 sg13g2_o21ai_1 _14460_ (.B1(_06167_),
    .Y(_06168_),
    .A1(_05788_),
    .A2(_06157_));
 sg13g2_and2_1 _14461_ (.A(_06077_),
    .B(_06095_),
    .X(_06169_));
 sg13g2_or2_1 _14462_ (.X(_06170_),
    .B(_06095_),
    .A(_06077_));
 sg13g2_o21ai_1 _14463_ (.B1(_06170_),
    .Y(_06171_),
    .A1(_06055_),
    .A2(_06169_));
 sg13g2_nor2_1 _14464_ (.A(_06055_),
    .B(_06170_),
    .Y(_06172_));
 sg13g2_a21oi_1 _14465_ (.A1(_06055_),
    .A2(_06170_),
    .Y(_06173_),
    .B1(_06169_));
 sg13g2_nand3_1 _14466_ (.B(_06051_),
    .C(_06169_),
    .A(_06055_),
    .Y(_06174_));
 sg13g2_o21ai_1 _14467_ (.B1(_06174_),
    .Y(_06175_),
    .A1(_06049_),
    .A2(_06173_));
 sg13g2_a221oi_1 _14468_ (.B2(_06049_),
    .C1(_06175_),
    .B1(_06172_),
    .A1(_06050_),
    .Y(_06176_),
    .A2(_06171_));
 sg13g2_nor2_1 _14469_ (.A(net89),
    .B(_06092_),
    .Y(_06177_));
 sg13g2_nor2b_1 _14470_ (.A(_06089_),
    .B_N(_06093_),
    .Y(_06178_));
 sg13g2_a21oi_2 _14471_ (.B1(_06178_),
    .Y(_06179_),
    .A2(_06177_),
    .A1(_06089_));
 sg13g2_buf_4 fanout859 (.X(net859),
    .A(net861));
 sg13g2_xor2_1 _14473_ (.B(_06056_),
    .A(net1329),
    .X(_06181_));
 sg13g2_buf_4 fanout858 (.X(net858),
    .A(net862));
 sg13g2_nor2_1 _14475_ (.A(net1321),
    .B(_06059_),
    .Y(_06183_));
 sg13g2_o21ai_1 _14476_ (.B1(_06183_),
    .Y(_06184_),
    .A1(net215),
    .A2(_06181_));
 sg13g2_a21oi_1 _14477_ (.A1(_04368_),
    .A2(net1321),
    .Y(_06185_),
    .B1(_06181_));
 sg13g2_nand2_1 _14478_ (.Y(_06186_),
    .A(net1321),
    .B(_06181_));
 sg13g2_o21ai_1 _14479_ (.B1(_06186_),
    .Y(_06187_),
    .A1(net1373),
    .A2(_06185_));
 sg13g2_nand2_1 _14480_ (.Y(_06188_),
    .A(_06059_),
    .B(_06187_));
 sg13g2_nand3_1 _14481_ (.B(net215),
    .C(_06181_),
    .A(_04368_),
    .Y(_06189_));
 sg13g2_nand3_1 _14482_ (.B(_06188_),
    .C(_06189_),
    .A(_06184_),
    .Y(_06190_));
 sg13g2_xnor2_1 _14483_ (.Y(_06191_),
    .A(_06179_),
    .B(_06190_));
 sg13g2_o21ai_1 _14484_ (.B1(_05566_),
    .Y(_06192_),
    .A1(_03950_),
    .A2(_05567_));
 sg13g2_nand2b_1 _14485_ (.Y(_06193_),
    .B(_06192_),
    .A_N(net269));
 sg13g2_a22oi_1 _14486_ (.Y(_06194_),
    .B1(net90),
    .B2(net254),
    .A2(net1258),
    .A1(net1473));
 sg13g2_buf_4 fanout857 (.X(net857),
    .A(net862));
 sg13g2_buf_4 fanout856 (.X(net856),
    .A(\register_file_i/_2885_ ));
 sg13g2_a22oi_1 _14489_ (.Y(_06197_),
    .B1(net135),
    .B2(_04608_),
    .A2(net1332),
    .A1(net252));
 sg13g2_xnor2_1 _14490_ (.Y(_06198_),
    .A(net1328),
    .B(_06197_));
 sg13g2_xor2_1 _14491_ (.B(_06198_),
    .A(_06194_),
    .X(_06199_));
 sg13g2_xnor2_1 _14492_ (.Y(_06200_),
    .A(_06193_),
    .B(_06199_));
 sg13g2_xor2_1 _14493_ (.B(_06070_),
    .A(net1337),
    .X(_06201_));
 sg13g2_xnor2_1 _14494_ (.Y(_06202_),
    .A(net159),
    .B(_06072_));
 sg13g2_xnor2_1 _14495_ (.Y(_06203_),
    .A(net1374),
    .B(_06073_));
 sg13g2_o21ai_1 _14496_ (.B1(_06203_),
    .Y(_06204_),
    .A1(_06201_),
    .A2(_06202_));
 sg13g2_nand2_1 _14497_ (.Y(_06205_),
    .A(_06201_),
    .B(_06202_));
 sg13g2_nand2_1 _14498_ (.Y(_06206_),
    .A(_06204_),
    .B(_06205_));
 sg13g2_a22oi_1 _14499_ (.Y(_06207_),
    .B1(net137),
    .B2(net1437),
    .A2(net1335),
    .A1(net248));
 sg13g2_xnor2_1 _14500_ (.Y(_06208_),
    .A(_05440_),
    .B(_06207_));
 sg13g2_buf_4 fanout855 (.X(net855),
    .A(net856));
 sg13g2_buf_4 fanout854 (.X(net854),
    .A(net856));
 sg13g2_a22oi_1 _14503_ (.Y(_06211_),
    .B1(net1322),
    .B2(net218),
    .A2(_05302_),
    .A1(net160));
 sg13g2_a22oi_1 _14504_ (.Y(_06212_),
    .B1(net1435),
    .B2(net1339),
    .A2(net247),
    .A1(net140));
 sg13g2_xnor2_1 _14505_ (.Y(_06213_),
    .A(_06211_),
    .B(_06212_));
 sg13g2_xnor2_1 _14506_ (.Y(_06214_),
    .A(_06208_),
    .B(_06213_));
 sg13g2_xnor2_1 _14507_ (.Y(_06215_),
    .A(_06206_),
    .B(_06214_));
 sg13g2_xnor2_1 _14508_ (.Y(_06216_),
    .A(_06200_),
    .B(_06215_));
 sg13g2_a22oi_1 _14509_ (.Y(_06217_),
    .B1(net213),
    .B2(net220),
    .A2(net244),
    .A1(net162));
 sg13g2_xnor2_1 _14510_ (.Y(_06218_),
    .A(net225),
    .B(_06217_));
 sg13g2_nand2_1 _14511_ (.Y(_06219_),
    .A(_06085_),
    .B(_06087_));
 sg13g2_nor2_1 _14512_ (.A(_06085_),
    .B(_06087_),
    .Y(_06220_));
 sg13g2_a21oi_1 _14513_ (.A1(_05924_),
    .A2(_06219_),
    .Y(_06221_),
    .B1(_06220_));
 sg13g2_xnor2_1 _14514_ (.Y(_06222_),
    .A(_06218_),
    .B(_06221_));
 sg13g2_nor2_1 _14515_ (.A(_06068_),
    .B(_06075_),
    .Y(_06223_));
 sg13g2_nand2_1 _14516_ (.Y(_06224_),
    .A(_06068_),
    .B(_06075_));
 sg13g2_o21ai_1 _14517_ (.B1(_06224_),
    .Y(_06225_),
    .A1(_06062_),
    .A2(_06223_));
 sg13g2_xor2_1 _14518_ (.B(_06225_),
    .A(_06222_),
    .X(_06226_));
 sg13g2_xnor2_1 _14519_ (.Y(_06227_),
    .A(_06216_),
    .B(_06226_));
 sg13g2_xnor2_1 _14520_ (.Y(_06228_),
    .A(_06191_),
    .B(_06227_));
 sg13g2_xor2_1 _14521_ (.B(_06228_),
    .A(_06176_),
    .X(_06229_));
 sg13g2_inv_1 _14522_ (.Y(_06230_),
    .A(_06112_));
 sg13g2_inv_1 _14523_ (.Y(_06231_),
    .A(_06098_));
 sg13g2_o21ai_1 _14524_ (.B1(_06113_),
    .Y(_06232_),
    .A1(_05941_),
    .A2(_06114_));
 sg13g2_o21ai_1 _14525_ (.B1(_06232_),
    .Y(_06233_),
    .A1(_06112_),
    .A2(_06231_));
 sg13g2_o21ai_1 _14526_ (.B1(_06233_),
    .Y(_06234_),
    .A1(_06230_),
    .A2(_06098_));
 sg13g2_xnor2_1 _14527_ (.Y(_06235_),
    .A(_06229_),
    .B(_06234_));
 sg13g2_xor2_1 _14528_ (.B(_06235_),
    .A(_06168_),
    .X(_06236_));
 sg13g2_xnor2_1 _14529_ (.Y(_06237_),
    .A(_06156_),
    .B(_06236_));
 sg13g2_xor2_1 _14530_ (.B(_06237_),
    .A(_06154_),
    .X(_06238_));
 sg13g2_mux2_1 _14531_ (.A0(_04393_),
    .A1(_06238_),
    .S(net1538),
    .X(_06239_));
 sg13g2_nand2_1 _14532_ (.Y(_06240_),
    .A(net1182),
    .B(_06239_));
 sg13g2_a21o_1 _14533_ (.A2(_06240_),
    .A1(net1478),
    .B1(net95),
    .X(_06241_));
 sg13g2_nand2_1 _14534_ (.Y(_06242_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .B(net1005));
 sg13g2_o21ai_1 _14535_ (.B1(_06242_),
    .Y(_06243_),
    .A1(_03274_),
    .A2(net1005));
 sg13g2_inv_1 _14536_ (.Y(_06244_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ));
 sg13g2_nor2_2 _14537_ (.A(_06244_),
    .B(_04331_),
    .Y(_06245_));
 sg13g2_a21oi_1 _14538_ (.A1(_04083_),
    .A2(_06245_),
    .Y(_06246_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_20_ ));
 sg13g2_nand2_1 _14539_ (.Y(_06247_),
    .A(net313),
    .B(_06246_));
 sg13g2_o21ai_1 _14540_ (.B1(_06247_),
    .Y(_06248_),
    .A1(net308),
    .A2(_06243_));
 sg13g2_nand2_1 _14541_ (.Y(_06249_),
    .A(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .B(net1218));
 sg13g2_o21ai_1 _14542_ (.B1(_06249_),
    .Y(_06250_),
    .A1(_03274_),
    .A2(net1218));
 sg13g2_o21ai_1 _14543_ (.B1(net1635),
    .Y(_06251_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ),
    .A2(net309));
 sg13g2_nand2_1 _14544_ (.Y(_06252_),
    .A(net1181),
    .B(_06251_));
 sg13g2_a221oi_1 _14545_ (.B2(net420),
    .C1(_06252_),
    .B1(_06250_),
    .A1(net1882),
    .Y(_06253_),
    .A2(_06136_));
 sg13g2_o21ai_1 _14546_ (.B1(_06253_),
    .Y(_06254_),
    .A1(net1708),
    .A2(_06248_));
 sg13g2_o21ai_1 _14547_ (.B1(_06254_),
    .Y(_06255_),
    .A1(net1578),
    .A2(net94));
 sg13g2_a22oi_1 _14548_ (.Y(_00143_),
    .B1(_06255_),
    .B2(_06240_),
    .A2(_06241_),
    .A1(_06147_));
 sg13g2_nand2_1 _14549_ (.Y(_06256_),
    .A(_06156_),
    .B(_06236_));
 sg13g2_nor2_1 _14550_ (.A(_06156_),
    .B(_06236_),
    .Y(_06257_));
 sg13g2_a21oi_1 _14551_ (.A1(_06154_),
    .A2(_06256_),
    .Y(_06258_),
    .B1(_06257_));
 sg13g2_nor2_1 _14552_ (.A(_05788_),
    .B(_06157_),
    .Y(_06259_));
 sg13g2_inv_1 _14553_ (.Y(_06260_),
    .A(_06229_));
 sg13g2_or2_1 _14554_ (.X(_06261_),
    .B(_06162_),
    .A(_06164_));
 sg13g2_a22oi_1 _14555_ (.Y(_06262_),
    .B1(_06261_),
    .B2(_06117_),
    .A2(_06162_),
    .A1(_06031_));
 sg13g2_a21o_1 _14556_ (.A2(_06234_),
    .A1(_06260_),
    .B1(_06262_),
    .X(_06263_));
 sg13g2_or2_1 _14557_ (.X(_06264_),
    .B(_06234_),
    .A(_06260_));
 sg13g2_a22oi_1 _14558_ (.Y(_06265_),
    .B1(_06263_),
    .B2(_06264_),
    .A2(_06235_),
    .A1(_06259_));
 sg13g2_nand2_1 _14559_ (.Y(_06266_),
    .A(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .B(net319));
 sg13g2_a21o_1 _14560_ (.A2(_06266_),
    .A1(net1568),
    .B1(net1565),
    .X(_06267_));
 sg13g2_a21oi_1 _14561_ (.A1(_06062_),
    .A2(_06224_),
    .Y(_06268_),
    .B1(_06223_));
 sg13g2_or2_1 _14562_ (.X(_06269_),
    .B(_06268_),
    .A(_06190_));
 sg13g2_inv_1 _14563_ (.Y(_06270_),
    .A(_06269_));
 sg13g2_nand2_1 _14564_ (.Y(_06271_),
    .A(_06190_),
    .B(_06225_));
 sg13g2_nand2_1 _14565_ (.Y(_06272_),
    .A(_06216_),
    .B(_06271_));
 sg13g2_a21oi_1 _14566_ (.A1(_06269_),
    .A2(_06272_),
    .Y(_06273_),
    .B1(_06222_));
 sg13g2_a21oi_1 _14567_ (.A1(_06216_),
    .A2(_06270_),
    .Y(_06274_),
    .B1(_06273_));
 sg13g2_and2_1 _14568_ (.A(_06190_),
    .B(_06225_),
    .X(_06275_));
 sg13g2_inv_1 _14569_ (.Y(_06276_),
    .A(_06179_));
 sg13g2_nor2b_1 _14570_ (.A(_06222_),
    .B_N(_06216_),
    .Y(_06277_));
 sg13g2_nand2b_1 _14571_ (.Y(_06278_),
    .B(_06222_),
    .A_N(_06216_));
 sg13g2_o21ai_1 _14572_ (.B1(_06278_),
    .Y(_06279_),
    .A1(_06276_),
    .A2(_06277_));
 sg13g2_nand2_1 _14573_ (.Y(_06280_),
    .A(_06179_),
    .B(_06269_));
 sg13g2_nor2_1 _14574_ (.A(_06278_),
    .B(_06280_),
    .Y(_06281_));
 sg13g2_a221oi_1 _14575_ (.B2(_06277_),
    .C1(_06281_),
    .B1(_06270_),
    .A1(_06275_),
    .Y(_06282_),
    .A2(_06279_));
 sg13g2_o21ai_1 _14576_ (.B1(_06282_),
    .Y(_06283_),
    .A1(_06179_),
    .A2(_06274_));
 sg13g2_a22oi_1 _14577_ (.Y(_06284_),
    .B1(net135),
    .B2(net251),
    .A2(net1332),
    .A1(net1437));
 sg13g2_xnor2_1 _14578_ (.Y(_06285_),
    .A(net1329),
    .B(_06284_));
 sg13g2_buf_4 fanout853 (.X(net853),
    .A(net856));
 sg13g2_buf_4 fanout852 (.X(net852),
    .A(net853));
 sg13g2_a22oi_1 _14581_ (.Y(_06288_),
    .B1(net91),
    .B2(net1473),
    .A2(net1258),
    .A1(net264));
 sg13g2_nor2_1 _14582_ (.A(net253),
    .B(_05686_),
    .Y(_06289_));
 sg13g2_xnor2_1 _14583_ (.Y(_06290_),
    .A(_06288_),
    .B(_06289_));
 sg13g2_xnor2_1 _14584_ (.Y(_06291_),
    .A(_06285_),
    .B(_06290_));
 sg13g2_xnor2_1 _14585_ (.Y(_06292_),
    .A(net1337),
    .B(_06212_));
 sg13g2_xnor2_1 _14586_ (.Y(_06293_),
    .A(net1374),
    .B(_06207_));
 sg13g2_xnor2_1 _14587_ (.Y(_06294_),
    .A(net158),
    .B(_06211_));
 sg13g2_a21oi_1 _14588_ (.A1(_06292_),
    .A2(_06293_),
    .Y(_06295_),
    .B1(_06294_));
 sg13g2_nor2_1 _14589_ (.A(_06292_),
    .B(_06293_),
    .Y(_06296_));
 sg13g2_nor2_2 _14590_ (.A(_06295_),
    .B(_06296_),
    .Y(_06297_));
 sg13g2_and2_1 _14591_ (.A(net246),
    .B(net1334),
    .X(_06298_));
 sg13g2_a21o_1 _14592_ (.A2(_05064_),
    .A1(net250),
    .B1(_06298_),
    .X(_06299_));
 sg13g2_xor2_1 _14593_ (.B(_06299_),
    .A(_05835_),
    .X(_06300_));
 sg13g2_a22oi_1 _14594_ (.Y(_06301_),
    .B1(_05302_),
    .B2(net1339),
    .A2(net1435),
    .A1(net140));
 sg13g2_a22oi_1 _14595_ (.Y(_06302_),
    .B1(net242),
    .B2(net218),
    .A2(net1322),
    .A1(net160));
 sg13g2_xnor2_1 _14596_ (.Y(_06303_),
    .A(_06301_),
    .B(_06302_));
 sg13g2_xnor2_1 _14597_ (.Y(_06304_),
    .A(_06300_),
    .B(_06303_));
 sg13g2_xor2_1 _14598_ (.B(_06304_),
    .A(_06297_),
    .X(_06305_));
 sg13g2_xnor2_1 _14599_ (.Y(_06306_),
    .A(_06291_),
    .B(_06305_));
 sg13g2_o21ai_1 _14600_ (.B1(_05806_),
    .Y(_06307_),
    .A1(_06085_),
    .A2(_06087_));
 sg13g2_a21oi_1 _14601_ (.A1(_06219_),
    .A2(_06307_),
    .Y(_06308_),
    .B1(_06218_));
 sg13g2_o21ai_1 _14602_ (.B1(_06198_),
    .Y(_06309_),
    .A1(net1326),
    .A2(_06194_));
 sg13g2_nor2_1 _14603_ (.A(net269),
    .B(net1372),
    .Y(_06310_));
 sg13g2_nor2_1 _14604_ (.A(_06194_),
    .B(_06198_),
    .Y(_06311_));
 sg13g2_a221oi_1 _14605_ (.B2(_06310_),
    .C1(_06311_),
    .B1(_06309_),
    .A1(net1326),
    .Y(_06312_),
    .A2(_06194_));
 sg13g2_nor3_1 _14606_ (.A(net1517),
    .B(net287),
    .C(net1521),
    .Y(_06313_));
 sg13g2_nand3_1 _14607_ (.B(net287),
    .C(net1521),
    .A(net1517),
    .Y(_06314_));
 sg13g2_nand2b_1 _14608_ (.Y(_06315_),
    .B(_06314_),
    .A_N(_06313_));
 sg13g2_or3_1 _14609_ (.A(net1506),
    .B(net1507),
    .C(net1510),
    .X(_06316_));
 sg13g2_nand3_1 _14610_ (.B(net1507),
    .C(net1510),
    .A(net1506),
    .Y(_06317_));
 sg13g2_nand3_1 _14611_ (.B(_06316_),
    .C(_06317_),
    .A(net1868),
    .Y(_06318_));
 sg13g2_o21ai_1 _14612_ (.B1(_06318_),
    .Y(_06319_),
    .A1(net1868),
    .A2(_06315_));
 sg13g2_and2_1 _14613_ (.A(net213),
    .B(_06319_),
    .X(_06320_));
 sg13g2_xnor2_1 _14614_ (.Y(_06321_),
    .A(net225),
    .B(_06320_));
 sg13g2_xnor2_1 _14615_ (.Y(_06322_),
    .A(_06312_),
    .B(_06321_));
 sg13g2_xnor2_1 _14616_ (.Y(_06323_),
    .A(_06308_),
    .B(_06322_));
 sg13g2_nand2_1 _14617_ (.Y(_06324_),
    .A(_06214_),
    .B(_06200_));
 sg13g2_nand2_1 _14618_ (.Y(_06325_),
    .A(_06206_),
    .B(_06324_));
 sg13g2_or2_1 _14619_ (.X(_06326_),
    .B(_06200_),
    .A(_06214_));
 sg13g2_nand3_1 _14620_ (.B(_06325_),
    .C(_06326_),
    .A(_06323_),
    .Y(_06327_));
 sg13g2_a21o_1 _14621_ (.A2(_06326_),
    .A1(_06325_),
    .B1(_06323_),
    .X(_06328_));
 sg13g2_nand2_1 _14622_ (.Y(_06329_),
    .A(_06327_),
    .B(_06328_));
 sg13g2_xnor2_1 _14623_ (.Y(_06330_),
    .A(_06306_),
    .B(_06329_));
 sg13g2_xnor2_1 _14624_ (.Y(_06331_),
    .A(_06283_),
    .B(_06330_));
 sg13g2_nand2_1 _14625_ (.Y(_06332_),
    .A(_06055_),
    .B(_06051_));
 sg13g2_nand3b_1 _14626_ (.B(_06049_),
    .C(_06332_),
    .Y(_06333_),
    .A_N(_06095_));
 sg13g2_nand2b_1 _14627_ (.Y(_06334_),
    .B(_06050_),
    .A_N(_06055_));
 sg13g2_a21oi_1 _14628_ (.A1(_06333_),
    .A2(_06334_),
    .Y(_06335_),
    .B1(_06077_));
 sg13g2_nor2_1 _14629_ (.A(_06095_),
    .B(_06334_),
    .Y(_06336_));
 sg13g2_nor2_1 _14630_ (.A(_06335_),
    .B(_06336_),
    .Y(_06337_));
 sg13g2_a21oi_2 _14631_ (.B1(_06175_),
    .Y(_06338_),
    .A2(_06337_),
    .A1(_06228_));
 sg13g2_xnor2_1 _14632_ (.Y(_06339_),
    .A(_06331_),
    .B(_06338_));
 sg13g2_xnor2_1 _14633_ (.Y(_06340_),
    .A(_06267_),
    .B(_06339_));
 sg13g2_xnor2_1 _14634_ (.Y(_06341_),
    .A(_06265_),
    .B(_06340_));
 sg13g2_xnor2_1 _14635_ (.Y(_06342_),
    .A(_06258_),
    .B(_06341_));
 sg13g2_nand2_1 _14636_ (.Y(_06343_),
    .A(net1541),
    .B(_06342_));
 sg13g2_or2_1 _14637_ (.X(_06344_),
    .B(_04479_),
    .A(net1541));
 sg13g2_nand4_1 _14638_ (.B(net1182),
    .C(_06343_),
    .A(net1188),
    .Y(_06345_),
    .D(_06344_));
 sg13g2_nor2_2 _14639_ (.A(_04487_),
    .B(_05891_),
    .Y(_06346_));
 sg13g2_a21oi_1 _14640_ (.A1(_04083_),
    .A2(_06346_),
    .Y(_06347_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_21_ ));
 sg13g2_mux2_1 _14641_ (.A0(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .A1(data_addr_o_21_),
    .S(net1009),
    .X(_06348_));
 sg13g2_nor2_1 _14642_ (.A(net307),
    .B(_06348_),
    .Y(_06349_));
 sg13g2_a21oi_1 _14643_ (.A1(net314),
    .A2(_06347_),
    .Y(_06350_),
    .B1(_06349_));
 sg13g2_nand2_1 _14644_ (.Y(_06351_),
    .A(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .B(net1219));
 sg13g2_o21ai_1 _14645_ (.B1(_06351_),
    .Y(_06352_),
    .A1(_02931_),
    .A2(net1219));
 sg13g2_nand2_1 _14646_ (.Y(_06353_),
    .A(net421),
    .B(_06352_));
 sg13g2_o21ai_1 _14647_ (.B1(net1638),
    .Y(_06354_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ),
    .A2(net310));
 sg13g2_nand3_1 _14648_ (.B(_06353_),
    .C(_06354_),
    .A(net1569),
    .Y(_06355_));
 sg13g2_a221oi_1 _14649_ (.B2(net1889),
    .C1(_06355_),
    .B1(_06350_),
    .A1(net1886),
    .Y(_06356_),
    .A2(_06243_));
 sg13g2_o21ai_1 _14650_ (.B1(net1188),
    .Y(_06357_),
    .A1(net337),
    .A2(_06356_));
 sg13g2_o21ai_1 _14651_ (.B1(_06357_),
    .Y(_06358_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .A2(_05153_));
 sg13g2_nand2_1 _14652_ (.Y(_00144_),
    .A(_06345_),
    .B(_06358_));
 sg13g2_buf_4 fanout851 (.X(net851),
    .A(\register_file_i/_2903_ ));
 sg13g2_nand2_1 _14654_ (.Y(_06360_),
    .A(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .B(net319));
 sg13g2_a21oi_1 _14655_ (.A1(net1568),
    .A2(_06360_),
    .Y(_06361_),
    .B1(net1566));
 sg13g2_inv_1 _14656_ (.Y(_06362_),
    .A(_06361_));
 sg13g2_inv_1 _14657_ (.Y(_06363_),
    .A(_06331_));
 sg13g2_nor2_1 _14658_ (.A(_06363_),
    .B(_06338_),
    .Y(_06364_));
 sg13g2_nor2b_1 _14659_ (.A(_06331_),
    .B_N(_06338_),
    .Y(_06365_));
 sg13g2_inv_1 _14660_ (.Y(_06366_),
    .A(_06365_));
 sg13g2_o21ai_1 _14661_ (.B1(_06366_),
    .Y(_06367_),
    .A1(_06265_),
    .A2(_06364_));
 sg13g2_a22oi_1 _14662_ (.Y(_06368_),
    .B1(net213),
    .B2(net218),
    .A2(net244),
    .A1(net160));
 sg13g2_xor2_1 _14663_ (.B(_06368_),
    .A(net157),
    .X(_06369_));
 sg13g2_a22oi_1 _14664_ (.Y(_06370_),
    .B1(net1435),
    .B2(net1334),
    .A2(_05064_),
    .A1(net246));
 sg13g2_a22oi_1 _14665_ (.Y(_06371_),
    .B1(net1322),
    .B2(net1339),
    .A2(_05302_),
    .A1(net139));
 sg13g2_xor2_1 _14666_ (.B(_06371_),
    .A(_05834_),
    .X(_06372_));
 sg13g2_xnor2_1 _14667_ (.Y(_06373_),
    .A(_06370_),
    .B(_06372_));
 sg13g2_xnor2_1 _14668_ (.Y(_06374_),
    .A(_06369_),
    .B(_06373_));
 sg13g2_a22oi_1 _14669_ (.Y(_06375_),
    .B1(net135),
    .B2(net1437),
    .A2(net1332),
    .A1(net248));
 sg13g2_xor2_1 _14670_ (.B(_06375_),
    .A(net1329),
    .X(_06376_));
 sg13g2_and2_1 _14671_ (.A(net252),
    .B(net1258),
    .X(_06377_));
 sg13g2_a21o_1 _14672_ (.A2(net92),
    .A1(net266),
    .B1(_06377_),
    .X(_06378_));
 sg13g2_nor2_1 _14673_ (.A(net1473),
    .B(_05686_),
    .Y(_06379_));
 sg13g2_xnor2_1 _14674_ (.Y(_06380_),
    .A(_06378_),
    .B(_06379_));
 sg13g2_xnor2_1 _14675_ (.Y(_06381_),
    .A(_06376_),
    .B(_06380_));
 sg13g2_xnor2_1 _14676_ (.Y(_06382_),
    .A(net158),
    .B(_06302_));
 sg13g2_xnor2_1 _14677_ (.Y(_06383_),
    .A(_05043_),
    .B(_06299_));
 sg13g2_xnor2_1 _14678_ (.Y(_06384_),
    .A(net1337),
    .B(_06301_));
 sg13g2_o21ai_1 _14679_ (.B1(_06384_),
    .Y(_06385_),
    .A1(_06382_),
    .A2(_06383_));
 sg13g2_nand2_1 _14680_ (.Y(_06386_),
    .A(_06382_),
    .B(_06383_));
 sg13g2_nand2_1 _14681_ (.Y(_06387_),
    .A(_06385_),
    .B(_06386_));
 sg13g2_nand2b_1 _14682_ (.Y(_06388_),
    .B(_06387_),
    .A_N(_06381_));
 sg13g2_nor2b_1 _14683_ (.A(_06387_),
    .B_N(_06381_),
    .Y(_06389_));
 sg13g2_inv_1 _14684_ (.Y(_06390_),
    .A(_06389_));
 sg13g2_nand2_1 _14685_ (.Y(_06391_),
    .A(_06388_),
    .B(_06390_));
 sg13g2_xnor2_1 _14686_ (.Y(_06392_),
    .A(_06374_),
    .B(_06391_));
 sg13g2_inv_1 _14687_ (.Y(_06393_),
    .A(_06291_));
 sg13g2_inv_1 _14688_ (.Y(_06394_),
    .A(_06297_));
 sg13g2_a21oi_1 _14689_ (.A1(_06394_),
    .A2(_06291_),
    .Y(_06395_),
    .B1(_06304_));
 sg13g2_a21oi_1 _14690_ (.A1(_06297_),
    .A2(_06393_),
    .Y(_06396_),
    .B1(_06395_));
 sg13g2_buf_4 fanout850 (.X(net850),
    .A(net851));
 sg13g2_o21ai_1 _14692_ (.B1(_06285_),
    .Y(_06398_),
    .A1(net1327),
    .A2(_06288_));
 sg13g2_nand3_1 _14693_ (.B(net216),
    .C(_06398_),
    .A(_04417_),
    .Y(_06399_));
 sg13g2_nor2_1 _14694_ (.A(_06288_),
    .B(_06285_),
    .Y(_06400_));
 sg13g2_a21oi_1 _14695_ (.A1(net1326),
    .A2(_06288_),
    .Y(_06401_),
    .B1(_06400_));
 sg13g2_nand2_2 _14696_ (.Y(_06402_),
    .A(_06399_),
    .B(_06401_));
 sg13g2_nand2_1 _14697_ (.Y(_06403_),
    .A(net1504),
    .B(_02283_));
 sg13g2_nor3_1 _14698_ (.A(net1876),
    .B(_06403_),
    .C(_05653_),
    .Y(_06404_));
 sg13g2_nand4_1 _14699_ (.B(_03897_),
    .C(net1877),
    .A(net1514),
    .Y(_06405_),
    .D(_05802_));
 sg13g2_nand2b_1 _14700_ (.Y(_06406_),
    .B(_06405_),
    .A_N(_06404_));
 sg13g2_a21oi_1 _14701_ (.A1(net162),
    .A2(net244),
    .Y(_06407_),
    .B1(net222));
 sg13g2_xnor2_1 _14702_ (.Y(_06408_),
    .A(net225),
    .B(_06407_));
 sg13g2_nand2b_1 _14703_ (.Y(_06409_),
    .B(_06408_),
    .A_N(_06406_));
 sg13g2_nand2_1 _14704_ (.Y(_06410_),
    .A(_04174_),
    .B(net166));
 sg13g2_buf_4 fanout849 (.X(net849),
    .A(\register_file_i/_2903_ ));
 sg13g2_nand2_1 _14706_ (.Y(_06412_),
    .A(net162),
    .B(net243));
 sg13g2_xnor2_1 _14707_ (.Y(_06413_),
    .A(net224),
    .B(_06412_));
 sg13g2_nand3_1 _14708_ (.B(_06410_),
    .C(_06413_),
    .A(_05658_),
    .Y(_06414_));
 sg13g2_o21ai_1 _14709_ (.B1(_06414_),
    .Y(_06415_),
    .A1(_05658_),
    .A2(_06409_));
 sg13g2_a21o_1 _14710_ (.A2(_03905_),
    .A1(_03911_),
    .B1(_04225_),
    .X(_06416_));
 sg13g2_nor3_1 _14711_ (.A(net1470),
    .B(net286),
    .C(net1515),
    .Y(_06417_));
 sg13g2_a21oi_1 _14712_ (.A1(net1517),
    .A2(_06416_),
    .Y(_06418_),
    .B1(_06417_));
 sg13g2_nor2_1 _14713_ (.A(net279),
    .B(net1502),
    .Y(_06419_));
 sg13g2_a221oi_1 _14714_ (.B2(_06419_),
    .C1(net1876),
    .B1(_06403_),
    .A1(net1505),
    .Y(_06420_),
    .A2(_04212_));
 sg13g2_a21o_1 _14715_ (.A2(_06418_),
    .A1(net1876),
    .B1(_06420_),
    .X(_06421_));
 sg13g2_nor2_1 _14716_ (.A(net1439),
    .B(net167),
    .Y(_06422_));
 sg13g2_nand2_1 _14717_ (.Y(_06423_),
    .A(_05658_),
    .B(_06422_));
 sg13g2_o21ai_1 _14718_ (.B1(_06423_),
    .Y(_06424_),
    .A1(net1371),
    .A2(_06421_));
 sg13g2_o21ai_1 _14719_ (.B1(_06321_),
    .Y(_06425_),
    .A1(_06415_),
    .A2(_06424_));
 sg13g2_xor2_1 _14720_ (.B(_06425_),
    .A(_06402_),
    .X(_06426_));
 sg13g2_xnor2_1 _14721_ (.Y(_06427_),
    .A(_06396_),
    .B(_06426_));
 sg13g2_xnor2_1 _14722_ (.Y(_06428_),
    .A(_06392_),
    .B(_06427_));
 sg13g2_buf_4 fanout848 (.X(net848),
    .A(net849));
 sg13g2_nand2b_1 _14724_ (.Y(_06430_),
    .B(_05206_),
    .A_N(_06422_));
 sg13g2_xnor2_1 _14725_ (.Y(_06431_),
    .A(net224),
    .B(_06319_));
 sg13g2_nand3_1 _14726_ (.B(_06421_),
    .C(_06431_),
    .A(net214),
    .Y(_06432_));
 sg13g2_o21ai_1 _14727_ (.B1(_06432_),
    .Y(_06433_),
    .A1(net214),
    .A2(_06430_));
 sg13g2_nand2b_1 _14728_ (.Y(_06434_),
    .B(_06433_),
    .A_N(_06415_));
 sg13g2_nand2_1 _14729_ (.Y(_06435_),
    .A(net1371),
    .B(_06410_));
 sg13g2_o21ai_1 _14730_ (.B1(_06435_),
    .Y(_06436_),
    .A1(net1371),
    .A2(_06406_));
 sg13g2_a21oi_1 _14731_ (.A1(_06088_),
    .A2(_06436_),
    .Y(_06437_),
    .B1(_06218_));
 sg13g2_o21ai_1 _14732_ (.B1(_06434_),
    .Y(_06438_),
    .A1(_06308_),
    .A2(_06321_));
 sg13g2_nand2_1 _14733_ (.Y(_06439_),
    .A(_06312_),
    .B(_06438_));
 sg13g2_o21ai_1 _14734_ (.B1(_06439_),
    .Y(_06440_),
    .A1(_06434_),
    .A2(_06437_));
 sg13g2_nand2b_1 _14735_ (.Y(_06441_),
    .B(_06327_),
    .A_N(_06306_));
 sg13g2_nand2_1 _14736_ (.Y(_06442_),
    .A(_06328_),
    .B(_06441_));
 sg13g2_xor2_1 _14737_ (.B(_06442_),
    .A(_06440_),
    .X(_06443_));
 sg13g2_xnor2_1 _14738_ (.Y(_06444_),
    .A(_06428_),
    .B(_06443_));
 sg13g2_o21ai_1 _14739_ (.B1(_06330_),
    .Y(_06445_),
    .A1(_06179_),
    .A2(_06269_));
 sg13g2_nand2_1 _14740_ (.Y(_06446_),
    .A(_06179_),
    .B(_06275_));
 sg13g2_a21oi_1 _14741_ (.A1(_06445_),
    .A2(_06446_),
    .Y(_06447_),
    .B1(_06277_));
 sg13g2_nand2_1 _14742_ (.Y(_06448_),
    .A(_06269_),
    .B(_06330_));
 sg13g2_a21oi_1 _14743_ (.A1(_06278_),
    .A2(_06448_),
    .Y(_06449_),
    .B1(_06271_));
 sg13g2_inv_1 _14744_ (.Y(_06450_),
    .A(_06330_));
 sg13g2_a21oi_1 _14745_ (.A1(_06278_),
    .A2(_06280_),
    .Y(_06451_),
    .B1(_06450_));
 sg13g2_nor4_2 _14746_ (.A(_06281_),
    .B(_06447_),
    .C(_06449_),
    .Y(_06452_),
    .D(_06451_));
 sg13g2_xnor2_1 _14747_ (.Y(_06453_),
    .A(_06444_),
    .B(_06452_));
 sg13g2_xnor2_1 _14748_ (.Y(_06454_),
    .A(_06367_),
    .B(_06453_));
 sg13g2_xnor2_1 _14749_ (.Y(_06455_),
    .A(_06362_),
    .B(_06454_));
 sg13g2_inv_1 _14750_ (.Y(_06456_),
    .A(_06153_));
 sg13g2_nand2_1 _14751_ (.Y(_06457_),
    .A(_05991_),
    .B(_06148_));
 sg13g2_inv_1 _14752_ (.Y(_06458_),
    .A(_05885_));
 sg13g2_nand3_1 _14753_ (.B(_05774_),
    .C(_06458_),
    .A(_05760_),
    .Y(_06459_));
 sg13g2_a21oi_1 _14754_ (.A1(_05756_),
    .A2(_05907_),
    .Y(_06460_),
    .B1(_05885_));
 sg13g2_nor3_1 _14755_ (.A(_06153_),
    .B(_06150_),
    .C(_06460_),
    .Y(_06461_));
 sg13g2_nand2b_1 _14756_ (.Y(_06462_),
    .B(_06341_),
    .A_N(_06237_));
 sg13g2_a221oi_1 _14757_ (.B2(_06461_),
    .C1(_06462_),
    .B1(_06459_),
    .A1(_06456_),
    .Y(_06463_),
    .A2(_06457_));
 sg13g2_nand2b_1 _14758_ (.Y(_06464_),
    .B(_06339_),
    .A_N(_06265_));
 sg13g2_inv_1 _14759_ (.Y(_06465_),
    .A(_06339_));
 sg13g2_a21oi_1 _14760_ (.A1(_06265_),
    .A2(_06465_),
    .Y(_06466_),
    .B1(_06267_));
 sg13g2_a22oi_1 _14761_ (.Y(_06467_),
    .B1(_06464_),
    .B2(_06466_),
    .A2(_06236_),
    .A1(_06156_));
 sg13g2_xnor2_1 _14762_ (.Y(_06468_),
    .A(_06265_),
    .B(_06465_));
 sg13g2_and2_1 _14763_ (.A(_06267_),
    .B(_06468_),
    .X(_06469_));
 sg13g2_nor2_1 _14764_ (.A(_06467_),
    .B(_06469_),
    .Y(_06470_));
 sg13g2_nor2_1 _14765_ (.A(_06463_),
    .B(_06470_),
    .Y(_06471_));
 sg13g2_xor2_1 _14766_ (.B(_06471_),
    .A(_06455_),
    .X(_06472_));
 sg13g2_nand2_1 _14767_ (.Y(_06473_),
    .A(net299),
    .B(_04558_));
 sg13g2_o21ai_1 _14768_ (.B1(_06473_),
    .Y(_06474_),
    .A1(net297),
    .A2(_06472_));
 sg13g2_nor2_1 _14769_ (.A(_03174_),
    .B(net1005),
    .Y(_06475_));
 sg13g2_a21oi_1 _14770_ (.A1(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .A2(net1005),
    .Y(_06476_),
    .B1(_06475_));
 sg13g2_a21oi_1 _14771_ (.A1(_04195_),
    .A2(_06245_),
    .Y(_06477_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_22_ ));
 sg13g2_mux2_1 _14772_ (.A0(_06476_),
    .A1(_06477_),
    .S(net306),
    .X(_06478_));
 sg13g2_nand2_1 _14773_ (.Y(_06479_),
    .A(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .B(net1219));
 sg13g2_o21ai_1 _14774_ (.B1(_06479_),
    .Y(_06480_),
    .A1(_03174_),
    .A2(net1219));
 sg13g2_o21ai_1 _14775_ (.B1(net1635),
    .Y(_06481_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ),
    .A2(net304));
 sg13g2_nand2_1 _14776_ (.Y(_06482_),
    .A(net1569),
    .B(_06481_));
 sg13g2_a221oi_1 _14777_ (.B2(net419),
    .C1(_06482_),
    .B1(_06480_),
    .A1(net1883),
    .Y(_06483_),
    .A2(_06348_));
 sg13g2_o21ai_1 _14778_ (.B1(_06483_),
    .Y(_06484_),
    .A1(net1708),
    .A2(_06478_));
 sg13g2_o21ai_1 _14779_ (.B1(_06484_),
    .Y(_06485_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .A2(net1572));
 sg13g2_a21oi_1 _14780_ (.A1(net1579),
    .A2(_06485_),
    .Y(_06486_),
    .B1(net376));
 sg13g2_o21ai_1 _14781_ (.B1(_06486_),
    .Y(_06487_),
    .A1(net1579),
    .A2(_06474_));
 sg13g2_nand2_1 _14782_ (.Y(_06488_),
    .A(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .B(net93));
 sg13g2_o21ai_1 _14783_ (.B1(_06488_),
    .Y(_00145_),
    .A1(net94),
    .A2(_06487_));
 sg13g2_nand2_1 _14784_ (.Y(_06489_),
    .A(net1185),
    .B(_04401_));
 sg13g2_o21ai_1 _14785_ (.B1(_06467_),
    .Y(_06490_),
    .A1(_06154_),
    .A2(_06257_));
 sg13g2_a21oi_1 _14786_ (.A1(_06265_),
    .A2(_06366_),
    .Y(_06491_),
    .B1(_06364_));
 sg13g2_xor2_1 _14787_ (.B(_06491_),
    .A(_06453_),
    .X(_06492_));
 sg13g2_a21oi_1 _14788_ (.A1(_06362_),
    .A2(_06492_),
    .Y(_06493_),
    .B1(_06469_));
 sg13g2_and2_1 _14789_ (.A(_06361_),
    .B(_06454_),
    .X(_06494_));
 sg13g2_a21oi_1 _14790_ (.A1(_06490_),
    .A2(_06493_),
    .Y(_06495_),
    .B1(_06494_));
 sg13g2_nand2_1 _14791_ (.Y(_06496_),
    .A(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .B(net319));
 sg13g2_buf_4 fanout847 (.X(net847),
    .A(net849));
 sg13g2_a21oi_2 _14793_ (.B1(net1565),
    .Y(_06498_),
    .A2(_06496_),
    .A1(net1567));
 sg13g2_nor2_1 _14794_ (.A(_06444_),
    .B(_06452_),
    .Y(_06499_));
 sg13g2_inv_1 _14795_ (.Y(_06500_),
    .A(_06499_));
 sg13g2_and2_1 _14796_ (.A(_06444_),
    .B(_06452_),
    .X(_06501_));
 sg13g2_a21oi_1 _14797_ (.A1(_06367_),
    .A2(_06500_),
    .Y(_06502_),
    .B1(_06501_));
 sg13g2_xnor2_1 _14798_ (.Y(_06503_),
    .A(net1374),
    .B(_06370_));
 sg13g2_xnor2_1 _14799_ (.Y(_06504_),
    .A(net1337),
    .B(_06371_));
 sg13g2_nor2_1 _14800_ (.A(_06503_),
    .B(_06504_),
    .Y(_06505_));
 sg13g2_nand2_1 _14801_ (.Y(_06506_),
    .A(_06503_),
    .B(_06504_));
 sg13g2_o21ai_1 _14802_ (.B1(_06506_),
    .Y(_06507_),
    .A1(_06369_),
    .A2(_06505_));
 sg13g2_a22oi_1 _14803_ (.Y(_06508_),
    .B1(net1433),
    .B2(net1334),
    .A2(net1435),
    .A1(net137));
 sg13g2_xnor2_1 _14804_ (.Y(_06509_),
    .A(_05835_),
    .B(_06508_));
 sg13g2_a22oi_1 _14805_ (.Y(_06510_),
    .B1(net242),
    .B2(net1339),
    .A2(net1322),
    .A1(net139));
 sg13g2_nand2_2 _14806_ (.Y(_06511_),
    .A(_04736_),
    .B(net213));
 sg13g2_xor2_1 _14807_ (.B(_06511_),
    .A(_06510_),
    .X(_06512_));
 sg13g2_xnor2_1 _14808_ (.Y(_06513_),
    .A(_06509_),
    .B(_06512_));
 sg13g2_and2_1 _14809_ (.A(net246),
    .B(net1332),
    .X(_06514_));
 sg13g2_a21o_1 _14810_ (.A2(net136),
    .A1(net250),
    .B1(_06514_),
    .X(_06515_));
 sg13g2_xnor2_1 _14811_ (.Y(_06516_),
    .A(_05532_),
    .B(_06515_));
 sg13g2_a22oi_1 _14812_ (.Y(_06517_),
    .B1(net91),
    .B2(net251),
    .A2(net1258),
    .A1(net1437));
 sg13g2_a21oi_1 _14813_ (.A1(net265),
    .A2(net1321),
    .Y(_06518_),
    .B1(net1373));
 sg13g2_xnor2_1 _14814_ (.Y(_06519_),
    .A(_06517_),
    .B(_06518_));
 sg13g2_xor2_1 _14815_ (.B(_06519_),
    .A(_06516_),
    .X(_06520_));
 sg13g2_xnor2_1 _14816_ (.Y(_06521_),
    .A(_06513_),
    .B(_06520_));
 sg13g2_xnor2_1 _14817_ (.Y(_06522_),
    .A(_06507_),
    .B(_06521_));
 sg13g2_nand2b_1 _14818_ (.Y(_06523_),
    .B(_06387_),
    .A_N(_06374_));
 sg13g2_nor2b_1 _14819_ (.A(_06387_),
    .B_N(_06374_),
    .Y(_06524_));
 sg13g2_a21oi_1 _14820_ (.A1(_06381_),
    .A2(_06523_),
    .Y(_06525_),
    .B1(_06524_));
 sg13g2_nand2b_1 _14821_ (.Y(_06526_),
    .B(_06431_),
    .A_N(_06421_));
 sg13g2_nand2_1 _14822_ (.Y(_06527_),
    .A(_05206_),
    .B(_06422_));
 sg13g2_mux2_2 _14823_ (.A0(_06526_),
    .A1(_06527_),
    .S(net1371),
    .X(_06528_));
 sg13g2_a21oi_1 _14824_ (.A1(net1321),
    .A2(_06378_),
    .Y(_06529_),
    .B1(_06376_));
 sg13g2_nor3_2 _14825_ (.A(net1473),
    .B(net1373),
    .C(_06529_),
    .Y(_06530_));
 sg13g2_nand2_1 _14826_ (.Y(_06531_),
    .A(_06376_),
    .B(_06378_));
 sg13g2_o21ai_1 _14827_ (.B1(_06531_),
    .Y(_06532_),
    .A1(net1321),
    .A2(_06378_));
 sg13g2_nor3_2 _14828_ (.A(_06528_),
    .B(_06530_),
    .C(_06532_),
    .Y(_06533_));
 sg13g2_o21ai_1 _14829_ (.B1(_06528_),
    .Y(_06534_),
    .A1(_06530_),
    .A2(_06532_));
 sg13g2_nor2b_1 _14830_ (.A(_06533_),
    .B_N(_06534_),
    .Y(_06535_));
 sg13g2_xnor2_1 _14831_ (.Y(_06536_),
    .A(_06525_),
    .B(_06535_));
 sg13g2_xnor2_1 _14832_ (.Y(_06537_),
    .A(_06522_),
    .B(_06536_));
 sg13g2_a21o_1 _14833_ (.A2(_06291_),
    .A1(_06304_),
    .B1(_06394_),
    .X(_06538_));
 sg13g2_o21ai_1 _14834_ (.B1(_06538_),
    .Y(_06539_),
    .A1(_06304_),
    .A2(_06291_));
 sg13g2_nand2b_1 _14835_ (.Y(_06540_),
    .B(_06539_),
    .A_N(_06402_));
 sg13g2_nor2b_1 _14836_ (.A(_06539_),
    .B_N(_06402_),
    .Y(_06541_));
 sg13g2_a21oi_1 _14837_ (.A1(_06392_),
    .A2(_06540_),
    .Y(_06542_),
    .B1(_06541_));
 sg13g2_nand2_2 _14838_ (.Y(_06543_),
    .A(_06415_),
    .B(_06433_));
 sg13g2_nor2_1 _14839_ (.A(_06402_),
    .B(_06543_),
    .Y(_06544_));
 sg13g2_and2_1 _14840_ (.A(_06392_),
    .B(_06543_),
    .X(_06545_));
 sg13g2_inv_1 _14841_ (.Y(_06546_),
    .A(_06528_));
 sg13g2_o21ai_1 _14842_ (.B1(_06543_),
    .Y(_06547_),
    .A1(_06402_),
    .A2(_06546_));
 sg13g2_a21oi_1 _14843_ (.A1(_06539_),
    .A2(_06547_),
    .Y(_06548_),
    .B1(_06544_));
 sg13g2_nor2_1 _14844_ (.A(_06392_),
    .B(_06548_),
    .Y(_06549_));
 sg13g2_a221oi_1 _14845_ (.B2(_06541_),
    .C1(_06549_),
    .B1(_06545_),
    .A1(_06539_),
    .Y(_06550_),
    .A2(_06544_));
 sg13g2_o21ai_1 _14846_ (.B1(_06550_),
    .Y(_06551_),
    .A1(_06528_),
    .A2(_06542_));
 sg13g2_xor2_1 _14847_ (.B(_06551_),
    .A(_06537_),
    .X(_06552_));
 sg13g2_nand2b_1 _14848_ (.Y(_06553_),
    .B(_06326_),
    .A_N(_06206_));
 sg13g2_nor2_1 _14849_ (.A(_06306_),
    .B(_06323_),
    .Y(_06554_));
 sg13g2_a21oi_1 _14850_ (.A1(_06324_),
    .A2(_06553_),
    .Y(_06555_),
    .B1(_06554_));
 sg13g2_a21oi_1 _14851_ (.A1(_06306_),
    .A2(_06323_),
    .Y(_06556_),
    .B1(_06555_));
 sg13g2_nand2_1 _14852_ (.Y(_06557_),
    .A(_06440_),
    .B(_06556_));
 sg13g2_nor2_1 _14853_ (.A(_06440_),
    .B(_06556_),
    .Y(_06558_));
 sg13g2_a21oi_2 _14854_ (.B1(_06558_),
    .Y(_06559_),
    .A2(_06557_),
    .A1(_06428_));
 sg13g2_xnor2_1 _14855_ (.Y(_06560_),
    .A(_06552_),
    .B(_06559_));
 sg13g2_xor2_1 _14856_ (.B(_06560_),
    .A(_06502_),
    .X(_06561_));
 sg13g2_xor2_1 _14857_ (.B(_06561_),
    .A(_06498_),
    .X(_06562_));
 sg13g2_xnor2_1 _14858_ (.Y(_06563_),
    .A(_06495_),
    .B(_06562_));
 sg13g2_nor2_1 _14859_ (.A(net1539),
    .B(_04656_),
    .Y(_06564_));
 sg13g2_a21oi_2 _14860_ (.B1(_06564_),
    .Y(_06565_),
    .A2(_06563_),
    .A1(net1539));
 sg13g2_a21oi_1 _14861_ (.A1(_04195_),
    .A2(_06346_),
    .Y(_06566_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_23_ ));
 sg13g2_nor2_1 _14862_ (.A(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .B(net1009),
    .Y(_06567_));
 sg13g2_a21oi_1 _14863_ (.A1(_03278_),
    .A2(net1009),
    .Y(_06568_),
    .B1(_06567_));
 sg13g2_nor2_1 _14864_ (.A(net309),
    .B(_06568_),
    .Y(_06569_));
 sg13g2_a21oi_1 _14865_ (.A1(net314),
    .A2(_06566_),
    .Y(_06570_),
    .B1(_06569_));
 sg13g2_nor2_1 _14866_ (.A(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .B(net1266),
    .Y(_06571_));
 sg13g2_a21oi_1 _14867_ (.A1(_03278_),
    .A2(net1266),
    .Y(_06572_),
    .B1(_06571_));
 sg13g2_nand2_1 _14868_ (.Y(_06573_),
    .A(net420),
    .B(_06572_));
 sg13g2_o21ai_1 _14869_ (.B1(net1635),
    .Y(_06574_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ),
    .A2(net311));
 sg13g2_nand2b_1 _14870_ (.Y(_06575_),
    .B(net1883),
    .A_N(_06476_));
 sg13g2_nand4_1 _14871_ (.B(_06573_),
    .C(_06574_),
    .A(net1569),
    .Y(_06576_),
    .D(_06575_));
 sg13g2_a21oi_1 _14872_ (.A1(net1891),
    .A2(_06570_),
    .Y(_06577_),
    .B1(_06576_));
 sg13g2_o21ai_1 _14873_ (.B1(net1187),
    .Y(_06578_),
    .A1(net337),
    .A2(_06577_));
 sg13g2_o21ai_1 _14874_ (.B1(_06578_),
    .Y(_06579_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .A2(net1181));
 sg13g2_o21ai_1 _14875_ (.B1(_06579_),
    .Y(_00146_),
    .A1(_06489_),
    .A2(_06565_));
 sg13g2_a21oi_1 _14876_ (.A1(_06455_),
    .A2(_06463_),
    .Y(_06580_),
    .B1(_06494_));
 sg13g2_o21ai_1 _14877_ (.B1(_06256_),
    .Y(_06581_),
    .A1(_06267_),
    .A2(_06468_));
 sg13g2_a22oi_1 _14878_ (.Y(_06582_),
    .B1(_06493_),
    .B2(_06581_),
    .A2(_06561_),
    .A1(_06498_));
 sg13g2_nor2_1 _14879_ (.A(_06498_),
    .B(_06561_),
    .Y(_06583_));
 sg13g2_a21oi_1 _14880_ (.A1(_06580_),
    .A2(_06582_),
    .Y(_06584_),
    .B1(_06583_));
 sg13g2_buf_4 fanout846 (.X(net846),
    .A(\register_file_i/_2907_ ));
 sg13g2_nand2_1 _14882_ (.Y(_06586_),
    .A(\ex_block_i.alu_i.imd_val_q_i_56_ ),
    .B(net321));
 sg13g2_a21oi_2 _14883_ (.B1(net1565),
    .Y(_06587_),
    .A2(_06586_),
    .A1(net1567));
 sg13g2_inv_1 _14884_ (.Y(_06588_),
    .A(_06587_));
 sg13g2_inv_1 _14885_ (.Y(_06589_),
    .A(_06392_));
 sg13g2_o21ai_1 _14886_ (.B1(_06537_),
    .Y(_06590_),
    .A1(_06392_),
    .A2(_06543_));
 sg13g2_o21ai_1 _14887_ (.B1(_06590_),
    .Y(_06591_),
    .A1(_06589_),
    .A2(_06528_));
 sg13g2_nor2_1 _14888_ (.A(_06537_),
    .B(_06541_),
    .Y(_06592_));
 sg13g2_nor2_1 _14889_ (.A(_06546_),
    .B(_06545_),
    .Y(_06593_));
 sg13g2_nor2_1 _14890_ (.A(_06592_),
    .B(_06593_),
    .Y(_06594_));
 sg13g2_a221oi_1 _14891_ (.B2(_06540_),
    .C1(_06594_),
    .B1(_06591_),
    .A1(_06537_),
    .Y(_06595_),
    .A2(_06541_));
 sg13g2_a22oi_1 _14892_ (.Y(_06596_),
    .B1(net135),
    .B2(net247),
    .A2(net1331),
    .A1(net1435));
 sg13g2_xnor2_1 _14893_ (.Y(_06597_),
    .A(net1328),
    .B(_06596_));
 sg13g2_a22oi_1 _14894_ (.Y(_06598_),
    .B1(net91),
    .B2(net1438),
    .A2(net1258),
    .A1(net248));
 sg13g2_nor2_1 _14895_ (.A(net252),
    .B(net1257),
    .Y(_06599_));
 sg13g2_xnor2_1 _14896_ (.Y(_06600_),
    .A(_06598_),
    .B(_06599_));
 sg13g2_xnor2_1 _14897_ (.Y(_06601_),
    .A(_06597_),
    .B(_06600_));
 sg13g2_a22oi_1 _14898_ (.Y(_06602_),
    .B1(net213),
    .B2(net1339),
    .A2(net245),
    .A1(net139));
 sg13g2_xnor2_1 _14899_ (.Y(_06603_),
    .A(net1337),
    .B(_06602_));
 sg13g2_a22oi_1 _14900_ (.Y(_06604_),
    .B1(net1322),
    .B2(net1334),
    .A2(net1433),
    .A1(net137));
 sg13g2_xnor2_1 _14901_ (.Y(_06605_),
    .A(net1374),
    .B(_06604_));
 sg13g2_xnor2_1 _14902_ (.Y(_06606_),
    .A(_06603_),
    .B(_06605_));
 sg13g2_xnor2_1 _14903_ (.Y(_06607_),
    .A(net1337),
    .B(_06510_));
 sg13g2_xnor2_1 _14904_ (.Y(_06608_),
    .A(net1374),
    .B(_06508_));
 sg13g2_nor2_1 _14905_ (.A(_06607_),
    .B(_06608_),
    .Y(_06609_));
 sg13g2_xnor2_1 _14906_ (.Y(_06610_),
    .A(net158),
    .B(_06511_));
 sg13g2_nand2_1 _14907_ (.Y(_06611_),
    .A(_06607_),
    .B(_06608_));
 sg13g2_nor2_1 _14908_ (.A(_06611_),
    .B(_06610_),
    .Y(_06612_));
 sg13g2_a21oi_1 _14909_ (.A1(_06609_),
    .A2(_06610_),
    .Y(_06613_),
    .B1(_06612_));
 sg13g2_xnor2_1 _14910_ (.Y(_06614_),
    .A(_06606_),
    .B(_06613_));
 sg13g2_xnor2_1 _14911_ (.Y(_06615_),
    .A(_06601_),
    .B(_06614_));
 sg13g2_xor2_1 _14912_ (.B(_06515_),
    .A(net1328),
    .X(_06616_));
 sg13g2_o21ai_1 _14913_ (.B1(_06616_),
    .Y(_06617_),
    .A1(net265),
    .A2(net1326));
 sg13g2_nor2_1 _14914_ (.A(net1326),
    .B(_06616_),
    .Y(_06618_));
 sg13g2_a21oi_1 _14915_ (.A1(_05684_),
    .A2(_06617_),
    .Y(_06619_),
    .B1(_06618_));
 sg13g2_nand2_1 _14916_ (.Y(_06620_),
    .A(net1326),
    .B(_06517_));
 sg13g2_a21oi_1 _14917_ (.A1(net1372),
    .A2(_06616_),
    .Y(_06621_),
    .B1(_06620_));
 sg13g2_nor3_1 _14918_ (.A(net265),
    .B(net1372),
    .C(_06616_),
    .Y(_06622_));
 sg13g2_nor2_1 _14919_ (.A(_06621_),
    .B(_06622_),
    .Y(_06623_));
 sg13g2_o21ai_1 _14920_ (.B1(_06623_),
    .Y(_06624_),
    .A1(_06517_),
    .A2(_06619_));
 sg13g2_a21oi_1 _14921_ (.A1(_06369_),
    .A2(_06506_),
    .Y(_06625_),
    .B1(_06505_));
 sg13g2_a21o_1 _14922_ (.A2(_06625_),
    .A1(_06513_),
    .B1(_06520_),
    .X(_06626_));
 sg13g2_o21ai_1 _14923_ (.B1(_06626_),
    .Y(_06627_),
    .A1(_06513_),
    .A2(_06625_));
 sg13g2_xor2_1 _14924_ (.B(_06627_),
    .A(_06624_),
    .X(_06628_));
 sg13g2_xnor2_1 _14925_ (.Y(_06629_),
    .A(_06615_),
    .B(_06628_));
 sg13g2_o21ai_1 _14926_ (.B1(_06388_),
    .Y(_06630_),
    .A1(_06374_),
    .A2(_06389_));
 sg13g2_a21o_1 _14927_ (.A2(_06534_),
    .A1(_06522_),
    .B1(_06533_),
    .X(_06631_));
 sg13g2_a21oi_1 _14928_ (.A1(_06374_),
    .A2(_06388_),
    .Y(_06632_),
    .B1(_06389_));
 sg13g2_nor3_1 _14929_ (.A(_06522_),
    .B(_06534_),
    .C(_06632_),
    .Y(_06633_));
 sg13g2_a221oi_1 _14930_ (.B2(_06631_),
    .C1(_06633_),
    .B1(_06630_),
    .A1(_06522_),
    .Y(_06634_),
    .A2(_06533_));
 sg13g2_xnor2_1 _14931_ (.Y(_06635_),
    .A(_06629_),
    .B(_06634_));
 sg13g2_xnor2_1 _14932_ (.Y(_06636_),
    .A(_06595_),
    .B(_06635_));
 sg13g2_or2_1 _14933_ (.X(_06637_),
    .B(_06491_),
    .A(_06501_));
 sg13g2_nor2_1 _14934_ (.A(_06552_),
    .B(_06559_),
    .Y(_06638_));
 sg13g2_nor2_1 _14935_ (.A(_06499_),
    .B(_06638_),
    .Y(_06639_));
 sg13g2_a22oi_1 _14936_ (.Y(_06640_),
    .B1(_06637_),
    .B2(_06639_),
    .A2(_06559_),
    .A1(_06552_));
 sg13g2_xnor2_1 _14937_ (.Y(_06641_),
    .A(_06636_),
    .B(_06640_));
 sg13g2_nand2_1 _14938_ (.Y(_06642_),
    .A(_06552_),
    .B(_06559_));
 sg13g2_xor2_1 _14939_ (.B(_06642_),
    .A(_06636_),
    .X(_06643_));
 sg13g2_a21oi_1 _14940_ (.A1(_06587_),
    .A2(_06643_),
    .Y(_06644_),
    .B1(_06637_));
 sg13g2_a21oi_1 _14941_ (.A1(_06499_),
    .A2(_06642_),
    .Y(_06645_),
    .B1(_06638_));
 sg13g2_xnor2_1 _14942_ (.Y(_06646_),
    .A(_06636_),
    .B(_06645_));
 sg13g2_nor2_1 _14943_ (.A(_06367_),
    .B(_06501_),
    .Y(_06647_));
 sg13g2_a21oi_1 _14944_ (.A1(_06587_),
    .A2(_06646_),
    .Y(_06648_),
    .B1(_06647_));
 sg13g2_nor2_2 _14945_ (.A(_06644_),
    .B(_06648_),
    .Y(_06649_));
 sg13g2_a21oi_1 _14946_ (.A1(_06588_),
    .A2(_06641_),
    .Y(_06650_),
    .B1(_06649_));
 sg13g2_xnor2_1 _14947_ (.Y(_06651_),
    .A(_06584_),
    .B(_06650_));
 sg13g2_nor2_1 _14948_ (.A(net1538),
    .B(_04756_),
    .Y(_06652_));
 sg13g2_a21oi_2 _14949_ (.B1(_06652_),
    .Y(_06653_),
    .A2(_06651_),
    .A1(net1539));
 sg13g2_nor2_1 _14950_ (.A(net556),
    .B(net1572),
    .Y(_06654_));
 sg13g2_a21oi_1 _14951_ (.A1(_04761_),
    .A2(_05632_),
    .Y(_06655_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_24_ ));
 sg13g2_mux2_1 _14952_ (.A0(net556),
    .A1(data_addr_o_24_),
    .S(net1007),
    .X(_06656_));
 sg13g2_nor2_1 _14953_ (.A(net306),
    .B(_06656_),
    .Y(_06657_));
 sg13g2_a21oi_1 _14954_ (.A1(net313),
    .A2(_06655_),
    .Y(_06658_),
    .B1(_06657_));
 sg13g2_mux2_1 _14955_ (.A0(net556),
    .A1(data_addr_o_24_),
    .S(net1260),
    .X(_06659_));
 sg13g2_nand2_1 _14956_ (.Y(_06660_),
    .A(net419),
    .B(_06659_));
 sg13g2_o21ai_1 _14957_ (.B1(net1634),
    .Y(_06661_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ),
    .A2(net306));
 sg13g2_nand3_1 _14958_ (.B(_06660_),
    .C(_06661_),
    .A(net1569),
    .Y(_06662_));
 sg13g2_a221oi_1 _14959_ (.B2(net1888),
    .C1(_06662_),
    .B1(_06658_),
    .A1(net1883),
    .Y(_06663_),
    .A2(_06568_));
 sg13g2_nor3_1 _14960_ (.A(net338),
    .B(_06654_),
    .C(_06663_),
    .Y(_06664_));
 sg13g2_a21oi_1 _14961_ (.A1(net342),
    .A2(_06653_),
    .Y(_06665_),
    .B1(_06664_));
 sg13g2_nor3_1 _14962_ (.A(net376),
    .B(net94),
    .C(_06665_),
    .Y(_06666_));
 sg13g2_a21o_1 _14963_ (.A2(net95),
    .A1(net556),
    .B1(_06666_),
    .X(_00147_));
 sg13g2_a221oi_1 _14964_ (.B2(_06641_),
    .C1(_06583_),
    .B1(_06588_),
    .A1(_06580_),
    .Y(_06667_),
    .A2(_06582_));
 sg13g2_nor2_1 _14965_ (.A(_06649_),
    .B(_06667_),
    .Y(_06668_));
 sg13g2_nand2_1 _14966_ (.Y(_06669_),
    .A(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .B(net321));
 sg13g2_a21o_2 _14967_ (.A2(_06669_),
    .A1(net1567),
    .B1(net1565),
    .X(_06670_));
 sg13g2_o21ai_1 _14968_ (.B1(_06611_),
    .Y(_06671_),
    .A1(_06601_),
    .A2(_06606_));
 sg13g2_inv_1 _14969_ (.Y(_06672_),
    .A(_06671_));
 sg13g2_a21oi_1 _14970_ (.A1(_06601_),
    .A2(_06606_),
    .Y(_06673_),
    .B1(_06672_));
 sg13g2_xor2_1 _14971_ (.B(_06511_),
    .A(net157),
    .X(_06674_));
 sg13g2_nor2_1 _14972_ (.A(_06601_),
    .B(_06609_),
    .Y(_06675_));
 sg13g2_nor3_1 _14973_ (.A(_06606_),
    .B(_06674_),
    .C(_06675_),
    .Y(_06676_));
 sg13g2_a21oi_1 _14974_ (.A1(_06601_),
    .A2(_06609_),
    .Y(_06677_),
    .B1(_06676_));
 sg13g2_o21ai_1 _14975_ (.B1(_06677_),
    .Y(_06678_),
    .A1(_06610_),
    .A2(_06673_));
 sg13g2_buf_4 fanout845 (.X(net845),
    .A(net846));
 sg13g2_o21ai_1 _14977_ (.B1(_06597_),
    .Y(_06680_),
    .A1(net1325),
    .A2(_06598_));
 sg13g2_nand3_1 _14978_ (.B(net216),
    .C(_06680_),
    .A(_04791_),
    .Y(_06681_));
 sg13g2_nor2_1 _14979_ (.A(_06598_),
    .B(_06597_),
    .Y(_06682_));
 sg13g2_a21oi_1 _14980_ (.A1(net1325),
    .A2(_06598_),
    .Y(_06683_),
    .B1(_06682_));
 sg13g2_nand2_2 _14981_ (.Y(_06684_),
    .A(_06681_),
    .B(_06683_));
 sg13g2_nand2_1 _14982_ (.Y(_06685_),
    .A(_06603_),
    .B(_06605_));
 sg13g2_nor2_1 _14983_ (.A(_06603_),
    .B(_06605_),
    .Y(_06686_));
 sg13g2_nand2_1 _14984_ (.Y(_06687_),
    .A(_06610_),
    .B(_06686_));
 sg13g2_o21ai_1 _14985_ (.B1(_06687_),
    .Y(_06688_),
    .A1(_06610_),
    .A2(_06685_));
 sg13g2_a22oi_1 _14986_ (.Y(_06689_),
    .B1(net135),
    .B2(net1435),
    .A2(net1433),
    .A1(net1331));
 sg13g2_xnor2_1 _14987_ (.Y(_06690_),
    .A(net1328),
    .B(_06689_));
 sg13g2_a22oi_1 _14988_ (.Y(_06691_),
    .B1(net91),
    .B2(net250),
    .A2(net1259),
    .A1(net246));
 sg13g2_nor2_1 _14989_ (.A(net1438),
    .B(net1257),
    .Y(_06692_));
 sg13g2_xnor2_1 _14990_ (.Y(_06693_),
    .A(_06691_),
    .B(_06692_));
 sg13g2_xnor2_1 _14991_ (.Y(_06694_),
    .A(_06690_),
    .B(_06693_));
 sg13g2_nor3_1 _14992_ (.A(net1493),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ),
    .C(net1495),
    .Y(_06695_));
 sg13g2_nor3_1 _14993_ (.A(_03882_),
    .B(_02058_),
    .C(_01990_),
    .Y(_06696_));
 sg13g2_nor3_1 _14994_ (.A(net1865),
    .B(_06695_),
    .C(_06696_),
    .Y(_06697_));
 sg13g2_nor3_1 _14995_ (.A(net281),
    .B(net1463),
    .C(net1464),
    .Y(_06698_));
 sg13g2_and3_1 _14996_ (.X(_06699_),
    .A(net281),
    .B(net1463),
    .C(net1464));
 sg13g2_nor3_1 _14997_ (.A(net1874),
    .B(_06698_),
    .C(_06699_),
    .Y(_06700_));
 sg13g2_o21ai_1 _14998_ (.B1(net214),
    .Y(_06701_),
    .A1(_06697_),
    .A2(_06700_));
 sg13g2_xor2_1 _14999_ (.B(_06701_),
    .A(net1338),
    .X(_06702_));
 sg13g2_a22oi_1 _15000_ (.Y(_06703_),
    .B1(net242),
    .B2(net1334),
    .A2(net1322),
    .A1(net137));
 sg13g2_xnor2_1 _15001_ (.Y(_06704_),
    .A(net1374),
    .B(_06703_));
 sg13g2_xor2_1 _15002_ (.B(_06704_),
    .A(_06702_),
    .X(_06705_));
 sg13g2_xnor2_1 _15003_ (.Y(_06706_),
    .A(_06694_),
    .B(_06705_));
 sg13g2_xnor2_1 _15004_ (.Y(_06707_),
    .A(_06688_),
    .B(_06706_));
 sg13g2_xnor2_1 _15005_ (.Y(_06708_),
    .A(_06684_),
    .B(_06707_));
 sg13g2_xnor2_1 _15006_ (.Y(_06709_),
    .A(_06678_),
    .B(_06708_));
 sg13g2_o21ai_1 _15007_ (.B1(_06513_),
    .Y(_06710_),
    .A1(_06520_),
    .A2(_06507_));
 sg13g2_nand2_1 _15008_ (.Y(_06711_),
    .A(_06520_),
    .B(_06507_));
 sg13g2_and2_1 _15009_ (.A(_06710_),
    .B(_06711_),
    .X(_06712_));
 sg13g2_or2_1 _15010_ (.X(_06713_),
    .B(_06712_),
    .A(_06624_));
 sg13g2_nand2_1 _15011_ (.Y(_06714_),
    .A(_06624_),
    .B(_06712_));
 sg13g2_mux2_1 _15012_ (.A0(_06713_),
    .A1(_06714_),
    .S(_06615_),
    .X(_06715_));
 sg13g2_xnor2_1 _15013_ (.Y(_06716_),
    .A(_06709_),
    .B(_06715_));
 sg13g2_inv_1 _15014_ (.Y(_06717_),
    .A(_06522_));
 sg13g2_xor2_1 _15015_ (.B(_06628_),
    .A(_06615_),
    .X(_06718_));
 sg13g2_a21o_1 _15016_ (.A2(_06718_),
    .A1(_06534_),
    .B1(_06630_),
    .X(_06719_));
 sg13g2_o21ai_1 _15017_ (.B1(_06719_),
    .Y(_06720_),
    .A1(_06533_),
    .A2(_06718_));
 sg13g2_o21ai_1 _15018_ (.B1(_06534_),
    .Y(_06721_),
    .A1(_06533_),
    .A2(_06630_));
 sg13g2_a22oi_1 _15019_ (.Y(_06722_),
    .B1(_06721_),
    .B2(_06629_),
    .A2(_06720_),
    .A1(_06717_));
 sg13g2_and2_2 _15020_ (.A(_06716_),
    .B(_06722_),
    .X(_06723_));
 sg13g2_nor2_1 _15021_ (.A(_06716_),
    .B(_06722_),
    .Y(_06724_));
 sg13g2_buf_4 fanout844 (.X(net844),
    .A(\register_file_i/_2907_ ));
 sg13g2_nor2_2 _15023_ (.A(_06723_),
    .B(net1076),
    .Y(_06726_));
 sg13g2_nor3_1 _15024_ (.A(_06453_),
    .B(_06560_),
    .C(_06636_),
    .Y(_06727_));
 sg13g2_nor2_1 _15025_ (.A(_06265_),
    .B(_06465_),
    .Y(_06728_));
 sg13g2_o21ai_1 _15026_ (.B1(_06444_),
    .Y(_06729_),
    .A1(_06365_),
    .A2(_06452_));
 sg13g2_nand2_1 _15027_ (.Y(_06730_),
    .A(_06365_),
    .B(_06452_));
 sg13g2_a21o_1 _15028_ (.A2(_06730_),
    .A1(_06729_),
    .B1(_06638_),
    .X(_06731_));
 sg13g2_nor2_1 _15029_ (.A(_06595_),
    .B(_06635_),
    .Y(_06732_));
 sg13g2_a21oi_1 _15030_ (.A1(_06642_),
    .A2(_06731_),
    .Y(_06733_),
    .B1(_06732_));
 sg13g2_a221oi_1 _15031_ (.B2(_06728_),
    .C1(_06733_),
    .B1(_06727_),
    .A1(_06595_),
    .Y(_06734_),
    .A2(_06635_));
 sg13g2_buf_4 fanout843 (.X(net843),
    .A(net844));
 sg13g2_xor2_1 _15033_ (.B(net808),
    .A(_06726_),
    .X(_06736_));
 sg13g2_xnor2_1 _15034_ (.Y(_06737_),
    .A(_06670_),
    .B(_06736_));
 sg13g2_xnor2_1 _15035_ (.Y(_06738_),
    .A(_06668_),
    .B(_06737_));
 sg13g2_nand3_1 _15036_ (.B(net1188),
    .C(_04144_),
    .A(net1615),
    .Y(_06739_));
 sg13g2_nor2_1 _15037_ (.A(net1578),
    .B(net1541),
    .Y(_06740_));
 sg13g2_a21oi_1 _15038_ (.A1(_04761_),
    .A2(_05892_),
    .Y(_06741_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_25_ ));
 sg13g2_mux2_1 _15039_ (.A0(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .A1(data_addr_o_25_),
    .S(net1007),
    .X(_06742_));
 sg13g2_nor2_1 _15040_ (.A(net309),
    .B(_06742_),
    .Y(_06743_));
 sg13g2_a21oi_1 _15041_ (.A1(net314),
    .A2(_06741_),
    .Y(_06744_),
    .B1(_06743_));
 sg13g2_nor2_1 _15042_ (.A(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .B(net1572),
    .Y(_06745_));
 sg13g2_nor3_1 _15043_ (.A(_04066_),
    .B(net341),
    .C(_06745_),
    .Y(_06746_));
 sg13g2_mux2_1 _15044_ (.A0(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .A1(data_addr_o_25_),
    .S(net1260),
    .X(_06747_));
 sg13g2_o21ai_1 _15045_ (.B1(net1634),
    .Y(_06748_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ),
    .A2(net304));
 sg13g2_nand2_1 _15046_ (.Y(_06749_),
    .A(net1569),
    .B(_06748_));
 sg13g2_a221oi_1 _15047_ (.B2(net419),
    .C1(_06749_),
    .B1(_06747_),
    .A1(net1882),
    .Y(_06750_),
    .A2(_06656_));
 sg13g2_nor3_1 _15048_ (.A(net337),
    .B(_06745_),
    .C(_06750_),
    .Y(_06751_));
 sg13g2_a221oi_1 _15049_ (.B2(_06746_),
    .C1(_06751_),
    .B1(_06744_),
    .A1(_04901_),
    .Y(_06752_),
    .A2(_06740_));
 sg13g2_nor3_1 _15050_ (.A(net375),
    .B(net94),
    .C(_06752_),
    .Y(_06753_));
 sg13g2_a21oi_1 _15051_ (.A1(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .A2(net95),
    .Y(_06754_),
    .B1(_06753_));
 sg13g2_o21ai_1 _15052_ (.B1(_06754_),
    .Y(_00148_),
    .A1(_06738_),
    .A2(_06739_));
 sg13g2_and2_1 _15053_ (.A(_06670_),
    .B(_06736_),
    .X(_06755_));
 sg13g2_or2_1 _15054_ (.X(_06756_),
    .B(_06736_),
    .A(_06670_));
 sg13g2_o21ai_1 _15055_ (.B1(_06756_),
    .Y(_06757_),
    .A1(_06668_),
    .A2(_06755_));
 sg13g2_nand2_1 _15056_ (.Y(_06758_),
    .A(_06716_),
    .B(_06722_));
 sg13g2_o21ai_1 _15057_ (.B1(_06758_),
    .Y(_06759_),
    .A1(net1076),
    .A2(net808));
 sg13g2_nand2_1 _15058_ (.Y(_06760_),
    .A(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .B(net319));
 sg13g2_a21oi_1 _15059_ (.A1(net1567),
    .A2(_06760_),
    .Y(_06761_),
    .B1(net1565));
 sg13g2_buf_4 fanout842 (.X(net842),
    .A(net844));
 sg13g2_inv_1 _15061_ (.Y(_06763_),
    .A(_06709_));
 sg13g2_a21oi_1 _15062_ (.A1(_06709_),
    .A2(_06713_),
    .Y(_06764_),
    .B1(_06615_));
 sg13g2_a21oi_2 _15063_ (.B1(_06764_),
    .Y(_06765_),
    .A2(_06714_),
    .A1(_06763_));
 sg13g2_o21ai_1 _15064_ (.B1(_06707_),
    .Y(_06766_),
    .A1(_06684_),
    .A2(_06678_));
 sg13g2_nand2_1 _15065_ (.Y(_06767_),
    .A(_06684_),
    .B(_06678_));
 sg13g2_nand2_2 _15066_ (.Y(_06768_),
    .A(_06766_),
    .B(_06767_));
 sg13g2_nand2_1 _15067_ (.Y(_06769_),
    .A(_06694_),
    .B(_06685_));
 sg13g2_nand3_1 _15068_ (.B(_06705_),
    .C(_06769_),
    .A(_06674_),
    .Y(_06770_));
 sg13g2_a21oi_1 _15069_ (.A1(_06694_),
    .A2(_06705_),
    .Y(_06771_),
    .B1(_06686_));
 sg13g2_nor2_1 _15070_ (.A(_06694_),
    .B(_06705_),
    .Y(_06772_));
 sg13g2_o21ai_1 _15071_ (.B1(_06610_),
    .Y(_06773_),
    .A1(_06771_),
    .A2(_06772_));
 sg13g2_or2_1 _15072_ (.X(_06774_),
    .B(_06685_),
    .A(_06694_));
 sg13g2_nand3_1 _15073_ (.B(_06773_),
    .C(_06774_),
    .A(_06770_),
    .Y(_06775_));
 sg13g2_o21ai_1 _15074_ (.B1(_06690_),
    .Y(_06776_),
    .A1(net1325),
    .A2(_06691_));
 sg13g2_nand3_1 _15075_ (.B(net215),
    .C(_06776_),
    .A(_04950_),
    .Y(_06777_));
 sg13g2_nor2_1 _15076_ (.A(_06691_),
    .B(_06690_),
    .Y(_06778_));
 sg13g2_a21oi_1 _15077_ (.A1(net1325),
    .A2(_06691_),
    .Y(_06779_),
    .B1(_06778_));
 sg13g2_nand2_1 _15078_ (.Y(_06780_),
    .A(_06777_),
    .B(_06779_));
 sg13g2_a22oi_1 _15079_ (.Y(_06781_),
    .B1(net1323),
    .B2(net1331),
    .A2(net136),
    .A1(net1434));
 sg13g2_xnor2_1 _15080_ (.Y(_06782_),
    .A(net1328),
    .B(_06781_));
 sg13g2_a22oi_1 _15081_ (.Y(_06783_),
    .B1(net91),
    .B2(net247),
    .A2(net1259),
    .A1(net1436));
 sg13g2_nor2_1 _15082_ (.A(net249),
    .B(net1257),
    .Y(_06784_));
 sg13g2_xnor2_1 _15083_ (.Y(_06785_),
    .A(_06783_),
    .B(_06784_));
 sg13g2_xnor2_1 _15084_ (.Y(_06786_),
    .A(_06782_),
    .B(_06785_));
 sg13g2_a22oi_1 _15085_ (.Y(_06787_),
    .B1(net213),
    .B2(net1334),
    .A2(net244),
    .A1(net137));
 sg13g2_xnor2_1 _15086_ (.Y(_06788_),
    .A(net1374),
    .B(_06787_));
 sg13g2_or2_1 _15087_ (.X(_06789_),
    .B(_06704_),
    .A(_06702_));
 sg13g2_nand3_1 _15088_ (.B(_06702_),
    .C(_06704_),
    .A(_06674_),
    .Y(_06790_));
 sg13g2_o21ai_1 _15089_ (.B1(_06790_),
    .Y(_06791_),
    .A1(_06674_),
    .A2(_06789_));
 sg13g2_xnor2_1 _15090_ (.Y(_06792_),
    .A(_06788_),
    .B(_06791_));
 sg13g2_xnor2_1 _15091_ (.Y(_06793_),
    .A(_06786_),
    .B(_06792_));
 sg13g2_xnor2_1 _15092_ (.Y(_06794_),
    .A(_06780_),
    .B(_06793_));
 sg13g2_xnor2_1 _15093_ (.Y(_06795_),
    .A(_06775_),
    .B(_06794_));
 sg13g2_xor2_1 _15094_ (.B(_06795_),
    .A(_06768_),
    .X(_06796_));
 sg13g2_xor2_1 _15095_ (.B(_06796_),
    .A(net1080),
    .X(_06797_));
 sg13g2_xnor2_1 _15096_ (.Y(_06798_),
    .A(net1369),
    .B(_06797_));
 sg13g2_xnor2_1 _15097_ (.Y(_06799_),
    .A(_06759_),
    .B(_06798_));
 sg13g2_xnor2_1 _15098_ (.Y(_06800_),
    .A(_06757_),
    .B(_06799_));
 sg13g2_nor2_1 _15099_ (.A(net1538),
    .B(_05012_),
    .Y(_06801_));
 sg13g2_a21oi_2 _15100_ (.B1(_06801_),
    .Y(_06802_),
    .A2(_06800_),
    .A1(net1538));
 sg13g2_nor2_1 _15101_ (.A(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .B(net1007),
    .Y(_06803_));
 sg13g2_a21oi_1 _15102_ (.A1(_03182_),
    .A2(net1007),
    .Y(_06804_),
    .B1(_06803_));
 sg13g2_a21oi_1 _15103_ (.A1(_05016_),
    .A2(_05632_),
    .Y(_06805_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_26_ ));
 sg13g2_nand2_1 _15104_ (.Y(_06806_),
    .A(net313),
    .B(_06805_));
 sg13g2_o21ai_1 _15105_ (.B1(_06806_),
    .Y(_06807_),
    .A1(net308),
    .A2(_06804_));
 sg13g2_nor3_1 _15106_ (.A(net1708),
    .B(net342),
    .C(_06807_),
    .Y(_06808_));
 sg13g2_nor2_1 _15107_ (.A(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .B(net1260),
    .Y(_06809_));
 sg13g2_a21oi_1 _15108_ (.A1(_03182_),
    .A2(net1260),
    .Y(_06810_),
    .B1(_06809_));
 sg13g2_o21ai_1 _15109_ (.B1(net1634),
    .Y(_06811_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ),
    .A2(net304));
 sg13g2_nand2_1 _15110_ (.Y(_06812_),
    .A(net1571),
    .B(_06811_));
 sg13g2_a221oi_1 _15111_ (.B2(net420),
    .C1(_06812_),
    .B1(_06810_),
    .A1(net1882),
    .Y(_06813_),
    .A2(_06742_));
 sg13g2_o21ai_1 _15112_ (.B1(net1187),
    .Y(_06814_),
    .A1(net339),
    .A2(_06813_));
 sg13g2_or2_1 _15113_ (.X(_06815_),
    .B(net1181),
    .A(\ex_block_i.alu_i.imd_val_q_i_58_ ));
 sg13g2_o21ai_1 _15114_ (.B1(_06815_),
    .Y(_06816_),
    .A1(_06808_),
    .A2(_06814_));
 sg13g2_o21ai_1 _15115_ (.B1(_06816_),
    .Y(_00149_),
    .A1(_06489_),
    .A2(_06802_));
 sg13g2_nor2_1 _15116_ (.A(net375),
    .B(net94),
    .Y(_06817_));
 sg13g2_a21oi_1 _15117_ (.A1(\ex_block_i.alu_i.imd_val_q_i_59_ ),
    .A2(net95),
    .Y(_06818_),
    .B1(_06817_));
 sg13g2_nand2_1 _15118_ (.Y(_06819_),
    .A(\ex_block_i.alu_i.imd_val_q_i_59_ ),
    .B(net319));
 sg13g2_a21oi_2 _15119_ (.B1(net1565),
    .Y(_06820_),
    .A2(_06819_),
    .A1(net1567));
 sg13g2_inv_1 _15120_ (.Y(_06821_),
    .A(_06820_));
 sg13g2_nand2b_1 _15121_ (.Y(_06822_),
    .B(_06788_),
    .A_N(_06786_));
 sg13g2_nand2b_1 _15122_ (.Y(_06823_),
    .B(_06786_),
    .A_N(_06788_));
 sg13g2_o21ai_1 _15123_ (.B1(_06823_),
    .Y(_06824_),
    .A1(_06674_),
    .A2(_06704_));
 sg13g2_a21oi_1 _15124_ (.A1(_06822_),
    .A2(_06824_),
    .Y(_06825_),
    .B1(_06702_));
 sg13g2_nand2_1 _15125_ (.Y(_06826_),
    .A(_06674_),
    .B(_06704_));
 sg13g2_nand2_1 _15126_ (.Y(_06827_),
    .A(_06786_),
    .B(_06826_));
 sg13g2_nand3b_1 _15127_ (.B(_06827_),
    .C(_06702_),
    .Y(_06828_),
    .A_N(_06788_));
 sg13g2_o21ai_1 _15128_ (.B1(_06828_),
    .Y(_06829_),
    .A1(_06786_),
    .A2(_06826_));
 sg13g2_or2_1 _15129_ (.X(_06830_),
    .B(_06829_),
    .A(_06825_));
 sg13g2_a22oi_1 _15130_ (.Y(_06831_),
    .B1(net90),
    .B2(net1436),
    .A2(net1259),
    .A1(net1434));
 sg13g2_xnor2_1 _15131_ (.Y(_06832_),
    .A(net1320),
    .B(_06831_));
 sg13g2_a22oi_1 _15132_ (.Y(_06833_),
    .B1(net243),
    .B2(net1331),
    .A2(net1323),
    .A1(net134));
 sg13g2_xnor2_1 _15133_ (.Y(_06834_),
    .A(net1330),
    .B(_06833_));
 sg13g2_o21ai_1 _15134_ (.B1(net216),
    .Y(_06835_),
    .A1(_05197_),
    .A2(net1324));
 sg13g2_xnor2_1 _15135_ (.Y(_06836_),
    .A(_06834_),
    .B(_06835_));
 sg13g2_xnor2_1 _15136_ (.Y(_06837_),
    .A(_06832_),
    .B(_06836_));
 sg13g2_o21ai_1 _15137_ (.B1(net214),
    .Y(_06838_),
    .A1(net1334),
    .A2(net137));
 sg13g2_xnor2_1 _15138_ (.Y(_06839_),
    .A(_05043_),
    .B(_06838_));
 sg13g2_nand3_1 _15139_ (.B(_06788_),
    .C(_06839_),
    .A(_06702_),
    .Y(_06840_));
 sg13g2_a21o_1 _15140_ (.A2(_06788_),
    .A1(_06702_),
    .B1(_06839_),
    .X(_06841_));
 sg13g2_nand2_1 _15141_ (.Y(_06842_),
    .A(_06840_),
    .B(_06841_));
 sg13g2_xor2_1 _15142_ (.B(_06842_),
    .A(_06837_),
    .X(_06843_));
 sg13g2_o21ai_1 _15143_ (.B1(_06782_),
    .Y(_06844_),
    .A1(net1324),
    .A2(_06783_));
 sg13g2_nand3b_1 _15144_ (.B(net216),
    .C(_06844_),
    .Y(_06845_),
    .A_N(net248));
 sg13g2_nor2_1 _15145_ (.A(_06783_),
    .B(_06782_),
    .Y(_06846_));
 sg13g2_a21oi_1 _15146_ (.A1(net1324),
    .A2(_06783_),
    .Y(_06847_),
    .B1(_06846_));
 sg13g2_nand2_1 _15147_ (.Y(_06848_),
    .A(_06845_),
    .B(_06847_));
 sg13g2_inv_1 _15148_ (.Y(_06849_),
    .A(_06848_));
 sg13g2_xnor2_1 _15149_ (.Y(_06850_),
    .A(_06843_),
    .B(_06849_));
 sg13g2_xnor2_1 _15150_ (.Y(_06851_),
    .A(_06830_),
    .B(_06850_));
 sg13g2_nand2b_1 _15151_ (.Y(_06852_),
    .B(_06780_),
    .A_N(_06793_));
 sg13g2_nor2b_1 _15152_ (.A(_06780_),
    .B_N(_06793_),
    .Y(_06853_));
 sg13g2_a21oi_2 _15153_ (.B1(_06853_),
    .Y(_06854_),
    .A2(_06852_),
    .A1(_06775_));
 sg13g2_xor2_1 _15154_ (.B(_06854_),
    .A(_06851_),
    .X(_06855_));
 sg13g2_or2_2 _15155_ (.X(_06856_),
    .B(_06795_),
    .A(_06768_));
 sg13g2_xor2_1 _15156_ (.B(_06856_),
    .A(_06855_),
    .X(_06857_));
 sg13g2_xnor2_1 _15157_ (.Y(_06858_),
    .A(_06821_),
    .B(_06857_));
 sg13g2_inv_1 _15158_ (.Y(_06859_),
    .A(net1369));
 sg13g2_inv_1 _15159_ (.Y(_06860_),
    .A(_06796_));
 sg13g2_nor2_2 _15160_ (.A(net1080),
    .B(_06860_),
    .Y(_06861_));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(\register_file_i/_2911_ ));
 sg13g2_inv_1 _15162_ (.Y(_06863_),
    .A(_06861_));
 sg13g2_nand2_2 _15163_ (.Y(_06864_),
    .A(net1080),
    .B(_06860_));
 sg13g2_inv_1 _15164_ (.Y(_06865_),
    .A(_06864_));
 sg13g2_a21oi_1 _15165_ (.A1(_06859_),
    .A2(_06863_),
    .Y(_06866_),
    .B1(_06865_));
 sg13g2_or2_1 _15166_ (.X(_06867_),
    .B(_06866_),
    .A(_06759_));
 sg13g2_nand2_1 _15167_ (.Y(_06868_),
    .A(_06859_),
    .B(_06865_));
 sg13g2_nand3_1 _15168_ (.B(net1370),
    .C(net1062),
    .A(_06759_),
    .Y(_06869_));
 sg13g2_nand3_1 _15169_ (.B(_06868_),
    .C(_06869_),
    .A(_06867_),
    .Y(_06870_));
 sg13g2_inv_1 _15170_ (.Y(_06871_),
    .A(_06756_));
 sg13g2_nor3_1 _15171_ (.A(_06649_),
    .B(_06667_),
    .C(_06871_),
    .Y(_06872_));
 sg13g2_or2_1 _15172_ (.X(_06873_),
    .B(_06872_),
    .A(_06755_));
 sg13g2_a21oi_1 _15173_ (.A1(net1369),
    .A2(_06864_),
    .Y(_06874_),
    .B1(net1062));
 sg13g2_and2_1 _15174_ (.A(_06758_),
    .B(net808),
    .X(_06875_));
 sg13g2_nor3_1 _15175_ (.A(net1076),
    .B(_06874_),
    .C(_06875_),
    .Y(_06876_));
 sg13g2_a21oi_1 _15176_ (.A1(net1369),
    .A2(net1062),
    .Y(_06877_),
    .B1(_06876_));
 sg13g2_o21ai_1 _15177_ (.B1(_06877_),
    .Y(_06878_),
    .A1(_06759_),
    .A2(_06868_));
 sg13g2_a22oi_1 _15178_ (.Y(_06879_),
    .B1(_06878_),
    .B2(_06757_),
    .A2(_06873_),
    .A1(_06870_));
 sg13g2_xnor2_1 _15179_ (.Y(_06880_),
    .A(_06858_),
    .B(_06879_));
 sg13g2_a21oi_1 _15180_ (.A1(_05016_),
    .A2(_05892_),
    .Y(_06881_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_27_ ));
 sg13g2_mux2_1 _15181_ (.A0(\ex_block_i.alu_i.imd_val_q_i_59_ ),
    .A1(data_addr_o_27_),
    .S(net1007),
    .X(_06882_));
 sg13g2_nor2_1 _15182_ (.A(net307),
    .B(_06882_),
    .Y(_06883_));
 sg13g2_a21oi_1 _15183_ (.A1(net314),
    .A2(_06881_),
    .Y(_06884_),
    .B1(_06883_));
 sg13g2_o21ai_1 _15184_ (.B1(net1635),
    .Y(_06885_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ),
    .A2(net311));
 sg13g2_nor2_1 _15185_ (.A(net2487),
    .B(net1218),
    .Y(_06886_));
 sg13g2_a21oi_1 _15186_ (.A1(_01899_),
    .A2(net1218),
    .Y(_06887_),
    .B1(_06886_));
 sg13g2_nand2_1 _15187_ (.Y(_06888_),
    .A(net422),
    .B(_06887_));
 sg13g2_nand3_1 _15188_ (.B(_06885_),
    .C(_06888_),
    .A(net1181),
    .Y(_06889_));
 sg13g2_a221oi_1 _15189_ (.B2(net1888),
    .C1(_06889_),
    .B1(_06884_),
    .A1(net1883),
    .Y(_06890_),
    .A2(_06804_));
 sg13g2_a221oi_1 _15190_ (.B2(_01899_),
    .C1(_06890_),
    .B1(net1478),
    .A1(net342),
    .Y(_06891_),
    .A2(net1188));
 sg13g2_a221oi_1 _15191_ (.B2(_04144_),
    .C1(_06891_),
    .B1(_06880_),
    .A1(_05128_),
    .Y(_06892_),
    .A2(_06740_));
 sg13g2_nor2_2 _15192_ (.A(_06818_),
    .B(_06892_),
    .Y(_00150_));
 sg13g2_mux2_1 _15193_ (.A0(net1511),
    .A1(data_addr_o_5_),
    .S(net1451),
    .X(_06893_));
 sg13g2_mux2_1 _15194_ (.A0(_06893_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_5_ ),
    .S(net1225),
    .X(_00151_));
 sg13g2_inv_2 _15195_ (.Y(_06894_),
    .A(\ex_block_i.alu_i.imd_val_q_i_60_ ));
 sg13g2_nand2_1 _15196_ (.Y(_06895_),
    .A(net299),
    .B(_05262_));
 sg13g2_nor2b_1 _15197_ (.A(net1076),
    .B_N(_06797_),
    .Y(_06896_));
 sg13g2_nor3_1 _15198_ (.A(_06716_),
    .B(_06722_),
    .C(net1062),
    .Y(_06897_));
 sg13g2_or2_1 _15199_ (.X(_06898_),
    .B(_06897_),
    .A(_06896_));
 sg13g2_inv_1 _15200_ (.Y(_06899_),
    .A(_06898_));
 sg13g2_nor2_1 _15201_ (.A(net1076),
    .B(net1369),
    .Y(_06900_));
 sg13g2_a22oi_1 _15202_ (.Y(_06901_),
    .B1(_06900_),
    .B2(net1062),
    .A2(_06899_),
    .A1(net1369));
 sg13g2_or3_1 _15203_ (.A(_06723_),
    .B(net1369),
    .C(_06797_),
    .X(_06902_));
 sg13g2_o21ai_1 _15204_ (.B1(_06902_),
    .Y(_06903_),
    .A1(_06859_),
    .A2(_06864_));
 sg13g2_a221oi_1 _15205_ (.B2(net1076),
    .C1(_06858_),
    .B1(_06903_),
    .A1(_06865_),
    .Y(_06904_),
    .A2(_06900_));
 sg13g2_a21o_1 _15206_ (.A2(_06901_),
    .A1(_06858_),
    .B1(_06904_),
    .X(_06905_));
 sg13g2_a21o_1 _15207_ (.A2(_06726_),
    .A1(_06670_),
    .B1(_06905_),
    .X(_06906_));
 sg13g2_xnor2_1 _15208_ (.Y(_06907_),
    .A(_06859_),
    .B(_06796_));
 sg13g2_and2_1 _15209_ (.A(_06758_),
    .B(net1080),
    .X(_06908_));
 sg13g2_nor2_1 _15210_ (.A(_06758_),
    .B(net1080),
    .Y(_06909_));
 sg13g2_mux2_1 _15211_ (.A0(_06908_),
    .A1(_06909_),
    .S(_06858_),
    .X(_06910_));
 sg13g2_nor2_1 _15212_ (.A(_06908_),
    .B(_06909_),
    .Y(_06911_));
 sg13g2_nor3_1 _15213_ (.A(net1370),
    .B(_06796_),
    .C(_06858_),
    .Y(_06912_));
 sg13g2_nand3_1 _15214_ (.B(_06796_),
    .C(_06858_),
    .A(net1370),
    .Y(_06913_));
 sg13g2_nand2b_1 _15215_ (.Y(_06914_),
    .B(_06913_),
    .A_N(_06912_));
 sg13g2_a22oi_1 _15216_ (.Y(_06915_),
    .B1(_06911_),
    .B2(_06914_),
    .A2(_06910_),
    .A1(_06907_));
 sg13g2_o21ai_1 _15217_ (.B1(_06670_),
    .Y(_06916_),
    .A1(_06723_),
    .A2(net1076));
 sg13g2_nand2b_1 _15218_ (.Y(_06917_),
    .B(_06916_),
    .A_N(_06915_));
 sg13g2_mux2_1 _15219_ (.A0(_06906_),
    .A1(_06917_),
    .S(net808),
    .X(_06918_));
 sg13g2_nor2_1 _15220_ (.A(_06668_),
    .B(_06918_),
    .Y(_06919_));
 sg13g2_nor2b_1 _15221_ (.A(_06915_),
    .B_N(_06726_),
    .Y(_06920_));
 sg13g2_nor3_1 _15222_ (.A(_06726_),
    .B(net808),
    .C(_06905_),
    .Y(_06921_));
 sg13g2_a21oi_1 _15223_ (.A1(net808),
    .A2(_06920_),
    .Y(_06922_),
    .B1(_06921_));
 sg13g2_o21ai_1 _15224_ (.B1(net1369),
    .Y(_06923_),
    .A1(_06759_),
    .A2(_06864_));
 sg13g2_nand2_1 _15225_ (.Y(_06924_),
    .A(net1370),
    .B(_06820_));
 sg13g2_o21ai_1 _15226_ (.B1(_06857_),
    .Y(_06925_),
    .A1(_06865_),
    .A2(_06924_));
 sg13g2_nor2b_1 _15227_ (.A(_06861_),
    .B_N(_06724_),
    .Y(_06926_));
 sg13g2_o21ai_1 _15228_ (.B1(_06857_),
    .Y(_06927_),
    .A1(_06724_),
    .A2(_06924_));
 sg13g2_and2_1 _15229_ (.A(_06820_),
    .B(_06857_),
    .X(_06928_));
 sg13g2_nand2b_1 _15230_ (.Y(_06929_),
    .B(_06924_),
    .A_N(_06857_));
 sg13g2_a22oi_1 _15231_ (.Y(_06930_),
    .B1(_06861_),
    .B2(_06929_),
    .A2(_06864_),
    .A1(_06928_));
 sg13g2_nand2_1 _15232_ (.Y(_06931_),
    .A(_06928_),
    .B(net1062));
 sg13g2_o21ai_1 _15233_ (.B1(_06931_),
    .Y(_06932_),
    .A1(_06724_),
    .A2(_06930_));
 sg13g2_a221oi_1 _15234_ (.B2(_06865_),
    .C1(_06932_),
    .B1(_06927_),
    .A1(_06925_),
    .Y(_06933_),
    .A2(_06926_));
 sg13g2_nand2_1 _15235_ (.Y(_06934_),
    .A(_06820_),
    .B(_06866_));
 sg13g2_mux2_1 _15236_ (.A0(net1062),
    .A1(_06934_),
    .S(_06857_),
    .X(_06935_));
 sg13g2_mux2_1 _15237_ (.A0(_06933_),
    .A1(_06935_),
    .S(_06875_),
    .X(_06936_));
 sg13g2_a21o_1 _15238_ (.A2(_06923_),
    .A1(_06821_),
    .B1(_06936_),
    .X(_06937_));
 sg13g2_o21ai_1 _15239_ (.B1(_06937_),
    .Y(_06938_),
    .A1(_06670_),
    .A2(_06922_));
 sg13g2_or2_1 _15240_ (.X(_06939_),
    .B(_06938_),
    .A(_06919_));
 sg13g2_nand2_1 _15241_ (.Y(_06940_),
    .A(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .B(net321));
 sg13g2_a21o_1 _15242_ (.A2(_06940_),
    .A1(net1567),
    .B1(net1565),
    .X(_06941_));
 sg13g2_inv_1 _15243_ (.Y(_06942_),
    .A(_06830_));
 sg13g2_o21ai_1 _15244_ (.B1(_06843_),
    .Y(_06943_),
    .A1(_06942_),
    .A2(_06848_));
 sg13g2_o21ai_1 _15245_ (.B1(_06943_),
    .Y(_06944_),
    .A1(_06830_),
    .A2(_06849_));
 sg13g2_o21ai_1 _15246_ (.B1(_06835_),
    .Y(_06945_),
    .A1(_06832_),
    .A2(_06834_));
 sg13g2_nand2_1 _15247_ (.Y(_06946_),
    .A(_06832_),
    .B(_06834_));
 sg13g2_nand2_1 _15248_ (.Y(_06947_),
    .A(_06945_),
    .B(_06946_));
 sg13g2_nor2_1 _15249_ (.A(_06702_),
    .B(_06839_),
    .Y(_06948_));
 sg13g2_inv_1 _15250_ (.Y(_06949_),
    .A(_06948_));
 sg13g2_a22oi_1 _15251_ (.Y(_06950_),
    .B1(net213),
    .B2(net1331),
    .A2(net244),
    .A1(net134));
 sg13g2_xnor2_1 _15252_ (.Y(_06951_),
    .A(net1330),
    .B(_06950_));
 sg13g2_a22oi_1 _15253_ (.Y(_06952_),
    .B1(net90),
    .B2(net1434),
    .A2(net1259),
    .A1(net1323));
 sg13g2_xnor2_1 _15254_ (.Y(_06953_),
    .A(net1320),
    .B(_06952_));
 sg13g2_o21ai_1 _15255_ (.B1(net216),
    .Y(_06954_),
    .A1(_05306_),
    .A2(net1324));
 sg13g2_xnor2_1 _15256_ (.Y(_06955_),
    .A(_06953_),
    .B(_06954_));
 sg13g2_xnor2_1 _15257_ (.Y(_06956_),
    .A(_06951_),
    .B(_06955_));
 sg13g2_xnor2_1 _15258_ (.Y(_06957_),
    .A(_06949_),
    .B(_06956_));
 sg13g2_o21ai_1 _15259_ (.B1(_06837_),
    .Y(_06958_),
    .A1(_06788_),
    .A2(_06839_));
 sg13g2_nand3_1 _15260_ (.B(_06949_),
    .C(_06958_),
    .A(_06840_),
    .Y(_06959_));
 sg13g2_xor2_1 _15261_ (.B(_06959_),
    .A(_06957_),
    .X(_06960_));
 sg13g2_xnor2_1 _15262_ (.Y(_06961_),
    .A(_06947_),
    .B(_06960_));
 sg13g2_xor2_1 _15263_ (.B(_06961_),
    .A(_06944_),
    .X(_06962_));
 sg13g2_nor2_1 _15264_ (.A(_06851_),
    .B(_06854_),
    .Y(_06963_));
 sg13g2_xnor2_1 _15265_ (.Y(_06964_),
    .A(_06962_),
    .B(_06963_));
 sg13g2_nor2_1 _15266_ (.A(_06716_),
    .B(_06722_),
    .Y(_06965_));
 sg13g2_nand2_1 _15267_ (.Y(_06966_),
    .A(net1080),
    .B(_06768_));
 sg13g2_nor2_1 _15268_ (.A(net1080),
    .B(_06768_),
    .Y(_06967_));
 sg13g2_nor2_1 _15269_ (.A(_06855_),
    .B(_06967_),
    .Y(_06968_));
 sg13g2_nor2_1 _15270_ (.A(_06795_),
    .B(_06968_),
    .Y(_06969_));
 sg13g2_a21oi_1 _15271_ (.A1(_06855_),
    .A2(_06966_),
    .Y(_06970_),
    .B1(_06969_));
 sg13g2_a21oi_1 _15272_ (.A1(net1080),
    .A2(_06768_),
    .Y(_06971_),
    .B1(_06795_));
 sg13g2_o21ai_1 _15273_ (.B1(_06855_),
    .Y(_06972_),
    .A1(_06967_),
    .A2(_06971_));
 sg13g2_o21ai_1 _15274_ (.B1(_06972_),
    .Y(_06973_),
    .A1(_06965_),
    .A2(_06970_));
 sg13g2_nor2b_1 _15275_ (.A(_06855_),
    .B_N(_06856_),
    .Y(_06974_));
 sg13g2_nand2_1 _15276_ (.Y(_06975_),
    .A(_06768_),
    .B(_06795_));
 sg13g2_nand2_1 _15277_ (.Y(_06976_),
    .A(_06855_),
    .B(_06975_));
 sg13g2_o21ai_1 _15278_ (.B1(_06976_),
    .Y(_06977_),
    .A1(_06765_),
    .A2(_06974_));
 sg13g2_inv_1 _15279_ (.Y(_06978_),
    .A(_06975_));
 sg13g2_o21ai_1 _15280_ (.B1(_06856_),
    .Y(_06979_),
    .A1(_06765_),
    .A2(_06978_));
 sg13g2_a22oi_1 _15281_ (.Y(_06980_),
    .B1(_06979_),
    .B2(_06855_),
    .A2(_06977_),
    .A1(_06723_));
 sg13g2_nand2_1 _15282_ (.Y(_06981_),
    .A(_06734_),
    .B(_06980_));
 sg13g2_o21ai_1 _15283_ (.B1(_06981_),
    .Y(_06982_),
    .A1(net808),
    .A2(_06973_));
 sg13g2_xor2_1 _15284_ (.B(_06982_),
    .A(_06964_),
    .X(_06983_));
 sg13g2_xnor2_1 _15285_ (.Y(_06984_),
    .A(_06941_),
    .B(_06983_));
 sg13g2_xor2_1 _15286_ (.B(_06984_),
    .A(_06939_),
    .X(_06985_));
 sg13g2_nand2_1 _15287_ (.Y(_06986_),
    .A(net1540),
    .B(_06985_));
 sg13g2_nand3_1 _15288_ (.B(_06895_),
    .C(_06986_),
    .A(net1182),
    .Y(_06987_));
 sg13g2_a21oi_1 _15289_ (.A1(_04761_),
    .A2(_06245_),
    .Y(_06988_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_28_ ));
 sg13g2_nand2_1 _15290_ (.Y(_06989_),
    .A(data_addr_o_28_),
    .B(net1007));
 sg13g2_o21ai_1 _15291_ (.B1(_06989_),
    .Y(_06990_),
    .A1(_06894_),
    .A2(net1007));
 sg13g2_nor2_1 _15292_ (.A(net311),
    .B(_06990_),
    .Y(_06991_));
 sg13g2_a21oi_1 _15293_ (.A1(net315),
    .A2(_06988_),
    .Y(_06992_),
    .B1(_06991_));
 sg13g2_o21ai_1 _15294_ (.B1(net1634),
    .Y(_06993_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_28_ ),
    .A2(net311));
 sg13g2_nand2_1 _15295_ (.Y(_06994_),
    .A(data_addr_o_28_),
    .B(net1260));
 sg13g2_o21ai_1 _15296_ (.B1(_06994_),
    .Y(_06995_),
    .A1(_06894_),
    .A2(net1260));
 sg13g2_nand2_1 _15297_ (.Y(_06996_),
    .A(net422),
    .B(_06995_));
 sg13g2_nand3_1 _15298_ (.B(_06993_),
    .C(_06996_),
    .A(net1571),
    .Y(_06997_));
 sg13g2_a221oi_1 _15299_ (.B2(net1888),
    .C1(_06997_),
    .B1(_06992_),
    .A1(net1882),
    .Y(_06998_),
    .A2(_06882_));
 sg13g2_o21ai_1 _15300_ (.B1(net1185),
    .Y(_06999_),
    .A1(net339),
    .A2(_06998_));
 sg13g2_o21ai_1 _15301_ (.B1(_06999_),
    .Y(_07000_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .A2(net1571));
 sg13g2_a22oi_1 _15302_ (.Y(_00152_),
    .B1(_06987_),
    .B2(_07000_),
    .A2(net95),
    .A1(_06894_));
 sg13g2_inv_1 _15303_ (.Y(_07001_),
    .A(\ex_block_i.alu_i.imd_val_q_i_61_ ));
 sg13g2_nor2_2 _15304_ (.A(net2093),
    .B(_04029_),
    .Y(_07002_));
 sg13g2_nand2_2 _15305_ (.Y(_07003_),
    .A(net341),
    .B(_07002_));
 sg13g2_nor2_1 _15306_ (.A(_06941_),
    .B(_06983_),
    .Y(_07004_));
 sg13g2_nand2_1 _15307_ (.Y(_07005_),
    .A(_06941_),
    .B(_06983_));
 sg13g2_o21ai_1 _15308_ (.B1(_07005_),
    .Y(_07006_),
    .A1(_06939_),
    .A2(_07004_));
 sg13g2_nand2_1 _15309_ (.Y(_07007_),
    .A(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .B(net321));
 sg13g2_a21oi_1 _15310_ (.A1(net1567),
    .A2(_07007_),
    .Y(_07008_),
    .B1(net1565));
 sg13g2_o21ai_1 _15311_ (.B1(_06834_),
    .Y(_07009_),
    .A1(_06832_),
    .A2(_06835_));
 sg13g2_nand2_1 _15312_ (.Y(_07010_),
    .A(_06832_),
    .B(_06835_));
 sg13g2_nand2_1 _15313_ (.Y(_07011_),
    .A(_07009_),
    .B(_07010_));
 sg13g2_xor2_1 _15314_ (.B(_07011_),
    .A(_06960_),
    .X(_07012_));
 sg13g2_nor2_2 _15315_ (.A(_06944_),
    .B(_07012_),
    .Y(_07013_));
 sg13g2_inv_1 _15316_ (.Y(_07014_),
    .A(_06959_));
 sg13g2_inv_1 _15317_ (.Y(_07015_),
    .A(_06957_));
 sg13g2_o21ai_1 _15318_ (.B1(_06947_),
    .Y(_07016_),
    .A1(_07015_),
    .A2(_06959_));
 sg13g2_o21ai_1 _15319_ (.B1(_07016_),
    .Y(_07017_),
    .A1(_06957_),
    .A2(_07014_));
 sg13g2_and2_2 _15320_ (.A(_06949_),
    .B(_06956_),
    .X(_07018_));
 sg13g2_inv_1 _15321_ (.Y(_07019_),
    .A(_07018_));
 sg13g2_o21ai_1 _15322_ (.B1(_06951_),
    .Y(_07020_),
    .A1(_06953_),
    .A2(_06954_));
 sg13g2_inv_1 _15323_ (.Y(_07021_),
    .A(_07020_));
 sg13g2_a21oi_2 _15324_ (.B1(_07021_),
    .Y(_07022_),
    .A2(_06954_),
    .A1(_06953_));
 sg13g2_o21ai_1 _15325_ (.B1(net214),
    .Y(_07023_),
    .A1(net1331),
    .A2(net134));
 sg13g2_xor2_1 _15326_ (.B(_07023_),
    .A(net1330),
    .X(_07024_));
 sg13g2_a22oi_1 _15327_ (.Y(_07025_),
    .B1(net90),
    .B2(net1323),
    .A2(net1259),
    .A1(net242));
 sg13g2_xnor2_1 _15328_ (.Y(_07026_),
    .A(net1320),
    .B(_07025_));
 sg13g2_a21oi_1 _15329_ (.A1(net1434),
    .A2(net1320),
    .Y(_07027_),
    .B1(net1372));
 sg13g2_inv_1 _15330_ (.Y(_07028_),
    .A(_07027_));
 sg13g2_xnor2_1 _15331_ (.Y(_07029_),
    .A(_07026_),
    .B(_07028_));
 sg13g2_xnor2_1 _15332_ (.Y(_07030_),
    .A(_07024_),
    .B(_07029_));
 sg13g2_inv_1 _15333_ (.Y(_07031_),
    .A(_07030_));
 sg13g2_xnor2_1 _15334_ (.Y(_07032_),
    .A(_07022_),
    .B(_07031_));
 sg13g2_xnor2_1 _15335_ (.Y(_07033_),
    .A(_07019_),
    .B(_07032_));
 sg13g2_xnor2_1 _15336_ (.Y(_07034_),
    .A(_07017_),
    .B(_07033_));
 sg13g2_xnor2_1 _15337_ (.Y(_07035_),
    .A(_07013_),
    .B(_07034_));
 sg13g2_a21o_1 _15338_ (.A2(_06856_),
    .A1(_06851_),
    .B1(_06854_),
    .X(_07036_));
 sg13g2_o21ai_1 _15339_ (.B1(_07036_),
    .Y(_07037_),
    .A1(_06851_),
    .A2(_06856_));
 sg13g2_nand2b_1 _15340_ (.Y(_07038_),
    .B(_07037_),
    .A_N(_06962_));
 sg13g2_inv_1 _15341_ (.Y(_07039_),
    .A(_07038_));
 sg13g2_nand2b_1 _15342_ (.Y(_07040_),
    .B(_06864_),
    .A_N(net1076));
 sg13g2_nor2_1 _15343_ (.A(_06723_),
    .B(net1062),
    .Y(_07041_));
 sg13g2_nand2b_1 _15344_ (.Y(_07042_),
    .B(_06964_),
    .A_N(_06857_));
 sg13g2_a221oi_1 _15345_ (.B2(net808),
    .C1(_07042_),
    .B1(_07041_),
    .A1(_06863_),
    .Y(_07043_),
    .A2(_07040_));
 sg13g2_or2_1 _15346_ (.X(_07044_),
    .B(_07043_),
    .A(_07039_));
 sg13g2_xor2_1 _15347_ (.B(_07044_),
    .A(_07035_),
    .X(_07045_));
 sg13g2_xnor2_1 _15348_ (.Y(_07046_),
    .A(_07008_),
    .B(_07045_));
 sg13g2_xnor2_1 _15349_ (.Y(_07047_),
    .A(_07006_),
    .B(_07046_));
 sg13g2_nand2_1 _15350_ (.Y(_07048_),
    .A(net299),
    .B(_05356_));
 sg13g2_o21ai_1 _15351_ (.B1(_07048_),
    .Y(_07049_),
    .A1(net297),
    .A2(_07047_));
 sg13g2_nor2_2 _15352_ (.A(_07003_),
    .B(_07049_),
    .Y(_07050_));
 sg13g2_o21ai_1 _15353_ (.B1(net1185),
    .Y(_07051_),
    .A1(net1571),
    .A2(_07050_));
 sg13g2_a21oi_1 _15354_ (.A1(_04761_),
    .A2(_06346_),
    .Y(_07052_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_29_ ));
 sg13g2_mux2_1 _15355_ (.A0(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .A1(data_addr_o_29_),
    .S(net1007),
    .X(_07053_));
 sg13g2_nor2_1 _15356_ (.A(net306),
    .B(_07053_),
    .Y(_07054_));
 sg13g2_a21oi_1 _15357_ (.A1(net313),
    .A2(_07052_),
    .Y(_07055_),
    .B1(_07054_));
 sg13g2_nand2_1 _15358_ (.Y(_07056_),
    .A(net1888),
    .B(_07055_));
 sg13g2_nor2_1 _15359_ (.A(data_addr_o_29_),
    .B(net1218),
    .Y(_07057_));
 sg13g2_a21oi_1 _15360_ (.A1(_07001_),
    .A2(net1218),
    .Y(_07058_),
    .B1(_07057_));
 sg13g2_o21ai_1 _15361_ (.B1(net1634),
    .Y(_07059_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ),
    .A2(net309));
 sg13g2_nand2_1 _15362_ (.Y(_07060_),
    .A(net1181),
    .B(_07059_));
 sg13g2_a221oi_1 _15363_ (.B2(net419),
    .C1(_07060_),
    .B1(_07058_),
    .A1(net1882),
    .Y(_07061_),
    .A2(_06990_));
 sg13g2_a22oi_1 _15364_ (.Y(_07062_),
    .B1(_07056_),
    .B2(_07061_),
    .A2(net1185),
    .A1(net337));
 sg13g2_nor2_1 _15365_ (.A(_07050_),
    .B(_07062_),
    .Y(_07063_));
 sg13g2_a21oi_1 _15366_ (.A1(_07001_),
    .A2(_07051_),
    .Y(_00153_),
    .B1(_07063_));
 sg13g2_nand2b_1 _15367_ (.Y(_07064_),
    .B(_07045_),
    .A_N(_07008_));
 sg13g2_o21ai_1 _15368_ (.B1(_06937_),
    .Y(_07065_),
    .A1(_06872_),
    .A2(_06918_));
 sg13g2_nor2b_1 _15369_ (.A(_06984_),
    .B_N(_07046_),
    .Y(_07066_));
 sg13g2_nor2b_1 _15370_ (.A(_07045_),
    .B_N(_07008_),
    .Y(_07067_));
 sg13g2_a221oi_1 _15371_ (.B2(_07066_),
    .C1(_07067_),
    .B1(_07065_),
    .A1(_07004_),
    .Y(_07068_),
    .A2(_07064_));
 sg13g2_nand2_1 _15372_ (.Y(_07069_),
    .A(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .B(net320));
 sg13g2_a21o_1 _15373_ (.A2(_07069_),
    .A1(net1568),
    .B1(net1566),
    .X(_07070_));
 sg13g2_inv_1 _15374_ (.Y(_07071_),
    .A(_07024_));
 sg13g2_inv_1 _15375_ (.Y(_07072_),
    .A(_07026_));
 sg13g2_a21oi_1 _15376_ (.A1(_07024_),
    .A2(_07026_),
    .Y(_07073_),
    .B1(_07028_));
 sg13g2_a21oi_1 _15377_ (.A1(_07071_),
    .A2(_07072_),
    .Y(_07074_),
    .B1(_07073_));
 sg13g2_o21ai_1 _15378_ (.B1(net216),
    .Y(_07075_),
    .A1(_05411_),
    .A2(net1324));
 sg13g2_a22oi_1 _15379_ (.Y(_07076_),
    .B1(net213),
    .B2(net1259),
    .A2(net92),
    .A1(net242));
 sg13g2_xnor2_1 _15380_ (.Y(_07077_),
    .A(net1320),
    .B(_07076_));
 sg13g2_xor2_1 _15381_ (.B(_07077_),
    .A(_07075_),
    .X(_07078_));
 sg13g2_xnor2_1 _15382_ (.Y(_07079_),
    .A(_07074_),
    .B(_07078_));
 sg13g2_nand2_2 _15383_ (.Y(_07080_),
    .A(_07022_),
    .B(_07031_));
 sg13g2_o21ai_1 _15384_ (.B1(_07013_),
    .Y(_07081_),
    .A1(_07018_),
    .A2(_07017_));
 sg13g2_nand2_1 _15385_ (.Y(_07082_),
    .A(_07018_),
    .B(_07017_));
 sg13g2_nand2_1 _15386_ (.Y(_07083_),
    .A(_07081_),
    .B(_07082_));
 sg13g2_nor2_1 _15387_ (.A(_07013_),
    .B(_07017_),
    .Y(_07084_));
 sg13g2_nor2_1 _15388_ (.A(_07018_),
    .B(_07080_),
    .Y(_07085_));
 sg13g2_nand2b_2 _15389_ (.Y(_07086_),
    .B(_07030_),
    .A_N(_07022_));
 sg13g2_a21oi_1 _15390_ (.A1(_07019_),
    .A2(_07084_),
    .Y(_07087_),
    .B1(_07086_));
 sg13g2_a221oi_1 _15391_ (.B2(_07085_),
    .C1(_07087_),
    .B1(_07084_),
    .A1(_07080_),
    .Y(_07088_),
    .A2(_07083_));
 sg13g2_xnor2_1 _15392_ (.Y(_07089_),
    .A(_07079_),
    .B(_07088_));
 sg13g2_nand2b_1 _15393_ (.Y(_07090_),
    .B(_07038_),
    .A_N(_07035_));
 sg13g2_nand2_1 _15394_ (.Y(_07091_),
    .A(_07019_),
    .B(_07086_));
 sg13g2_a21oi_1 _15395_ (.A1(_07080_),
    .A2(_07091_),
    .Y(_07092_),
    .B1(_07017_));
 sg13g2_nor2_1 _15396_ (.A(_07082_),
    .B(_07086_),
    .Y(_07093_));
 sg13g2_nor3_1 _15397_ (.A(_07085_),
    .B(_07092_),
    .C(_07093_),
    .Y(_07094_));
 sg13g2_xnor2_1 _15398_ (.Y(_07095_),
    .A(_07079_),
    .B(_07094_));
 sg13g2_xnor2_1 _15399_ (.Y(_07096_),
    .A(_07043_),
    .B(_07095_));
 sg13g2_nor2_1 _15400_ (.A(_07096_),
    .B(_07090_),
    .Y(_07097_));
 sg13g2_a21oi_2 _15401_ (.B1(_07097_),
    .Y(_07098_),
    .A2(_07090_),
    .A1(_07089_));
 sg13g2_xor2_1 _15402_ (.B(_07098_),
    .A(_07070_),
    .X(_07099_));
 sg13g2_xnor2_1 _15403_ (.Y(_07100_),
    .A(_07068_),
    .B(_07099_));
 sg13g2_nor2_1 _15404_ (.A(net1538),
    .B(_05470_),
    .Y(_07101_));
 sg13g2_a21oi_1 _15405_ (.A1(net1538),
    .A2(_07100_),
    .Y(_07102_),
    .B1(_07101_));
 sg13g2_nand2_2 _15406_ (.Y(_07103_),
    .A(_06016_),
    .B(_07102_));
 sg13g2_mux2_1 _15407_ (.A0(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .A1(data_addr_o_30_),
    .S(net1008),
    .X(_07104_));
 sg13g2_a21oi_1 _15408_ (.A1(_05016_),
    .A2(_06245_),
    .Y(_07105_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_30_ ));
 sg13g2_nand2_1 _15409_ (.Y(_07106_),
    .A(net313),
    .B(_07105_));
 sg13g2_o21ai_1 _15410_ (.B1(_07106_),
    .Y(_07107_),
    .A1(net308),
    .A2(_07104_));
 sg13g2_mux2_1 _15411_ (.A0(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .A1(data_addr_o_30_),
    .S(net1260),
    .X(_07108_));
 sg13g2_o21ai_1 _15412_ (.B1(net1635),
    .Y(_07109_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ),
    .A2(net307));
 sg13g2_nand2_1 _15413_ (.Y(_07110_),
    .A(net1181),
    .B(_07109_));
 sg13g2_a221oi_1 _15414_ (.B2(net419),
    .C1(_07110_),
    .B1(_07108_),
    .A1(net1883),
    .Y(_07111_),
    .A2(_07053_));
 sg13g2_o21ai_1 _15415_ (.B1(_07111_),
    .Y(_07112_),
    .A1(net1708),
    .A2(_07107_));
 sg13g2_o21ai_1 _15416_ (.B1(_07112_),
    .Y(_07113_),
    .A1(net1579),
    .A2(net94));
 sg13g2_a21oi_1 _15417_ (.A1(net1478),
    .A2(_07103_),
    .Y(_07114_),
    .B1(net94));
 sg13g2_nor2_1 _15418_ (.A(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .B(_07114_),
    .Y(_07115_));
 sg13g2_a21oi_1 _15419_ (.A1(_07103_),
    .A2(_07113_),
    .Y(_00154_),
    .B1(_07115_));
 sg13g2_nand2_1 _15420_ (.Y(_07116_),
    .A(net299),
    .B(_05616_));
 sg13g2_nand2_1 _15421_ (.Y(_07117_),
    .A(_07070_),
    .B(_07068_));
 sg13g2_nor2_1 _15422_ (.A(_07070_),
    .B(_07068_),
    .Y(_07118_));
 sg13g2_a21oi_1 _15423_ (.A1(_07098_),
    .A2(_07117_),
    .Y(_07119_),
    .B1(_07118_));
 sg13g2_nand2_1 _15424_ (.Y(_07120_),
    .A(\ex_block_i.alu_i.imd_val_q_i_63_ ),
    .B(net320));
 sg13g2_a21oi_2 _15425_ (.B1(net1566),
    .Y(_07121_),
    .A2(_07120_),
    .A1(net1567));
 sg13g2_nand2_1 _15426_ (.Y(_07122_),
    .A(_07018_),
    .B(_07080_));
 sg13g2_nand2_1 _15427_ (.Y(_07123_),
    .A(_07086_),
    .B(_07122_));
 sg13g2_and2_2 _15428_ (.A(_07079_),
    .B(_07123_),
    .X(_07124_));
 sg13g2_buf_4 fanout840 (.X(net840),
    .A(net841));
 sg13g2_o21ai_1 _15430_ (.B1(_07024_),
    .Y(_07126_),
    .A1(_07026_),
    .A2(_07028_));
 sg13g2_o21ai_1 _15431_ (.B1(_07126_),
    .Y(_07127_),
    .A1(_07072_),
    .A2(_07027_));
 sg13g2_nor2_1 _15432_ (.A(_07078_),
    .B(_07127_),
    .Y(_07128_));
 sg13g2_a21oi_2 _15433_ (.B1(_07128_),
    .Y(_07129_),
    .A2(_07078_),
    .A1(_07024_));
 sg13g2_a21oi_1 _15434_ (.A1(_07075_),
    .A2(_07077_),
    .Y(_07130_),
    .B1(_07024_));
 sg13g2_nor2_1 _15435_ (.A(_07075_),
    .B(_07077_),
    .Y(_07131_));
 sg13g2_nor2_1 _15436_ (.A(_07130_),
    .B(_07131_),
    .Y(_07132_));
 sg13g2_o21ai_1 _15437_ (.B1(net214),
    .Y(_07133_),
    .A1(net1259),
    .A2(net90));
 sg13g2_xnor2_1 _15438_ (.Y(_07134_),
    .A(net1324),
    .B(_07133_));
 sg13g2_a21oi_1 _15439_ (.A1(net243),
    .A2(net1320),
    .Y(_07135_),
    .B1(net1372));
 sg13g2_xor2_1 _15440_ (.B(_07135_),
    .A(_07134_),
    .X(_07136_));
 sg13g2_xnor2_1 _15441_ (.Y(_07137_),
    .A(_07132_),
    .B(_07136_));
 sg13g2_xnor2_1 _15442_ (.Y(_07138_),
    .A(_07129_),
    .B(_07137_));
 sg13g2_xnor2_1 _15443_ (.Y(_07139_),
    .A(_07124_),
    .B(_07138_));
 sg13g2_nor2_1 _15444_ (.A(_07035_),
    .B(_07095_),
    .Y(_07140_));
 sg13g2_mux2_1 _15445_ (.A0(_07086_),
    .A1(_07080_),
    .S(_07079_),
    .X(_07141_));
 sg13g2_nand2b_1 _15446_ (.Y(_07142_),
    .B(_07079_),
    .A_N(_07032_));
 sg13g2_mux2_1 _15447_ (.A0(_07141_),
    .A1(_07142_),
    .S(_07019_),
    .X(_07143_));
 sg13g2_nor2_1 _15448_ (.A(_07018_),
    .B(_07030_),
    .Y(_07144_));
 sg13g2_mux2_1 _15449_ (.A0(_07123_),
    .A1(_07144_),
    .S(_07079_),
    .X(_07145_));
 sg13g2_nand3_1 _15450_ (.B(_07017_),
    .C(_07145_),
    .A(_07013_),
    .Y(_07146_));
 sg13g2_o21ai_1 _15451_ (.B1(_07146_),
    .Y(_07147_),
    .A1(_07084_),
    .A2(_07143_));
 sg13g2_a21oi_2 _15452_ (.B1(_07147_),
    .Y(_07148_),
    .A2(_07140_),
    .A1(_07044_));
 sg13g2_xnor2_1 _15453_ (.Y(_07149_),
    .A(_07139_),
    .B(_07148_));
 sg13g2_xnor2_1 _15454_ (.Y(_07150_),
    .A(_07121_),
    .B(_07149_));
 sg13g2_xnor2_1 _15455_ (.Y(_07151_),
    .A(_07119_),
    .B(_07150_));
 sg13g2_nand2_1 _15456_ (.Y(_07152_),
    .A(net1539),
    .B(_07151_));
 sg13g2_nand3_1 _15457_ (.B(_07116_),
    .C(_07152_),
    .A(net1182),
    .Y(_07153_));
 sg13g2_a21oi_1 _15458_ (.A1(_05016_),
    .A2(_06346_),
    .Y(_07154_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_31_ ));
 sg13g2_a21oi_1 _15459_ (.A1(\ex_block_i.alu_i.imd_val_q_i_63_ ),
    .A2(net37),
    .Y(_07155_),
    .B1(net310));
 sg13g2_a21oi_1 _15460_ (.A1(net315),
    .A2(_07154_),
    .Y(_07156_),
    .B1(_07155_));
 sg13g2_nand2_1 _15461_ (.Y(_07157_),
    .A(net36),
    .B(net1261));
 sg13g2_o21ai_1 _15462_ (.B1(_07157_),
    .Y(_07158_),
    .A1(_01846_),
    .A2(net1262));
 sg13g2_nand2_1 _15463_ (.Y(_07159_),
    .A(net422),
    .B(_07158_));
 sg13g2_o21ai_1 _15464_ (.B1(net1636),
    .Y(_07160_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .A2(net304));
 sg13g2_nand3_1 _15465_ (.B(_07159_),
    .C(_07160_),
    .A(net1575),
    .Y(_07161_));
 sg13g2_a221oi_1 _15466_ (.B2(net1890),
    .C1(_07161_),
    .B1(_07156_),
    .A1(net1884),
    .Y(_07162_),
    .A2(_07104_));
 sg13g2_nand2_1 _15467_ (.Y(_07163_),
    .A(net360),
    .B(net1579));
 sg13g2_o21ai_1 _15468_ (.B1(net1186),
    .Y(_07164_),
    .A1(_07162_),
    .A2(_07163_));
 sg13g2_o21ai_1 _15469_ (.B1(_07164_),
    .Y(_07165_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_63_ ),
    .A2(net1575));
 sg13g2_a22oi_1 _15470_ (.Y(_00155_),
    .B1(_07153_),
    .B2(_07165_),
    .A2(net95),
    .A1(_01846_));
 sg13g2_mux2_1 _15471_ (.A0(net1513),
    .A1(data_addr_o_6_),
    .S(net1451),
    .X(_07166_));
 sg13g2_mux2_1 _15472_ (.A0(_07166_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_6_ ),
    .S(net1223),
    .X(_00156_));
 sg13g2_mux2_1 _15473_ (.A0(net283),
    .A1(data_addr_o_7_),
    .S(_03951_),
    .X(_07167_));
 sg13g2_mux2_1 _15474_ (.A0(_07167_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_7_ ),
    .S(net1230),
    .X(_00157_));
 sg13g2_nand2_1 _15475_ (.Y(_07168_),
    .A(_03914_),
    .B(net1449));
 sg13g2_o21ai_1 _15476_ (.B1(_07168_),
    .Y(_07169_),
    .A1(data_addr_o_8_),
    .A2(net1449));
 sg13g2_nand2_1 _15477_ (.Y(_07170_),
    .A(\ex_block_i.alu_i.imd_val_q_i_8_ ),
    .B(net1228));
 sg13g2_o21ai_1 _15478_ (.B1(_07170_),
    .Y(_00158_),
    .A1(net1228),
    .A2(_07169_));
 sg13g2_mux2_1 _15479_ (.A0(net1466),
    .A1(data_addr_o_9_),
    .S(net1451),
    .X(_07171_));
 sg13g2_mux2_1 _15480_ (.A0(_07171_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_9_ ),
    .S(net1225),
    .X(_00159_));
 sg13g2_nand3_1 _15481_ (.B(net308),
    .C(net1634),
    .A(_03957_),
    .Y(_07172_));
 sg13g2_nand2_1 _15482_ (.Y(_07173_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .B(_07172_));
 sg13g2_o21ai_1 _15483_ (.B1(_07173_),
    .Y(_00160_),
    .A1(_03184_),
    .A2(_07172_));
 sg13g2_buf_4 fanout839 (.X(net839),
    .A(\register_file_i/_2911_ ));
 sg13g2_nand2_1 _15485_ (.Y(_07175_),
    .A(net2111),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ));
 sg13g2_a21oi_1 _15486_ (.A1(_04129_),
    .A2(_07175_),
    .Y(_07176_),
    .B1(_01535_));
 sg13g2_nor2_2 _15487_ (.A(net2105),
    .B(_07176_),
    .Y(_07177_));
 sg13g2_nor3_1 _15488_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .B(net142),
    .C(_07177_),
    .Y(_07178_));
 sg13g2_a21oi_1 _15489_ (.A1(_04486_),
    .A2(net143),
    .Y(_00161_),
    .B1(_07178_));
 sg13g2_xor2_1 _15490_ (.B(net2113),
    .A(net554),
    .X(_07179_));
 sg13g2_nor3_1 _15491_ (.A(net142),
    .B(_07177_),
    .C(_07179_),
    .Y(_07180_));
 sg13g2_a21oi_1 _15492_ (.A1(_04194_),
    .A2(net143),
    .Y(_00162_),
    .B1(_07180_));
 sg13g2_nor3_1 _15493_ (.A(net142),
    .B(_04101_),
    .C(_07177_),
    .Y(_07181_));
 sg13g2_a21oi_1 _15494_ (.A1(_04487_),
    .A2(net143),
    .Y(_00163_),
    .B1(_07181_));
 sg13g2_nor3_1 _15495_ (.A(net142),
    .B(_04104_),
    .C(_07177_),
    .Y(_07182_));
 sg13g2_a21oi_1 _15496_ (.A1(_04112_),
    .A2(net143),
    .Y(_00164_),
    .B1(_07182_));
 sg13g2_nor3_1 _15497_ (.A(net142),
    .B(_04114_),
    .C(_07177_),
    .Y(_07183_));
 sg13g2_a21oi_1 _15498_ (.A1(_06244_),
    .A2(net143),
    .Y(_00165_),
    .B1(_07183_));
 sg13g2_inv_1 _15499_ (.Y(_07184_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ));
 sg13g2_nor3_1 _15500_ (.A(_04035_),
    .B(net323),
    .C(_05912_),
    .Y(_07185_));
 sg13g2_a21oi_1 _15501_ (.A1(_07184_),
    .A2(_04035_),
    .Y(_00166_),
    .B1(_07185_));
 sg13g2_inv_1 _15502_ (.Y(_07186_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ));
 sg13g2_nor2_1 _15503_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ),
    .Y(_07187_));
 sg13g2_nor3_1 _15504_ (.A(_04035_),
    .B(net322),
    .C(_07187_),
    .Y(_07188_));
 sg13g2_a21oi_1 _15505_ (.A1(_07186_),
    .A2(_04035_),
    .Y(_00167_),
    .B1(_07188_));
 sg13g2_nor2_1 _15506_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ),
    .B(_05153_),
    .Y(_07189_));
 sg13g2_nand3_1 _15507_ (.B(net1885),
    .C(net36),
    .A(\ex_block_i.alu_i.imd_val_q_i_63_ ),
    .Y(_07190_));
 sg13g2_and2_1 _15508_ (.A(net419),
    .B(net1220),
    .X(_07191_));
 sg13g2_a221oi_1 _15509_ (.B2(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ),
    .C1(_04134_),
    .B1(_07191_),
    .A1(net313),
    .Y(_07192_),
    .A2(net1638));
 sg13g2_a21oi_1 _15510_ (.A1(_07190_),
    .A2(_07192_),
    .Y(_07193_),
    .B1(net337));
 sg13g2_nor2_1 _15511_ (.A(net93),
    .B(_07193_),
    .Y(_07194_));
 sg13g2_nor2_1 _15512_ (.A(net297),
    .B(_07003_),
    .Y(_07195_));
 sg13g2_nand2_1 _15513_ (.Y(_07196_),
    .A(_07121_),
    .B(_07149_));
 sg13g2_o21ai_1 _15514_ (.B1(_07117_),
    .Y(_07197_),
    .A1(_07098_),
    .A2(_07118_));
 sg13g2_nor2_1 _15515_ (.A(_07121_),
    .B(_07149_),
    .Y(_07198_));
 sg13g2_a21oi_1 _15516_ (.A1(_07196_),
    .A2(_07197_),
    .Y(_07199_),
    .B1(_07198_));
 sg13g2_nand2_1 _15517_ (.Y(_07200_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ),
    .B(net320));
 sg13g2_a21oi_1 _15518_ (.A1(_05910_),
    .A2(_07200_),
    .Y(_07201_),
    .B1(_05912_));
 sg13g2_nand2_1 _15519_ (.Y(_07202_),
    .A(_07024_),
    .B(_07077_));
 sg13g2_nand3_1 _15520_ (.B(net215),
    .C(_07202_),
    .A(_05411_),
    .Y(_07203_));
 sg13g2_o21ai_1 _15521_ (.B1(_07203_),
    .Y(_07204_),
    .A1(_07024_),
    .A2(_07077_));
 sg13g2_o21ai_1 _15522_ (.B1(net216),
    .Y(_07205_),
    .A1(net1324),
    .A2(net1371));
 sg13g2_nor2b_1 _15523_ (.A(_07134_),
    .B_N(_07205_),
    .Y(_07206_));
 sg13g2_a21oi_1 _15524_ (.A1(net243),
    .A2(net1320),
    .Y(_07207_),
    .B1(_07134_));
 sg13g2_nor3_1 _15525_ (.A(_07130_),
    .B(_07131_),
    .C(_07207_),
    .Y(_07208_));
 sg13g2_and3_1 _15526_ (.X(_07209_),
    .A(net242),
    .B(net1320),
    .C(_07134_));
 sg13g2_o21ai_1 _15527_ (.B1(net1371),
    .Y(_07210_),
    .A1(_07208_),
    .A2(_07209_));
 sg13g2_nand3_1 _15528_ (.B(_07132_),
    .C(_07134_),
    .A(net1324),
    .Y(_07211_));
 sg13g2_a21oi_2 _15529_ (.B1(net1372),
    .Y(_07212_),
    .A2(_07211_),
    .A1(_07210_));
 sg13g2_a21oi_2 _15530_ (.B1(_07212_),
    .Y(_07213_),
    .A2(_07206_),
    .A1(_07204_));
 sg13g2_a21o_1 _15531_ (.A2(_07129_),
    .A1(_07124_),
    .B1(_07137_),
    .X(_07214_));
 sg13g2_o21ai_1 _15532_ (.B1(_07214_),
    .Y(_07215_),
    .A1(_07124_),
    .A2(_07129_));
 sg13g2_or2_1 _15533_ (.X(_07216_),
    .B(_07137_),
    .A(_07129_));
 sg13g2_and2_1 _15534_ (.A(_07129_),
    .B(_07137_),
    .X(_07217_));
 sg13g2_nand3b_1 _15535_ (.B(_07217_),
    .C(_07124_),
    .Y(_07218_),
    .A_N(_07148_));
 sg13g2_o21ai_1 _15536_ (.B1(_07218_),
    .Y(_07219_),
    .A1(_07124_),
    .A2(_07216_));
 sg13g2_a21oi_1 _15537_ (.A1(_07148_),
    .A2(_07215_),
    .Y(_07220_),
    .B1(_07219_));
 sg13g2_xnor2_1 _15538_ (.Y(_07221_),
    .A(_07213_),
    .B(_07220_));
 sg13g2_xor2_1 _15539_ (.B(_07221_),
    .A(_07201_),
    .X(_07222_));
 sg13g2_xnor2_1 _15540_ (.Y(_07223_),
    .A(_07199_),
    .B(_07222_));
 sg13g2_nand3_1 _15541_ (.B(net1472),
    .C(_07223_),
    .A(net1188),
    .Y(_07224_));
 sg13g2_o21ai_1 _15542_ (.B1(_07224_),
    .Y(_00168_),
    .A1(_07189_),
    .A2(_07194_));
 sg13g2_nand2b_1 _15543_ (.Y(_07225_),
    .B(_07221_),
    .A_N(_07201_));
 sg13g2_o21ai_1 _15544_ (.B1(_07196_),
    .Y(_07226_),
    .A1(_07119_),
    .A2(_07198_));
 sg13g2_nor2b_1 _15545_ (.A(_07221_),
    .B_N(_07201_),
    .Y(_07227_));
 sg13g2_a21oi_1 _15546_ (.A1(_07225_),
    .A2(_07226_),
    .Y(_07228_),
    .B1(_07227_));
 sg13g2_or2_1 _15547_ (.X(_07229_),
    .B(_07217_),
    .A(_07213_));
 sg13g2_a22oi_1 _15548_ (.Y(_07230_),
    .B1(_07229_),
    .B2(_07124_),
    .A2(_07216_),
    .A1(_07213_));
 sg13g2_a21oi_1 _15549_ (.A1(_07124_),
    .A2(_07216_),
    .Y(_07231_),
    .B1(_07217_));
 sg13g2_nand2b_1 _15550_ (.Y(_07232_),
    .B(_07213_),
    .A_N(_07231_));
 sg13g2_o21ai_1 _15551_ (.B1(_07232_),
    .Y(_07233_),
    .A1(_07148_),
    .A2(_07230_));
 sg13g2_nand2_1 _15552_ (.Y(_07234_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ),
    .B(net320));
 sg13g2_a21oi_1 _15553_ (.A1(net1568),
    .A2(_07234_),
    .Y(_07235_),
    .B1(net1566));
 sg13g2_xnor2_1 _15554_ (.Y(_07236_),
    .A(_07212_),
    .B(_07235_));
 sg13g2_xnor2_1 _15555_ (.Y(_07237_),
    .A(_07233_),
    .B(_07236_));
 sg13g2_xnor2_1 _15556_ (.Y(_07238_),
    .A(_07228_),
    .B(_07237_));
 sg13g2_nand3_1 _15557_ (.B(net1543),
    .C(net1182),
    .A(net1188),
    .Y(_07239_));
 sg13g2_nor2_1 _15558_ (.A(net375),
    .B(net341),
    .Y(_07240_));
 sg13g2_nand2_1 _15559_ (.Y(_07241_),
    .A(net315),
    .B(net1638));
 sg13g2_o21ai_1 _15560_ (.B1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ),
    .Y(_07242_),
    .A1(_04134_),
    .A2(_07191_));
 sg13g2_o21ai_1 _15561_ (.B1(_07242_),
    .Y(_07243_),
    .A1(net93),
    .A2(_07241_));
 sg13g2_a22oi_1 _15562_ (.Y(_07244_),
    .B1(_07240_),
    .B2(_07243_),
    .A2(net97),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ));
 sg13g2_o21ai_1 _15563_ (.B1(_07244_),
    .Y(_00169_),
    .A1(_07238_),
    .A2(_07239_));
 sg13g2_a21oi_1 _15564_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .A2(net2110),
    .Y(_07245_),
    .B1(net2105));
 sg13g2_o21ai_1 _15565_ (.B1(_07175_),
    .Y(_07246_),
    .A1(_04065_),
    .A2(_07245_));
 sg13g2_nor3_1 _15566_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .B(net2112),
    .C(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .Y(_07247_));
 sg13g2_and2_1 _15567_ (.A(_04084_),
    .B(_07247_),
    .X(_07248_));
 sg13g2_o21ai_1 _15568_ (.B1(net2111),
    .Y(_07249_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ),
    .A2(_07248_));
 sg13g2_a221oi_1 _15569_ (.B2(_04130_),
    .C1(net1888),
    .B1(_07249_),
    .A1(_03184_),
    .Y(_07250_),
    .A2(net1634));
 sg13g2_nor3_1 _15570_ (.A(net142),
    .B(_07246_),
    .C(_07250_),
    .Y(_07251_));
 sg13g2_a21o_1 _15571_ (.A2(net143),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0_ ),
    .B1(_07251_),
    .X(_00170_));
 sg13g2_nand2_2 _15572_ (.Y(_07252_),
    .A(_03848_),
    .B(net1634));
 sg13g2_a21oi_1 _15573_ (.A1(_04130_),
    .A2(_07249_),
    .Y(_07253_),
    .B1(net1710));
 sg13g2_a21oi_2 _15574_ (.B1(_07246_),
    .Y(_07254_),
    .A2(_07253_),
    .A1(_07252_));
 sg13g2_mux2_1 _15575_ (.A0(net2110),
    .A1(_07254_),
    .S(_03957_),
    .X(_00171_));
 sg13g2_or2_1 _15576_ (.X(_07255_),
    .B(net419),
    .A(net1888));
 sg13g2_a21oi_1 _15577_ (.A1(net1882),
    .A2(_07248_),
    .Y(_07256_),
    .B1(_07255_));
 sg13g2_a21oi_2 _15578_ (.B1(_07246_),
    .Y(_07257_),
    .A2(_07256_),
    .A1(_07252_));
 sg13g2_mux2_1 _15579_ (.A0(net2105),
    .A1(_07257_),
    .S(_03957_),
    .X(_00172_));
 sg13g2_and2_1 _15580_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .B(_04118_),
    .X(_07258_));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(net839));
 sg13g2_nand2_1 _15582_ (.Y(_07260_),
    .A(net1145),
    .B(net1431));
 sg13g2_o21ai_1 _15583_ (.B1(_07260_),
    .Y(_07261_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ),
    .A2(net1431));
 sg13g2_nand3_1 _15584_ (.B(net1893),
    .C(_03957_),
    .A(net1881),
    .Y(_07262_));
 sg13g2_buf_4 fanout837 (.X(net837),
    .A(net839));
 sg13g2_buf_2 fanout836 (.A(\register_file_i/_2913_ ),
    .X(net836));
 sg13g2_nand2_1 _15587_ (.Y(_07265_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_0_ ),
    .B(net1254));
 sg13g2_o21ai_1 _15588_ (.B1(_07265_),
    .Y(_00173_),
    .A1(_07261_),
    .A2(net1254));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(\register_file_i/_2913_ ));
 sg13g2_buf_2 fanout834 (.A(\register_file_i/_2913_ ),
    .X(net834));
 sg13g2_nand2_1 _15591_ (.Y(_07268_),
    .A(_02895_),
    .B(net1430));
 sg13g2_o21ai_1 _15592_ (.B1(_07268_),
    .Y(_07269_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ),
    .A2(net1428));
 sg13g2_nand2_1 _15593_ (.Y(_07270_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_10_ ),
    .B(net1254));
 sg13g2_o21ai_1 _15594_ (.B1(_07270_),
    .Y(_00174_),
    .A1(net1254),
    .A2(_07269_));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(net834));
 sg13g2_buf_4 fanout832 (.X(net832),
    .A(net834));
 sg13g2_nand2b_1 _15597_ (.Y(_07273_),
    .B(net1442),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_o21ai_1 _15598_ (.B1(_07273_),
    .Y(_07274_),
    .A1(data_addr_o_11_),
    .A2(net1442));
 sg13g2_nand2_1 _15599_ (.Y(_07275_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_11_ ),
    .B(net1254));
 sg13g2_o21ai_1 _15600_ (.B1(_07275_),
    .Y(_00175_),
    .A1(net1253),
    .A2(_07274_));
 sg13g2_nor3_1 _15601_ (.A(net2105),
    .B(_01839_),
    .C(net142),
    .Y(_07276_));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(\register_file_i/_2927_ ));
 sg13g2_buf_2 fanout830 (.A(net831),
    .X(net830));
 sg13g2_and2_1 _15604_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ),
    .B(net1441),
    .X(_07279_));
 sg13g2_a21oi_1 _15605_ (.A1(data_addr_o_12_),
    .A2(net1429),
    .Y(_07280_),
    .B1(_07279_));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(net831));
 sg13g2_nor2_1 _15607_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_12_ ),
    .B(net1212),
    .Y(_07282_));
 sg13g2_a21oi_1 _15608_ (.A1(net1212),
    .A2(_07280_),
    .Y(_00176_),
    .B1(_07282_));
 sg13g2_nand2b_1 _15609_ (.Y(_07283_),
    .B(net1445),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_o21ai_1 _15610_ (.B1(_07283_),
    .Y(_07284_),
    .A1(data_addr_o_13_),
    .A2(net1445));
 sg13g2_nand2_1 _15611_ (.Y(_07285_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_13_ ),
    .B(net1252));
 sg13g2_o21ai_1 _15612_ (.B1(_07285_),
    .Y(_00177_),
    .A1(net1252),
    .A2(_07284_));
 sg13g2_nand2_1 _15613_ (.Y(_07286_),
    .A(_03265_),
    .B(net1432));
 sg13g2_o21ai_1 _15614_ (.B1(_07286_),
    .Y(_07287_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ),
    .A2(net1431));
 sg13g2_buf_4 fanout828 (.X(net828),
    .A(net831));
 sg13g2_nand2_1 _15616_ (.Y(_07289_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_14_ ),
    .B(net1252));
 sg13g2_o21ai_1 _15617_ (.B1(_07289_),
    .Y(_00178_),
    .A1(net1252),
    .A2(_07287_));
 sg13g2_nand2b_1 _15618_ (.Y(_07290_),
    .B(net1441),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_o21ai_1 _15619_ (.B1(_07290_),
    .Y(_07291_),
    .A1(data_addr_o_15_),
    .A2(net1441));
 sg13g2_nand2_1 _15620_ (.Y(_07292_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_15_ ),
    .B(net1252));
 sg13g2_o21ai_1 _15621_ (.B1(_07292_),
    .Y(_00179_),
    .A1(net1252),
    .A2(_07291_));
 sg13g2_nand2b_1 _15622_ (.Y(_07293_),
    .B(net1442),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ));
 sg13g2_o21ai_1 _15623_ (.B1(_07293_),
    .Y(_07294_),
    .A1(data_addr_o_16_),
    .A2(net1442));
 sg13g2_nand2_1 _15624_ (.Y(_07295_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_16_ ),
    .B(net1255));
 sg13g2_o21ai_1 _15625_ (.B1(_07295_),
    .Y(_00180_),
    .A1(net1254),
    .A2(_07294_));
 sg13g2_nor2_1 _15626_ (.A(_04296_),
    .B(net1428),
    .Y(_07296_));
 sg13g2_a21oi_1 _15627_ (.A1(data_addr_o_17_),
    .A2(net1428),
    .Y(_07297_),
    .B1(_07296_));
 sg13g2_nor2_1 _15628_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_17_ ),
    .B(net1215),
    .Y(_07298_));
 sg13g2_a21oi_1 _15629_ (.A1(net1217),
    .A2(_07297_),
    .Y(_00181_),
    .B1(_07298_));
 sg13g2_nor2_1 _15630_ (.A(_04216_),
    .B(net1428),
    .Y(_07299_));
 sg13g2_a21oi_1 _15631_ (.A1(data_addr_o_18_),
    .A2(net1428),
    .Y(_07300_),
    .B1(_07299_));
 sg13g2_nor2_1 _15632_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_18_ ),
    .B(net1215),
    .Y(_07301_));
 sg13g2_a21oi_1 _15633_ (.A1(net1215),
    .A2(_07300_),
    .Y(_00182_),
    .B1(_07301_));
 sg13g2_and2_1 _15634_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ),
    .B(net1446),
    .X(_07302_));
 sg13g2_a21oi_1 _15635_ (.A1(data_addr_o_19_),
    .A2(net1431),
    .Y(_07303_),
    .B1(_07302_));
 sg13g2_nor2_1 _15636_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_19_ ),
    .B(net1215),
    .Y(_07304_));
 sg13g2_a21oi_1 _15637_ (.A1(net1217),
    .A2(_07303_),
    .Y(_00183_),
    .B1(_07304_));
 sg13g2_nor2_1 _15638_ (.A(_02293_),
    .B(net1432),
    .Y(_07305_));
 sg13g2_a21oi_2 _15639_ (.B1(_07305_),
    .Y(_07306_),
    .A2(net1431),
    .A1(net1111));
 sg13g2_buf_4 fanout827 (.X(net827),
    .A(net828));
 sg13g2_nor2_1 _15641_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_1_ ),
    .B(net1214),
    .Y(_07308_));
 sg13g2_a21oi_1 _15642_ (.A1(net1214),
    .A2(_07306_),
    .Y(_00184_),
    .B1(_07308_));
 sg13g2_nor2_1 _15643_ (.A(_03274_),
    .B(net1446),
    .Y(_07309_));
 sg13g2_a21oi_1 _15644_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ),
    .A2(net1445),
    .Y(_07310_),
    .B1(_07309_));
 sg13g2_nor2_1 _15645_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_20_ ),
    .B(_07276_),
    .Y(_07311_));
 sg13g2_a21oi_1 _15646_ (.A1(net1217),
    .A2(_07310_),
    .Y(_00185_),
    .B1(_07311_));
 sg13g2_nor2_1 _15647_ (.A(_04416_),
    .B(net1432),
    .Y(_07312_));
 sg13g2_a21oi_1 _15648_ (.A1(data_addr_o_21_),
    .A2(net1431),
    .Y(_07313_),
    .B1(_07312_));
 sg13g2_nor2_1 _15649_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_21_ ),
    .B(net1217),
    .Y(_07314_));
 sg13g2_a21oi_1 _15650_ (.A1(net1217),
    .A2(_07313_),
    .Y(_00186_),
    .B1(_07314_));
 sg13g2_nor2_1 _15651_ (.A(_03174_),
    .B(net1445),
    .Y(_07315_));
 sg13g2_a21oi_1 _15652_ (.A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ),
    .A2(net1445),
    .Y(_07316_),
    .B1(_07315_));
 sg13g2_nor2_1 _15653_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_22_ ),
    .B(net1217),
    .Y(_07317_));
 sg13g2_a21oi_1 _15654_ (.A1(net1217),
    .A2(_07316_),
    .Y(_00187_),
    .B1(_07317_));
 sg13g2_nand2_1 _15655_ (.Y(_07318_),
    .A(_03278_),
    .B(net1430));
 sg13g2_o21ai_1 _15656_ (.B1(_07318_),
    .Y(_07319_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ),
    .A2(net1430));
 sg13g2_nand2_1 _15657_ (.Y(_07320_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_23_ ),
    .B(net1256));
 sg13g2_o21ai_1 _15658_ (.B1(_07320_),
    .Y(_00188_),
    .A1(net1255),
    .A2(_07319_));
 sg13g2_nand2b_1 _15659_ (.Y(_07321_),
    .B(net1443),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ));
 sg13g2_o21ai_1 _15660_ (.B1(_07321_),
    .Y(_07322_),
    .A1(data_addr_o_24_),
    .A2(net1443));
 sg13g2_nand2_1 _15661_ (.Y(_07323_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_24_ ),
    .B(net1256));
 sg13g2_o21ai_1 _15662_ (.B1(_07323_),
    .Y(_00189_),
    .A1(net1255),
    .A2(_07322_));
 sg13g2_nand2b_1 _15663_ (.Y(_07324_),
    .B(net1443),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_o21ai_1 _15664_ (.B1(_07324_),
    .Y(_07325_),
    .A1(data_addr_o_25_),
    .A2(net1442));
 sg13g2_nand2_1 _15665_ (.Y(_07326_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_25_ ),
    .B(net1255));
 sg13g2_o21ai_1 _15666_ (.B1(_07326_),
    .Y(_00190_),
    .A1(net1255),
    .A2(_07325_));
 sg13g2_nand2_1 _15667_ (.Y(_07327_),
    .A(_03182_),
    .B(net1430));
 sg13g2_o21ai_1 _15668_ (.B1(_07327_),
    .Y(_07328_),
    .A1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ),
    .A2(net1430));
 sg13g2_nand2_1 _15669_ (.Y(_07329_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_26_ ),
    .B(net1256));
 sg13g2_o21ai_1 _15670_ (.B1(_07329_),
    .Y(_00191_),
    .A1(net1253),
    .A2(_07328_));
 sg13g2_nand2_1 _15671_ (.Y(_07330_),
    .A(_01907_),
    .B(net1444));
 sg13g2_o21ai_1 _15672_ (.B1(_07330_),
    .Y(_07331_),
    .A1(net2487),
    .A2(net1441));
 sg13g2_nand2_1 _15673_ (.Y(_07332_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_27_ ),
    .B(net1255));
 sg13g2_o21ai_1 _15674_ (.B1(_07332_),
    .Y(_00192_),
    .A1(net1253),
    .A2(_07331_));
 sg13g2_nor2_1 _15675_ (.A(_01281_),
    .B(net1429),
    .Y(_07333_));
 sg13g2_a21oi_1 _15676_ (.A1(data_addr_o_28_),
    .A2(net1429),
    .Y(_07334_),
    .B1(_07333_));
 sg13g2_nor2_1 _15677_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_28_ ),
    .B(net1213),
    .Y(_07335_));
 sg13g2_a21oi_1 _15678_ (.A1(net1213),
    .A2(_07334_),
    .Y(_00193_),
    .B1(_07335_));
 sg13g2_nand2b_1 _15679_ (.Y(_07336_),
    .B(net1444),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_o21ai_1 _15680_ (.B1(_07336_),
    .Y(_07337_),
    .A1(data_addr_o_29_),
    .A2(net1441));
 sg13g2_nand2_1 _15681_ (.Y(_07338_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_29_ ),
    .B(net1252));
 sg13g2_o21ai_1 _15682_ (.B1(_07338_),
    .Y(_00194_),
    .A1(net1252),
    .A2(_07337_));
 sg13g2_nor2_1 _15683_ (.A(_04215_),
    .B(net1431),
    .Y(_07339_));
 sg13g2_a21oi_1 _15684_ (.A1(data_addr_o_2_),
    .A2(net1431),
    .Y(_07340_),
    .B1(_07339_));
 sg13g2_nor2_1 _15685_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_2_ ),
    .B(net1214),
    .Y(_07341_));
 sg13g2_a21oi_1 _15686_ (.A1(net1214),
    .A2(_07340_),
    .Y(_00195_),
    .B1(_07341_));
 sg13g2_nand2b_1 _15687_ (.Y(_07342_),
    .B(net1444),
    .A_N(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ));
 sg13g2_o21ai_1 _15688_ (.B1(_07342_),
    .Y(_07343_),
    .A1(net2494),
    .A2(net1441));
 sg13g2_nand2_1 _15689_ (.Y(_07344_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_30_ ),
    .B(net1253));
 sg13g2_o21ai_1 _15690_ (.B1(_07344_),
    .Y(_00196_),
    .A1(net1253),
    .A2(_07343_));
 sg13g2_inv_1 _15691_ (.Y(_07345_),
    .A(_04118_));
 sg13g2_o21ai_1 _15692_ (.B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ),
    .Y(_07346_),
    .A1(net36),
    .A2(_07345_));
 sg13g2_nand2_1 _15693_ (.Y(_07347_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31_ ),
    .B(net1253));
 sg13g2_o21ai_1 _15694_ (.B1(_07347_),
    .Y(_00197_),
    .A1(net1253),
    .A2(_07346_));
 sg13g2_and2_1 _15695_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ),
    .B(net1442),
    .X(_07348_));
 sg13g2_a21oi_1 _15696_ (.A1(data_addr_o_3_),
    .A2(net1428),
    .Y(_07349_),
    .B1(_07348_));
 sg13g2_nor2_1 _15697_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_3_ ),
    .B(net1214),
    .Y(_07350_));
 sg13g2_a21oi_1 _15698_ (.A1(net1214),
    .A2(_07349_),
    .Y(_00198_),
    .B1(_07350_));
 sg13g2_nor2_1 _15699_ (.A(_02263_),
    .B(net1429),
    .Y(_07351_));
 sg13g2_a21oi_1 _15700_ (.A1(data_addr_o_4_),
    .A2(net1429),
    .Y(_07352_),
    .B1(_07351_));
 sg13g2_nor2_1 _15701_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_4_ ),
    .B(net1212),
    .Y(_07353_));
 sg13g2_a21oi_1 _15702_ (.A1(net1212),
    .A2(_07352_),
    .Y(_00199_),
    .B1(_07353_));
 sg13g2_nor2_1 _15703_ (.A(_04415_),
    .B(net1430),
    .Y(_07354_));
 sg13g2_a21oi_1 _15704_ (.A1(data_addr_o_5_),
    .A2(net1428),
    .Y(_07355_),
    .B1(_07354_));
 sg13g2_nor2_1 _15705_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_5_ ),
    .B(net1212),
    .Y(_07356_));
 sg13g2_a21oi_1 _15706_ (.A1(net1212),
    .A2(_07355_),
    .Y(_00200_),
    .B1(_07356_));
 sg13g2_and2_1 _15707_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ),
    .B(net1442),
    .X(_07357_));
 sg13g2_a21oi_1 _15708_ (.A1(data_addr_o_6_),
    .A2(net1428),
    .Y(_07358_),
    .B1(_07357_));
 sg13g2_nor2_1 _15709_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_6_ ),
    .B(net1214),
    .Y(_07359_));
 sg13g2_a21oi_1 _15710_ (.A1(net1214),
    .A2(_07358_),
    .Y(_00201_),
    .B1(_07359_));
 sg13g2_and2_1 _15711_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ),
    .B(net1441),
    .X(_07360_));
 sg13g2_a21oi_1 _15712_ (.A1(data_addr_o_7_),
    .A2(net1429),
    .Y(_07361_),
    .B1(_07360_));
 sg13g2_nor2_1 _15713_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_7_ ),
    .B(net1212),
    .Y(_07362_));
 sg13g2_a21oi_1 _15714_ (.A1(net1212),
    .A2(_07361_),
    .Y(_00202_),
    .B1(_07362_));
 sg13g2_nand2_1 _15715_ (.Y(_07363_),
    .A(_02175_),
    .B(net1443));
 sg13g2_o21ai_1 _15716_ (.B1(_07363_),
    .Y(_07364_),
    .A1(data_addr_o_8_),
    .A2(net1442));
 sg13g2_nand2_1 _15717_ (.Y(_07365_),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_8_ ),
    .B(net1254));
 sg13g2_o21ai_1 _15718_ (.B1(_07365_),
    .Y(_00203_),
    .A1(net1254),
    .A2(_07364_));
 sg13g2_and2_1 _15719_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ),
    .B(net1441),
    .X(_07366_));
 sg13g2_a21oi_1 _15720_ (.A1(data_addr_o_9_),
    .A2(net1429),
    .Y(_07367_),
    .B1(_07366_));
 sg13g2_nor2_1 _15721_ (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_9_ ),
    .B(net1213),
    .Y(_07368_));
 sg13g2_a21oi_1 _15722_ (.A1(net1213),
    .A2(_07367_),
    .Y(_00204_),
    .B1(_07368_));
 sg13g2_nor2_1 _15723_ (.A(_01831_),
    .B(net1255),
    .Y(_07369_));
 sg13g2_buf_4 fanout826 (.X(net826),
    .A(net828));
 sg13g2_nand2_2 _15725_ (.Y(_07371_),
    .A(net1883),
    .B(_03957_));
 sg13g2_nor4_2 _15726_ (.A(net2112),
    .B(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .C(net1006),
    .Y(_07372_),
    .D(_07371_));
 sg13g2_a21oi_1 _15727_ (.A1(_04085_),
    .A2(_07372_),
    .Y(_07373_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_0_ ));
 sg13g2_nor2_1 _15728_ (.A(net1209),
    .B(_07373_),
    .Y(_00205_));
 sg13g2_nor4_2 _15729_ (.A(_04112_),
    .B(_04194_),
    .C(net1006),
    .Y(_07374_),
    .D(_07371_));
 sg13g2_a21oi_1 _15730_ (.A1(_04085_),
    .A2(_07374_),
    .Y(_07375_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_10_ ));
 sg13g2_nor2_1 _15731_ (.A(net1209),
    .B(_07375_),
    .Y(_00206_));
 sg13g2_a21oi_1 _15732_ (.A1(_04151_),
    .A2(_07374_),
    .Y(_07376_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_11_ ));
 sg13g2_nor2_1 _15733_ (.A(net1209),
    .B(_07376_),
    .Y(_00207_));
 sg13g2_nor3_2 _15734_ (.A(net1005),
    .B(_04760_),
    .C(_07371_),
    .Y(_07377_));
 sg13g2_a21oi_1 _15735_ (.A1(_04332_),
    .A2(_07377_),
    .Y(_07378_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_12_ ));
 sg13g2_nor2_1 _15736_ (.A(net1210),
    .B(_07378_),
    .Y(_00208_));
 sg13g2_a21oi_1 _15737_ (.A1(_04488_),
    .A2(_07377_),
    .Y(_07379_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_13_ ));
 sg13g2_nor2_1 _15738_ (.A(net1208),
    .B(_07379_),
    .Y(_00209_));
 sg13g2_a21oi_1 _15739_ (.A1(_04332_),
    .A2(_07374_),
    .Y(_07380_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_14_ ));
 sg13g2_nor2_1 _15740_ (.A(net1210),
    .B(_07380_),
    .Y(_00210_));
 sg13g2_a21oi_1 _15741_ (.A1(_04488_),
    .A2(_07374_),
    .Y(_07381_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_15_ ));
 sg13g2_nor2_1 _15742_ (.A(net1208),
    .B(_07381_),
    .Y(_00211_));
 sg13g2_a21oi_1 _15743_ (.A1(_05632_),
    .A2(_07372_),
    .Y(_07382_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_16_ ));
 sg13g2_nor2_1 _15744_ (.A(net1209),
    .B(_07382_),
    .Y(_00212_));
 sg13g2_a21oi_1 _15745_ (.A1(_05892_),
    .A2(_07372_),
    .Y(_07383_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_17_ ));
 sg13g2_nor2_1 _15746_ (.A(net1210),
    .B(_07383_),
    .Y(_00213_));
 sg13g2_nor4_2 _15747_ (.A(net2112),
    .B(_04194_),
    .C(net1005),
    .Y(_07384_),
    .D(_07371_));
 sg13g2_a21oi_1 _15748_ (.A1(_05632_),
    .A2(_07384_),
    .Y(_07385_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_18_ ));
 sg13g2_nor2_1 _15749_ (.A(net1209),
    .B(_07385_),
    .Y(_00214_));
 sg13g2_buf_2 fanout825 (.A(\register_file_i/_2932_ ),
    .X(net825));
 sg13g2_a21oi_1 _15751_ (.A1(_05892_),
    .A2(_07384_),
    .Y(_07387_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_19_ ));
 sg13g2_nor2_1 _15752_ (.A(net1207),
    .B(_07387_),
    .Y(_00215_));
 sg13g2_a21oi_1 _15753_ (.A1(_04151_),
    .A2(_07372_),
    .Y(_07388_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_1_ ));
 sg13g2_nor2_1 _15754_ (.A(net1210),
    .B(_07388_),
    .Y(_00216_));
 sg13g2_a21oi_1 _15755_ (.A1(_06245_),
    .A2(_07372_),
    .Y(_07389_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_20_ ));
 sg13g2_nor2_1 _15756_ (.A(net1208),
    .B(_07389_),
    .Y(_00217_));
 sg13g2_a21oi_1 _15757_ (.A1(_06346_),
    .A2(_07372_),
    .Y(_07390_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_21_ ));
 sg13g2_nor2_1 _15758_ (.A(net1207),
    .B(_07390_),
    .Y(_00218_));
 sg13g2_a21oi_1 _15759_ (.A1(_06245_),
    .A2(_07384_),
    .Y(_07391_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_22_ ));
 sg13g2_nor2_1 _15760_ (.A(net1207),
    .B(_07391_),
    .Y(_00219_));
 sg13g2_a21oi_1 _15761_ (.A1(_06346_),
    .A2(_07384_),
    .Y(_07392_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_23_ ));
 sg13g2_nor2_1 _15762_ (.A(net1207),
    .B(_07392_),
    .Y(_00220_));
 sg13g2_a21oi_1 _15763_ (.A1(_05632_),
    .A2(_07377_),
    .Y(_07393_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_24_ ));
 sg13g2_nor2_1 _15764_ (.A(net1208),
    .B(_07393_),
    .Y(_00221_));
 sg13g2_a21oi_1 _15765_ (.A1(_05892_),
    .A2(_07377_),
    .Y(_07394_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_25_ ));
 sg13g2_nor2_1 _15766_ (.A(net1207),
    .B(_07394_),
    .Y(_00222_));
 sg13g2_a21oi_1 _15767_ (.A1(_05632_),
    .A2(_07374_),
    .Y(_07395_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_26_ ));
 sg13g2_nor2_1 _15768_ (.A(net1208),
    .B(_07395_),
    .Y(_00223_));
 sg13g2_a21oi_1 _15769_ (.A1(_05892_),
    .A2(_07374_),
    .Y(_07396_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_27_ ));
 sg13g2_nor2_1 _15770_ (.A(net1207),
    .B(_07396_),
    .Y(_00224_));
 sg13g2_buf_2 fanout824 (.A(net825),
    .X(net824));
 sg13g2_a21oi_1 _15772_ (.A1(_06245_),
    .A2(_07377_),
    .Y(_07398_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_28_ ));
 sg13g2_nor2_1 _15773_ (.A(net1208),
    .B(_07398_),
    .Y(_00225_));
 sg13g2_a21oi_1 _15774_ (.A1(_06346_),
    .A2(_07377_),
    .Y(_07399_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_29_ ));
 sg13g2_nor2_1 _15775_ (.A(net1208),
    .B(_07399_),
    .Y(_00226_));
 sg13g2_a21oi_1 _15776_ (.A1(_04085_),
    .A2(_07384_),
    .Y(_07400_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_2_ ));
 sg13g2_nor2_1 _15777_ (.A(net1209),
    .B(_07400_),
    .Y(_00227_));
 sg13g2_a21oi_1 _15778_ (.A1(_06245_),
    .A2(_07374_),
    .Y(_07401_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_30_ ));
 sg13g2_nor2_1 _15779_ (.A(net1208),
    .B(_07401_),
    .Y(_00228_));
 sg13g2_a21oi_1 _15780_ (.A1(_06346_),
    .A2(_07374_),
    .Y(_07402_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_31_ ));
 sg13g2_nor2_1 _15781_ (.A(net1211),
    .B(_07402_),
    .Y(_00229_));
 sg13g2_a21oi_1 _15782_ (.A1(_04151_),
    .A2(_07384_),
    .Y(_07403_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_3_ ));
 sg13g2_nor2_1 _15783_ (.A(net1210),
    .B(_07403_),
    .Y(_00230_));
 sg13g2_a21oi_1 _15784_ (.A1(_04332_),
    .A2(_07372_),
    .Y(_07404_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_4_ ));
 sg13g2_nor2_1 _15785_ (.A(net1210),
    .B(_07404_),
    .Y(_00231_));
 sg13g2_a21oi_1 _15786_ (.A1(_04488_),
    .A2(_07372_),
    .Y(_07405_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_5_ ));
 sg13g2_nor2_1 _15787_ (.A(net1207),
    .B(_07405_),
    .Y(_00232_));
 sg13g2_a21oi_1 _15788_ (.A1(_04332_),
    .A2(_07384_),
    .Y(_07406_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_6_ ));
 sg13g2_nor2_1 _15789_ (.A(net1210),
    .B(_07406_),
    .Y(_00233_));
 sg13g2_a21oi_1 _15790_ (.A1(_04488_),
    .A2(_07384_),
    .Y(_07407_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_7_ ));
 sg13g2_nor2_1 _15791_ (.A(net1207),
    .B(_07407_),
    .Y(_00234_));
 sg13g2_a21oi_1 _15792_ (.A1(_04085_),
    .A2(_07377_),
    .Y(_07408_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_8_ ));
 sg13g2_nor2_1 _15793_ (.A(net1209),
    .B(_07408_),
    .Y(_00235_));
 sg13g2_a21oi_1 _15794_ (.A1(_04151_),
    .A2(_07377_),
    .Y(_07409_),
    .B1(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_9_ ));
 sg13g2_nor2_1 _15795_ (.A(net1209),
    .B(_07409_),
    .Y(_00236_));
 sg13g2_inv_1 _15796_ (.Y(exc_cause_4_),
    .A(_03440_));
 sg13g2_and3_1 _15797_ (.X(_07410_),
    .A(_01631_),
    .B(_01520_),
    .C(_01632_));
 sg13g2_o21ai_1 _15798_ (.B1(_07410_),
    .Y(_07411_),
    .A1(\id_stage_i.branch_jump_set_done_q ),
    .A2(_01437_));
 sg13g2_nor2b_1 _15799_ (.A(_07411_),
    .B_N(_03194_),
    .Y(\id_stage_i.branch_jump_set_done_d ));
 sg13g2_nor2b_2 _15800_ (.A(_03849_),
    .B_N(_03846_),
    .Y(_07412_));
 sg13g2_nor2b_1 _15801_ (.A(_07412_),
    .B_N(\id_stage_i.perf_branch_o ),
    .Y(\id_stage_i.branch_set_raw_d ));
 sg13g2_nor2_1 _15802_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .B(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .Y(_07413_));
 sg13g2_nor2_1 _15803_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .B(net2104),
    .Y(_07414_));
 sg13g2_nand2b_1 _15804_ (.Y(_07415_),
    .B(_07414_),
    .A_N(fetch_enable_i));
 sg13g2_o21ai_1 _15805_ (.B1(_07415_),
    .Y(_07416_),
    .A1(\id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ),
    .A2(_01493_));
 sg13g2_nand2_1 _15806_ (.Y(_07417_),
    .A(_07413_),
    .B(_07416_));
 sg13g2_and2_1 _15807_ (.A(_01462_),
    .B(_07414_),
    .X(_07418_));
 sg13g2_and2_1 _15808_ (.A(_01577_),
    .B(_07418_),
    .X(_07419_));
 sg13g2_nand3_1 _15809_ (.B(_03195_),
    .C(_07419_),
    .A(_01466_),
    .Y(_07420_));
 sg13g2_and2_2 _15810_ (.A(_07417_),
    .B(_07420_),
    .X(_07421_));
 sg13g2_a21oi_1 _15811_ (.A1(net2102),
    .A2(net2104),
    .Y(_07422_),
    .B1(\id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ));
 sg13g2_o21ai_1 _15812_ (.B1(_07413_),
    .Y(_07423_),
    .A1(_07414_),
    .A2(_07422_));
 sg13g2_nand2b_1 _15813_ (.Y(_07424_),
    .B(_07423_),
    .A_N(_01488_));
 sg13g2_inv_1 _15814_ (.Y(_07425_),
    .A(\id_in_ready_$_AND__Y_A_$_AND__Y_A_$_AND__A_Y_$_AND__A_B ));
 sg13g2_or2_1 _15815_ (.X(_07426_),
    .B(_03193_),
    .A(_07425_));
 sg13g2_nor2_2 _15816_ (.A(_01577_),
    .B(_07426_),
    .Y(_07427_));
 sg13g2_a21oi_1 _15817_ (.A1(_03189_),
    .A2(_03184_),
    .Y(_07428_),
    .B1(_03849_));
 sg13g2_o21ai_1 _15818_ (.B1(_02865_),
    .Y(_07429_),
    .A1(_02863_),
    .A2(_07428_));
 sg13g2_and2_1 _15819_ (.A(_01601_),
    .B(_07429_),
    .X(_07430_));
 sg13g2_nand2_1 _15820_ (.Y(_07431_),
    .A(_01329_),
    .B(_07430_));
 sg13g2_and3_1 _15821_ (.X(\id_stage_i.controller_i.wfi_insn_i ),
    .A(_01449_),
    .B(_01450_),
    .C(_01585_));
 sg13g2_and4_1 _15822_ (.A(net436),
    .B(_01443_),
    .C(_01584_),
    .D(\id_stage_i.controller_i.wfi_insn_i ),
    .X(_07432_));
 sg13g2_o21ai_1 _15823_ (.B1(\id_stage_i.controller_i.enter_debug_mode_prio_q ),
    .Y(_07433_),
    .A1(_01455_),
    .A2(_03853_));
 sg13g2_and2_1 _15824_ (.A(net395),
    .B(_07433_),
    .X(_07434_));
 sg13g2_nand2b_1 _15825_ (.Y(_07435_),
    .B(_07434_),
    .A_N(_07432_));
 sg13g2_inv_1 _15826_ (.Y(_07436_),
    .A(_07435_));
 sg13g2_o21ai_1 _15827_ (.B1(_07413_),
    .Y(_07437_),
    .A1(_01476_),
    .A2(_01461_));
 sg13g2_nor2_1 _15828_ (.A(_03298_),
    .B(_07419_),
    .Y(_07438_));
 sg13g2_o21ai_1 _15829_ (.B1(_07438_),
    .Y(_07439_),
    .A1(net2104),
    .A2(_07437_));
 sg13g2_nor2_1 _15830_ (.A(_07436_),
    .B(_07439_),
    .Y(_07440_));
 sg13g2_o21ai_1 _15831_ (.B1(_07440_),
    .Y(_07441_),
    .A1(_07427_),
    .A2(_07431_));
 sg13g2_nand2_1 _15832_ (.Y(_07442_),
    .A(_07424_),
    .B(_07441_));
 sg13g2_o21ai_1 _15833_ (.B1(_07440_),
    .Y(_07443_),
    .A1(_01466_),
    .A2(_07426_));
 sg13g2_nand2_2 _15834_ (.Y(_07444_),
    .A(_07421_),
    .B(_07443_));
 sg13g2_a22oi_1 _15835_ (.Y(_00237_),
    .B1(_07444_),
    .B2(_01460_),
    .A2(_07442_),
    .A1(_07421_));
 sg13g2_nor2_1 _15836_ (.A(_01466_),
    .B(_07426_),
    .Y(_07445_));
 sg13g2_nor3_1 _15837_ (.A(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .B(_03186_),
    .C(_07445_),
    .Y(_07446_));
 sg13g2_nor2b_1 _15838_ (.A(_01466_),
    .B_N(_07419_),
    .Y(_07447_));
 sg13g2_a221oi_1 _15839_ (.B2(_07434_),
    .C1(_07447_),
    .B1(_07432_),
    .A1(_01460_),
    .Y(_07448_),
    .A2(_01496_));
 sg13g2_o21ai_1 _15840_ (.B1(_07448_),
    .Y(_07449_),
    .A1(net1715),
    .A2(_07446_));
 sg13g2_nand3_1 _15841_ (.B(_07430_),
    .C(_07448_),
    .A(_07427_),
    .Y(_07450_));
 sg13g2_nand4_1 _15842_ (.B(_07424_),
    .C(_07449_),
    .A(_07421_),
    .Y(_07451_),
    .D(_07450_));
 sg13g2_o21ai_1 _15843_ (.B1(_07451_),
    .Y(_00238_),
    .A1(_01476_),
    .A2(_07421_));
 sg13g2_inv_1 _15844_ (.Y(_07452_),
    .A(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ));
 sg13g2_o21ai_1 _15845_ (.B1(_07438_),
    .Y(_07453_),
    .A1(net2102),
    .A2(_07437_));
 sg13g2_a21oi_1 _15846_ (.A1(_01457_),
    .A2(_07436_),
    .Y(_07454_),
    .B1(_07453_));
 sg13g2_nand2b_1 _15847_ (.Y(_07455_),
    .B(_07454_),
    .A_N(_03186_));
 sg13g2_o21ai_1 _15848_ (.B1(_07420_),
    .Y(_07456_),
    .A1(_07445_),
    .A2(_07455_));
 sg13g2_inv_1 _15849_ (.Y(_07457_),
    .A(_07455_));
 sg13g2_o21ai_1 _15850_ (.B1(_07457_),
    .Y(_07458_),
    .A1(net1715),
    .A2(_07427_));
 sg13g2_nand3_1 _15851_ (.B(_07424_),
    .C(_07458_),
    .A(_07417_),
    .Y(_07459_));
 sg13g2_a22oi_1 _15852_ (.Y(_00239_),
    .B1(_07459_),
    .B2(_07420_),
    .A2(_07456_),
    .A1(_07452_));
 sg13g2_nand3_1 _15853_ (.B(_07427_),
    .C(_07430_),
    .A(_01329_),
    .Y(_07460_));
 sg13g2_inv_1 _15854_ (.Y(_07461_),
    .A(_01577_));
 sg13g2_nand2_1 _15855_ (.Y(_07462_),
    .A(_01457_),
    .B(_07433_));
 sg13g2_a22oi_1 _15856_ (.Y(_07463_),
    .B1(_07462_),
    .B2(_01582_),
    .A2(_07418_),
    .A1(_07461_));
 sg13g2_inv_1 _15857_ (.Y(_07464_),
    .A(_07424_));
 sg13g2_a21oi_1 _15858_ (.A1(_07460_),
    .A2(_07463_),
    .Y(_07465_),
    .B1(_07464_));
 sg13g2_mux2_1 _15859_ (.A0(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .A1(_07465_),
    .S(_07421_),
    .X(_00240_));
 sg13g2_a21oi_1 _15860_ (.A1(_01583_),
    .A2(_01588_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ),
    .B1(net395));
 sg13g2_nor2b_1 _15861_ (.A(net1984),
    .B_N(instr_rdata_i_16_),
    .Y(_07466_));
 sg13g2_a21oi_1 _15862_ (.A1(net1984),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16_ ),
    .Y(_07467_),
    .B1(_07466_));
 sg13g2_mux2_1 _15863_ (.A0(instr_rdata_i_0_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0_ ),
    .S(net1983),
    .X(_07468_));
 sg13g2_nor2_1 _15864_ (.A(net559),
    .B(_07468_),
    .Y(_07469_));
 sg13g2_a21oi_1 _15865_ (.A1(net558),
    .A2(_07467_),
    .Y(_07470_),
    .B1(_07469_));
 sg13g2_buf_8 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_4 fanout822 (.X(net822),
    .A(\register_file_i/_2932_ ));
 sg13g2_mux2_1 _15868_ (.A0(\id_stage_i.controller_i.instr_compressed_i_0_ ),
    .A1(net1537),
    .S(net762),
    .X(_00241_));
 sg13g2_mux2_1 _15869_ (.A0(instr_rdata_i_26_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_26_ ),
    .S(net1980),
    .X(_07473_));
 sg13g2_mux2_1 _15870_ (.A0(instr_rdata_i_10_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_10_ ),
    .S(net1978),
    .X(_07474_));
 sg13g2_inv_1 _15871_ (.Y(_07475_),
    .A(net557));
 sg13g2_mux2_1 _15872_ (.A0(_07473_),
    .A1(_07474_),
    .S(net1861),
    .X(_07476_));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(net822));
 sg13g2_mux2_1 _15874_ (.A0(\id_stage_i.controller_i.instr_compressed_i_10_ ),
    .A1(net394),
    .S(net763),
    .X(_00242_));
 sg13g2_mux2_1 _15875_ (.A0(instr_rdata_i_27_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_27_ ),
    .S(net1980),
    .X(_07478_));
 sg13g2_mux2_1 _15876_ (.A0(instr_rdata_i_11_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_11_ ),
    .S(net1978),
    .X(_07479_));
 sg13g2_mux2_1 _15877_ (.A0(_07478_),
    .A1(_07479_),
    .S(net1862),
    .X(_07480_));
 sg13g2_buf_4 fanout820 (.X(net820),
    .A(net822));
 sg13g2_mux2_1 _15879_ (.A0(\id_stage_i.controller_i.instr_compressed_i_11_ ),
    .A1(net391),
    .S(net757),
    .X(_00243_));
 sg13g2_nor2b_1 _15880_ (.A(net1982),
    .B_N(instr_rdata_i_28_),
    .Y(_07482_));
 sg13g2_a21oi_2 _15881_ (.B1(_07482_),
    .Y(_07483_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_28_ ),
    .A1(net1982));
 sg13g2_mux2_1 _15882_ (.A0(instr_rdata_i_12_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_12_ ),
    .S(net1979),
    .X(_07484_));
 sg13g2_nor2_1 _15883_ (.A(net558),
    .B(_07484_),
    .Y(_07485_));
 sg13g2_a21oi_2 _15884_ (.B1(_07485_),
    .Y(_07486_),
    .A2(_07483_),
    .A1(net557));
 sg13g2_buf_2 fanout819 (.A(\register_file_i/_2936_ ),
    .X(net819));
 sg13g2_buf_2 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_8 fanout817 (.A(net819),
    .X(net817));
 sg13g2_mux2_1 _15888_ (.A0(\id_stage_i.controller_i.instr_compressed_i_12_ ),
    .A1(net336),
    .S(net763),
    .X(_00244_));
 sg13g2_nor2b_1 _15889_ (.A(net1981),
    .B_N(instr_rdata_i_29_),
    .Y(_07490_));
 sg13g2_a21oi_2 _15890_ (.B1(_07490_),
    .Y(_07491_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_29_ ),
    .A1(net1981));
 sg13g2_mux2_1 _15891_ (.A0(instr_rdata_i_13_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_13_ ),
    .S(net1978),
    .X(_07492_));
 sg13g2_nor2_1 _15892_ (.A(net557),
    .B(_07492_),
    .Y(_07493_));
 sg13g2_a21oi_1 _15893_ (.A1(net558),
    .A2(_07491_),
    .Y(_07494_),
    .B1(_07493_));
 sg13g2_buf_4 fanout816 (.X(net816),
    .A(\register_file_i/_2936_ ));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(net816));
 sg13g2_mux2_1 _15896_ (.A0(\id_stage_i.controller_i.instr_compressed_i_13_ ),
    .A1(net1673),
    .S(net764),
    .X(_00245_));
 sg13g2_nor2b_1 _15897_ (.A(net1980),
    .B_N(instr_rdata_i_30_),
    .Y(_07497_));
 sg13g2_a21oi_2 _15898_ (.B1(_07497_),
    .Y(_07498_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_30_ ),
    .A1(net1980));
 sg13g2_mux2_1 _15899_ (.A0(instr_rdata_i_14_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_14_ ),
    .S(net1978),
    .X(_07499_));
 sg13g2_nor2_1 _15900_ (.A(net557),
    .B(_07499_),
    .Y(_07500_));
 sg13g2_a21oi_1 _15901_ (.A1(net557),
    .A2(_07498_),
    .Y(_07501_),
    .B1(_07500_));
 sg13g2_buf_4 fanout814 (.X(net814),
    .A(net816));
 sg13g2_buf_4 fanout813 (.X(net813),
    .A(\register_file_i/_2995_ ));
 sg13g2_mux2_1 _15904_ (.A0(\id_stage_i.controller_i.instr_compressed_i_14_ ),
    .A1(net1669),
    .S(net757),
    .X(_00246_));
 sg13g2_nor2b_1 _15905_ (.A(net1981),
    .B_N(instr_rdata_i_31_),
    .Y(_07504_));
 sg13g2_a21oi_2 _15906_ (.B1(_07504_),
    .Y(_07505_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_31_ ),
    .A1(net1981));
 sg13g2_mux2_1 _15907_ (.A0(instr_rdata_i_15_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_15_ ),
    .S(net1979),
    .X(_07506_));
 sg13g2_nor2_1 _15908_ (.A(net557),
    .B(_07506_),
    .Y(_07507_));
 sg13g2_a21oi_2 _15909_ (.B1(_07507_),
    .Y(_07508_),
    .A2(_07505_),
    .A1(net557));
 sg13g2_buf_4 fanout812 (.X(net812),
    .A(net813));
 sg13g2_mux2_1 _15911_ (.A0(\id_stage_i.controller_i.instr_compressed_i_15_ ),
    .A1(net1630),
    .S(net762),
    .X(_00247_));
 sg13g2_nor2b_1 _15912_ (.A(net1985),
    .B_N(instr_rdata_i_17_),
    .Y(_07510_));
 sg13g2_a21oi_2 _15913_ (.B1(_07510_),
    .Y(_07511_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17_ ),
    .A1(net1985));
 sg13g2_mux2_1 _15914_ (.A0(instr_rdata_i_1_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1_ ),
    .S(net1985),
    .X(_07512_));
 sg13g2_nor2_1 _15915_ (.A(net558),
    .B(_07512_),
    .Y(_07513_));
 sg13g2_a21oi_1 _15916_ (.A1(net559),
    .A2(_07511_),
    .Y(_07514_),
    .B1(_07513_));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(\register_file_i/_2995_ ));
 sg13g2_mux2_1 _15918_ (.A0(\id_stage_i.controller_i.instr_compressed_i_1_ ),
    .A1(net1530),
    .S(net764),
    .X(_00248_));
 sg13g2_mux2_1 _15919_ (.A0(instr_rdata_i_18_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_18_ ),
    .S(net1980),
    .X(_07516_));
 sg13g2_mux2_1 _15920_ (.A0(instr_rdata_i_2_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_2_ ),
    .S(net1978),
    .X(_07517_));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(net811));
 sg13g2_mux2_1 _15922_ (.A0(_07516_),
    .A1(_07517_),
    .S(net1862),
    .X(_07519_));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(net811));
 sg13g2_mux2_1 _15924_ (.A0(\id_stage_i.controller_i.instr_compressed_i_2_ ),
    .A1(net1610),
    .S(net765),
    .X(_00249_));
 sg13g2_mux2_1 _15925_ (.A0(instr_rdata_i_19_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_19_ ),
    .S(net1981),
    .X(_07521_));
 sg13g2_mux2_1 _15926_ (.A0(instr_rdata_i_3_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_3_ ),
    .S(net1978),
    .X(_07522_));
 sg13g2_mux2_2 _15927_ (.A0(_07521_),
    .A1(_07522_),
    .S(net1862),
    .X(_07523_));
 sg13g2_buf_2 fanout808 (.A(_06734_),
    .X(net808));
 sg13g2_mux2_1 _15929_ (.A0(\id_stage_i.controller_i.instr_compressed_i_3_ ),
    .A1(net1609),
    .S(net765),
    .X(_00250_));
 sg13g2_mux2_1 _15930_ (.A0(instr_rdata_i_20_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_20_ ),
    .S(net1981),
    .X(_07525_));
 sg13g2_mux2_1 _15931_ (.A0(instr_rdata_i_4_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_4_ ),
    .S(net1979),
    .X(_07526_));
 sg13g2_mux2_1 _15932_ (.A0(_07525_),
    .A1(_07526_),
    .S(net1862),
    .X(_07527_));
 sg13g2_buf_2 fanout807 (.A(rf_wdata_wb_9_),
    .X(net807));
 sg13g2_mux2_1 _15934_ (.A0(\id_stage_i.controller_i.instr_compressed_i_4_ ),
    .A1(net1607),
    .S(net757),
    .X(_00251_));
 sg13g2_mux2_1 _15935_ (.A0(instr_rdata_i_21_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_21_ ),
    .S(net1980),
    .X(_07529_));
 sg13g2_mux2_1 _15936_ (.A0(instr_rdata_i_5_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_5_ ),
    .S(net1978),
    .X(_07530_));
 sg13g2_mux2_1 _15937_ (.A0(_07529_),
    .A1(_07530_),
    .S(net1861),
    .X(_07531_));
 sg13g2_buf_2 fanout806 (.A(net807),
    .X(net806));
 sg13g2_mux2_1 _15939_ (.A0(\id_stage_i.controller_i.instr_compressed_i_5_ ),
    .A1(net1627),
    .S(net762),
    .X(_00252_));
 sg13g2_mux2_2 _15940_ (.A0(instr_rdata_i_22_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_22_ ),
    .S(net1980),
    .X(_07533_));
 sg13g2_mux2_1 _15941_ (.A0(instr_rdata_i_6_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_6_ ),
    .S(net1978),
    .X(_07534_));
 sg13g2_mux2_1 _15942_ (.A0(_07533_),
    .A1(_07534_),
    .S(net1861),
    .X(_07535_));
 sg13g2_buf_2 fanout805 (.A(rf_wdata_wb_9_),
    .X(net805));
 sg13g2_mux2_1 _15944_ (.A0(\id_stage_i.controller_i.instr_compressed_i_6_ ),
    .A1(net1625),
    .S(net762),
    .X(_00253_));
 sg13g2_mux4_1 _15945_ (.S0(net1985),
    .A0(instr_rdata_i_7_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_7_ ),
    .A2(instr_rdata_i_23_),
    .A3(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23_ ),
    .S1(crash_dump_o_65_),
    .X(_07537_));
 sg13g2_buf_2 fanout804 (.A(rf_wdata_wb_9_),
    .X(net804));
 sg13g2_buf_2 fanout803 (.A(rf_wdata_wb_12_),
    .X(net803));
 sg13g2_mux2_1 _15948_ (.A0(\id_stage_i.controller_i.instr_compressed_i_7_ ),
    .A1(net1662),
    .S(net762),
    .X(_00254_));
 sg13g2_mux2_1 _15949_ (.A0(instr_rdata_i_24_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_24_ ),
    .S(net1980),
    .X(_07540_));
 sg13g2_mux2_1 _15950_ (.A0(instr_rdata_i_8_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_8_ ),
    .S(net1979),
    .X(_07541_));
 sg13g2_mux2_1 _15951_ (.A0(_07540_),
    .A1(_07541_),
    .S(net1862),
    .X(_07542_));
 sg13g2_buf_2 fanout802 (.A(net803),
    .X(net802));
 sg13g2_mux2_1 _15953_ (.A0(\id_stage_i.controller_i.instr_compressed_i_8_ ),
    .A1(net386),
    .S(net769),
    .X(_00255_));
 sg13g2_mux2_1 _15954_ (.A0(instr_rdata_i_25_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_25_ ),
    .S(net1981),
    .X(_07544_));
 sg13g2_mux2_1 _15955_ (.A0(instr_rdata_i_9_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_9_ ),
    .S(net1979),
    .X(_07545_));
 sg13g2_mux2_2 _15956_ (.A0(_07544_),
    .A1(_07545_),
    .S(net1862),
    .X(_07546_));
 sg13g2_mux2_1 _15957_ (.A0(\id_stage_i.controller_i.instr_compressed_i_9_ ),
    .A1(net1661),
    .S(net758),
    .X(_00256_));
 sg13g2_buf_2 fanout801 (.A(net803),
    .X(net801));
 sg13g2_buf_2 fanout800 (.A(net803),
    .X(net800));
 sg13g2_buf_2 fanout799 (.A(net800),
    .X(net799));
 sg13g2_nor3_1 _15961_ (.A(instr_err_i),
    .B(net434),
    .C(_01513_),
    .Y(_07550_));
 sg13g2_nor3_1 _15962_ (.A(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ),
    .B(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ),
    .C(_01472_),
    .Y(_07551_));
 sg13g2_nand2_1 _15963_ (.Y(_07552_),
    .A(_01512_),
    .B(_01472_));
 sg13g2_a221oi_1 _15964_ (.B2(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ),
    .C1(_01517_),
    .B1(_07552_),
    .A1(_01472_),
    .Y(_07553_),
    .A2(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_0_ ));
 sg13g2_nor4_1 _15965_ (.A(net1864),
    .B(_07550_),
    .C(_07551_),
    .D(_07553_),
    .Y(_07554_));
 sg13g2_a21oi_2 _15966_ (.B1(_07554_),
    .Y(_07555_),
    .A2(_01514_),
    .A1(net1863));
 sg13g2_nor2_2 _15967_ (.A(\id_stage_i.controller_i.instr_fetch_err_i ),
    .B(net767),
    .Y(_07556_));
 sg13g2_a21oi_1 _15968_ (.A1(net767),
    .A2(_07555_),
    .Y(_00257_),
    .B1(_07556_));
 sg13g2_inv_1 _15969_ (.Y(_07557_),
    .A(\id_stage_i.controller_i.instr_fetch_err_plus2_i ));
 sg13g2_buf_2 fanout798 (.A(rf_wdata_wb_10_),
    .X(net798));
 sg13g2_nor2b_1 _15971_ (.A(net435),
    .B_N(instr_err_i),
    .Y(_07559_));
 sg13g2_a22oi_1 _15972_ (.Y(_07560_),
    .B1(_07559_),
    .B2(net1983),
    .A2(net435),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ));
 sg13g2_inv_1 _15973_ (.Y(_07561_),
    .A(_07560_));
 sg13g2_nand4_1 _15974_ (.B(\if_stage_i.prefetch_buffer_i.fifo_i.err_plus2_$_AND__Y_B ),
    .C(net768),
    .A(net560),
    .Y(_07562_),
    .D(_07561_));
 sg13g2_o21ai_1 _15975_ (.B1(_07562_),
    .Y(_00258_),
    .A1(_07557_),
    .A2(net768));
 sg13g2_a21o_1 _15976_ (.A2(_07467_),
    .A1(net560),
    .B1(_07469_),
    .X(_07563_));
 sg13g2_buf_2 fanout797 (.A(net798),
    .X(net797));
 sg13g2_buf_2 fanout796 (.A(rf_wdata_wb_10_),
    .X(net796));
 sg13g2_a21o_1 _15979_ (.A2(_07511_),
    .A1(net560),
    .B1(_07513_),
    .X(_07566_));
 sg13g2_nand2_2 _15980_ (.Y(_07567_),
    .A(net1633),
    .B(net1524));
 sg13g2_a21o_1 _15981_ (.A2(_07491_),
    .A1(net560),
    .B1(_07493_),
    .X(_07568_));
 sg13g2_buf_2 fanout795 (.A(rf_wdata_wb_10_),
    .X(net795));
 sg13g2_buf_8 fanout794 (.A(rf_wdata_wb_11_),
    .X(net794));
 sg13g2_o21ai_1 _15984_ (.B1(net1658),
    .Y(_07571_),
    .A1(net1665),
    .A2(_07567_));
 sg13g2_nand2_1 _15985_ (.Y(_07572_),
    .A(net1527),
    .B(_07571_));
 sg13g2_mux2_1 _15986_ (.A0(\id_stage_i.controller_i.instr_i_0_ ),
    .A1(_07572_),
    .S(net765),
    .X(_00259_));
 sg13g2_buf_8 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_8 fanout792 (.A(net794),
    .X(net792));
 sg13g2_a21o_1 _15989_ (.A2(_07505_),
    .A1(net560),
    .B1(_07507_),
    .X(_07575_));
 sg13g2_nor2_2 _15990_ (.A(net1668),
    .B(net1623),
    .Y(_07576_));
 sg13g2_nor2_1 _15991_ (.A(net1526),
    .B(net1670),
    .Y(_07577_));
 sg13g2_inv_2 _15992_ (.Y(_07578_),
    .A(net392));
 sg13g2_buf_8 fanout791 (.A(net794),
    .X(net791));
 sg13g2_nand2_2 _15994_ (.Y(_07580_),
    .A(net1659),
    .B(net1623));
 sg13g2_a21oi_1 _15995_ (.A1(_07578_),
    .A2(_07580_),
    .Y(_07581_),
    .B1(net1536));
 sg13g2_a21o_1 _15996_ (.A2(_07577_),
    .A1(_07576_),
    .B1(_07581_),
    .X(_07582_));
 sg13g2_nor2_2 _15997_ (.A(net1672),
    .B(net1666),
    .Y(_07583_));
 sg13g2_or2_1 _15998_ (.X(_07584_),
    .B(net1625),
    .A(net1627));
 sg13g2_nor4_2 _15999_ (.A(net1610),
    .B(net1609),
    .C(net1607),
    .Y(_07585_),
    .D(_07584_));
 sg13g2_a21o_1 _16000_ (.A2(_07498_),
    .A1(net560),
    .B1(_07500_),
    .X(_07586_));
 sg13g2_nand2_2 _16001_ (.Y(_07587_),
    .A(net1658),
    .B(net388));
 sg13g2_nor2_2 _16002_ (.A(net1623),
    .B(_07587_),
    .Y(_07588_));
 sg13g2_and2_2 _16003_ (.A(_07585_),
    .B(_07588_),
    .X(_07589_));
 sg13g2_nand2_2 _16004_ (.Y(_07590_),
    .A(net1528),
    .B(net1530));
 sg13g2_a21oi_1 _16005_ (.A1(_07583_),
    .A2(_07589_),
    .Y(_07591_),
    .B1(_07590_));
 sg13g2_nor2_2 _16006_ (.A(net1656),
    .B(net1664),
    .Y(_07592_));
 sg13g2_buf_8 fanout790 (.A(net794),
    .X(net790));
 sg13g2_buf_2 fanout789 (.A(rf_wdata_wb_13_),
    .X(net789));
 sg13g2_nand2_1 _16009_ (.Y(_07595_),
    .A(net1533),
    .B(net394));
 sg13g2_a21oi_1 _16010_ (.A1(net1523),
    .A2(net1606),
    .Y(_07596_),
    .B1(_07595_));
 sg13g2_a221oi_1 _16011_ (.B2(net392),
    .C1(_07596_),
    .B1(_07591_),
    .A1(net1523),
    .Y(_07597_),
    .A2(_07582_));
 sg13g2_nor2_2 _16012_ (.A(net2099),
    .B(net763),
    .Y(_07598_));
 sg13g2_a21oi_1 _16013_ (.A1(net763),
    .A2(_07597_),
    .Y(_00260_),
    .B1(_07598_));
 sg13g2_buf_2 fanout788 (.A(rf_wdata_wb_13_),
    .X(net788));
 sg13g2_and2_2 _16015_ (.A(net392),
    .B(net391),
    .X(_07600_));
 sg13g2_nand2_2 _16016_ (.Y(_07601_),
    .A(net335),
    .B(_07600_));
 sg13g2_a21oi_1 _16017_ (.A1(net1629),
    .A2(_07601_),
    .Y(_07602_),
    .B1(net1670));
 sg13g2_buf_2 fanout787 (.A(rf_wdata_wb_13_),
    .X(net787));
 sg13g2_nand2_2 _16019_ (.Y(_07604_),
    .A(net389),
    .B(net1524));
 sg13g2_nor2_1 _16020_ (.A(_07602_),
    .B(_07604_),
    .Y(_07605_));
 sg13g2_nor2_1 _16021_ (.A(net1526),
    .B(_07605_),
    .Y(_07606_));
 sg13g2_buf_8 fanout786 (.A(net787),
    .X(net786));
 sg13g2_nor2_2 _16023_ (.A(net1671),
    .B(net1630),
    .Y(_07608_));
 sg13g2_nor3_1 _16024_ (.A(net1533),
    .B(net1529),
    .C(_07608_),
    .Y(_07609_));
 sg13g2_nor3_1 _16025_ (.A(_07591_),
    .B(_07606_),
    .C(_07609_),
    .Y(_07610_));
 sg13g2_nor2b_1 _16026_ (.A(_07610_),
    .B_N(net391),
    .Y(_07611_));
 sg13g2_mux2_1 _16027_ (.A0(net553),
    .A1(_07611_),
    .S(net758),
    .X(_00261_));
 sg13g2_nor2_2 _16028_ (.A(net1535),
    .B(net1522),
    .Y(_07612_));
 sg13g2_buf_8 fanout785 (.A(net787),
    .X(net785));
 sg13g2_nor2_2 _16030_ (.A(net1630),
    .B(_07587_),
    .Y(_07614_));
 sg13g2_a21oi_1 _16031_ (.A1(net1523),
    .A2(_07576_),
    .Y(_07615_),
    .B1(net1670));
 sg13g2_nand2_1 _16032_ (.Y(_07616_),
    .A(net1533),
    .B(net1529));
 sg13g2_o21ai_1 _16033_ (.B1(_07616_),
    .Y(_07617_),
    .A1(net1534),
    .A2(_07615_));
 sg13g2_nor4_1 _16034_ (.A(net392),
    .B(net390),
    .C(net1662),
    .D(net1661),
    .Y(_07618_));
 sg13g2_and2_1 _16035_ (.A(net385),
    .B(_07618_),
    .X(_07619_));
 sg13g2_buf_2 fanout784 (.A(rf_wdata_wb_15_),
    .X(net784));
 sg13g2_nor3_2 _16037_ (.A(net1659),
    .B(net388),
    .C(net1632),
    .Y(_07621_));
 sg13g2_nor2b_2 _16038_ (.A(_07619_),
    .B_N(_07621_),
    .Y(_07622_));
 sg13g2_buf_2 fanout783 (.A(net784),
    .X(net783));
 sg13g2_nand2_1 _16040_ (.Y(_07624_),
    .A(net1627),
    .B(net1625));
 sg13g2_a21oi_1 _16041_ (.A1(_07600_),
    .A2(_07624_),
    .Y(_07625_),
    .B1(net1670));
 sg13g2_o21ai_1 _16042_ (.B1(_07580_),
    .Y(_07626_),
    .A1(net334),
    .A2(_07625_));
 sg13g2_nand3_1 _16043_ (.B(net1664),
    .C(net1629),
    .A(net1670),
    .Y(_07627_));
 sg13g2_o21ai_1 _16044_ (.B1(_07627_),
    .Y(_07628_),
    .A1(net1664),
    .A2(_07626_));
 sg13g2_a21oi_1 _16045_ (.A1(net1610),
    .A2(_07622_),
    .Y(_07629_),
    .B1(_07628_));
 sg13g2_nand2_2 _16046_ (.Y(_07630_),
    .A(net1533),
    .B(net1523));
 sg13g2_nor2_1 _16047_ (.A(_07630_),
    .B(_07614_),
    .Y(_07631_));
 sg13g2_nor2b_1 _16048_ (.A(_07629_),
    .B_N(_07631_),
    .Y(_07632_));
 sg13g2_a221oi_1 _16049_ (.B2(net335),
    .C1(_07632_),
    .B1(_07617_),
    .A1(_07612_),
    .Y(_07633_),
    .A2(_07614_));
 sg13g2_nor2_2 _16050_ (.A(net2097),
    .B(net761),
    .Y(_07634_));
 sg13g2_a21oi_2 _16051_ (.B1(_07634_),
    .Y(_00262_),
    .A2(_07633_),
    .A1(net761));
 sg13g2_nand3_1 _16052_ (.B(net1609),
    .C(_07622_),
    .A(net1522),
    .Y(_07635_));
 sg13g2_and2_1 _16053_ (.A(net390),
    .B(_07588_),
    .X(_07636_));
 sg13g2_a21o_1 _16054_ (.A2(_07483_),
    .A1(net560),
    .B1(_07485_),
    .X(_07637_));
 sg13g2_buf_2 fanout782 (.A(net784),
    .X(net782));
 sg13g2_a21oi_1 _16056_ (.A1(net1604),
    .A2(net1626),
    .Y(_07639_),
    .B1(_07578_));
 sg13g2_nor2_1 _16057_ (.A(net1530),
    .B(_07639_),
    .Y(_07640_));
 sg13g2_buf_2 fanout781 (.A(net784),
    .X(net781));
 sg13g2_buf_2 fanout780 (.A(net784),
    .X(net780));
 sg13g2_o21ai_1 _16060_ (.B1(net1525),
    .Y(_07643_),
    .A1(net1605),
    .A2(net1668));
 sg13g2_a221oi_1 _16061_ (.B2(net1673),
    .C1(net1527),
    .B1(_07643_),
    .A1(_07636_),
    .Y(_07644_),
    .A2(_07640_));
 sg13g2_nand2_1 _16062_ (.Y(_07645_),
    .A(net1536),
    .B(net1633));
 sg13g2_a22oi_1 _16063_ (.Y(_07646_),
    .B1(_07645_),
    .B2(_07583_),
    .A2(_07644_),
    .A1(_07635_));
 sg13g2_mux2_1 _16064_ (.A0(net551),
    .A1(_07646_),
    .S(net761),
    .X(_00263_));
 sg13g2_nand2_2 _16065_ (.Y(_07647_),
    .A(net393),
    .B(net390));
 sg13g2_a21oi_1 _16066_ (.A1(net1605),
    .A2(_07584_),
    .Y(_07648_),
    .B1(_07647_));
 sg13g2_nand2_1 _16067_ (.Y(_07649_),
    .A(net1607),
    .B(_07622_));
 sg13g2_o21ai_1 _16068_ (.B1(_07649_),
    .Y(_07650_),
    .A1(_07587_),
    .A2(_07648_));
 sg13g2_nor3_1 _16069_ (.A(net1603),
    .B(net1656),
    .C(_07604_),
    .Y(_07651_));
 sg13g2_a21oi_1 _16070_ (.A1(net1664),
    .A2(net1529),
    .Y(_07652_),
    .B1(_07651_));
 sg13g2_a21oi_1 _16071_ (.A1(net1670),
    .A2(net1664),
    .Y(_07653_),
    .B1(net1533));
 sg13g2_a21oi_1 _16072_ (.A1(net1533),
    .A2(_07652_),
    .Y(_07654_),
    .B1(_07653_));
 sg13g2_a21oi_2 _16073_ (.B1(_07654_),
    .Y(_07655_),
    .A2(_07650_),
    .A1(_07631_));
 sg13g2_nor2_2 _16074_ (.A(net2089),
    .B(net759),
    .Y(_07656_));
 sg13g2_a21oi_2 _16075_ (.B1(_07656_),
    .Y(_00264_),
    .A2(_07655_),
    .A1(net760));
 sg13g2_buf_8 fanout779 (.A(_03196_),
    .X(net779));
 sg13g2_nand2_1 _16077_ (.Y(_07658_),
    .A(net1656),
    .B(_07647_));
 sg13g2_a22oi_1 _16078_ (.Y(_07659_),
    .B1(_07658_),
    .B2(net336),
    .A2(net1662),
    .A1(net1656));
 sg13g2_nand3_1 _16079_ (.B(net1629),
    .C(net1662),
    .A(net1664),
    .Y(_07660_));
 sg13g2_o21ai_1 _16080_ (.B1(_07660_),
    .Y(_07661_),
    .A1(net1664),
    .A2(_07659_));
 sg13g2_a21oi_1 _16081_ (.A1(net1627),
    .A2(_07622_),
    .Y(_07662_),
    .B1(_07661_));
 sg13g2_nand2_2 _16082_ (.Y(_07663_),
    .A(net1624),
    .B(_07583_));
 sg13g2_nor2_1 _16083_ (.A(net1526),
    .B(net1529),
    .Y(_07664_));
 sg13g2_buf_8 fanout778 (.A(_03196_),
    .X(net778));
 sg13g2_o21ai_1 _16085_ (.B1(net1426),
    .Y(_07666_),
    .A1(net1662),
    .A2(_07663_));
 sg13g2_nor2_2 _16086_ (.A(net1536),
    .B(net1672),
    .Y(_07667_));
 sg13g2_nor3_1 _16087_ (.A(net334),
    .B(net1624),
    .C(_07585_),
    .Y(_07668_));
 sg13g2_nor2_2 _16088_ (.A(_07587_),
    .B(_07668_),
    .Y(_07669_));
 sg13g2_nand3_1 _16089_ (.B(net1662),
    .C(_07669_),
    .A(net1526),
    .Y(_07670_));
 sg13g2_o21ai_1 _16090_ (.B1(_07670_),
    .Y(_07671_),
    .A1(net1623),
    .A2(_07667_));
 sg13g2_nor2_2 _16091_ (.A(net1672),
    .B(net388),
    .Y(_07672_));
 sg13g2_nor2_1 _16092_ (.A(net1623),
    .B(net1622),
    .Y(_07673_));
 sg13g2_a21oi_1 _16093_ (.A1(net1662),
    .A2(net1622),
    .Y(_07674_),
    .B1(_07673_));
 sg13g2_nor3_1 _16094_ (.A(net1534),
    .B(net1529),
    .C(_07674_),
    .Y(_07675_));
 sg13g2_a21oi_1 _16095_ (.A1(net1529),
    .A2(_07671_),
    .Y(_07676_),
    .B1(_07675_));
 sg13g2_o21ai_1 _16096_ (.B1(_07676_),
    .Y(_07677_),
    .A1(_07662_),
    .A2(_07666_));
 sg13g2_mux2_1 _16097_ (.A0(net2050),
    .A1(_07677_),
    .S(net763),
    .X(_00265_));
 sg13g2_nand2_2 _16098_ (.Y(_07678_),
    .A(net1666),
    .B(net1624));
 sg13g2_inv_1 _16099_ (.Y(_07679_),
    .A(_07678_));
 sg13g2_o21ai_1 _16100_ (.B1(_07679_),
    .Y(_07680_),
    .A1(net1626),
    .A2(net333));
 sg13g2_o21ai_1 _16101_ (.B1(_07680_),
    .Y(_07681_),
    .A1(net1604),
    .A2(net1667));
 sg13g2_nor2_1 _16102_ (.A(net1603),
    .B(_07647_),
    .Y(_07682_));
 sg13g2_mux2_1 _16103_ (.A0(instr_rdata_i_0_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_32_ ),
    .S(net431),
    .X(_07683_));
 sg13g2_nor2_1 _16104_ (.A(net1863),
    .B(_07683_),
    .Y(_07684_));
 sg13g2_a21oi_1 _16105_ (.A1(net1863),
    .A2(_07467_),
    .Y(_07685_),
    .B1(_07684_));
 sg13g2_and2_1 _16106_ (.A(_07583_),
    .B(_07685_),
    .X(_07686_));
 sg13g2_a22oi_1 _16107_ (.Y(_07687_),
    .B1(net296),
    .B2(_07686_),
    .A2(net386),
    .A1(net1667));
 sg13g2_nand2_1 _16108_ (.Y(_07688_),
    .A(net1633),
    .B(net296));
 sg13g2_nand3_1 _16109_ (.B(_07583_),
    .C(_07688_),
    .A(net386),
    .Y(_07689_));
 sg13g2_o21ai_1 _16110_ (.B1(_07689_),
    .Y(_07690_),
    .A1(net1624),
    .A2(_07687_));
 sg13g2_a21oi_1 _16111_ (.A1(net1672),
    .A2(_07681_),
    .Y(_07691_),
    .B1(_07690_));
 sg13g2_nand2_2 _16112_ (.Y(_07692_),
    .A(net388),
    .B(net1629));
 sg13g2_nand2_2 _16113_ (.Y(_07693_),
    .A(net1656),
    .B(_07692_));
 sg13g2_nor2_2 _16114_ (.A(net1536),
    .B(net1530),
    .Y(_07694_));
 sg13g2_nor2_2 _16115_ (.A(net1528),
    .B(net1524),
    .Y(_07695_));
 sg13g2_a21o_1 _16116_ (.A2(_07694_),
    .A1(net1563),
    .B1(_07695_),
    .X(_07696_));
 sg13g2_nand2_1 _16117_ (.Y(_07697_),
    .A(net1660),
    .B(net1667));
 sg13g2_nand2_1 _16118_ (.Y(_07698_),
    .A(net385),
    .B(_07669_));
 sg13g2_a21oi_1 _16119_ (.A1(net1672),
    .A2(_07685_),
    .Y(_07699_),
    .B1(net1524));
 sg13g2_nand3_1 _16120_ (.B(_07698_),
    .C(_07699_),
    .A(_07697_),
    .Y(_07700_));
 sg13g2_nor2_1 _16121_ (.A(net1622),
    .B(net1563),
    .Y(_07701_));
 sg13g2_a21oi_1 _16122_ (.A1(net385),
    .A2(net1622),
    .Y(_07702_),
    .B1(_07701_));
 sg13g2_a21oi_1 _16123_ (.A1(net1525),
    .A2(_07702_),
    .Y(_07703_),
    .B1(net1537));
 sg13g2_a22oi_1 _16124_ (.Y(_07704_),
    .B1(_07700_),
    .B2(_07703_),
    .A2(_07696_),
    .A1(_07685_));
 sg13g2_o21ai_1 _16125_ (.B1(_07704_),
    .Y(_07705_),
    .A1(_07630_),
    .A2(_07691_));
 sg13g2_mux2_1 _16126_ (.A0(net536),
    .A1(_07705_),
    .S(net757),
    .X(_00266_));
 sg13g2_inv_1 _16127_ (.Y(_07706_),
    .A(net1661));
 sg13g2_mux2_1 _16128_ (.A0(instr_rdata_i_1_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_33_ ),
    .S(net430),
    .X(_07707_));
 sg13g2_nor2_1 _16129_ (.A(net1863),
    .B(_07707_),
    .Y(_07708_));
 sg13g2_a21oi_2 _16130_ (.B1(_07708_),
    .Y(_07709_),
    .A2(_07511_),
    .A1(net1863));
 sg13g2_nand2_1 _16131_ (.Y(_07710_),
    .A(net296),
    .B(_07709_));
 sg13g2_o21ai_1 _16132_ (.B1(_07710_),
    .Y(_07711_),
    .A1(_07706_),
    .A2(net296));
 sg13g2_nor2_1 _16133_ (.A(net1606),
    .B(_07622_),
    .Y(_07712_));
 sg13g2_nor2_2 _16134_ (.A(net1604),
    .B(_07712_),
    .Y(_07713_));
 sg13g2_a21oi_1 _16135_ (.A1(_07588_),
    .A2(_07711_),
    .Y(_07714_),
    .B1(_07713_));
 sg13g2_nor2_2 _16136_ (.A(net388),
    .B(net1623),
    .Y(_07715_));
 sg13g2_o21ai_1 _16137_ (.B1(net1661),
    .Y(_07716_),
    .A1(_07614_),
    .A2(_07715_));
 sg13g2_o21ai_1 _16138_ (.B1(_07716_),
    .Y(_07717_),
    .A1(_07614_),
    .A2(_07714_));
 sg13g2_a21oi_1 _16139_ (.A1(net1661),
    .A2(net1622),
    .Y(_07718_),
    .B1(net1531));
 sg13g2_a21oi_1 _16140_ (.A1(net1528),
    .A2(net1563),
    .Y(_07719_),
    .B1(net1530));
 sg13g2_nand2b_1 _16141_ (.Y(_07720_),
    .B(_07709_),
    .A_N(_07719_));
 sg13g2_o21ai_1 _16142_ (.B1(_07720_),
    .Y(_07721_),
    .A1(net1536),
    .A2(_07718_));
 sg13g2_a221oi_1 _16143_ (.B2(net1672),
    .C1(_07590_),
    .B1(_07709_),
    .A1(net1661),
    .Y(_07722_),
    .A2(_07669_));
 sg13g2_inv_1 _16144_ (.Y(_07723_),
    .A(_07722_));
 sg13g2_a22oi_1 _16145_ (.Y(_07724_),
    .B1(_07721_),
    .B2(_07723_),
    .A2(_07717_),
    .A1(net1427));
 sg13g2_buf_16 fanout777 (.X(net777),
    .A(net778));
 sg13g2_nor2_2 _16147_ (.A(net525),
    .B(net757),
    .Y(_07726_));
 sg13g2_a21oi_2 _16148_ (.B1(_07726_),
    .Y(_00267_),
    .A2(_07724_),
    .A1(net757));
 sg13g2_mux2_1 _16149_ (.A0(instr_rdata_i_2_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_34_ ),
    .S(net432),
    .X(_07727_));
 sg13g2_mux2_2 _16150_ (.A0(_07516_),
    .A1(_07727_),
    .S(net559),
    .X(_07728_));
 sg13g2_nand3_1 _16151_ (.B(net391),
    .C(net334),
    .A(net393),
    .Y(_07729_));
 sg13g2_nor3_1 _16152_ (.A(net1624),
    .B(_07728_),
    .C(_07729_),
    .Y(_07730_));
 sg13g2_o21ai_1 _16153_ (.B1(net389),
    .Y(_07731_),
    .A1(net1671),
    .A2(_07730_));
 sg13g2_a21oi_1 _16154_ (.A1(_07678_),
    .A2(_07731_),
    .Y(_07732_),
    .B1(_07713_));
 sg13g2_o21ai_1 _16155_ (.B1(net1427),
    .Y(_07733_),
    .A1(net392),
    .A2(_07663_));
 sg13g2_nor2_1 _16156_ (.A(_07578_),
    .B(_07590_),
    .Y(_07734_));
 sg13g2_nand2_1 _16157_ (.Y(_07735_),
    .A(net1660),
    .B(_07567_));
 sg13g2_a22oi_1 _16158_ (.Y(_07736_),
    .B1(_07728_),
    .B2(_07735_),
    .A2(net1622),
    .A1(net1524));
 sg13g2_nor2_1 _16159_ (.A(net1537),
    .B(_07736_),
    .Y(_07737_));
 sg13g2_a221oi_1 _16160_ (.B2(_07669_),
    .C1(_07737_),
    .B1(_07734_),
    .A1(_07695_),
    .Y(_07738_),
    .A2(_07728_));
 sg13g2_o21ai_1 _16161_ (.B1(_07738_),
    .Y(_07739_),
    .A1(_07732_),
    .A2(_07733_));
 sg13g2_mux2_1 _16162_ (.A0(net2009),
    .A1(_07739_),
    .S(net758),
    .X(_00268_));
 sg13g2_a21oi_1 _16163_ (.A1(net1534),
    .A2(net296),
    .Y(_07740_),
    .B1(_07694_));
 sg13g2_nor2_1 _16164_ (.A(_07692_),
    .B(_07740_),
    .Y(_07741_));
 sg13g2_o21ai_1 _16165_ (.B1(_07616_),
    .Y(_07742_),
    .A1(net1533),
    .A2(net1656));
 sg13g2_mux2_1 _16166_ (.A0(instr_rdata_i_3_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_35_ ),
    .S(net432),
    .X(_07743_));
 sg13g2_mux2_2 _16167_ (.A0(_07521_),
    .A1(_07743_),
    .S(net559),
    .X(_07744_));
 sg13g2_o21ai_1 _16168_ (.B1(_07744_),
    .Y(_07745_),
    .A1(_07741_),
    .A2(_07742_));
 sg13g2_o21ai_1 _16169_ (.B1(net1668),
    .Y(_07746_),
    .A1(net1629),
    .A2(net333));
 sg13g2_nand4_1 _16170_ (.B(net1670),
    .C(net1426),
    .A(net336),
    .Y(_07747_),
    .D(_07746_));
 sg13g2_a22oi_1 _16171_ (.Y(_07748_),
    .B1(_07669_),
    .B2(_07612_),
    .A2(_07614_),
    .A1(net1426));
 sg13g2_nand2b_1 _16172_ (.Y(_07749_),
    .B(net390),
    .A_N(_07748_));
 sg13g2_nand3_1 _16173_ (.B(_07747_),
    .C(_07749_),
    .A(_07745_),
    .Y(_07750_));
 sg13g2_mux2_1 _16174_ (.A0(\id_stage_i.controller_i.instr_i_19_ ),
    .A1(_07750_),
    .S(net762),
    .X(_00269_));
 sg13g2_buf_16 fanout776 (.X(net776),
    .A(net777));
 sg13g2_o21ai_1 _16176_ (.B1(net1535),
    .Y(_07752_),
    .A1(net1673),
    .A2(_07729_));
 sg13g2_nand4_1 _16177_ (.B(net1522),
    .C(net1564),
    .A(net764),
    .Y(_07753_),
    .D(_07752_));
 sg13g2_o21ai_1 _16178_ (.B1(_07753_),
    .Y(_07754_),
    .A1(\id_stage_i.controller_i.instr_i_1_ ),
    .A2(net766));
 sg13g2_inv_1 _16179_ (.Y(_00270_),
    .A(_07754_));
 sg13g2_nand2_2 _16180_ (.Y(_07755_),
    .A(net1528),
    .B(net1659));
 sg13g2_mux2_1 _16181_ (.A0(instr_rdata_i_4_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_36_ ),
    .S(net430),
    .X(_07756_));
 sg13g2_mux2_1 _16182_ (.A0(_07525_),
    .A1(_07756_),
    .S(net558),
    .X(_07757_));
 sg13g2_nand2b_1 _16183_ (.Y(_07758_),
    .B(_07618_),
    .A_N(net385));
 sg13g2_nor2_1 _16184_ (.A(net1603),
    .B(_07758_),
    .Y(_07759_));
 sg13g2_a22oi_1 _16185_ (.Y(_07760_),
    .B1(_07759_),
    .B2(_07589_),
    .A2(_07678_),
    .A1(net1610));
 sg13g2_nor3_1 _16186_ (.A(net1666),
    .B(net1632),
    .C(net1611),
    .Y(_07761_));
 sg13g2_nor3_1 _16187_ (.A(_07755_),
    .B(_07760_),
    .C(_07761_),
    .Y(_07762_));
 sg13g2_a21oi_1 _16188_ (.A1(_07755_),
    .A2(_07757_),
    .Y(_07763_),
    .B1(_07762_));
 sg13g2_nand2_1 _16189_ (.Y(_07764_),
    .A(net1563),
    .B(_07757_));
 sg13g2_nand3_1 _16190_ (.B(net1611),
    .C(net1622),
    .A(net1632),
    .Y(_07765_));
 sg13g2_a21oi_1 _16191_ (.A1(_07764_),
    .A2(_07765_),
    .Y(_07766_),
    .B1(net1536));
 sg13g2_nand2_1 _16192_ (.Y(_07767_),
    .A(net1624),
    .B(net1610));
 sg13g2_and2_1 _16193_ (.A(net296),
    .B(_07757_),
    .X(_07768_));
 sg13g2_a21oi_1 _16194_ (.A1(net1611),
    .A2(_07601_),
    .Y(_07769_),
    .B1(_07768_));
 sg13g2_a221oi_1 _16195_ (.B2(net1633),
    .C1(net1672),
    .B1(_07769_),
    .A1(net1666),
    .Y(_07770_),
    .A2(_07767_));
 sg13g2_nor2_1 _16196_ (.A(_07713_),
    .B(_07770_),
    .Y(_07771_));
 sg13g2_nor2_1 _16197_ (.A(net1611),
    .B(_07663_),
    .Y(_07772_));
 sg13g2_nor3_1 _16198_ (.A(net1528),
    .B(_07771_),
    .C(_07772_),
    .Y(_07773_));
 sg13g2_nor3_1 _16199_ (.A(net1531),
    .B(_07766_),
    .C(_07773_),
    .Y(_07774_));
 sg13g2_a21oi_2 _16200_ (.B1(_07774_),
    .Y(_07775_),
    .A2(_07763_),
    .A1(net1531));
 sg13g2_mux2_1 _16201_ (.A0(net513),
    .A1(_07775_),
    .S(net764),
    .X(_00271_));
 sg13g2_mux2_1 _16202_ (.A0(instr_rdata_i_5_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_37_ ),
    .S(net431),
    .X(_07776_));
 sg13g2_mux2_1 _16203_ (.A0(_07529_),
    .A1(_07776_),
    .S(net559),
    .X(_07777_));
 sg13g2_nor2_1 _16204_ (.A(net1672),
    .B(_07601_),
    .Y(_07778_));
 sg13g2_o21ai_1 _16205_ (.B1(_07580_),
    .Y(_07779_),
    .A1(net1666),
    .A2(_07778_));
 sg13g2_nand2b_1 _16206_ (.Y(_07780_),
    .B(_07621_),
    .A_N(net333));
 sg13g2_nand3_1 _16207_ (.B(_07600_),
    .C(_07777_),
    .A(_07588_),
    .Y(_07781_));
 sg13g2_o21ai_1 _16208_ (.B1(net336),
    .Y(_07782_),
    .A1(_07523_),
    .A2(_07663_));
 sg13g2_a21oi_1 _16209_ (.A1(_07780_),
    .A2(_07781_),
    .Y(_07783_),
    .B1(_07782_));
 sg13g2_a21o_1 _16210_ (.A2(_07779_),
    .A1(_07523_),
    .B1(_07783_),
    .X(_07784_));
 sg13g2_and4_1 _16211_ (.A(_07523_),
    .B(_07604_),
    .C(_07667_),
    .D(_07678_),
    .X(_07785_));
 sg13g2_a221oi_1 _16212_ (.B2(net1427),
    .C1(_07785_),
    .B1(_07784_),
    .A1(_07617_),
    .Y(_07786_),
    .A2(_07777_));
 sg13g2_nor2_1 _16213_ (.A(net448),
    .B(net766),
    .Y(_07787_));
 sg13g2_a21oi_2 _16214_ (.B1(_07787_),
    .Y(_00272_),
    .A2(_07786_),
    .A1(net765));
 sg13g2_mux2_1 _16215_ (.A0(instr_rdata_i_6_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_38_ ),
    .S(net431),
    .X(_07788_));
 sg13g2_mux2_1 _16216_ (.A0(_07533_),
    .A1(_07788_),
    .S(net559),
    .X(_07789_));
 sg13g2_nand3_1 _16217_ (.B(_07600_),
    .C(_07789_),
    .A(_07588_),
    .Y(_07790_));
 sg13g2_nand2_1 _16218_ (.Y(_07791_),
    .A(_07780_),
    .B(_07790_));
 sg13g2_a22oi_1 _16219_ (.Y(_07792_),
    .B1(_07791_),
    .B2(net335),
    .A2(_07779_),
    .A1(net1608));
 sg13g2_o21ai_1 _16220_ (.B1(net1427),
    .Y(_07793_),
    .A1(net1608),
    .A2(_07663_));
 sg13g2_inv_1 _16221_ (.Y(_07794_),
    .A(_07789_));
 sg13g2_inv_1 _16222_ (.Y(_07795_),
    .A(net1607));
 sg13g2_nand3_1 _16223_ (.B(_07508_),
    .C(_07795_),
    .A(net1667),
    .Y(_07796_));
 sg13g2_o21ai_1 _16224_ (.B1(_07796_),
    .Y(_07797_),
    .A1(net1633),
    .A2(net1626));
 sg13g2_a221oi_1 _16225_ (.B2(net1659),
    .C1(net1536),
    .B1(_07797_),
    .A1(net1563),
    .Y(_07798_),
    .A2(_07794_));
 sg13g2_nand2_1 _16226_ (.Y(_07799_),
    .A(net1608),
    .B(_07667_));
 sg13g2_nand2_1 _16227_ (.Y(_07800_),
    .A(_07755_),
    .B(_07789_));
 sg13g2_nand3_1 _16228_ (.B(_07799_),
    .C(_07800_),
    .A(net1531),
    .Y(_07801_));
 sg13g2_o21ai_1 _16229_ (.B1(_07801_),
    .Y(_07802_),
    .A1(net1531),
    .A2(_07798_));
 sg13g2_o21ai_1 _16230_ (.B1(_07802_),
    .Y(_07803_),
    .A1(_07792_),
    .A2(_07793_));
 sg13g2_mux2_1 _16231_ (.A0(net447),
    .A1(_07803_),
    .S(net759),
    .X(_00273_));
 sg13g2_o21ai_1 _16232_ (.B1(net1631),
    .Y(_07804_),
    .A1(net1668),
    .A2(_07600_));
 sg13g2_mux2_1 _16233_ (.A0(instr_rdata_i_7_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_39_ ),
    .S(net430),
    .X(_07805_));
 sg13g2_nand2_1 _16234_ (.Y(_07806_),
    .A(_01512_),
    .B(instr_rdata_i_23_));
 sg13g2_nand2_1 _16235_ (.Y(_07807_),
    .A(net1985),
    .B(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23_ ));
 sg13g2_nand3_1 _16236_ (.B(_07806_),
    .C(_07807_),
    .A(net1864),
    .Y(_07808_));
 sg13g2_o21ai_1 _16237_ (.B1(_07808_),
    .Y(_07809_),
    .A1(net1864),
    .A2(_07805_));
 sg13g2_a21oi_1 _16238_ (.A1(net335),
    .A2(_07809_),
    .Y(_07810_),
    .B1(_07647_));
 sg13g2_a22oi_1 _16239_ (.Y(_07811_),
    .B1(_07810_),
    .B2(_07576_),
    .A2(_07804_),
    .A1(net1628));
 sg13g2_and2_1 _16240_ (.A(net388),
    .B(net1627),
    .X(_07812_));
 sg13g2_nor4_1 _16241_ (.A(net1603),
    .B(net389),
    .C(net1629),
    .D(net333),
    .Y(_07813_));
 sg13g2_nor3_1 _16242_ (.A(net1657),
    .B(_07812_),
    .C(_07813_),
    .Y(_07814_));
 sg13g2_a21oi_1 _16243_ (.A1(net1657),
    .A2(_07811_),
    .Y(_07815_),
    .B1(_07814_));
 sg13g2_a21oi_1 _16244_ (.A1(net393),
    .A2(net1668),
    .Y(_07816_),
    .B1(_07812_));
 sg13g2_a221oi_1 _16245_ (.B2(_07608_),
    .C1(net1534),
    .B1(_07816_),
    .A1(net1564),
    .Y(_07817_),
    .A2(_07809_));
 sg13g2_a21oi_1 _16246_ (.A1(net1534),
    .A2(_07815_),
    .Y(_07818_),
    .B1(_07817_));
 sg13g2_nand2_1 _16247_ (.Y(_07819_),
    .A(net1627),
    .B(_07667_));
 sg13g2_o21ai_1 _16248_ (.B1(_07819_),
    .Y(_07820_),
    .A1(_07667_),
    .A2(_07809_));
 sg13g2_nor2_1 _16249_ (.A(net1523),
    .B(_07820_),
    .Y(_07821_));
 sg13g2_a21oi_1 _16250_ (.A1(net1523),
    .A2(_07818_),
    .Y(_07822_),
    .B1(_07821_));
 sg13g2_mux2_1 _16251_ (.A0(net2007),
    .A1(_07822_),
    .S(net763),
    .X(_00274_));
 sg13g2_mux2_1 _16252_ (.A0(instr_rdata_i_8_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_40_ ),
    .S(net430),
    .X(_07823_));
 sg13g2_mux2_2 _16253_ (.A0(_07540_),
    .A1(_07823_),
    .S(net558),
    .X(_07824_));
 sg13g2_a221oi_1 _16254_ (.B2(_07824_),
    .C1(net1529),
    .B1(net1564),
    .A1(net391),
    .Y(_07825_),
    .A2(_07608_));
 sg13g2_a21oi_1 _16255_ (.A1(net1656),
    .A2(net1625),
    .Y(_07826_),
    .B1(net1523));
 sg13g2_nor2_1 _16256_ (.A(net1533),
    .B(_07826_),
    .Y(_07827_));
 sg13g2_a21oi_1 _16257_ (.A1(_07742_),
    .A2(_07824_),
    .Y(_07828_),
    .B1(_07827_));
 sg13g2_o21ai_1 _16258_ (.B1(net1426),
    .Y(_07829_),
    .A1(net1625),
    .A2(_07663_));
 sg13g2_nand2_1 _16259_ (.Y(_07830_),
    .A(net1626),
    .B(_07647_));
 sg13g2_nand3_1 _16260_ (.B(_07600_),
    .C(_07824_),
    .A(net335),
    .Y(_07831_));
 sg13g2_nand3_1 _16261_ (.B(_07830_),
    .C(_07831_),
    .A(net1629),
    .Y(_07832_));
 sg13g2_a22oi_1 _16262_ (.Y(_07833_),
    .B1(_07832_),
    .B2(net389),
    .A2(net1626),
    .A1(net1623));
 sg13g2_nand2_1 _16263_ (.Y(_07834_),
    .A(net1626),
    .B(net333));
 sg13g2_o21ai_1 _16264_ (.B1(_07834_),
    .Y(_07835_),
    .A1(net1604),
    .A2(net333));
 sg13g2_a22oi_1 _16265_ (.Y(_07836_),
    .B1(_07621_),
    .B2(_07835_),
    .A2(_07592_),
    .A1(net390));
 sg13g2_o21ai_1 _16266_ (.B1(_07836_),
    .Y(_07837_),
    .A1(net1671),
    .A2(_07833_));
 sg13g2_nand2b_1 _16267_ (.Y(_07838_),
    .B(_07837_),
    .A_N(_07829_));
 sg13g2_o21ai_1 _16268_ (.B1(_07838_),
    .Y(_07839_),
    .A1(_07825_),
    .A2(_07828_));
 sg13g2_mux2_1 _16269_ (.A0(\id_stage_i.controller_i.instr_i_24_ ),
    .A1(_07839_),
    .S(net759),
    .X(_00275_));
 sg13g2_nand2_1 _16270_ (.Y(_07840_),
    .A(net335),
    .B(net1667));
 sg13g2_mux2_1 _16271_ (.A0(instr_rdata_i_9_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_41_ ),
    .S(net430),
    .X(_07841_));
 sg13g2_mux2_2 _16272_ (.A0(_07544_),
    .A1(_07841_),
    .S(net558),
    .X(_07842_));
 sg13g2_nand2_1 _16273_ (.Y(_07843_),
    .A(_07755_),
    .B(_07842_));
 sg13g2_o21ai_1 _16274_ (.B1(_07843_),
    .Y(_07844_),
    .A1(_07755_),
    .A2(_07840_));
 sg13g2_nand2_1 _16275_ (.Y(_07845_),
    .A(_07697_),
    .B(net1563));
 sg13g2_a221oi_1 _16276_ (.B2(net334),
    .C1(net1537),
    .B1(_07845_),
    .A1(_07693_),
    .Y(_07846_),
    .A2(_07842_));
 sg13g2_and2_1 _16277_ (.A(net334),
    .B(_07636_),
    .X(_07847_));
 sg13g2_nand2b_1 _16278_ (.Y(_07848_),
    .B(net392),
    .A_N(_07842_));
 sg13g2_nand2_1 _16279_ (.Y(_07849_),
    .A(net335),
    .B(net1659));
 sg13g2_nor2_1 _16280_ (.A(_07678_),
    .B(_07849_),
    .Y(_07850_));
 sg13g2_a21oi_1 _16281_ (.A1(_07847_),
    .A2(_07848_),
    .Y(_07851_),
    .B1(_07850_));
 sg13g2_nand2b_1 _16282_ (.Y(_07852_),
    .B(_07851_),
    .A_N(_07715_));
 sg13g2_o21ai_1 _16283_ (.B1(_07852_),
    .Y(_07853_),
    .A1(net1667),
    .A2(net1633));
 sg13g2_o21ai_1 _16284_ (.B1(net1611),
    .Y(_07854_),
    .A1(net333),
    .A2(_07678_));
 sg13g2_a22oi_1 _16285_ (.Y(_07855_),
    .B1(_07854_),
    .B2(_07851_),
    .A2(_07853_),
    .A1(net1659));
 sg13g2_a21oi_1 _16286_ (.A1(_07780_),
    .A2(_07663_),
    .Y(_07856_),
    .B1(net1604));
 sg13g2_nor3_1 _16287_ (.A(_07563_),
    .B(_07855_),
    .C(_07856_),
    .Y(_07857_));
 sg13g2_nor3_1 _16288_ (.A(net1530),
    .B(_07846_),
    .C(_07857_),
    .Y(_07858_));
 sg13g2_a21oi_2 _16289_ (.B1(_07858_),
    .Y(_07859_),
    .A2(_07844_),
    .A1(net1530));
 sg13g2_nor2_2 _16290_ (.A(net2005),
    .B(net759),
    .Y(_07860_));
 sg13g2_a21oi_2 _16291_ (.B1(_07860_),
    .Y(_00276_),
    .A2(_07859_),
    .A1(net759));
 sg13g2_mux2_1 _16292_ (.A0(instr_rdata_i_10_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_42_ ),
    .S(net431),
    .X(_07861_));
 sg13g2_mux2_2 _16293_ (.A0(_07473_),
    .A1(_07861_),
    .S(net559),
    .X(_07862_));
 sg13g2_o21ai_1 _16294_ (.B1(_07847_),
    .Y(_07863_),
    .A1(_07578_),
    .A2(_07862_));
 sg13g2_and2_1 _16295_ (.A(net333),
    .B(_07621_),
    .X(_07864_));
 sg13g2_nand2_1 _16296_ (.Y(_07865_),
    .A(net1628),
    .B(_07864_));
 sg13g2_nand2_1 _16297_ (.Y(_07866_),
    .A(net1632),
    .B(net1628));
 sg13g2_o21ai_1 _16298_ (.B1(_07866_),
    .Y(_07867_),
    .A1(net1632),
    .A2(_07849_));
 sg13g2_a22oi_1 _16299_ (.Y(_07868_),
    .B1(_07867_),
    .B2(net1666),
    .A2(_07592_),
    .A1(net1662));
 sg13g2_nand3_1 _16300_ (.B(_07865_),
    .C(_07868_),
    .A(_07863_),
    .Y(_07869_));
 sg13g2_a21oi_1 _16301_ (.A1(_07663_),
    .A2(_07869_),
    .Y(_07870_),
    .B1(_07856_));
 sg13g2_nand2_1 _16302_ (.Y(_07871_),
    .A(net1663),
    .B(_07701_));
 sg13g2_a22oi_1 _16303_ (.Y(_07872_),
    .B1(net1563),
    .B2(_07862_),
    .A2(_07672_),
    .A1(net1628));
 sg13g2_a21oi_1 _16304_ (.A1(_07871_),
    .A2(_07872_),
    .Y(_07873_),
    .B1(net1536));
 sg13g2_nand2_1 _16305_ (.Y(_07874_),
    .A(net1632),
    .B(net1663));
 sg13g2_nand2_1 _16306_ (.Y(_07875_),
    .A(_07874_),
    .B(_07767_));
 sg13g2_nand3_1 _16307_ (.B(_07672_),
    .C(_07875_),
    .A(net1528),
    .Y(_07876_));
 sg13g2_a21oi_1 _16308_ (.A1(_07755_),
    .A2(_07862_),
    .Y(_07877_),
    .B1(net1524));
 sg13g2_nand2_1 _16309_ (.Y(_07878_),
    .A(_07876_),
    .B(_07877_));
 sg13g2_o21ai_1 _16310_ (.B1(_07878_),
    .Y(_07879_),
    .A1(net1531),
    .A2(_07873_));
 sg13g2_o21ai_1 _16311_ (.B1(_07879_),
    .Y(_07880_),
    .A1(_07630_),
    .A2(_07870_));
 sg13g2_mux2_1 _16312_ (.A0(net2003),
    .A1(_07880_),
    .S(net759),
    .X(_00277_));
 sg13g2_nand2_1 _16313_ (.Y(_07881_),
    .A(net385),
    .B(_07697_));
 sg13g2_mux2_1 _16314_ (.A0(instr_rdata_i_11_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_43_ ),
    .S(net431),
    .X(_07882_));
 sg13g2_mux2_2 _16315_ (.A0(_07478_),
    .A1(_07882_),
    .S(net559),
    .X(_07883_));
 sg13g2_nand2_1 _16316_ (.Y(_07884_),
    .A(_07693_),
    .B(_07883_));
 sg13g2_o21ai_1 _16317_ (.B1(_07884_),
    .Y(_07885_),
    .A1(net1563),
    .A2(_07881_));
 sg13g2_nand2b_1 _16318_ (.Y(_07886_),
    .B(net392),
    .A_N(_07883_));
 sg13g2_o21ai_1 _16319_ (.B1(net1626),
    .Y(_07887_),
    .A1(_07592_),
    .A2(_07715_));
 sg13g2_nand2b_1 _16320_ (.Y(_07888_),
    .B(_07887_),
    .A_N(_07850_));
 sg13g2_a221oi_1 _16321_ (.B2(_07847_),
    .C1(_07888_),
    .B1(_07886_),
    .A1(net1609),
    .Y(_07889_),
    .A2(_07864_));
 sg13g2_inv_1 _16322_ (.Y(_07890_),
    .A(_07856_));
 sg13g2_o21ai_1 _16323_ (.B1(_07890_),
    .Y(_07891_),
    .A1(_07614_),
    .A2(_07889_));
 sg13g2_nand2_1 _16324_ (.Y(_07892_),
    .A(_07755_),
    .B(_07883_));
 sg13g2_mux2_1 _16325_ (.A0(net1609),
    .A1(net386),
    .S(net1632),
    .X(_07893_));
 sg13g2_nand3_1 _16326_ (.B(_07667_),
    .C(_07893_),
    .A(net1666),
    .Y(_07894_));
 sg13g2_a21oi_1 _16327_ (.A1(_07892_),
    .A2(_07894_),
    .Y(_07895_),
    .B1(net1524));
 sg13g2_a221oi_1 _16328_ (.B2(net1427),
    .C1(_07895_),
    .B1(_07891_),
    .A1(_07694_),
    .Y(_07896_),
    .A2(_07885_));
 sg13g2_nor2_2 _16329_ (.A(\id_stage_i.controller_i.instr_i_27_ ),
    .B(net759),
    .Y(_07897_));
 sg13g2_a21oi_1 _16330_ (.A1(net759),
    .A2(_07896_),
    .Y(_00278_),
    .B1(_07897_));
 sg13g2_mux2_1 _16331_ (.A0(instr_rdata_i_12_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_44_ ),
    .S(net430),
    .X(_07898_));
 sg13g2_nor2_1 _16332_ (.A(net1863),
    .B(_07898_),
    .Y(_07899_));
 sg13g2_a21oi_2 _16333_ (.B1(_07899_),
    .Y(_07900_),
    .A2(_07483_),
    .A1(net1863));
 sg13g2_nand2b_1 _16334_ (.Y(_07901_),
    .B(net392),
    .A_N(_07900_));
 sg13g2_nor2_1 _16335_ (.A(net1659),
    .B(net1633),
    .Y(_07902_));
 sg13g2_nand2_1 _16336_ (.Y(_07903_),
    .A(net1661),
    .B(net1606));
 sg13g2_o21ai_1 _16337_ (.B1(_07903_),
    .Y(_07904_),
    .A1(_07902_),
    .A2(_07840_));
 sg13g2_a221oi_1 _16338_ (.B2(_07847_),
    .C1(_07904_),
    .B1(_07901_),
    .A1(net1608),
    .Y(_07905_),
    .A2(_07864_));
 sg13g2_o21ai_1 _16339_ (.B1(_07890_),
    .Y(_07906_),
    .A1(_07614_),
    .A2(_07905_));
 sg13g2_nand2_1 _16340_ (.Y(_07907_),
    .A(net1427),
    .B(_07906_));
 sg13g2_and2_1 _16341_ (.A(_07694_),
    .B(_07701_),
    .X(_07908_));
 sg13g2_a22oi_1 _16342_ (.Y(_07909_),
    .B1(_07908_),
    .B2(_07546_),
    .A2(_07900_),
    .A1(_07617_));
 sg13g2_nand3_1 _16343_ (.B(_07907_),
    .C(_07909_),
    .A(net764),
    .Y(_07910_));
 sg13g2_o21ai_1 _16344_ (.B1(_07910_),
    .Y(_07911_),
    .A1(\id_stage_i.controller_i.instr_i_28_ ),
    .A2(net765));
 sg13g2_inv_1 _16345_ (.Y(_00279_),
    .A(_07911_));
 sg13g2_mux2_1 _16346_ (.A0(instr_rdata_i_13_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_45_ ),
    .S(net431),
    .X(_07912_));
 sg13g2_nor2_1 _16347_ (.A(net1861),
    .B(_07912_),
    .Y(_07913_));
 sg13g2_a21oi_2 _16348_ (.B1(_07913_),
    .Y(_07914_),
    .A2(_07491_),
    .A1(net1861));
 sg13g2_a21oi_1 _16349_ (.A1(net393),
    .A2(net1670),
    .Y(_07915_),
    .B1(_07608_));
 sg13g2_mux2_1 _16350_ (.A0(net1604),
    .A1(_07915_),
    .S(net389),
    .X(_07916_));
 sg13g2_o21ai_1 _16351_ (.B1(_07847_),
    .Y(_07917_),
    .A1(_07578_),
    .A2(_07914_));
 sg13g2_a221oi_1 _16352_ (.B2(_07917_),
    .C1(_07630_),
    .B1(_07916_),
    .A1(net1604),
    .Y(_07918_),
    .A2(_07614_));
 sg13g2_a221oi_1 _16353_ (.B2(_07617_),
    .C1(_07918_),
    .B1(_07914_),
    .A1(net393),
    .Y(_07919_),
    .A2(_07908_));
 sg13g2_nor2_1 _16354_ (.A(\id_stage_i.controller_i.instr_i_29_ ),
    .B(net766),
    .Y(_07920_));
 sg13g2_a21oi_2 _16355_ (.B1(_07920_),
    .Y(_00280_),
    .A2(_07919_),
    .A1(net765));
 sg13g2_a21oi_1 _16356_ (.A1(_07577_),
    .A2(net296),
    .Y(_07921_),
    .B1(_07694_));
 sg13g2_a21oi_1 _16357_ (.A1(net1673),
    .A2(_07694_),
    .Y(_07922_),
    .B1(_07695_));
 sg13g2_o21ai_1 _16358_ (.B1(_07922_),
    .Y(_07923_),
    .A1(_07692_),
    .A2(_07921_));
 sg13g2_inv_1 _16359_ (.Y(_07924_),
    .A(_07759_));
 sg13g2_a22oi_1 _16360_ (.Y(_07925_),
    .B1(_07589_),
    .B2(_07924_),
    .A2(net1610),
    .A1(net1671));
 sg13g2_o21ai_1 _16361_ (.B1(_07631_),
    .Y(_07926_),
    .A1(net1606),
    .A2(_07622_));
 sg13g2_o21ai_1 _16362_ (.B1(_07926_),
    .Y(_07927_),
    .A1(_07590_),
    .A2(_07925_));
 sg13g2_a21oi_1 _16363_ (.A1(net1610),
    .A2(_07923_),
    .Y(_07928_),
    .B1(_07927_));
 sg13g2_nor2_2 _16364_ (.A(\id_stage_i.controller_i.instr_i_2_ ),
    .B(net767),
    .Y(_07929_));
 sg13g2_a21oi_1 _16365_ (.A1(net767),
    .A2(_07928_),
    .Y(_00281_),
    .B1(_07929_));
 sg13g2_mux2_1 _16366_ (.A0(instr_rdata_i_14_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_46_ ),
    .S(net430),
    .X(_07930_));
 sg13g2_nor2_1 _16367_ (.A(net1861),
    .B(_07930_),
    .Y(_07931_));
 sg13g2_a21oi_2 _16368_ (.B1(_07931_),
    .Y(_07932_),
    .A2(_07498_),
    .A1(net1861));
 sg13g2_nand2_1 _16369_ (.Y(_07933_),
    .A(net389),
    .B(_07580_));
 sg13g2_o21ai_1 _16370_ (.B1(net390),
    .Y(_07934_),
    .A1(net334),
    .A2(_07584_));
 sg13g2_nor2b_1 _16371_ (.A(net393),
    .B_N(net390),
    .Y(_07935_));
 sg13g2_a21oi_1 _16372_ (.A1(net393),
    .A2(_07932_),
    .Y(_07936_),
    .B1(_07935_));
 sg13g2_o21ai_1 _16373_ (.B1(net1629),
    .Y(_07937_),
    .A1(net1603),
    .A2(_07936_));
 sg13g2_a21oi_1 _16374_ (.A1(net393),
    .A2(_07934_),
    .Y(_07938_),
    .B1(_07937_));
 sg13g2_nand2_1 _16375_ (.Y(_07939_),
    .A(net1657),
    .B(_07938_));
 sg13g2_o21ai_1 _16376_ (.B1(_07939_),
    .Y(_07940_),
    .A1(net1657),
    .A2(net385));
 sg13g2_a221oi_1 _16377_ (.B2(net389),
    .C1(_07630_),
    .B1(_07940_),
    .A1(net1605),
    .Y(_07941_),
    .A2(_07933_));
 sg13g2_a21oi_2 _16378_ (.B1(_07941_),
    .Y(_07942_),
    .A2(_07932_),
    .A1(_07617_));
 sg13g2_nor2_2 _16379_ (.A(net441),
    .B(net761),
    .Y(_07943_));
 sg13g2_a21oi_2 _16380_ (.B1(_07943_),
    .Y(_00282_),
    .A2(_07942_),
    .A1(net761));
 sg13g2_mux2_1 _16381_ (.A0(instr_rdata_i_15_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_47_ ),
    .S(net431),
    .X(_07944_));
 sg13g2_nor2_1 _16382_ (.A(net1861),
    .B(_07944_),
    .Y(_07945_));
 sg13g2_a21oi_1 _16383_ (.A1(net1863),
    .A2(_07505_),
    .Y(_07946_),
    .B1(_07945_));
 sg13g2_o21ai_1 _16384_ (.B1(net390),
    .Y(_07947_),
    .A1(_07578_),
    .A2(_07946_));
 sg13g2_nand2_1 _16385_ (.Y(_07948_),
    .A(net335),
    .B(net1426));
 sg13g2_a21oi_1 _16386_ (.A1(_07588_),
    .A2(_07947_),
    .Y(_07949_),
    .B1(_07948_));
 sg13g2_a21oi_1 _16387_ (.A1(_07617_),
    .A2(_07946_),
    .Y(_07950_),
    .B1(_07949_));
 sg13g2_nor2_2 _16388_ (.A(net2002),
    .B(net763),
    .Y(_07951_));
 sg13g2_a21oi_1 _16389_ (.A1(net763),
    .A2(_07950_),
    .Y(_00283_),
    .B1(_07951_));
 sg13g2_nand3_1 _16390_ (.B(net296),
    .C(net1426),
    .A(_07588_),
    .Y(_07952_));
 sg13g2_nand2b_1 _16391_ (.Y(_07953_),
    .B(_07952_),
    .A_N(_07617_));
 sg13g2_a22oi_1 _16392_ (.Y(_07954_),
    .B1(_07953_),
    .B2(net1609),
    .A2(net1426),
    .A1(net1606));
 sg13g2_nor2_2 _16393_ (.A(net1998),
    .B(net765),
    .Y(_07955_));
 sg13g2_a21oi_1 _16394_ (.A1(net765),
    .A2(_07954_),
    .Y(_00284_),
    .B1(_07955_));
 sg13g2_nand3_1 _16395_ (.B(_07585_),
    .C(_07924_),
    .A(net1631),
    .Y(_07956_));
 sg13g2_nand3_1 _16396_ (.B(net388),
    .C(_07956_),
    .A(net1658),
    .Y(_07957_));
 sg13g2_o21ai_1 _16397_ (.B1(_07957_),
    .Y(_07958_),
    .A1(net1658),
    .A2(_07795_));
 sg13g2_o21ai_1 _16398_ (.B1(net388),
    .Y(_07959_),
    .A1(net1607),
    .A2(_07729_));
 sg13g2_a21oi_1 _16399_ (.A1(net1631),
    .A2(_07959_),
    .Y(_07960_),
    .B1(net1606));
 sg13g2_a22oi_1 _16400_ (.Y(_07961_),
    .B1(_07795_),
    .B2(net1564),
    .A2(net1668),
    .A1(net1658));
 sg13g2_mux4_1 _16401_ (.S0(net1527),
    .A0(net1607),
    .A1(_07958_),
    .A2(_07960_),
    .A3(_07961_),
    .S1(net1522),
    .X(_07962_));
 sg13g2_mux2_1 _16402_ (.A0(net1997),
    .A1(_07962_),
    .S(net760),
    .X(_00285_));
 sg13g2_a21oi_1 _16403_ (.A1(net1656),
    .A2(_07604_),
    .Y(_07963_),
    .B1(net1627));
 sg13g2_or2_1 _16404_ (.X(_07964_),
    .B(_07963_),
    .A(_07608_));
 sg13g2_a21oi_1 _16405_ (.A1(net1666),
    .A2(_07780_),
    .Y(_07965_),
    .B1(_07583_));
 sg13g2_o21ai_1 _16406_ (.B1(_07600_),
    .Y(_07966_),
    .A1(net1604),
    .A2(net1628));
 sg13g2_nand2_1 _16407_ (.Y(_07967_),
    .A(_07583_),
    .B(_07966_));
 sg13g2_o21ai_1 _16408_ (.B1(_07967_),
    .Y(_07968_),
    .A1(net1632),
    .A2(_07965_));
 sg13g2_nor3_1 _16409_ (.A(net1526),
    .B(net1523),
    .C(net1627),
    .Y(_07969_));
 sg13g2_a221oi_1 _16410_ (.B2(net1426),
    .C1(_07969_),
    .B1(_07968_),
    .A1(net1526),
    .Y(_07970_),
    .A2(_07964_));
 sg13g2_mux2_1 _16411_ (.A0(net1996),
    .A1(_07970_),
    .S(net760),
    .X(_00286_));
 sg13g2_a21o_1 _16412_ (.A2(_07682_),
    .A1(net1625),
    .B1(net1665),
    .X(_07971_));
 sg13g2_a21oi_1 _16413_ (.A1(net1630),
    .A2(_07971_),
    .Y(_07972_),
    .B1(net1606));
 sg13g2_a22oi_1 _16414_ (.Y(_07973_),
    .B1(_07617_),
    .B2(net1625),
    .A2(_07612_),
    .A1(_07589_));
 sg13g2_o21ai_1 _16415_ (.B1(_07973_),
    .Y(_07974_),
    .A1(_07630_),
    .A2(_07972_));
 sg13g2_mux2_1 _16416_ (.A0(net1995),
    .A1(_07974_),
    .S(net760),
    .X(_00287_));
 sg13g2_a22oi_1 _16417_ (.Y(_07975_),
    .B1(_07902_),
    .B2(net1525),
    .A2(net1663),
    .A1(net1659));
 sg13g2_nor2_1 _16418_ (.A(_07567_),
    .B(_07840_),
    .Y(_07976_));
 sg13g2_a21oi_1 _16419_ (.A1(net1663),
    .A2(_07567_),
    .Y(_07977_),
    .B1(_07976_));
 sg13g2_o21ai_1 _16420_ (.B1(_07977_),
    .Y(_07978_),
    .A1(net1667),
    .A2(_07975_));
 sg13g2_nor2_1 _16421_ (.A(net1671),
    .B(net1623),
    .Y(_07979_));
 sg13g2_o21ai_1 _16422_ (.B1(_07979_),
    .Y(_07980_),
    .A1(net1668),
    .A2(_07585_));
 sg13g2_and2_1 _16423_ (.A(net334),
    .B(_07758_),
    .X(_07981_));
 sg13g2_a221oi_1 _16424_ (.B2(_07589_),
    .C1(net1525),
    .B1(_07981_),
    .A1(net1663),
    .Y(_07982_),
    .A2(_07980_));
 sg13g2_a221oi_1 _16425_ (.B2(net1663),
    .C1(net1532),
    .B1(net1564),
    .A1(net1610),
    .Y(_07983_),
    .A2(_07608_));
 sg13g2_nor3_1 _16426_ (.A(net1535),
    .B(_07982_),
    .C(_07983_),
    .Y(_07984_));
 sg13g2_a21oi_1 _16427_ (.A1(net1535),
    .A2(_07978_),
    .Y(_07985_),
    .B1(_07984_));
 sg13g2_nor2_2 _16428_ (.A(net1994),
    .B(net762),
    .Y(_07986_));
 sg13g2_a21oi_1 _16429_ (.A1(net762),
    .A2(_07985_),
    .Y(_00288_),
    .B1(_07986_));
 sg13g2_a21oi_1 _16430_ (.A1(net1609),
    .A2(_07715_),
    .Y(_07987_),
    .B1(net1527));
 sg13g2_o21ai_1 _16431_ (.B1(net1524),
    .Y(_07988_),
    .A1(net1606),
    .A2(_07715_));
 sg13g2_nand2_1 _16432_ (.Y(_07989_),
    .A(net385),
    .B(_07988_));
 sg13g2_o21ai_1 _16433_ (.B1(_07989_),
    .Y(_07990_),
    .A1(net1530),
    .A2(_07987_));
 sg13g2_nor2_1 _16434_ (.A(net1525),
    .B(_07980_),
    .Y(_07991_));
 sg13g2_a221oi_1 _16435_ (.B2(net385),
    .C1(net1532),
    .B1(net1564),
    .A1(net1609),
    .Y(_07992_),
    .A2(_07608_));
 sg13g2_o21ai_1 _16436_ (.B1(net1526),
    .Y(_07993_),
    .A1(_07991_),
    .A2(_07992_));
 sg13g2_nand3_1 _16437_ (.B(_07990_),
    .C(_07993_),
    .A(net764),
    .Y(_07994_));
 sg13g2_o21ai_1 _16438_ (.B1(_07994_),
    .Y(_00289_),
    .A1(_02333_),
    .A2(net760));
 sg13g2_nand3_1 _16439_ (.B(net1522),
    .C(net1607),
    .A(net1630),
    .Y(_07995_));
 sg13g2_o21ai_1 _16440_ (.B1(_07995_),
    .Y(_07996_),
    .A1(net1630),
    .A2(_07706_));
 sg13g2_nand2_1 _16441_ (.Y(_07997_),
    .A(net1522),
    .B(_07587_));
 sg13g2_a22oi_1 _16442_ (.Y(_07998_),
    .B1(_07997_),
    .B2(net1661),
    .A2(_07996_),
    .A1(net1665));
 sg13g2_nand3b_1 _16443_ (.B(net1630),
    .C(net1664),
    .Y(_07999_),
    .A_N(net1625));
 sg13g2_o21ai_1 _16444_ (.B1(_07999_),
    .Y(_08000_),
    .A1(net1630),
    .A2(net1607));
 sg13g2_a221oi_1 _16445_ (.B2(net1658),
    .C1(net1529),
    .B1(_08000_),
    .A1(_07706_),
    .Y(_08001_),
    .A2(net1564));
 sg13g2_nor3_1 _16446_ (.A(net1522),
    .B(_07706_),
    .C(_07589_),
    .Y(_08002_));
 sg13g2_nor3_1 _16447_ (.A(net1535),
    .B(_08001_),
    .C(_08002_),
    .Y(_08003_));
 sg13g2_a21oi_1 _16448_ (.A1(net1535),
    .A2(_07998_),
    .Y(_08004_),
    .B1(_08003_));
 sg13g2_mux2_1 _16449_ (.A0(net1991),
    .A1(_08004_),
    .S(net758),
    .X(_00290_));
 sg13g2_nor2_2 _16450_ (.A(net438),
    .B(net766),
    .Y(_08005_));
 sg13g2_a21oi_2 _16451_ (.B1(_08005_),
    .Y(_00291_),
    .A2(_07695_),
    .A1(net766));
 sg13g2_o21ai_1 _16452_ (.B1(_01494_),
    .Y(_08006_),
    .A1(net2102),
    .A2(_01466_));
 sg13g2_nor2b_1 _16453_ (.A(_01467_),
    .B_N(_08006_),
    .Y(_08007_));
 sg13g2_a21oi_1 _16454_ (.A1(_01463_),
    .A2(exc_cause_5_),
    .Y(_08008_),
    .B1(\id_stage_i.controller_i.nmi_mode_o ));
 sg13g2_a21oi_1 _16455_ (.A1(net344),
    .A2(_08007_),
    .Y(_00292_),
    .B1(_08008_));
 sg13g2_and4_1 _16456_ (.A(\id_stage_i.branch_set_$_AND__Y_B ),
    .B(net1904),
    .C(_01435_),
    .D(_02862_),
    .X(\id_stage_i.controller_i.perf_jump_o ));
 sg13g2_and3_1 _16457_ (.X(\id_stage_i.controller_i.perf_tbranch_o ),
    .A(\id_stage_i.branch_set_raw ),
    .B(\id_stage_i.branch_set_$_AND__Y_B ),
    .C(net1904));
 sg13g2_and4_1 _16458_ (.A(net1603),
    .B(net1671),
    .C(_07585_),
    .D(_07679_),
    .X(_08009_));
 sg13g2_nor3_1 _16459_ (.A(_07692_),
    .B(_07935_),
    .C(_07849_),
    .Y(_08010_));
 sg13g2_nor3_1 _16460_ (.A(net1526),
    .B(_08009_),
    .C(_08010_),
    .Y(_08011_));
 sg13g2_nor4_1 _16461_ (.A(net334),
    .B(_07584_),
    .C(net1622),
    .D(_07758_),
    .Y(_08012_));
 sg13g2_nor3_1 _16462_ (.A(net1537),
    .B(net1564),
    .C(_08012_),
    .Y(_08013_));
 sg13g2_nor2_1 _16463_ (.A(_08011_),
    .B(_08013_),
    .Y(_08014_));
 sg13g2_nand3_1 _16464_ (.B(_07576_),
    .C(_07585_),
    .A(net1603),
    .Y(_08015_));
 sg13g2_a21oi_1 _16465_ (.A1(_07678_),
    .A2(_08015_),
    .Y(_08016_),
    .B1(_07758_));
 sg13g2_nor3_1 _16466_ (.A(net1603),
    .B(net1665),
    .C(net1631),
    .Y(_08017_));
 sg13g2_or3_1 _16467_ (.A(net1671),
    .B(_08016_),
    .C(_08017_),
    .X(_08018_));
 sg13g2_a22oi_1 _16468_ (.Y(_08019_),
    .B1(_08018_),
    .B2(_07612_),
    .A2(_08014_),
    .A1(net1522));
 sg13g2_nor2_2 _16469_ (.A(\id_stage_i.decoder_i.illegal_c_insn_i ),
    .B(net757),
    .Y(_08020_));
 sg13g2_a21oi_2 _16470_ (.B1(_08020_),
    .Y(_00293_),
    .A2(_08019_),
    .A1(net757));
 sg13g2_nand2_1 _16471_ (.Y(_08021_),
    .A(net358),
    .B(_01552_));
 sg13g2_or2_1 _16472_ (.X(_08022_),
    .B(_07412_),
    .A(_01624_));
 sg13g2_nand4_1 _16473_ (.B(_01433_),
    .C(_08021_),
    .A(_01162_),
    .Y(_08023_),
    .D(_08022_));
 sg13g2_a21oi_1 _16474_ (.A1(_01569_),
    .A2(_08023_),
    .Y(_08024_),
    .B1(\id_stage_i.id_fsm_q ));
 sg13g2_nor3_1 _16475_ (.A(_01429_),
    .B(_01434_),
    .C(_01567_),
    .Y(_08025_));
 sg13g2_nor2_1 _16476_ (.A(_08024_),
    .B(_08025_),
    .Y(_00294_));
 sg13g2_nand2_1 _16477_ (.Y(_08026_),
    .A(\id_stage_i.id_fsm_q ),
    .B(_01566_));
 sg13g2_nand2_1 _16478_ (.Y(_08027_),
    .A(_01552_),
    .B(_08026_));
 sg13g2_o21ai_1 _16479_ (.B1(_08027_),
    .Y(_08028_),
    .A1(_01626_),
    .A2(_08026_));
 sg13g2_and3_1 _16480_ (.X(\id_stage_i.perf_div_wait_o ),
    .A(net355),
    .B(_03957_),
    .C(_08028_));
 sg13g2_nor3_1 _16481_ (.A(_01434_),
    .B(_03216_),
    .C(_01626_),
    .Y(\id_stage_i.perf_dside_wait_o ));
 sg13g2_nor4_2 _16482_ (.A(net105),
    .B(_01519_),
    .C(_01580_),
    .Y(_08029_),
    .D(_03194_));
 sg13g2_nand3_1 _16483_ (.B(_07410_),
    .C(_03194_),
    .A(net437),
    .Y(_08030_));
 sg13g2_nand2b_1 _16484_ (.Y(\if_stage_i.instr_valid_id_d ),
    .B(_08030_),
    .A_N(_08029_));
 sg13g2_inv_1 _16485_ (.Y(_08031_),
    .A(\if_stage_i.prefetch_buffer_i.discard_req_q ));
 sg13g2_inv_1 _16486_ (.Y(_08032_),
    .A(\if_stage_i.prefetch_buffer_i.valid_req_q ));
 sg13g2_buf_16 fanout775 (.X(net775),
    .A(net776));
 sg13g2_a21oi_2 _16488_ (.B1(net1965),
    .Y(\if_stage_i.prefetch_buffer_i.discard_req_d ),
    .A2(net117),
    .A1(_08031_));
 sg13g2_and2_1 _16489_ (.A(instr_gnt_i),
    .B(instr_req_o),
    .X(_08034_));
 sg13g2_and2_1 _16490_ (.A(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .B(_08034_),
    .X(_08035_));
 sg13g2_a221oi_1 _16491_ (.B2(_08035_),
    .C1(\if_stage_i.prefetch_buffer_i.branch_discard_q_1_ ),
    .B1(\if_stage_i.prefetch_buffer_i.discard_req_d ),
    .A1(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ),
    .Y(_08036_),
    .A2(_03283_));
 sg13g2_or2_1 _16492_ (.X(_08037_),
    .B(instr_rvalid_i),
    .A(\if_stage_i.prefetch_buffer_i.branch_discard_q_0_ ));
 sg13g2_a221oi_1 _16493_ (.B2(_08034_),
    .C1(_08037_),
    .B1(\if_stage_i.prefetch_buffer_i.discard_req_d ),
    .A1(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .Y(_08038_),
    .A2(_03283_));
 sg13g2_a21oi_1 _16494_ (.A1(instr_rvalid_i),
    .A2(_08036_),
    .Y(\if_stage_i.prefetch_buffer_i.branch_discard_s_0_ ),
    .B1(_08038_));
 sg13g2_nor2_1 _16495_ (.A(instr_rvalid_i),
    .B(_08036_),
    .Y(\if_stage_i.prefetch_buffer_i.branch_discard_s_1_ ));
 sg13g2_and2_2 _16496_ (.A(\if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__A_B ),
    .B(_01490_),
    .X(_08039_));
 sg13g2_nand2_1 _16497_ (.Y(_08040_),
    .A(net114),
    .B(_08039_));
 sg13g2_nor2_1 _16498_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_10_ ),
    .B(_08040_),
    .Y(_08041_));
 sg13g2_a21oi_2 _16499_ (.B1(_03470_),
    .Y(_08042_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_9_ ));
 sg13g2_nand2_2 _16500_ (.Y(_08043_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_7_ ),
    .B(net111));
 sg13g2_nor2b_2 _16501_ (.A(_03451_),
    .B_N(_08043_),
    .Y(_08044_));
 sg13g2_inv_1 _16502_ (.Y(_08045_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_6_ ));
 sg13g2_nand2_1 _16503_ (.Y(_08046_),
    .A(net107),
    .B(_03444_));
 sg13g2_o21ai_1 _16504_ (.B1(_08046_),
    .Y(_08047_),
    .A1(_08045_),
    .A2(net103));
 sg13g2_mux2_2 _16505_ (.A0(\if_stage_i.prefetch_buffer_i.fetch_addr_q_5_ ),
    .A1(_03436_),
    .S(net103),
    .X(_08048_));
 sg13g2_a21o_2 _16506_ (.A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ),
    .B1(_03420_),
    .X(_08049_));
 sg13g2_nand2_1 _16507_ (.Y(_08050_),
    .A(\if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__A_B ),
    .B(_01490_));
 sg13g2_nor3_1 _16508_ (.A(net1396),
    .B(_03368_),
    .C(_03405_),
    .Y(_08051_));
 sg13g2_nor2_1 _16509_ (.A(net111),
    .B(_08051_),
    .Y(_08052_));
 sg13g2_nor2b_1 _16510_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ),
    .B_N(net1099),
    .Y(_08053_));
 sg13g2_nor2_1 _16511_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ),
    .B(_03406_),
    .Y(_08054_));
 sg13g2_nor4_2 _16512_ (.A(net1170),
    .B(_08052_),
    .C(_08053_),
    .Y(_08055_),
    .D(_08054_));
 sg13g2_and2_1 _16513_ (.A(_08049_),
    .B(_08055_),
    .X(_08056_));
 sg13g2_nand3_1 _16514_ (.B(_08048_),
    .C(_08056_),
    .A(_08047_),
    .Y(_08057_));
 sg13g2_or2_1 _16515_ (.X(_08058_),
    .B(_08057_),
    .A(_08044_));
 sg13g2_inv_1 _16516_ (.Y(_08059_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_8_ ));
 sg13g2_nand2_2 _16517_ (.Y(_08060_),
    .A(net107),
    .B(_03462_));
 sg13g2_o21ai_1 _16518_ (.B1(_08060_),
    .Y(_08061_),
    .A1(_08059_),
    .A2(net103));
 sg13g2_nor2b_1 _16519_ (.A(_08058_),
    .B_N(_08061_),
    .Y(_08062_));
 sg13g2_nor2b_2 _16520_ (.A(_08042_),
    .B_N(_08062_),
    .Y(_08063_));
 sg13g2_o21ai_1 _16521_ (.B1(_08063_),
    .Y(_08064_),
    .A1(_03479_),
    .A2(_08041_));
 sg13g2_inv_1 _16522_ (.Y(_08065_),
    .A(_08063_));
 sg13g2_nand2_1 _16523_ (.Y(_08066_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_10_ ),
    .B(net111));
 sg13g2_o21ai_1 _16524_ (.B1(_08066_),
    .Y(_08067_),
    .A1(net111),
    .A2(_03478_));
 sg13g2_nor2_1 _16525_ (.A(net104),
    .B(_08039_),
    .Y(_08068_));
 sg13g2_buf_16 fanout774 (.X(net774),
    .A(net775));
 sg13g2_a22oi_1 _16527_ (.Y(_08070_),
    .B1(net49),
    .B2(\if_stage_i.prefetch_buffer_i.fetch_addr_q_10_ ),
    .A2(_08067_),
    .A1(_08065_));
 sg13g2_nand2_1 _16528_ (.Y(_00295_),
    .A(_08064_),
    .B(_08070_));
 sg13g2_nand2_2 _16529_ (.Y(_08071_),
    .A(net114),
    .B(net1170));
 sg13g2_nand2_1 _16530_ (.Y(_08072_),
    .A(_03488_),
    .B(net1121));
 sg13g2_nand3_1 _16531_ (.B(net114),
    .C(_08039_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_11_ ),
    .Y(_08073_));
 sg13g2_nand2_1 _16532_ (.Y(_08074_),
    .A(_08063_),
    .B(_08067_));
 sg13g2_a21oi_1 _16533_ (.A1(_08072_),
    .A2(_08073_),
    .Y(_08075_),
    .B1(_08074_));
 sg13g2_a21o_1 _16534_ (.A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_11_ ),
    .B1(_03488_),
    .X(_08076_));
 sg13g2_a21oi_1 _16535_ (.A1(_08063_),
    .A2(_08067_),
    .Y(_08077_),
    .B1(_08076_));
 sg13g2_buf_16 fanout773 (.X(net773),
    .A(net777));
 sg13g2_nor2_1 _16537_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_11_ ),
    .B(net1122),
    .Y(_08079_));
 sg13g2_nor3_1 _16538_ (.A(_08075_),
    .B(_08077_),
    .C(_08079_),
    .Y(_00296_));
 sg13g2_a21oi_2 _16539_ (.B1(_03496_),
    .Y(_08080_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_12_ ));
 sg13g2_nand3_1 _16540_ (.B(_08067_),
    .C(_08076_),
    .A(_08063_),
    .Y(_08081_));
 sg13g2_nor2_2 _16541_ (.A(_08080_),
    .B(_08081_),
    .Y(_08082_));
 sg13g2_nand2_1 _16542_ (.Y(_08083_),
    .A(_08080_),
    .B(_08081_));
 sg13g2_o21ai_1 _16543_ (.B1(_08083_),
    .Y(_08084_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_12_ ),
    .A2(net1122));
 sg13g2_a21oi_2 _16544_ (.B1(_08084_),
    .Y(_00297_),
    .A2(_08082_),
    .A1(net1122));
 sg13g2_a21o_2 _16545_ (.A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ),
    .B1(_03505_),
    .X(_08085_));
 sg13g2_nor2_1 _16546_ (.A(_08082_),
    .B(_08085_),
    .Y(_08086_));
 sg13g2_nor2_2 _16547_ (.A(net104),
    .B(net1170),
    .Y(_08087_));
 sg13g2_a22oi_1 _16548_ (.Y(_08088_),
    .B1(net1121),
    .B2(_03505_),
    .A2(_08087_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ));
 sg13g2_nor3_1 _16549_ (.A(_08080_),
    .B(_08081_),
    .C(_08088_),
    .Y(_08089_));
 sg13g2_nor2_1 _16550_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ),
    .B(net1121),
    .Y(_08090_));
 sg13g2_nor3_1 _16551_ (.A(_08086_),
    .B(_08089_),
    .C(_08090_),
    .Y(_00298_));
 sg13g2_inv_1 _16552_ (.Y(_08091_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ));
 sg13g2_buf_16 fanout772 (.X(net772),
    .A(net773));
 sg13g2_nand2_2 _16554_ (.Y(_08093_),
    .A(_08082_),
    .B(_08085_));
 sg13g2_a21o_1 _16555_ (.A2(net121),
    .A1(_08091_),
    .B1(_03518_),
    .X(_08094_));
 sg13g2_nor2_1 _16556_ (.A(net111),
    .B(_03517_),
    .Y(_08095_));
 sg13g2_a21oi_1 _16557_ (.A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ),
    .A2(_08087_),
    .Y(_08096_),
    .B1(_08095_));
 sg13g2_nor2_1 _16558_ (.A(_08096_),
    .B(_08093_),
    .Y(_08097_));
 sg13g2_a221oi_1 _16559_ (.B2(_08094_),
    .C1(_08097_),
    .B1(_08093_),
    .A1(_08091_),
    .Y(_00299_),
    .A2(_08068_));
 sg13g2_nand2_1 _16560_ (.Y(_08098_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_15_ ),
    .B(net111));
 sg13g2_a21o_2 _16561_ (.A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ),
    .B1(_08095_),
    .X(_08099_));
 sg13g2_nand2_1 _16562_ (.Y(_08100_),
    .A(_03505_),
    .B(_08099_));
 sg13g2_nand3_1 _16563_ (.B(\if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ),
    .C(net111),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ),
    .Y(_08101_));
 sg13g2_nand2_1 _16564_ (.Y(_08102_),
    .A(_08100_),
    .B(_08101_));
 sg13g2_nand2_1 _16565_ (.Y(_08103_),
    .A(_08082_),
    .B(_08102_));
 sg13g2_xnor2_1 _16566_ (.Y(_08104_),
    .A(_03527_),
    .B(_08103_));
 sg13g2_nand4_1 _16567_ (.B(_08039_),
    .C(_08082_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_15_ ),
    .Y(_08105_),
    .D(_08102_));
 sg13g2_o21ai_1 _16568_ (.B1(_08105_),
    .Y(_08106_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_15_ ),
    .A2(_08039_));
 sg13g2_a22oi_1 _16569_ (.Y(_00300_),
    .B1(_08106_),
    .B2(net118),
    .A2(_08104_),
    .A1(_08098_));
 sg13g2_inv_1 _16570_ (.Y(_08107_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_16_ ));
 sg13g2_nand2_2 _16571_ (.Y(_08108_),
    .A(_03527_),
    .B(_08098_));
 sg13g2_nand3_1 _16572_ (.B(_08102_),
    .C(_08108_),
    .A(_08082_),
    .Y(_08109_));
 sg13g2_inv_2 _16573_ (.Y(_08110_),
    .A(_03536_));
 sg13g2_a21oi_2 _16574_ (.B1(_08110_),
    .Y(_08111_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_16_ ));
 sg13g2_a22oi_1 _16575_ (.Y(_08112_),
    .B1(net1121),
    .B2(_08110_),
    .A2(_08087_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_16_ ));
 sg13g2_nor2_1 _16576_ (.A(_08109_),
    .B(_08112_),
    .Y(_08113_));
 sg13g2_a221oi_1 _16577_ (.B2(_08111_),
    .C1(_08113_),
    .B1(_08109_),
    .A1(_08107_),
    .Y(_00301_),
    .A2(_08068_));
 sg13g2_mux2_1 _16578_ (.A0(\if_stage_i.prefetch_buffer_i.fetch_addr_q_17_ ),
    .A1(_03542_),
    .S(net103),
    .X(_08114_));
 sg13g2_o21ai_1 _16579_ (.B1(_08114_),
    .Y(_08115_),
    .A1(_03325_),
    .A2(_03541_));
 sg13g2_nor2_1 _16580_ (.A(_08109_),
    .B(_08111_),
    .Y(_08116_));
 sg13g2_xor2_1 _16581_ (.B(_08116_),
    .A(_08115_),
    .X(_08117_));
 sg13g2_nor2_1 _16582_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_17_ ),
    .B(_08071_),
    .Y(_08118_));
 sg13g2_a21oi_1 _16583_ (.A1(_08071_),
    .A2(_08117_),
    .Y(_00302_),
    .B1(_08118_));
 sg13g2_mux2_1 _16584_ (.A0(\if_stage_i.prefetch_buffer_i.fetch_addr_q_18_ ),
    .A1(_03551_),
    .S(net103),
    .X(_08119_));
 sg13g2_or2_1 _16585_ (.X(_08120_),
    .B(_03550_),
    .A(_03325_));
 sg13g2_nand2_2 _16586_ (.Y(_08121_),
    .A(_08119_),
    .B(_08120_));
 sg13g2_inv_1 _16587_ (.Y(_08122_),
    .A(_08121_));
 sg13g2_nor3_2 _16588_ (.A(_08109_),
    .B(_08111_),
    .C(_08115_),
    .Y(_08123_));
 sg13g2_xnor2_1 _16589_ (.Y(_08124_),
    .A(_08122_),
    .B(_08123_));
 sg13g2_nor2_1 _16590_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_18_ ),
    .B(_08071_),
    .Y(_08125_));
 sg13g2_a21oi_1 _16591_ (.A1(net1122),
    .A2(_08124_),
    .Y(_00303_),
    .B1(_08125_));
 sg13g2_a22oi_1 _16592_ (.Y(_08126_),
    .B1(_03564_),
    .B2(_08120_),
    .A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_19_ ));
 sg13g2_nor2b_1 _16593_ (.A(_08126_),
    .B_N(_08119_),
    .Y(_08127_));
 sg13g2_and2_1 _16594_ (.A(_08123_),
    .B(_08127_),
    .X(_08128_));
 sg13g2_a21o_1 _16595_ (.A2(net119),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_19_ ),
    .B1(_03564_),
    .X(_08129_));
 sg13g2_a21oi_1 _16596_ (.A1(_08122_),
    .A2(_08123_),
    .Y(_08130_),
    .B1(_08129_));
 sg13g2_nor3_1 _16597_ (.A(net48),
    .B(_08128_),
    .C(_08130_),
    .Y(_08131_));
 sg13g2_a21o_1 _16598_ (.A2(net50),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_19_ ),
    .B1(_08131_),
    .X(_00304_));
 sg13g2_nor2_1 _16599_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_20_ ),
    .B(_08040_),
    .Y(_08132_));
 sg13g2_or2_1 _16600_ (.X(_08133_),
    .B(_08132_),
    .A(_03573_));
 sg13g2_inv_1 _16601_ (.Y(_08134_),
    .A(_03325_));
 sg13g2_and3_1 _16602_ (.X(_08135_),
    .A(boot_addr_i_20_),
    .B(net107),
    .C(net1396));
 sg13g2_a221oi_1 _16603_ (.B2(_03570_),
    .C1(_08135_),
    .B1(_08134_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_20_ ),
    .Y(_08136_),
    .A2(net119));
 sg13g2_nor2_1 _16604_ (.A(_08128_),
    .B(_08136_),
    .Y(_08137_));
 sg13g2_a221oi_1 _16605_ (.B2(_08133_),
    .C1(_08137_),
    .B1(_08128_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_20_ ),
    .Y(_08138_),
    .A2(net50));
 sg13g2_inv_1 _16606_ (.Y(_00305_),
    .A(_08138_));
 sg13g2_and2_1 _16607_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_21_ ),
    .B(net112),
    .X(_08139_));
 sg13g2_nor2_2 _16608_ (.A(_03581_),
    .B(_08139_),
    .Y(_08140_));
 sg13g2_nor3_1 _16609_ (.A(_08111_),
    .B(_08115_),
    .C(_08136_),
    .Y(_08141_));
 sg13g2_nand3b_1 _16610_ (.B(_08127_),
    .C(_08141_),
    .Y(_08142_),
    .A_N(_08109_));
 sg13g2_xnor2_1 _16611_ (.Y(_08143_),
    .A(_08140_),
    .B(_08142_));
 sg13g2_nand2_1 _16612_ (.Y(_08144_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_21_ ),
    .B(net49));
 sg13g2_o21ai_1 _16613_ (.B1(_08144_),
    .Y(_00306_),
    .A1(net49),
    .A2(_08143_));
 sg13g2_nor2_1 _16614_ (.A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ),
    .B(_08040_),
    .Y(_08145_));
 sg13g2_nor2_2 _16615_ (.A(_08140_),
    .B(_08142_),
    .Y(_08146_));
 sg13g2_o21ai_1 _16616_ (.B1(_08146_),
    .Y(_08147_),
    .A1(_03590_),
    .A2(_08145_));
 sg13g2_inv_1 _16617_ (.Y(_08148_),
    .A(_08146_));
 sg13g2_mux2_2 _16618_ (.A0(\if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ),
    .A1(_03589_),
    .S(net103),
    .X(_08149_));
 sg13g2_a22oi_1 _16619_ (.Y(_08150_),
    .B1(_08148_),
    .B2(_08149_),
    .A2(net50),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ));
 sg13g2_nand2_1 _16620_ (.Y(_00307_),
    .A(_08147_),
    .B(_08150_));
 sg13g2_inv_1 _16621_ (.Y(_08151_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_23_ ));
 sg13g2_a22oi_1 _16622_ (.Y(_08152_),
    .B1(_08149_),
    .B2(_03581_),
    .A2(_08139_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ));
 sg13g2_nor2_2 _16623_ (.A(_08142_),
    .B(_08152_),
    .Y(_08153_));
 sg13g2_buf_16 fanout771 (.X(net771),
    .A(net772));
 sg13g2_nand2_2 _16625_ (.Y(_08155_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_23_ ),
    .B(net112));
 sg13g2_nand2_1 _16626_ (.Y(_08156_),
    .A(_03595_),
    .B(net1122));
 sg13g2_o21ai_1 _16627_ (.B1(_08156_),
    .Y(_08157_),
    .A1(_08050_),
    .A2(_08155_));
 sg13g2_nor2b_2 _16628_ (.A(_03595_),
    .B_N(_08155_),
    .Y(_08158_));
 sg13g2_nor2b_1 _16629_ (.A(_08153_),
    .B_N(_08158_),
    .Y(_08159_));
 sg13g2_a221oi_1 _16630_ (.B2(_08157_),
    .C1(_08159_),
    .B1(_08153_),
    .A1(_08151_),
    .Y(_00308_),
    .A2(net50));
 sg13g2_a21oi_2 _16631_ (.B1(_03605_),
    .Y(_08160_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_24_ ));
 sg13g2_nand2b_1 _16632_ (.Y(_08161_),
    .B(_08153_),
    .A_N(_08158_));
 sg13g2_xnor2_1 _16633_ (.Y(_08162_),
    .A(_08160_),
    .B(_08161_));
 sg13g2_nand2_1 _16634_ (.Y(_08163_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_24_ ),
    .B(net48));
 sg13g2_o21ai_1 _16635_ (.B1(_08163_),
    .Y(_00309_),
    .A1(net48),
    .A2(_08162_));
 sg13g2_nor2_1 _16636_ (.A(net112),
    .B(_03610_),
    .Y(_08164_));
 sg13g2_a21oi_2 _16637_ (.B1(_08164_),
    .Y(_08165_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_25_ ));
 sg13g2_or2_1 _16638_ (.X(_08166_),
    .B(_08158_),
    .A(_08152_));
 sg13g2_nor3_2 _16639_ (.A(_08142_),
    .B(_08160_),
    .C(_08166_),
    .Y(_08167_));
 sg13g2_xor2_1 _16640_ (.B(_08167_),
    .A(_08165_),
    .X(_08168_));
 sg13g2_nand2_1 _16641_ (.Y(_08169_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_25_ ),
    .B(net48));
 sg13g2_o21ai_1 _16642_ (.B1(_08169_),
    .Y(_00310_),
    .A1(net48),
    .A2(_08168_));
 sg13g2_nor4_2 _16643_ (.A(_08142_),
    .B(_08160_),
    .C(_08165_),
    .Y(_08170_),
    .D(_08166_));
 sg13g2_a22oi_1 _16644_ (.Y(_08171_),
    .B1(_03622_),
    .B2(net1121),
    .A2(net121),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ));
 sg13g2_nand3_1 _16645_ (.B(net116),
    .C(net1170),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ),
    .Y(_08172_));
 sg13g2_o21ai_1 _16646_ (.B1(_08172_),
    .Y(_08173_),
    .A1(_08170_),
    .A2(_08171_));
 sg13g2_o21ai_1 _16647_ (.B1(net116),
    .Y(_08174_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ),
    .A2(net1170));
 sg13g2_nand3b_1 _16648_ (.B(_08170_),
    .C(_08174_),
    .Y(_08175_),
    .A_N(_03622_));
 sg13g2_nand2b_1 _16649_ (.Y(_00311_),
    .B(_08175_),
    .A_N(_08173_));
 sg13g2_a21oi_2 _16650_ (.B1(_03622_),
    .Y(_08176_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ));
 sg13g2_nor2b_2 _16651_ (.A(_08176_),
    .B_N(_08170_),
    .Y(_08177_));
 sg13g2_o21ai_1 _16652_ (.B1(net114),
    .Y(_08178_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_27_ ),
    .A2(net1171));
 sg13g2_and3_1 _16653_ (.X(_08179_),
    .A(_03630_),
    .B(_08177_),
    .C(_08178_));
 sg13g2_nand2_1 _16654_ (.Y(_08180_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_27_ ),
    .B(net112));
 sg13g2_a21oi_2 _16655_ (.B1(_08180_),
    .Y(_08181_),
    .A2(_08177_),
    .A1(_08039_));
 sg13g2_nor3_1 _16656_ (.A(_03630_),
    .B(net49),
    .C(_08177_),
    .Y(_08182_));
 sg13g2_or3_1 _16657_ (.A(_08179_),
    .B(_08181_),
    .C(_08182_),
    .X(_00312_));
 sg13g2_inv_1 _16658_ (.Y(_08183_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_28_ ));
 sg13g2_nand2_1 _16659_ (.Y(_08184_),
    .A(_03630_),
    .B(_08180_));
 sg13g2_and2_2 _16660_ (.A(_08177_),
    .B(_08184_),
    .X(_08185_));
 sg13g2_nand2_1 _16661_ (.Y(_08186_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_28_ ),
    .B(_08087_));
 sg13g2_o21ai_1 _16662_ (.B1(_08186_),
    .Y(_08187_),
    .A1(net113),
    .A2(_03638_));
 sg13g2_o21ai_1 _16663_ (.B1(_03639_),
    .Y(_08188_),
    .A1(_08183_),
    .A2(net103));
 sg13g2_nor2_1 _16664_ (.A(_08185_),
    .B(_08188_),
    .Y(_08189_));
 sg13g2_a221oi_1 _16665_ (.B2(_08187_),
    .C1(_08189_),
    .B1(_08185_),
    .A1(_08183_),
    .Y(_00313_),
    .A2(net50));
 sg13g2_inv_1 _16666_ (.Y(_08190_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_29_ ));
 sg13g2_o21ai_1 _16667_ (.B1(_03646_),
    .Y(_08191_),
    .A1(_08190_),
    .A2(net103));
 sg13g2_nand3_1 _16668_ (.B(_08185_),
    .C(_08188_),
    .A(net1122),
    .Y(_08192_));
 sg13g2_xnor2_1 _16669_ (.Y(_00314_),
    .A(_08191_),
    .B(_08192_));
 sg13g2_nand2_1 _16670_ (.Y(_08193_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ),
    .B(net112));
 sg13g2_nand2_2 _16671_ (.Y(_08194_),
    .A(net1099),
    .B(_08193_));
 sg13g2_o21ai_1 _16672_ (.B1(_08193_),
    .Y(_08195_),
    .A1(net113),
    .A2(net1099));
 sg13g2_nand2_1 _16673_ (.Y(_08196_),
    .A(net1171),
    .B(_08195_));
 sg13g2_o21ai_1 _16674_ (.B1(_08196_),
    .Y(_00315_),
    .A1(net1171),
    .A2(_08194_));
 sg13g2_nand4_1 _16675_ (.B(_08185_),
    .C(_08188_),
    .A(net1122),
    .Y(_08197_),
    .D(_08191_));
 sg13g2_inv_1 _16676_ (.Y(_08198_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_30_ ));
 sg13g2_o21ai_1 _16677_ (.B1(_03657_),
    .Y(_08199_),
    .A1(_08198_),
    .A2(net104));
 sg13g2_xnor2_1 _16678_ (.Y(_00316_),
    .A(_08197_),
    .B(_08199_));
 sg13g2_a21oi_1 _16679_ (.A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_31_ ),
    .A2(net1171),
    .Y(_08200_),
    .B1(net104));
 sg13g2_o21ai_1 _16680_ (.B1(_08200_),
    .Y(_08201_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_31_ ),
    .A2(net1171));
 sg13g2_and2_1 _16681_ (.A(net2491),
    .B(_08201_),
    .X(_08202_));
 sg13g2_inv_1 _16682_ (.Y(_08203_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_31_ ));
 sg13g2_o21ai_1 _16683_ (.B1(net2491),
    .Y(_08204_),
    .A1(_08203_),
    .A2(net104));
 sg13g2_nand4_1 _16684_ (.B(_08188_),
    .C(_08191_),
    .A(_08185_),
    .Y(_08205_),
    .D(_08199_));
 sg13g2_mux2_1 _16685_ (.A0(_08202_),
    .A1(_08204_),
    .S(_08205_),
    .X(_00317_));
 sg13g2_a21oi_2 _16686_ (.B1(_03406_),
    .Y(_08206_),
    .A2(net117),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ));
 sg13g2_nand4_1 _16687_ (.B(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ),
    .C(net1099),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ),
    .Y(_08207_),
    .D(_03407_));
 sg13g2_o21ai_1 _16688_ (.B1(_08207_),
    .Y(_08208_),
    .A1(net1099),
    .A2(_08206_));
 sg13g2_o21ai_1 _16689_ (.B1(net114),
    .Y(_08209_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ),
    .A2(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ));
 sg13g2_a22oi_1 _16690_ (.Y(_08210_),
    .B1(_08209_),
    .B2(net1099),
    .A2(net1170),
    .A1(net108));
 sg13g2_nand2b_1 _16691_ (.Y(_08211_),
    .B(net49),
    .A_N(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ));
 sg13g2_o21ai_1 _16692_ (.B1(_08211_),
    .Y(_08212_),
    .A1(_03406_),
    .A2(_08210_));
 sg13g2_a21oi_1 _16693_ (.A1(_08039_),
    .A2(_08208_),
    .Y(_00318_),
    .B1(_08212_));
 sg13g2_a22oi_1 _16694_ (.Y(_08213_),
    .B1(_03420_),
    .B2(net1121),
    .A2(net121),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ));
 sg13g2_nand3_1 _16695_ (.B(net114),
    .C(net1170),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ),
    .Y(_08214_));
 sg13g2_o21ai_1 _16696_ (.B1(_08214_),
    .Y(_08215_),
    .A1(_08055_),
    .A2(_08213_));
 sg13g2_o21ai_1 _16697_ (.B1(net116),
    .Y(_08216_),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ),
    .A2(net1170));
 sg13g2_nand3b_1 _16698_ (.B(_08055_),
    .C(_08216_),
    .Y(_08217_),
    .A_N(_03420_));
 sg13g2_nand2b_1 _16699_ (.Y(_00319_),
    .B(_08217_),
    .A_N(_08215_));
 sg13g2_nand2_1 _16700_ (.Y(_08218_),
    .A(_08049_),
    .B(_08055_));
 sg13g2_inv_1 _16701_ (.Y(_08219_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_5_ ));
 sg13g2_a21oi_1 _16702_ (.A1(_08219_),
    .A2(_08087_),
    .Y(_08220_),
    .B1(_03437_));
 sg13g2_a22oi_1 _16703_ (.Y(_08221_),
    .B1(net49),
    .B2(\if_stage_i.prefetch_buffer_i.fetch_addr_q_5_ ),
    .A2(_08218_),
    .A1(_08048_));
 sg13g2_o21ai_1 _16704_ (.B1(_08221_),
    .Y(_00320_),
    .A1(_08218_),
    .A2(_08220_));
 sg13g2_a21o_1 _16705_ (.A2(_08056_),
    .A1(_08048_),
    .B1(_08047_),
    .X(_08222_));
 sg13g2_nand3_1 _16706_ (.B(net1121),
    .C(_08222_),
    .A(_08057_),
    .Y(_08223_));
 sg13g2_o21ai_1 _16707_ (.B1(_08223_),
    .Y(_00321_),
    .A1(_08045_),
    .A2(net1121));
 sg13g2_nor2b_1 _16708_ (.A(_03451_),
    .B_N(_08057_),
    .Y(_08224_));
 sg13g2_o21ai_1 _16709_ (.B1(_08043_),
    .Y(_08225_),
    .A1(net48),
    .A2(_08224_));
 sg13g2_a22oi_1 _16710_ (.Y(_08226_),
    .B1(_08225_),
    .B2(_08058_),
    .A2(net50),
    .A1(\if_stage_i.prefetch_buffer_i.fetch_addr_q_7_ ));
 sg13g2_inv_1 _16711_ (.Y(_00322_),
    .A(_08226_));
 sg13g2_a21oi_1 _16712_ (.A1(_08059_),
    .A2(_08087_),
    .Y(_08227_),
    .B1(_03463_));
 sg13g2_a22oi_1 _16713_ (.Y(_08228_),
    .B1(net49),
    .B2(\if_stage_i.prefetch_buffer_i.fetch_addr_q_8_ ),
    .A2(_08058_),
    .A1(_08061_));
 sg13g2_o21ai_1 _16714_ (.B1(_08228_),
    .Y(_00323_),
    .A1(_08058_),
    .A2(_08227_));
 sg13g2_xor2_1 _16715_ (.B(_08062_),
    .A(_08042_),
    .X(_08229_));
 sg13g2_nand2_1 _16716_ (.Y(_08230_),
    .A(\if_stage_i.prefetch_buffer_i.fetch_addr_q_9_ ),
    .B(net48));
 sg13g2_o21ai_1 _16717_ (.B1(_08230_),
    .Y(_00324_),
    .A1(net48),
    .A2(_08229_));
 sg13g2_buf_8 fanout770 (.A(_03196_),
    .X(net770));
 sg13g2_a21o_1 _16719_ (.A2(net435),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ),
    .B1(_07559_),
    .X(_08232_));
 sg13g2_nor3_2 _16720_ (.A(_01519_),
    .B(_03195_),
    .C(_03295_),
    .Y(_08233_));
 sg13g2_nand3_1 _16721_ (.B(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_1__$_AND__Y_A ),
    .C(_01506_),
    .A(net1983),
    .Y(_08234_));
 sg13g2_and2_1 _16722_ (.A(_01472_),
    .B(_08234_),
    .X(_08235_));
 sg13g2_a21oi_2 _16723_ (.B1(_08233_),
    .Y(_08236_),
    .A2(_01506_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_0_ ));
 sg13g2_a21o_1 _16724_ (.A2(_08235_),
    .A1(_08233_),
    .B1(_08236_),
    .X(_08237_));
 sg13g2_buf_16 fanout769 (.X(net769),
    .A(net770));
 sg13g2_buf_16 fanout768 (.X(net768),
    .A(net769));
 sg13g2_mux2_1 _16727_ (.A0(_08232_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ),
    .S(net732),
    .X(_00325_));
 sg13g2_buf_16 fanout767 (.X(net767),
    .A(net768));
 sg13g2_mux2_1 _16729_ (.A0(instr_err_i),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_2_ ),
    .S(net1990),
    .X(_08241_));
 sg13g2_nand3_1 _16730_ (.B(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_2__$_AND__Y_A ),
    .C(_01506_),
    .A(net434),
    .Y(_08242_));
 sg13g2_buf_16 fanout766 (.X(net766),
    .A(net767));
 sg13g2_nor2b_1 _16732_ (.A(net1990),
    .B_N(net1860),
    .Y(_08244_));
 sg13g2_mux2_1 _16733_ (.A0(_08234_),
    .A1(_08244_),
    .S(_08233_),
    .X(_08245_));
 sg13g2_buf_16 fanout765 (.X(net765),
    .A(net766));
 sg13g2_buf_16 fanout764 (.X(net764),
    .A(net769));
 sg13g2_mux2_1 _16736_ (.A0(_08241_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ),
    .S(net746),
    .X(_00326_));
 sg13g2_buf_16 fanout763 (.X(net763),
    .A(net764));
 sg13g2_mux2_1 _16738_ (.A0(instr_err_i),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_2_ ),
    .S(net1860),
    .X(_00327_));
 sg13g2_mux2_1 _16739_ (.A0(_07683_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0_ ),
    .S(net732),
    .X(_00328_));
 sg13g2_mux2_1 _16740_ (.A0(_07861_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_10_ ),
    .S(net728),
    .X(_00329_));
 sg13g2_mux2_1 _16741_ (.A0(_07882_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_11_ ),
    .S(net728),
    .X(_00330_));
 sg13g2_mux2_1 _16742_ (.A0(_07898_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_12_ ),
    .S(net729),
    .X(_00331_));
 sg13g2_mux2_1 _16743_ (.A0(_07912_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_13_ ),
    .S(net729),
    .X(_00332_));
 sg13g2_mux2_1 _16744_ (.A0(_07930_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_14_ ),
    .S(net729),
    .X(_00333_));
 sg13g2_mux2_1 _16745_ (.A0(_07944_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_15_ ),
    .S(net729),
    .X(_00334_));
 sg13g2_mux2_1 _16746_ (.A0(instr_rdata_i_16_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_48_ ),
    .S(net434),
    .X(_08249_));
 sg13g2_mux2_1 _16747_ (.A0(_08249_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16_ ),
    .S(net732),
    .X(_00335_));
 sg13g2_mux2_1 _16748_ (.A0(instr_rdata_i_17_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_49_ ),
    .S(net434),
    .X(_08250_));
 sg13g2_mux2_1 _16749_ (.A0(_08250_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17_ ),
    .S(net732),
    .X(_00336_));
 sg13g2_mux2_1 _16750_ (.A0(instr_rdata_i_18_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_50_ ),
    .S(net433),
    .X(_08251_));
 sg13g2_buf_16 fanout762 (.X(net762),
    .A(net764));
 sg13g2_mux2_1 _16752_ (.A0(_08251_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_18_ ),
    .S(net730),
    .X(_00337_));
 sg13g2_mux2_1 _16753_ (.A0(instr_rdata_i_19_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_51_ ),
    .S(net433),
    .X(_08253_));
 sg13g2_mux2_1 _16754_ (.A0(_08253_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_19_ ),
    .S(net730),
    .X(_00338_));
 sg13g2_mux2_1 _16755_ (.A0(_07707_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1_ ),
    .S(_08237_),
    .X(_00339_));
 sg13g2_mux2_1 _16756_ (.A0(instr_rdata_i_20_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_52_ ),
    .S(net433),
    .X(_08254_));
 sg13g2_mux2_1 _16757_ (.A0(_08254_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_20_ ),
    .S(net730),
    .X(_00340_));
 sg13g2_mux2_1 _16758_ (.A0(instr_rdata_i_21_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_53_ ),
    .S(net433),
    .X(_08255_));
 sg13g2_mux2_1 _16759_ (.A0(_08255_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_21_ ),
    .S(net730),
    .X(_00341_));
 sg13g2_mux2_1 _16760_ (.A0(instr_rdata_i_22_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_54_ ),
    .S(net433),
    .X(_08256_));
 sg13g2_mux2_1 _16761_ (.A0(_08256_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_22_ ),
    .S(net730),
    .X(_00342_));
 sg13g2_mux2_1 _16762_ (.A0(instr_rdata_i_23_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_55_ ),
    .S(net433),
    .X(_08257_));
 sg13g2_mux2_1 _16763_ (.A0(_08257_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23_ ),
    .S(net731),
    .X(_00343_));
 sg13g2_mux2_1 _16764_ (.A0(instr_rdata_i_24_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_56_ ),
    .S(net433),
    .X(_08258_));
 sg13g2_mux2_1 _16765_ (.A0(_08258_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_24_ ),
    .S(net730),
    .X(_00344_));
 sg13g2_mux2_1 _16766_ (.A0(instr_rdata_i_25_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_57_ ),
    .S(net433),
    .X(_08259_));
 sg13g2_mux2_1 _16767_ (.A0(_08259_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_25_ ),
    .S(net731),
    .X(_00345_));
 sg13g2_mux2_1 _16768_ (.A0(instr_rdata_i_26_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_58_ ),
    .S(net432),
    .X(_08260_));
 sg13g2_mux2_1 _16769_ (.A0(_08260_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_26_ ),
    .S(net730),
    .X(_00346_));
 sg13g2_mux2_1 _16770_ (.A0(instr_rdata_i_27_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_59_ ),
    .S(net432),
    .X(_08261_));
 sg13g2_buf_16 fanout761 (.X(net761),
    .A(net769));
 sg13g2_mux2_1 _16772_ (.A0(_08261_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_27_ ),
    .S(net731),
    .X(_00347_));
 sg13g2_mux2_1 _16773_ (.A0(instr_rdata_i_28_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_60_ ),
    .S(net432),
    .X(_08263_));
 sg13g2_mux2_1 _16774_ (.A0(_08263_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_28_ ),
    .S(net731),
    .X(_00348_));
 sg13g2_mux2_1 _16775_ (.A0(instr_rdata_i_29_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_61_ ),
    .S(net432),
    .X(_08264_));
 sg13g2_mux2_1 _16776_ (.A0(_08264_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_29_ ),
    .S(net731),
    .X(_00349_));
 sg13g2_mux2_1 _16777_ (.A0(_07727_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_2_ ),
    .S(net728),
    .X(_00350_));
 sg13g2_mux2_1 _16778_ (.A0(instr_rdata_i_30_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_62_ ),
    .S(net432),
    .X(_08265_));
 sg13g2_mux2_1 _16779_ (.A0(_08265_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_30_ ),
    .S(net730),
    .X(_00351_));
 sg13g2_mux2_1 _16780_ (.A0(instr_rdata_i_31_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_63_ ),
    .S(net432),
    .X(_08266_));
 sg13g2_mux2_1 _16781_ (.A0(_08266_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_31_ ),
    .S(net731),
    .X(_00352_));
 sg13g2_mux2_1 _16782_ (.A0(instr_rdata_i_0_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_64_ ),
    .S(net1987),
    .X(_08267_));
 sg13g2_mux2_1 _16783_ (.A0(_08267_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_32_ ),
    .S(net746),
    .X(_00353_));
 sg13g2_mux2_1 _16784_ (.A0(instr_rdata_i_1_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_65_ ),
    .S(net1987),
    .X(_08268_));
 sg13g2_mux2_1 _16785_ (.A0(_08268_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_33_ ),
    .S(net746),
    .X(_00354_));
 sg13g2_mux2_1 _16786_ (.A0(instr_rdata_i_2_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_66_ ),
    .S(net1987),
    .X(_08269_));
 sg13g2_mux2_1 _16787_ (.A0(_08269_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_34_ ),
    .S(net741),
    .X(_00355_));
 sg13g2_mux2_1 _16788_ (.A0(instr_rdata_i_3_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_67_ ),
    .S(net1987),
    .X(_08270_));
 sg13g2_mux2_1 _16789_ (.A0(_08270_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_35_ ),
    .S(net741),
    .X(_00356_));
 sg13g2_mux2_1 _16790_ (.A0(instr_rdata_i_4_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_68_ ),
    .S(net1986),
    .X(_08271_));
 sg13g2_mux2_1 _16791_ (.A0(_08271_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_36_ ),
    .S(net742),
    .X(_00357_));
 sg13g2_mux2_1 _16792_ (.A0(instr_rdata_i_5_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_69_ ),
    .S(net1986),
    .X(_08272_));
 sg13g2_mux2_1 _16793_ (.A0(_08272_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_37_ ),
    .S(net741),
    .X(_00358_));
 sg13g2_mux2_1 _16794_ (.A0(instr_rdata_i_6_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_70_ ),
    .S(net1986),
    .X(_08273_));
 sg13g2_mux2_1 _16795_ (.A0(_08273_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_38_ ),
    .S(net741),
    .X(_00359_));
 sg13g2_mux2_1 _16796_ (.A0(instr_rdata_i_7_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_71_ ),
    .S(net1989),
    .X(_08274_));
 sg13g2_mux2_1 _16797_ (.A0(_08274_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_39_ ),
    .S(net746),
    .X(_00360_));
 sg13g2_mux2_1 _16798_ (.A0(_07743_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_3_ ),
    .S(net728),
    .X(_00361_));
 sg13g2_mux2_1 _16799_ (.A0(instr_rdata_i_8_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_72_ ),
    .S(net1986),
    .X(_08275_));
 sg13g2_mux2_1 _16800_ (.A0(_08275_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_40_ ),
    .S(net741),
    .X(_00362_));
 sg13g2_buf_16 fanout760 (.X(net760),
    .A(net761));
 sg13g2_mux2_1 _16802_ (.A0(instr_rdata_i_9_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_73_ ),
    .S(net1989),
    .X(_08277_));
 sg13g2_buf_16 fanout759 (.X(net759),
    .A(net761));
 sg13g2_mux2_1 _16804_ (.A0(_08277_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_41_ ),
    .S(net744),
    .X(_00363_));
 sg13g2_mux2_1 _16805_ (.A0(instr_rdata_i_10_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_74_ ),
    .S(net1986),
    .X(_08279_));
 sg13g2_mux2_1 _16806_ (.A0(_08279_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_42_ ),
    .S(net741),
    .X(_00364_));
 sg13g2_mux2_1 _16807_ (.A0(instr_rdata_i_11_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_75_ ),
    .S(net1986),
    .X(_08280_));
 sg13g2_mux2_1 _16808_ (.A0(_08280_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_43_ ),
    .S(net741),
    .X(_00365_));
 sg13g2_mux2_1 _16809_ (.A0(instr_rdata_i_12_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_76_ ),
    .S(net1990),
    .X(_08281_));
 sg13g2_mux2_1 _16810_ (.A0(_08281_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_44_ ),
    .S(net742),
    .X(_00366_));
 sg13g2_mux2_1 _16811_ (.A0(instr_rdata_i_13_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_77_ ),
    .S(net1986),
    .X(_08282_));
 sg13g2_mux2_1 _16812_ (.A0(_08282_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_45_ ),
    .S(net742),
    .X(_00367_));
 sg13g2_mux2_1 _16813_ (.A0(instr_rdata_i_14_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_78_ ),
    .S(net1986),
    .X(_08283_));
 sg13g2_mux2_1 _16814_ (.A0(_08283_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_46_ ),
    .S(net742),
    .X(_00368_));
 sg13g2_mux2_1 _16815_ (.A0(instr_rdata_i_15_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_79_ ),
    .S(net1987),
    .X(_08284_));
 sg13g2_mux2_1 _16816_ (.A0(_08284_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_47_ ),
    .S(net742),
    .X(_00369_));
 sg13g2_mux2_1 _16817_ (.A0(instr_rdata_i_16_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_80_ ),
    .S(net1990),
    .X(_08285_));
 sg13g2_mux2_1 _16818_ (.A0(_08285_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_48_ ),
    .S(net746),
    .X(_00370_));
 sg13g2_mux2_1 _16819_ (.A0(instr_rdata_i_17_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_81_ ),
    .S(net1987),
    .X(_08286_));
 sg13g2_mux2_1 _16820_ (.A0(_08286_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_49_ ),
    .S(net746),
    .X(_00371_));
 sg13g2_mux2_1 _16821_ (.A0(_07756_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_4_ ),
    .S(net729),
    .X(_00372_));
 sg13g2_mux2_1 _16822_ (.A0(instr_rdata_i_18_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_82_ ),
    .S(net1988),
    .X(_08287_));
 sg13g2_mux2_1 _16823_ (.A0(_08287_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_50_ ),
    .S(net743),
    .X(_00373_));
 sg13g2_buf_16 fanout758 (.X(net758),
    .A(net769));
 sg13g2_mux2_1 _16825_ (.A0(instr_rdata_i_19_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_83_ ),
    .S(net1989),
    .X(_08289_));
 sg13g2_buf_16 fanout757 (.X(net757),
    .A(net758));
 sg13g2_mux2_1 _16827_ (.A0(_08289_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_51_ ),
    .S(net743),
    .X(_00374_));
 sg13g2_mux2_1 _16828_ (.A0(instr_rdata_i_20_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_84_ ),
    .S(net1989),
    .X(_08291_));
 sg13g2_mux2_1 _16829_ (.A0(_08291_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_52_ ),
    .S(net743),
    .X(_00375_));
 sg13g2_mux2_1 _16830_ (.A0(instr_rdata_i_21_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_85_ ),
    .S(net1988),
    .X(_08292_));
 sg13g2_mux2_1 _16831_ (.A0(_08292_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_53_ ),
    .S(net743),
    .X(_00376_));
 sg13g2_mux2_1 _16832_ (.A0(instr_rdata_i_22_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_86_ ),
    .S(net1989),
    .X(_08293_));
 sg13g2_mux2_1 _16833_ (.A0(_08293_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_54_ ),
    .S(net743),
    .X(_00377_));
 sg13g2_mux2_1 _16834_ (.A0(instr_rdata_i_23_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_87_ ),
    .S(net1989),
    .X(_08294_));
 sg13g2_mux2_1 _16835_ (.A0(_08294_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_55_ ),
    .S(net744),
    .X(_00378_));
 sg13g2_mux2_1 _16836_ (.A0(instr_rdata_i_24_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_88_ ),
    .S(net1988),
    .X(_08295_));
 sg13g2_mux2_1 _16837_ (.A0(_08295_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_56_ ),
    .S(net744),
    .X(_00379_));
 sg13g2_mux2_1 _16838_ (.A0(instr_rdata_i_25_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_89_ ),
    .S(net1989),
    .X(_08296_));
 sg13g2_mux2_1 _16839_ (.A0(_08296_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_57_ ),
    .S(net744),
    .X(_00380_));
 sg13g2_mux2_1 _16840_ (.A0(instr_rdata_i_26_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_90_ ),
    .S(net1987),
    .X(_08297_));
 sg13g2_mux2_1 _16841_ (.A0(_08297_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_58_ ),
    .S(net741),
    .X(_00381_));
 sg13g2_mux2_1 _16842_ (.A0(instr_rdata_i_27_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_91_ ),
    .S(net1988),
    .X(_08298_));
 sg13g2_mux2_1 _16843_ (.A0(_08298_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_59_ ),
    .S(net743),
    .X(_00382_));
 sg13g2_mux2_1 _16844_ (.A0(_07776_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_5_ ),
    .S(net728),
    .X(_00383_));
 sg13g2_mux2_1 _16845_ (.A0(instr_rdata_i_28_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_92_ ),
    .S(net1988),
    .X(_08299_));
 sg13g2_mux2_1 _16846_ (.A0(_08299_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_60_ ),
    .S(net744),
    .X(_00384_));
 sg13g2_mux2_1 _16847_ (.A0(instr_rdata_i_29_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_93_ ),
    .S(net1988),
    .X(_08300_));
 sg13g2_mux2_1 _16848_ (.A0(_08300_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_61_ ),
    .S(net744),
    .X(_00385_));
 sg13g2_mux2_1 _16849_ (.A0(instr_rdata_i_30_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_94_ ),
    .S(net1988),
    .X(_08301_));
 sg13g2_mux2_1 _16850_ (.A0(_08301_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_62_ ),
    .S(net743),
    .X(_00386_));
 sg13g2_mux2_1 _16851_ (.A0(instr_rdata_i_31_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_95_ ),
    .S(net1988),
    .X(_08302_));
 sg13g2_mux2_1 _16852_ (.A0(_08302_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_63_ ),
    .S(net743),
    .X(_00387_));
 sg13g2_mux2_1 _16853_ (.A0(instr_rdata_i_0_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_64_ ),
    .S(net1860),
    .X(_00388_));
 sg13g2_mux2_1 _16854_ (.A0(instr_rdata_i_1_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_65_ ),
    .S(net1860),
    .X(_00389_));
 sg13g2_mux2_1 _16855_ (.A0(instr_rdata_i_2_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_66_ ),
    .S(net1855),
    .X(_00390_));
 sg13g2_mux2_1 _16856_ (.A0(instr_rdata_i_3_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_67_ ),
    .S(net1855),
    .X(_00391_));
 sg13g2_mux2_1 _16857_ (.A0(instr_rdata_i_4_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_68_ ),
    .S(net1856),
    .X(_00392_));
 sg13g2_mux2_1 _16858_ (.A0(instr_rdata_i_5_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_69_ ),
    .S(net1855),
    .X(_00393_));
 sg13g2_mux2_1 _16859_ (.A0(_07788_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_6_ ),
    .S(net728),
    .X(_00394_));
 sg13g2_mux2_1 _16860_ (.A0(instr_rdata_i_6_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_70_ ),
    .S(net1855),
    .X(_00395_));
 sg13g2_mux2_1 _16861_ (.A0(instr_rdata_i_7_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_71_ ),
    .S(net1860),
    .X(_00396_));
 sg13g2_mux2_1 _16862_ (.A0(instr_rdata_i_8_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_72_ ),
    .S(net1855),
    .X(_00397_));
 sg13g2_buf_8 fanout756 (.A(rf_wdata_wb_0_),
    .X(net756));
 sg13g2_mux2_1 _16864_ (.A0(instr_rdata_i_9_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_73_ ),
    .S(net1856),
    .X(_00398_));
 sg13g2_mux2_1 _16865_ (.A0(instr_rdata_i_10_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_74_ ),
    .S(net1855),
    .X(_00399_));
 sg13g2_mux2_1 _16866_ (.A0(instr_rdata_i_11_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_75_ ),
    .S(net1855),
    .X(_00400_));
 sg13g2_mux2_1 _16867_ (.A0(instr_rdata_i_12_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_76_ ),
    .S(net1856),
    .X(_00401_));
 sg13g2_mux2_1 _16868_ (.A0(instr_rdata_i_13_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_77_ ),
    .S(net1856),
    .X(_00402_));
 sg13g2_mux2_1 _16869_ (.A0(instr_rdata_i_14_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_78_ ),
    .S(net1856),
    .X(_00403_));
 sg13g2_mux2_1 _16870_ (.A0(instr_rdata_i_15_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_79_ ),
    .S(net1856),
    .X(_00404_));
 sg13g2_mux2_1 _16871_ (.A0(_07805_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_7_ ),
    .S(net732),
    .X(_00405_));
 sg13g2_mux2_1 _16872_ (.A0(instr_rdata_i_16_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_80_ ),
    .S(net1860),
    .X(_00406_));
 sg13g2_mux2_1 _16873_ (.A0(instr_rdata_i_17_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_81_ ),
    .S(net1860),
    .X(_00407_));
 sg13g2_mux2_1 _16874_ (.A0(instr_rdata_i_18_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_82_ ),
    .S(net1857),
    .X(_00408_));
 sg13g2_buf_8 fanout755 (.A(rf_wdata_wb_0_),
    .X(net755));
 sg13g2_mux2_1 _16876_ (.A0(instr_rdata_i_19_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_83_ ),
    .S(net1857),
    .X(_00409_));
 sg13g2_mux2_1 _16877_ (.A0(instr_rdata_i_20_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_84_ ),
    .S(net1857),
    .X(_00410_));
 sg13g2_mux2_1 _16878_ (.A0(instr_rdata_i_21_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_85_ ),
    .S(net1857),
    .X(_00411_));
 sg13g2_mux2_1 _16879_ (.A0(instr_rdata_i_22_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_86_ ),
    .S(net1857),
    .X(_00412_));
 sg13g2_mux2_1 _16880_ (.A0(instr_rdata_i_23_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_87_ ),
    .S(net1858),
    .X(_00413_));
 sg13g2_mux2_1 _16881_ (.A0(instr_rdata_i_24_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_88_ ),
    .S(net1858),
    .X(_00414_));
 sg13g2_mux2_1 _16882_ (.A0(instr_rdata_i_25_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_89_ ),
    .S(net1858),
    .X(_00415_));
 sg13g2_mux2_1 _16883_ (.A0(_07823_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_8_ ),
    .S(net728),
    .X(_00416_));
 sg13g2_mux2_1 _16884_ (.A0(instr_rdata_i_26_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_90_ ),
    .S(net1855),
    .X(_00417_));
 sg13g2_mux2_1 _16885_ (.A0(instr_rdata_i_27_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_91_ ),
    .S(net1857),
    .X(_00418_));
 sg13g2_mux2_1 _16886_ (.A0(instr_rdata_i_28_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_92_ ),
    .S(net1858),
    .X(_00419_));
 sg13g2_mux2_1 _16887_ (.A0(instr_rdata_i_29_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_93_ ),
    .S(net1858),
    .X(_00420_));
 sg13g2_mux2_1 _16888_ (.A0(instr_rdata_i_30_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_94_ ),
    .S(net1857),
    .X(_00421_));
 sg13g2_mux2_1 _16889_ (.A0(instr_rdata_i_31_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_95_ ),
    .S(net1857),
    .X(_00422_));
 sg13g2_mux2_1 _16890_ (.A0(_07841_),
    .A1(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_9_ ),
    .S(net728),
    .X(_00423_));
 sg13g2_a221oi_1 _16891_ (.B2(_08233_),
    .C1(net105),
    .B1(_08235_),
    .A1(_01512_),
    .Y(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_0_ ),
    .A2(_08236_));
 sg13g2_inv_1 _16892_ (.Y(_08305_),
    .A(_08235_));
 sg13g2_o21ai_1 _16893_ (.B1(net114),
    .Y(_08306_),
    .A1(_08233_),
    .A2(_08305_));
 sg13g2_a21oi_1 _16894_ (.A1(_08233_),
    .A2(_08244_),
    .Y(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_1_ ),
    .B1(_08306_));
 sg13g2_nor3_1 _16895_ (.A(net104),
    .B(_08233_),
    .C(_08244_),
    .Y(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_2_ ));
 sg13g2_inv_1 _16896_ (.Y(_08307_),
    .A(_08034_));
 sg13g2_nand2_1 _16897_ (.Y(_08308_),
    .A(_01471_),
    .B(instr_rvalid_i));
 sg13g2_o21ai_1 _16898_ (.B1(_08308_),
    .Y(_08309_),
    .A1(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .A2(instr_rvalid_i));
 sg13g2_a22oi_1 _16899_ (.Y(\if_stage_i.prefetch_buffer_i.rdata_outstanding_s_0_ ),
    .B1(_08307_),
    .B2(_08309_),
    .A2(_01497_),
    .A1(instr_rvalid_i));
 sg13g2_nor2_1 _16900_ (.A(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ),
    .B(_08035_),
    .Y(_08310_));
 sg13g2_nor2_1 _16901_ (.A(instr_rvalid_i),
    .B(_08310_),
    .Y(\if_stage_i.prefetch_buffer_i.rdata_outstanding_s_1_ ));
 sg13g2_buf_8 fanout754 (.A(rf_wdata_wb_0_),
    .X(net754));
 sg13g2_mux2_2 _16903_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_10_ ),
    .A1(_08067_),
    .S(net1968),
    .X(instr_addr_o_10_));
 sg13g2_nor2_1 _16904_ (.A(instr_gnt_i),
    .B(net1171),
    .Y(_08312_));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_8 fanout752 (.A(net754),
    .X(net752));
 sg13g2_mux2_1 _16907_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_10_ ),
    .A1(instr_addr_o_10_),
    .S(net1143),
    .X(_00424_));
 sg13g2_mux2_2 _16908_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_11_ ),
    .A1(_08076_),
    .S(net1965),
    .X(instr_addr_o_11_));
 sg13g2_mux2_1 _16909_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_11_ ),
    .A1(instr_addr_o_11_),
    .S(net1140),
    .X(_00425_));
 sg13g2_buf_2 fanout751 (.A(rf_wdata_wb_14_),
    .X(net751));
 sg13g2_buf_2 fanout750 (.A(rf_wdata_wb_14_),
    .X(net750));
 sg13g2_nor2_1 _16912_ (.A(net1967),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_12_ ),
    .Y(_08317_));
 sg13g2_a21oi_2 _16913_ (.B1(_08317_),
    .Y(instr_addr_o_12_),
    .A2(_08080_),
    .A1(net1967));
 sg13g2_mux2_1 _16914_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_12_ ),
    .A1(instr_addr_o_12_),
    .S(net1142),
    .X(_00426_));
 sg13g2_mux2_2 _16915_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_13_ ),
    .A1(_08085_),
    .S(net1968),
    .X(instr_addr_o_13_));
 sg13g2_mux2_1 _16916_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_13_ ),
    .A1(instr_addr_o_13_),
    .S(net1143),
    .X(_00427_));
 sg13g2_mux2_2 _16917_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_14_ ),
    .A1(_08099_),
    .S(net1968),
    .X(instr_addr_o_14_));
 sg13g2_mux2_1 _16918_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_14_ ),
    .A1(instr_addr_o_14_),
    .S(net1143),
    .X(_00428_));
 sg13g2_mux2_2 _16919_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_15_ ),
    .A1(_08108_),
    .S(net1965),
    .X(instr_addr_o_15_));
 sg13g2_mux2_1 _16920_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_15_ ),
    .A1(instr_addr_o_15_),
    .S(net1140),
    .X(_00429_));
 sg13g2_nor2_1 _16921_ (.A(net1966),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_16_ ),
    .Y(_08318_));
 sg13g2_a21oi_2 _16922_ (.B1(_08318_),
    .Y(instr_addr_o_16_),
    .A2(_08111_),
    .A1(net1966));
 sg13g2_mux2_1 _16923_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_16_ ),
    .A1(instr_addr_o_16_),
    .S(net1142),
    .X(_00430_));
 sg13g2_nand2_1 _16924_ (.Y(_08319_),
    .A(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_17_ ));
 sg13g2_o21ai_1 _16925_ (.B1(_08319_),
    .Y(instr_addr_o_17_),
    .A1(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .A2(_08115_));
 sg13g2_mux2_1 _16926_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_17_ ),
    .A1(instr_addr_o_17_),
    .S(net1141),
    .X(_00431_));
 sg13g2_nand2_1 _16927_ (.Y(_08320_),
    .A(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_18_ ));
 sg13g2_o21ai_1 _16928_ (.B1(_08320_),
    .Y(instr_addr_o_18_),
    .A1(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .A2(_08121_));
 sg13g2_mux2_1 _16929_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_18_ ),
    .A1(instr_addr_o_18_),
    .S(net1141),
    .X(_00432_));
 sg13g2_mux2_2 _16930_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_19_ ),
    .A1(_08129_),
    .S(net1966),
    .X(instr_addr_o_19_));
 sg13g2_mux2_1 _16931_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_19_ ),
    .A1(instr_addr_o_19_),
    .S(net1142),
    .X(_00433_));
 sg13g2_nor2_1 _16932_ (.A(net1964),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_20_ ),
    .Y(_08321_));
 sg13g2_a21oi_2 _16933_ (.B1(_08321_),
    .Y(instr_addr_o_20_),
    .A2(_08136_),
    .A1(net1964));
 sg13g2_buf_2 fanout749 (.A(rf_wdata_wb_14_),
    .X(net749));
 sg13g2_mux2_1 _16935_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_20_ ),
    .A1(instr_addr_o_20_),
    .S(net1141),
    .X(_00434_));
 sg13g2_nor2_1 _16936_ (.A(net1969),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_21_ ),
    .Y(_08323_));
 sg13g2_a21oi_2 _16937_ (.B1(_08323_),
    .Y(instr_addr_o_21_),
    .A2(_08140_),
    .A1(net1968));
 sg13g2_mux2_1 _16938_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_21_ ),
    .A1(instr_addr_o_21_),
    .S(net1143),
    .X(_00435_));
 sg13g2_mux2_2 _16939_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_22_ ),
    .A1(_08149_),
    .S(net1966),
    .X(instr_addr_o_22_));
 sg13g2_mux2_1 _16940_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_22_ ),
    .A1(instr_addr_o_22_),
    .S(net1142),
    .X(_00436_));
 sg13g2_nor2_1 _16941_ (.A(net1967),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_23_ ),
    .Y(_08324_));
 sg13g2_a21oi_2 _16942_ (.B1(_08324_),
    .Y(instr_addr_o_23_),
    .A2(_08158_),
    .A1(net1967));
 sg13g2_mux2_1 _16943_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_23_ ),
    .A1(instr_addr_o_23_),
    .S(net1142),
    .X(_00437_));
 sg13g2_nor2_1 _16944_ (.A(net1970),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_24_ ),
    .Y(_08325_));
 sg13g2_a21oi_2 _16945_ (.B1(_08325_),
    .Y(instr_addr_o_24_),
    .A2(_08160_),
    .A1(net1964));
 sg13g2_nor3_2 _16946_ (.A(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .B(instr_gnt_i),
    .C(net1171),
    .Y(_08326_));
 sg13g2_nor2_1 _16947_ (.A(\if_stage_i.prefetch_buffer_i.stored_addr_q_24_ ),
    .B(_08326_),
    .Y(_08327_));
 sg13g2_a21oi_1 _16948_ (.A1(_08160_),
    .A2(_08326_),
    .Y(_00438_),
    .B1(_08327_));
 sg13g2_nor2_1 _16949_ (.A(net1967),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_25_ ),
    .Y(_08328_));
 sg13g2_a21oi_2 _16950_ (.B1(_08328_),
    .Y(instr_addr_o_25_),
    .A2(_08165_),
    .A1(net1966));
 sg13g2_mux2_1 _16951_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_25_ ),
    .A1(instr_addr_o_25_),
    .S(net1142),
    .X(_00439_));
 sg13g2_nor2_1 _16952_ (.A(net1966),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_26_ ),
    .Y(_08329_));
 sg13g2_a21oi_2 _16953_ (.B1(_08329_),
    .Y(instr_addr_o_26_),
    .A2(_08176_),
    .A1(net1966));
 sg13g2_mux2_1 _16954_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_26_ ),
    .A1(instr_addr_o_26_),
    .S(net1142),
    .X(_00440_));
 sg13g2_mux2_2 _16955_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_27_ ),
    .A1(_08184_),
    .S(net1965),
    .X(instr_addr_o_27_));
 sg13g2_mux2_1 _16956_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_27_ ),
    .A1(instr_addr_o_27_),
    .S(net1140),
    .X(_00441_));
 sg13g2_mux2_2 _16957_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_28_ ),
    .A1(_08188_),
    .S(net1964),
    .X(instr_addr_o_28_));
 sg13g2_mux2_1 _16958_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_28_ ),
    .A1(_08188_),
    .S(_08326_),
    .X(_00442_));
 sg13g2_mux2_2 _16959_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_29_ ),
    .A1(_08191_),
    .S(net1966),
    .X(instr_addr_o_29_));
 sg13g2_mux2_1 _16960_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_29_ ),
    .A1(instr_addr_o_29_),
    .S(net1142),
    .X(_00443_));
 sg13g2_mux2_2 _16961_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_2_ ),
    .A1(_08194_),
    .S(net1964),
    .X(instr_addr_o_2_));
 sg13g2_mux2_1 _16962_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_2_ ),
    .A1(instr_addr_o_2_),
    .S(net1141),
    .X(_00444_));
 sg13g2_mux2_2 _16963_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_30_ ),
    .A1(_08199_),
    .S(net1968),
    .X(instr_addr_o_30_));
 sg13g2_mux2_1 _16964_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_30_ ),
    .A1(instr_addr_o_30_),
    .S(net1143),
    .X(_00445_));
 sg13g2_mux2_2 _16965_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_31_ ),
    .A1(_08204_),
    .S(net1964),
    .X(instr_addr_o_31_));
 sg13g2_mux2_1 _16966_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_31_ ),
    .A1(instr_addr_o_31_),
    .S(net1140),
    .X(_00446_));
 sg13g2_nor2_1 _16967_ (.A(net1965),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_3_ ),
    .Y(_08330_));
 sg13g2_a21oi_2 _16968_ (.B1(_08330_),
    .Y(instr_addr_o_3_),
    .A2(_08206_),
    .A1(net1965));
 sg13g2_mux2_1 _16969_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_3_ ),
    .A1(instr_addr_o_3_),
    .S(net1140),
    .X(_00447_));
 sg13g2_mux2_2 _16970_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_4_ ),
    .A1(_08049_),
    .S(net1968),
    .X(instr_addr_o_4_));
 sg13g2_mux2_1 _16971_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_4_ ),
    .A1(instr_addr_o_4_),
    .S(net1143),
    .X(_00448_));
 sg13g2_mux2_2 _16972_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_5_ ),
    .A1(_08048_),
    .S(net1964),
    .X(instr_addr_o_5_));
 sg13g2_mux2_1 _16973_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_5_ ),
    .A1(instr_addr_o_5_),
    .S(net1140),
    .X(_00449_));
 sg13g2_mux2_2 _16974_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_6_ ),
    .A1(_08047_),
    .S(net1968),
    .X(instr_addr_o_6_));
 sg13g2_mux2_1 _16975_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_6_ ),
    .A1(instr_addr_o_6_),
    .S(net1143),
    .X(_00450_));
 sg13g2_nor2_1 _16976_ (.A(net1964),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_7_ ),
    .Y(_08331_));
 sg13g2_a21oi_2 _16977_ (.B1(_08331_),
    .Y(instr_addr_o_7_),
    .A2(_08044_),
    .A1(net1970));
 sg13g2_mux2_1 _16978_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_7_ ),
    .A1(instr_addr_o_7_),
    .S(net1140),
    .X(_00451_));
 sg13g2_mux2_2 _16979_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_8_ ),
    .A1(_08061_),
    .S(net1968),
    .X(instr_addr_o_8_));
 sg13g2_mux2_1 _16980_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_8_ ),
    .A1(instr_addr_o_8_),
    .S(net1143),
    .X(_00452_));
 sg13g2_nor2_1 _16981_ (.A(net1965),
    .B(\if_stage_i.prefetch_buffer_i.stored_addr_q_9_ ),
    .Y(_08332_));
 sg13g2_a21oi_2 _16982_ (.B1(_08332_),
    .Y(instr_addr_o_9_),
    .A2(_08042_),
    .A1(net1965));
 sg13g2_mux2_1 _16983_ (.A0(\if_stage_i.prefetch_buffer_i.stored_addr_q_9_ ),
    .A1(instr_addr_o_9_),
    .S(net1140),
    .X(_00453_));
 sg13g2_nor2b_1 _16984_ (.A(instr_gnt_i),
    .B_N(instr_req_o),
    .Y(\if_stage_i.prefetch_buffer_i.valid_req_d ));
 sg13g2_inv_1 _16985_ (.Y(_08333_),
    .A(\load_store_unit_i.data_sign_ext_q ));
 sg13g2_nor2b_1 _16986_ (.A(_03230_),
    .B_N(_03221_),
    .Y(_08334_));
 sg13g2_a21o_2 _16987_ (.A2(_03218_),
    .A1(data_gnt_i),
    .B1(_08334_),
    .X(_08335_));
 sg13g2_buf_1 fanout748 (.A(net749),
    .X(net748));
 sg13g2_nand4_1 _16989_ (.B(_01139_),
    .C(net1906),
    .A(net2087),
    .Y(_08337_),
    .D(_08335_));
 sg13g2_o21ai_1 _16990_ (.B1(_08337_),
    .Y(_00454_),
    .A1(_08333_),
    .A2(_08335_));
 sg13g2_nor2_2 _16991_ (.A(_01162_),
    .B(_01373_),
    .Y(_08338_));
 sg13g2_mux2_1 _16992_ (.A0(\load_store_unit_i.data_type_q_0_ ),
    .A1(_08338_),
    .S(_08335_),
    .X(_00455_));
 sg13g2_mux2_1 _16993_ (.A0(\load_store_unit_i.data_type_q_1_ ),
    .A1(_03872_),
    .S(_08335_),
    .X(_00456_));
 sg13g2_mux2_1 _16994_ (.A0(\load_store_unit_i.data_we_q ),
    .A1(data_we_o),
    .S(_08335_),
    .X(_00457_));
 sg13g2_inv_1 _16995_ (.Y(_08339_),
    .A(_03222_));
 sg13g2_o21ai_1 _16996_ (.B1(net1147),
    .Y(_08340_),
    .A1(_03239_),
    .A2(_08338_));
 sg13g2_nor2_1 _16997_ (.A(_01373_),
    .B(net1113),
    .Y(_08341_));
 sg13g2_o21ai_1 _16998_ (.B1(_03859_),
    .Y(_08342_),
    .A1(_03858_),
    .A2(_08341_));
 sg13g2_nand2_2 _16999_ (.Y(_08343_),
    .A(_08340_),
    .B(_08342_));
 sg13g2_nand2_1 _17000_ (.Y(_08344_),
    .A(_03876_),
    .B(_03230_));
 sg13g2_nor2_1 _17001_ (.A(\load_store_unit_i.ls_fsm_cs_1_ ),
    .B(_03220_),
    .Y(_08345_));
 sg13g2_nand2b_2 _17002_ (.Y(_08346_),
    .B(_01770_),
    .A_N(net1977));
 sg13g2_nor3_1 _17003_ (.A(data_gnt_i),
    .B(_01564_),
    .C(_08346_),
    .Y(_08347_));
 sg13g2_a21oi_1 _17004_ (.A1(_08344_),
    .A2(_08345_),
    .Y(_08348_),
    .B1(_08347_));
 sg13g2_o21ai_1 _17005_ (.B1(_08348_),
    .Y(_08349_),
    .A1(_08339_),
    .A2(_08343_));
 sg13g2_nor4_1 _17006_ (.A(data_rvalid_i),
    .B(\load_store_unit_i.pmp_err_q ),
    .C(data_gnt_i),
    .D(_08346_),
    .Y(_08350_));
 sg13g2_nor2_1 _17007_ (.A(_01625_),
    .B(_03217_),
    .Y(_08351_));
 sg13g2_nor3_1 _17008_ (.A(net1976),
    .B(\load_store_unit_i.ls_fsm_cs_0__$_NOT__A_Y ),
    .C(_01141_),
    .Y(_08352_));
 sg13g2_o21ai_1 _17009_ (.B1(_03224_),
    .Y(_08353_),
    .A1(_01495_),
    .A2(_08352_));
 sg13g2_o21ai_1 _17010_ (.B1(_08353_),
    .Y(_08354_),
    .A1(_01495_),
    .A2(_08339_));
 sg13g2_nor3_1 _17011_ (.A(_08350_),
    .B(_08351_),
    .C(_08354_),
    .Y(_08355_));
 sg13g2_mux2_1 _17012_ (.A0(\load_store_unit_i.handle_misaligned_q ),
    .A1(_08349_),
    .S(_08355_),
    .X(_00458_));
 sg13g2_o21ai_1 _17013_ (.B1(_01625_),
    .Y(_08356_),
    .A1(_01564_),
    .A2(_08346_));
 sg13g2_nand2_1 _17014_ (.Y(_08357_),
    .A(_03224_),
    .B(_08356_));
 sg13g2_nor2_1 _17015_ (.A(net2466),
    .B(_01144_),
    .Y(_08358_));
 sg13g2_and2_1 _17016_ (.A(_03230_),
    .B(_03221_),
    .X(_08359_));
 sg13g2_or4_2 _17017_ (.A(_08350_),
    .B(_08351_),
    .C(_08358_),
    .D(_08359_),
    .X(_08360_));
 sg13g2_nand2_1 _17018_ (.Y(_08361_),
    .A(net1977),
    .B(_08360_));
 sg13g2_o21ai_1 _17019_ (.B1(_08361_),
    .Y(_00459_),
    .A1(_08357_),
    .A2(_08360_));
 sg13g2_xnor2_1 _17020_ (.Y(_08362_),
    .A(data_gnt_i),
    .B(_08343_));
 sg13g2_nor2_1 _17021_ (.A(_08347_),
    .B(_08345_),
    .Y(_08363_));
 sg13g2_o21ai_1 _17022_ (.B1(_08363_),
    .Y(_08364_),
    .A1(_01625_),
    .A2(_08362_));
 sg13g2_mux2_1 _17023_ (.A0(_08364_),
    .A1(\load_store_unit_i.ls_fsm_cs_1_ ),
    .S(_08360_),
    .X(_00460_));
 sg13g2_nor4_1 _17024_ (.A(net2466),
    .B(net1976),
    .C(_08346_),
    .D(_08360_),
    .Y(_08365_));
 sg13g2_a21o_1 _17025_ (.A2(_08360_),
    .A1(\load_store_unit_i.ls_fsm_cs_2_ ),
    .B1(_08365_),
    .X(_00461_));
 sg13g2_a22oi_1 _17026_ (.Y(_08366_),
    .B1(_01595_),
    .B2(_03219_),
    .A2(_01771_),
    .A1(data_err_i));
 sg13g2_a21oi_1 _17027_ (.A1(_01144_),
    .A2(_03225_),
    .Y(_08367_),
    .B1(net2466));
 sg13g2_and2_1 _17028_ (.A(_08346_),
    .B(_03223_),
    .X(_08368_));
 sg13g2_nor3_1 _17029_ (.A(_08351_),
    .B(_08367_),
    .C(_08368_),
    .Y(_08369_));
 sg13g2_nor2_1 _17030_ (.A(\load_store_unit_i.lsu_err_q ),
    .B(_08369_),
    .Y(_08370_));
 sg13g2_a21oi_1 _17031_ (.A1(_08366_),
    .A2(_08369_),
    .Y(_00462_),
    .B1(_08370_));
 sg13g2_nor2b_1 _17032_ (.A(data_we_o),
    .B_N(_03218_),
    .Y(\load_store_unit_i.perf_load_o ));
 sg13g2_and2_1 _17033_ (.A(_03218_),
    .B(data_we_o),
    .X(\load_store_unit_i.perf_store_o ));
 sg13g2_o21ai_1 _17034_ (.B1(net1976),
    .Y(_08371_),
    .A1(_08358_),
    .A2(_08368_));
 sg13g2_inv_1 _17035_ (.Y(_00463_),
    .A(_08371_));
 sg13g2_nor2_1 _17036_ (.A(\load_store_unit_i.rdata_offset_q_0_ ),
    .B(_08335_),
    .Y(_08372_));
 sg13g2_a21oi_1 _17037_ (.A1(net1147),
    .A2(_08335_),
    .Y(_00464_),
    .B1(_08372_));
 sg13g2_mux2_1 _17038_ (.A0(\load_store_unit_i.rdata_offset_q_1_ ),
    .A1(net1113),
    .S(_08335_),
    .X(_00465_));
 sg13g2_a21oi_1 _17039_ (.A1(net1976),
    .A2(_01144_),
    .Y(_08373_),
    .B1(net2466));
 sg13g2_o21ai_1 _17040_ (.B1(\load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ),
    .Y(_08374_),
    .A1(_01771_),
    .A2(_03219_));
 sg13g2_nor2_1 _17041_ (.A(_08373_),
    .B(_08374_),
    .Y(_08375_));
 sg13g2_buf_2 fanout747 (.A(net749),
    .X(net747));
 sg13g2_mux2_1 _17043_ (.A0(\load_store_unit_i.rdata_q_0_ ),
    .A1(data_rdata_i_8_),
    .S(net1653),
    .X(_00466_));
 sg13g2_mux2_1 _17044_ (.A0(\load_store_unit_i.rdata_q_10_ ),
    .A1(data_rdata_i_18_),
    .S(net1652),
    .X(_00467_));
 sg13g2_mux2_1 _17045_ (.A0(\load_store_unit_i.rdata_q_11_ ),
    .A1(data_rdata_i_19_),
    .S(net1654),
    .X(_00468_));
 sg13g2_mux2_1 _17046_ (.A0(\load_store_unit_i.rdata_q_12_ ),
    .A1(data_rdata_i_20_),
    .S(net1654),
    .X(_00469_));
 sg13g2_mux2_1 _17047_ (.A0(\load_store_unit_i.rdata_q_13_ ),
    .A1(data_rdata_i_21_),
    .S(net1654),
    .X(_00470_));
 sg13g2_mux2_1 _17048_ (.A0(\load_store_unit_i.rdata_q_14_ ),
    .A1(data_rdata_i_22_),
    .S(net1653),
    .X(_00471_));
 sg13g2_mux2_1 _17049_ (.A0(\load_store_unit_i.rdata_q_15_ ),
    .A1(data_rdata_i_23_),
    .S(net1652),
    .X(_00472_));
 sg13g2_mux2_1 _17050_ (.A0(\load_store_unit_i.rdata_q_16_ ),
    .A1(data_rdata_i_24_),
    .S(net1653),
    .X(_00473_));
 sg13g2_mux2_1 _17051_ (.A0(\load_store_unit_i.rdata_q_17_ ),
    .A1(data_rdata_i_25_),
    .S(net1654),
    .X(_00474_));
 sg13g2_mux2_1 _17052_ (.A0(\load_store_unit_i.rdata_q_18_ ),
    .A1(data_rdata_i_26_),
    .S(net1652),
    .X(_00475_));
 sg13g2_buf_8 fanout746 (.A(_08245_),
    .X(net746));
 sg13g2_mux2_1 _17054_ (.A0(\load_store_unit_i.rdata_q_19_ ),
    .A1(data_rdata_i_27_),
    .S(net1654),
    .X(_00476_));
 sg13g2_mux2_1 _17055_ (.A0(\load_store_unit_i.rdata_q_1_ ),
    .A1(data_rdata_i_9_),
    .S(net1655),
    .X(_00477_));
 sg13g2_mux2_1 _17056_ (.A0(\load_store_unit_i.rdata_q_20_ ),
    .A1(data_rdata_i_28_),
    .S(net1655),
    .X(_00478_));
 sg13g2_mux2_1 _17057_ (.A0(\load_store_unit_i.rdata_q_21_ ),
    .A1(data_rdata_i_29_),
    .S(net1655),
    .X(_00479_));
 sg13g2_mux2_1 _17058_ (.A0(\load_store_unit_i.rdata_q_22_ ),
    .A1(data_rdata_i_30_),
    .S(net1653),
    .X(_00480_));
 sg13g2_mux2_1 _17059_ (.A0(\load_store_unit_i.rdata_q_23_ ),
    .A1(data_rdata_i_31_),
    .S(net1652),
    .X(_00481_));
 sg13g2_mux2_1 _17060_ (.A0(\load_store_unit_i.rdata_q_2_ ),
    .A1(data_rdata_i_10_),
    .S(net1652),
    .X(_00482_));
 sg13g2_mux2_1 _17061_ (.A0(\load_store_unit_i.rdata_q_3_ ),
    .A1(data_rdata_i_11_),
    .S(net1654),
    .X(_00483_));
 sg13g2_mux2_1 _17062_ (.A0(\load_store_unit_i.rdata_q_4_ ),
    .A1(data_rdata_i_12_),
    .S(net1654),
    .X(_00484_));
 sg13g2_mux2_1 _17063_ (.A0(\load_store_unit_i.rdata_q_5_ ),
    .A1(data_rdata_i_13_),
    .S(net1653),
    .X(_00485_));
 sg13g2_mux2_1 _17064_ (.A0(\load_store_unit_i.rdata_q_6_ ),
    .A1(data_rdata_i_14_),
    .S(net1652),
    .X(_00486_));
 sg13g2_mux2_1 _17065_ (.A0(\load_store_unit_i.rdata_q_7_ ),
    .A1(data_rdata_i_15_),
    .S(net1652),
    .X(_00487_));
 sg13g2_mux2_1 _17066_ (.A0(\load_store_unit_i.rdata_q_8_ ),
    .A1(data_rdata_i_16_),
    .S(net1652),
    .X(_00488_));
 sg13g2_mux2_1 _17067_ (.A0(\load_store_unit_i.rdata_q_9_ ),
    .A1(data_rdata_i_17_),
    .S(net1654),
    .X(_00489_));
 sg13g2_nor3_1 _17068_ (.A(_01573_),
    .B(_01403_),
    .C(_01584_),
    .Y(_08378_));
 sg13g2_nor2_1 _17069_ (.A(_01401_),
    .B(_01419_),
    .Y(_08379_));
 sg13g2_o21ai_1 _17070_ (.B1(_01450_),
    .Y(_08380_),
    .A1(_08378_),
    .A2(_08379_));
 sg13g2_nand2_1 _17071_ (.Y(_08381_),
    .A(_01626_),
    .B(_01599_));
 sg13g2_nor2_1 _17072_ (.A(\id_stage_i.illegal_csr_insn_i ),
    .B(_01568_),
    .Y(_08382_));
 sg13g2_nand4_1 _17073_ (.B(_08380_),
    .C(_08381_),
    .A(\id_stage_i.instr_perf_count_id_o_$_AND__Y_B ),
    .Y(_08383_),
    .D(_08382_));
 sg13g2_nor3_2 _17074_ (.A(_01633_),
    .B(_03193_),
    .C(_08383_),
    .Y(perf_instr_ret_wb));
 sg13g2_and2_1 _17075_ (.A(net438),
    .B(perf_instr_ret_wb),
    .X(perf_instr_ret_compressed_wb));
 sg13g2_nor2_1 _17076_ (.A(_07425_),
    .B(_03195_),
    .Y(perf_iside_wait));
 sg13g2_and4_1 _17077_ (.A(net2466),
    .B(\load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ),
    .C(_01495_),
    .D(_01596_),
    .X(_08384_));
 sg13g2_buf_16 fanout745 (.X(net745),
    .A(net746));
 sg13g2_a21oi_1 _17079_ (.A1(\load_store_unit_i.data_type_q_0_ ),
    .A2(\load_store_unit_i.data_type_q_0__$_NOT__A_Y ),
    .Y(_08386_),
    .B1(\load_store_unit_i.data_type_q_1__$_NOT__A_Y ));
 sg13g2_buf_16 fanout744 (.X(net744),
    .A(net745));
 sg13g2_or2_1 _17081_ (.X(_08388_),
    .B(\load_store_unit_i.data_type_q_1_ ),
    .A(\load_store_unit_i.data_type_q_0__$_NOT__A_Y ));
 sg13g2_buf_16 fanout743 (.X(net743),
    .A(net745));
 sg13g2_nand2b_1 _17083_ (.Y(_08390_),
    .B(net1959),
    .A_N(net1961));
 sg13g2_buf_16 fanout742 (.X(net742),
    .A(net745));
 sg13g2_nor2_1 _17085_ (.A(\load_store_unit_i.rdata_offset_q_0__$_NOT__A_Y ),
    .B(\load_store_unit_i.rdata_offset_q_1_ ),
    .Y(_08392_));
 sg13g2_buf_16 fanout741 (.X(net741),
    .A(net745));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(rf_wdata_wb_20_));
 sg13g2_nor2_1 _17088_ (.A(\load_store_unit_i.rdata_offset_q_0__$_NOT__A_Y ),
    .B(\load_store_unit_i.rdata_offset_q_1__$_NOT__A_Y ),
    .Y(_08395_));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_1 fanout738 (.A(net739),
    .X(net738));
 sg13g2_nor2_1 _17091_ (.A(\load_store_unit_i.rdata_offset_q_0_ ),
    .B(\load_store_unit_i.rdata_offset_q_1__$_NOT__A_Y ),
    .Y(_08398_));
 sg13g2_buf_1 fanout737 (.A(net738),
    .X(net737));
 sg13g2_buf_2 fanout736 (.A(net737),
    .X(net736));
 sg13g2_and2_1 _17094_ (.A(\load_store_unit_i.rdata_q_8_ ),
    .B(net1937),
    .X(_08401_));
 sg13g2_a221oi_1 _17095_ (.B2(\load_store_unit_i.rdata_q_16_ ),
    .C1(_08401_),
    .B1(net1945),
    .A1(\load_store_unit_i.rdata_q_0_ ),
    .Y(_08402_),
    .A2(net1953));
 sg13g2_nor2_1 _17096_ (.A(\load_store_unit_i.data_type_q_0__$_NOT__A_Y ),
    .B(\load_store_unit_i.data_type_q_1_ ),
    .Y(_08403_));
 sg13g2_nor2_2 _17097_ (.A(net1960),
    .B(net1931),
    .Y(_08404_));
 sg13g2_a22oi_1 _17098_ (.Y(_08405_),
    .B1(net1953),
    .B2(data_rdata_i_8_),
    .A2(net1937),
    .A1(data_rdata_i_16_));
 sg13g2_a22oi_1 _17099_ (.Y(_08406_),
    .B1(net1933),
    .B2(\load_store_unit_i.rdata_q_16_ ),
    .A2(net1962),
    .A1(data_rdata_i_24_));
 sg13g2_nand2b_1 _17100_ (.Y(_08407_),
    .B(net1945),
    .A_N(_08406_));
 sg13g2_o21ai_1 _17101_ (.B1(_08407_),
    .Y(_08408_),
    .A1(net1704),
    .A2(_08405_));
 sg13g2_nor3_1 _17102_ (.A(net1938),
    .B(net1954),
    .C(net1946),
    .Y(_08409_));
 sg13g2_buf_8 fanout735 (.A(\cs_registers_i/_2062_ ),
    .X(net735));
 sg13g2_buf_1 fanout734 (.A(net735),
    .X(net734));
 sg13g2_nand2b_1 _17105_ (.Y(_08412_),
    .B(net414),
    .A_N(data_rdata_i_0_));
 sg13g2_o21ai_1 _17106_ (.B1(_08412_),
    .Y(_08413_),
    .A1(_08408_),
    .A2(net413));
 sg13g2_o21ai_1 _17107_ (.B1(_08413_),
    .Y(_08414_),
    .A1(net1707),
    .A2(_08402_));
 sg13g2_nand4_1 _17108_ (.B(net1581),
    .C(_01682_),
    .A(_01719_),
    .Y(_08415_),
    .D(_01738_));
 sg13g2_and2_1 _17109_ (.A(_01752_),
    .B(_08415_),
    .X(_08416_));
 sg13g2_and2_1 _17110_ (.A(_01732_),
    .B(_02840_),
    .X(_08417_));
 sg13g2_inv_1 _17111_ (.Y(_08418_),
    .A(_08417_));
 sg13g2_nor2_1 _17112_ (.A(_01703_),
    .B(_08418_),
    .Y(_08419_));
 sg13g2_a21oi_1 _17113_ (.A1(_08416_),
    .A2(_08419_),
    .Y(_08420_),
    .B1(_01742_));
 sg13g2_a21oi_1 _17114_ (.A1(_01719_),
    .A2(_01682_),
    .Y(_08421_),
    .B1(_01697_));
 sg13g2_a22oi_1 _17115_ (.Y(_08422_),
    .B1(_08421_),
    .B2(_01663_),
    .A2(_01697_),
    .A1(_01662_));
 sg13g2_and2_1 _17116_ (.A(_01724_),
    .B(_02840_),
    .X(_08423_));
 sg13g2_nand2_1 _17117_ (.Y(_08424_),
    .A(_01722_),
    .B(_08423_));
 sg13g2_nor2_1 _17118_ (.A(_08422_),
    .B(_08424_),
    .Y(_08425_));
 sg13g2_buf_8 fanout733 (.A(net735),
    .X(net733));
 sg13g2_buf_8 fanout732 (.A(_08237_),
    .X(net732));
 sg13g2_a21oi_1 _17121_ (.A1(net1247),
    .A2(net1457),
    .Y(_08428_),
    .B1(_01187_));
 sg13g2_xnor2_1 _17122_ (.Y(_08429_),
    .A(_02328_),
    .B(_08428_));
 sg13g2_buf_16 fanout731 (.X(net731),
    .A(net732));
 sg13g2_buf_16 fanout730 (.X(net730),
    .A(net731));
 sg13g2_buf_16 fanout729 (.X(net729),
    .A(net732));
 sg13g2_nor2_1 _17126_ (.A(_01187_),
    .B(net1460),
    .Y(_08433_));
 sg13g2_xnor2_1 _17127_ (.Y(_08434_),
    .A(net1247),
    .B(_08433_));
 sg13g2_buf_16 fanout728 (.X(net728),
    .A(net732));
 sg13g2_buf_2 fanout727 (.A(rf_wdata_wb_17_),
    .X(net727));
 sg13g2_buf_2 fanout726 (.A(net727),
    .X(net726));
 sg13g2_and3_2 _17131_ (.X(_08438_),
    .A(_01662_),
    .B(_01722_),
    .C(_08421_));
 sg13g2_nand3_1 _17132_ (.B(_02840_),
    .C(_08438_),
    .A(_01744_),
    .Y(_08439_));
 sg13g2_buf_2 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_2 fanout724 (.A(net727),
    .X(net724));
 sg13g2_mux4_1 _17135_ (.S0(net1462),
    .A0(net1201),
    .A1(net1199),
    .A2(net1408),
    .A3(net1409),
    .S1(net211),
    .X(_08442_));
 sg13g2_and3_1 _17136_ (.X(_08443_),
    .A(_01744_),
    .B(_02840_),
    .C(_08438_));
 sg13g2_buf_2 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout722 (.A(\cs_registers_i/_0580_ ),
    .X(net722));
 sg13g2_buf_8 fanout721 (.A(\cs_registers_i/_1926_ ),
    .X(net721));
 sg13g2_mux4_1 _17140_ (.S0(net201),
    .A0(net1411),
    .A1(net1190),
    .A2(net198),
    .A3(alu_operand_a_ex_31_),
    .S1(net1458),
    .X(_08447_));
 sg13g2_nor2b_1 _17141_ (.A(net1178),
    .B_N(_08447_),
    .Y(_08448_));
 sg13g2_a21oi_1 _17142_ (.A1(net1178),
    .A2(_08442_),
    .Y(_08449_),
    .B1(_08448_));
 sg13g2_buf_8 fanout720 (.A(\cs_registers_i/_1934_ ),
    .X(net720));
 sg13g2_mux4_1 _17144_ (.S0(net1461),
    .A0(net87),
    .A1(net124),
    .A2(net1404),
    .A3(net1407),
    .S1(net211),
    .X(_08451_));
 sg13g2_mux4_1 _17145_ (.S0(net1461),
    .A0(net125),
    .A1(net1202),
    .A2(net148),
    .A3(net1350),
    .S1(net211),
    .X(_08452_));
 sg13g2_buf_8 fanout719 (.A(\cs_registers_i/_2068_ ),
    .X(net719));
 sg13g2_buf_1 fanout718 (.A(net719),
    .X(net718));
 sg13g2_mux2_1 _17148_ (.A0(_08451_),
    .A1(_08452_),
    .S(net1179),
    .X(_08455_));
 sg13g2_nor2_1 _17149_ (.A(net1164),
    .B(_08455_),
    .Y(_08456_));
 sg13g2_a21oi_1 _17150_ (.A1(net1164),
    .A2(_08449_),
    .Y(_08457_),
    .B1(_08456_));
 sg13g2_and3_1 _17151_ (.X(_08458_),
    .A(_02412_),
    .B(net1247),
    .C(net1457));
 sg13g2_nor2_1 _17152_ (.A(_01187_),
    .B(_08458_),
    .Y(_08459_));
 sg13g2_xnor2_1 _17153_ (.Y(_08460_),
    .A(_02287_),
    .B(_08459_));
 sg13g2_buf_2 fanout717 (.A(net719),
    .X(net717));
 sg13g2_mux4_1 _17155_ (.S0(net1460),
    .A0(net195),
    .A1(net150),
    .A2(net194),
    .A3(net1279),
    .S1(net210),
    .X(_08462_));
 sg13g2_mux4_1 _17156_ (.S0(_03067_),
    .A0(net151),
    .A1(net1415),
    .A2(net126),
    .A3(net1281),
    .S1(net205),
    .X(_08463_));
 sg13g2_mux2_1 _17157_ (.A0(_08462_),
    .A1(_08463_),
    .S(net1177),
    .X(_08464_));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(\cs_registers_i/_2109_ ));
 sg13g2_buf_2 fanout715 (.A(net716),
    .X(net715));
 sg13g2_mux4_1 _17160_ (.S0(_03067_),
    .A0(net1413),
    .A1(net1352),
    .A2(_01248_),
    .A3(net1203),
    .S1(net205),
    .X(_08467_));
 sg13g2_mux4_1 _17161_ (.S0(net200),
    .A0(net1351),
    .A1(alu_operand_a_ex_16_),
    .A2(net1283),
    .A3(net1250),
    .S1(net1460),
    .X(_08468_));
 sg13g2_mux2_1 _17162_ (.A0(_08467_),
    .A1(_08468_),
    .S(net1177),
    .X(_08469_));
 sg13g2_nor2b_1 _17163_ (.A(net1164),
    .B_N(_08469_),
    .Y(_08470_));
 sg13g2_a21oi_1 _17164_ (.A1(_08464_),
    .A2(net1164),
    .Y(_08471_),
    .B1(_08470_));
 sg13g2_nor2_1 _17165_ (.A(_08471_),
    .B(net1137),
    .Y(_08472_));
 sg13g2_a21oi_1 _17166_ (.A1(_08457_),
    .A2(net1137),
    .Y(_08473_),
    .B1(_08472_));
 sg13g2_a21oi_1 _17167_ (.A1(_03244_),
    .A2(_08458_),
    .Y(_08474_),
    .B1(_01187_));
 sg13g2_xnor2_1 _17168_ (.Y(_08475_),
    .A(_02261_),
    .B(_08474_));
 sg13g2_buf_8 fanout714 (.A(\cs_registers_i/_2125_ ),
    .X(net714));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(\cs_registers_i/_2166_ ));
 sg13g2_mux4_1 _17171_ (.S0(net1460),
    .A0(net1283),
    .A1(net1351),
    .A2(net1250),
    .A3(alu_operand_a_ex_16_),
    .S1(net210),
    .X(_08478_));
 sg13g2_mux4_1 _17172_ (.S0(net1460),
    .A0(net1413),
    .A1(net1352),
    .A2(_01248_),
    .A3(net1203),
    .S1(net210),
    .X(_08479_));
 sg13g2_mux2_1 _17173_ (.A0(_08478_),
    .A1(_08479_),
    .S(net1177),
    .X(_08480_));
 sg13g2_mux4_1 _17174_ (.S0(net1460),
    .A0(net151),
    .A1(net1415),
    .A2(net127),
    .A3(net1281),
    .S1(net210),
    .X(_08481_));
 sg13g2_mux4_1 _17175_ (.S0(net200),
    .A0(net149),
    .A1(net1279),
    .A2(net196),
    .A3(net194),
    .S1(net1461),
    .X(_08482_));
 sg13g2_mux2_1 _17176_ (.A0(_08481_),
    .A1(_08482_),
    .S(net1177),
    .X(_08483_));
 sg13g2_nor2b_1 _17177_ (.A(net1164),
    .B_N(_08483_),
    .Y(_08484_));
 sg13g2_a21oi_1 _17178_ (.A1(net1164),
    .A2(_08480_),
    .Y(_08485_),
    .B1(_08484_));
 sg13g2_mux4_1 _17179_ (.S0(net199),
    .A0(net1199),
    .A1(net1409),
    .A2(net1201),
    .A3(net1408),
    .S1(net1461),
    .X(_08486_));
 sg13g2_nand2b_1 _17180_ (.Y(_08487_),
    .B(net199),
    .A_N(net197));
 sg13g2_o21ai_1 _17181_ (.B1(_08487_),
    .Y(_08488_),
    .A1(net81),
    .A2(net199));
 sg13g2_nor2_1 _17182_ (.A(net1190),
    .B(net203),
    .Y(_08489_));
 sg13g2_a21oi_1 _17183_ (.A1(_02331_),
    .A2(net203),
    .Y(_08490_),
    .B1(_08489_));
 sg13g2_nand2_1 _17184_ (.Y(_08491_),
    .A(net1458),
    .B(_08490_));
 sg13g2_o21ai_1 _17185_ (.B1(_08491_),
    .Y(_08492_),
    .A1(net1458),
    .A2(_08488_));
 sg13g2_mux2_2 _17186_ (.A0(_08486_),
    .A1(_08492_),
    .S(net1179),
    .X(_08493_));
 sg13g2_mux4_1 _17187_ (.S0(net200),
    .A0(net1202),
    .A1(net1350),
    .A2(net125),
    .A3(net148),
    .S1(net1461),
    .X(_08494_));
 sg13g2_mux4_1 _17188_ (.S0(net199),
    .A0(net123),
    .A1(net1407),
    .A2(net88),
    .A3(net1404),
    .S1(net1461),
    .X(_08495_));
 sg13g2_mux2_1 _17189_ (.A0(_08494_),
    .A1(_08495_),
    .S(net1179),
    .X(_08496_));
 sg13g2_mux2_1 _17190_ (.A0(_08493_),
    .A1(_08496_),
    .S(net1168),
    .X(_08497_));
 sg13g2_nor2_1 _17191_ (.A(net1137),
    .B(_08497_),
    .Y(_08498_));
 sg13g2_a21oi_1 _17192_ (.A1(net1137),
    .A2(_08485_),
    .Y(_08499_),
    .B1(_08498_));
 sg13g2_nand2_1 _17193_ (.Y(_08500_),
    .A(_08499_),
    .B(net1135));
 sg13g2_o21ai_1 _17194_ (.B1(_08500_),
    .Y(_08501_),
    .A1(_08473_),
    .A2(net1134));
 sg13g2_xnor2_1 _17195_ (.Y(_08502_),
    .A(_03244_),
    .B(_08459_));
 sg13g2_nor2_2 _17196_ (.A(net45),
    .B(net1134),
    .Y(_08503_));
 sg13g2_buf_8 fanout712 (.A(net713),
    .X(net712));
 sg13g2_nand2_2 _17198_ (.Y(_08505_),
    .A(_08423_),
    .B(_08438_));
 sg13g2_nor2b_1 _17199_ (.A(net1180),
    .B_N(net1165),
    .Y(_08506_));
 sg13g2_nand2_1 _17200_ (.Y(_08507_),
    .A(net1462),
    .B(_08506_));
 sg13g2_a21oi_1 _17201_ (.A1(_08505_),
    .A2(_08507_),
    .Y(_08508_),
    .B1(_08488_));
 sg13g2_or2_2 _17202_ (.X(_08509_),
    .B(_08505_),
    .A(_08488_));
 sg13g2_nor2_2 _17203_ (.A(_08509_),
    .B(net1120),
    .Y(_08510_));
 sg13g2_a21o_1 _17204_ (.A2(_08508_),
    .A1(net1120),
    .B1(_08510_),
    .X(_08511_));
 sg13g2_buf_8 fanout711 (.A(rf_wdata_wb_16_),
    .X(net711));
 sg13g2_mux2_1 _17206_ (.A0(_08501_),
    .A1(_08511_),
    .S(net201),
    .X(_08513_));
 sg13g2_nor2_1 _17207_ (.A(_01722_),
    .B(_01758_),
    .Y(_08514_));
 sg13g2_nor3_1 _17208_ (.A(_01704_),
    .B(_08514_),
    .C(_08418_),
    .Y(_08515_));
 sg13g2_buf_16 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_8 fanout709 (.A(rf_wdata_wb_16_),
    .X(net709));
 sg13g2_or2_1 _17211_ (.X(_08518_),
    .B(_02841_),
    .A(_01702_));
 sg13g2_or3_1 _17212_ (.A(_01685_),
    .B(_01722_),
    .C(_08518_),
    .X(_08519_));
 sg13g2_buf_8 fanout708 (.A(rf_wdata_wb_16_),
    .X(net708));
 sg13g2_xnor2_1 _17214_ (.Y(_08521_),
    .A(_01715_),
    .B(net1562));
 sg13g2_or3_1 _17215_ (.A(_01724_),
    .B(_08518_),
    .C(_08521_),
    .X(_08522_));
 sg13g2_nand2b_1 _17216_ (.Y(_08523_),
    .B(net1424),
    .A_N(net1358));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(rf_wdata_wb_18_));
 sg13g2_buf_2 fanout706 (.A(net707),
    .X(net706));
 sg13g2_a21oi_1 _17219_ (.A1(net197),
    .A2(net131),
    .Y(_08526_),
    .B1(_03067_));
 sg13g2_buf_2 fanout705 (.A(net707),
    .X(net705));
 sg13g2_buf_2 fanout704 (.A(net707),
    .X(net704));
 sg13g2_buf_2 fanout703 (.A(net707),
    .X(net703));
 sg13g2_buf_2 fanout702 (.A(rf_wdata_wb_19_),
    .X(net702));
 sg13g2_buf_2 fanout701 (.A(net702),
    .X(net701));
 sg13g2_buf_2 fanout700 (.A(net702),
    .X(net700));
 sg13g2_nand2_1 _17226_ (.Y(_08533_),
    .A(_02346_),
    .B(net1354));
 sg13g2_o21ai_1 _17227_ (.B1(_08533_),
    .Y(_08534_),
    .A1(net197),
    .A2(net1354));
 sg13g2_a21o_1 _17228_ (.A2(_01724_),
    .A1(_01715_),
    .B1(_08518_),
    .X(_08535_));
 sg13g2_buf_2 fanout699 (.A(net702),
    .X(net699));
 sg13g2_buf_2 fanout698 (.A(net699),
    .X(net698));
 sg13g2_a21o_1 _17231_ (.A2(_08534_),
    .A1(net1421),
    .B1(net1417),
    .X(_08538_));
 sg13g2_nand2_1 _17232_ (.Y(_08539_),
    .A(_04144_),
    .B(_04064_));
 sg13g2_o21ai_1 _17233_ (.B1(_08539_),
    .Y(_08540_),
    .A1(_02304_),
    .A2(_04144_));
 sg13g2_a21oi_2 _17234_ (.B1(net1680),
    .Y(_08541_),
    .A2(_08540_),
    .A1(net360));
 sg13g2_o21ai_1 _17235_ (.B1(_08541_),
    .Y(_08542_),
    .A1(_08526_),
    .A2(_08538_));
 sg13g2_a221oi_1 _17236_ (.B2(net1368),
    .C1(_08542_),
    .B1(_08513_),
    .A1(net1128),
    .Y(_08543_),
    .A2(net1319));
 sg13g2_o21ai_1 _17237_ (.B1(_08543_),
    .Y(_08544_),
    .A1(_07412_),
    .A2(_08420_));
 sg13g2_inv_1 _17238_ (.Y(_08545_),
    .A(net1419));
 sg13g2_inv_1 _17239_ (.Y(_08546_),
    .A(_08420_));
 sg13g2_nor4_2 _17240_ (.A(net1364),
    .B(_08545_),
    .C(net1315),
    .Y(_08547_),
    .D(_08546_));
 sg13g2_or2_2 _17241_ (.X(_08548_),
    .B(net1194),
    .A(net355));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(rf_wdata_wb_22_));
 sg13g2_nand4_1 _17243_ (.B(_01365_),
    .C(_01659_),
    .A(net397),
    .Y(_08550_),
    .D(_01796_));
 sg13g2_nand3_1 _17244_ (.B(_08382_),
    .C(_08550_),
    .A(_08021_),
    .Y(_08551_));
 sg13g2_inv_1 _17245_ (.Y(_08552_),
    .A(net1075));
 sg13g2_o21ai_1 _17246_ (.B1(_08552_),
    .Y(_08553_),
    .A1(csr_rdata_0_),
    .A2(net397));
 sg13g2_a21oi_2 _17247_ (.B1(_08553_),
    .Y(_08554_),
    .A2(_08548_),
    .A1(_08541_));
 sg13g2_a22oi_1 _17248_ (.Y(_08555_),
    .B1(_08544_),
    .B2(_08554_),
    .A2(_08414_),
    .A1(net1651));
 sg13g2_inv_2 _17249_ (.Y(rf_wdata_wb_0_),
    .A(_08555_));
 sg13g2_buf_1 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout695 (.A(net697),
    .X(net695));
 sg13g2_buf_2 fanout694 (.A(net697),
    .X(net694));
 sg13g2_buf_2 fanout693 (.A(net697),
    .X(net693));
 sg13g2_buf_2 fanout692 (.A(rf_wdata_wb_23_),
    .X(net692));
 sg13g2_mux2_1 _17255_ (.A0(_08479_),
    .A1(_08481_),
    .S(net1177),
    .X(_08561_));
 sg13g2_mux2_1 _17256_ (.A0(_08482_),
    .A1(_08494_),
    .S(net1180),
    .X(_08562_));
 sg13g2_nor2b_1 _17257_ (.A(net1167),
    .B_N(_08562_),
    .Y(_08563_));
 sg13g2_a21oi_1 _17258_ (.A1(net1166),
    .A2(_08561_),
    .Y(_08564_),
    .B1(_08563_));
 sg13g2_nor2_2 _17259_ (.A(_08488_),
    .B(_08505_),
    .Y(_08565_));
 sg13g2_mux2_1 _17260_ (.A0(_08492_),
    .A1(net1133),
    .S(net1180),
    .X(_08566_));
 sg13g2_nor2b_1 _17261_ (.A(net1179),
    .B_N(_08495_),
    .Y(_08567_));
 sg13g2_a21oi_1 _17262_ (.A1(net1179),
    .A2(_08486_),
    .Y(_08568_),
    .B1(_08567_));
 sg13g2_nand2_1 _17263_ (.Y(_08569_),
    .A(net1167),
    .B(_08568_));
 sg13g2_o21ai_1 _17264_ (.B1(_08569_),
    .Y(_08570_),
    .A1(net1167),
    .A2(_08566_));
 sg13g2_mux2_1 _17265_ (.A0(_08463_),
    .A1(_08467_),
    .S(net1177),
    .X(_08571_));
 sg13g2_mux2_1 _17266_ (.A0(_08468_),
    .A1(_08478_),
    .S(net1177),
    .X(_08572_));
 sg13g2_nor2b_1 _17267_ (.A(net1166),
    .B_N(_08572_),
    .Y(_08573_));
 sg13g2_a21oi_1 _17268_ (.A1(net1166),
    .A2(_08571_),
    .Y(_08574_),
    .B1(_08573_));
 sg13g2_xnor2_1 _17269_ (.Y(_08575_),
    .A(net1399),
    .B(_08474_));
 sg13g2_mux4_1 _17270_ (.S0(net41),
    .A0(_08509_),
    .A1(_08564_),
    .A2(_08570_),
    .A3(_08574_),
    .S1(net1138),
    .X(_08576_));
 sg13g2_buf_2 fanout691 (.A(net692),
    .X(net691));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_mux4_1 _17273_ (.S0(net200),
    .A0(net88),
    .A1(net1404),
    .A2(net1202),
    .A3(net1350),
    .S1(net1459),
    .X(_08579_));
 sg13g2_mux4_1 _17274_ (.S0(net200),
    .A0(net1201),
    .A1(net1408),
    .A2(net124),
    .A3(net1407),
    .S1(net1458),
    .X(_08580_));
 sg13g2_mux2_1 _17275_ (.A0(_08579_),
    .A1(_08580_),
    .S(net1175),
    .X(_08581_));
 sg13g2_mux4_1 _17276_ (.S0(net206),
    .A0(net151),
    .A1(net127),
    .A2(net194),
    .A3(net196),
    .S1(_03067_),
    .X(_08582_));
 sg13g2_mux4_1 _17277_ (.S0(net199),
    .A0(net125),
    .A1(alu_operand_a_ex_7_),
    .A2(net150),
    .A3(net1279),
    .S1(net1459),
    .X(_08583_));
 sg13g2_mux2_1 _17278_ (.A0(_08582_),
    .A1(_08583_),
    .S(net1175),
    .X(_08584_));
 sg13g2_mux2_1 _17279_ (.A0(_08581_),
    .A1(_08584_),
    .S(net1163),
    .X(_08585_));
 sg13g2_buf_2 fanout689 (.A(net691),
    .X(net689));
 sg13g2_mux4_1 _17281_ (.S0(net1459),
    .A0(net1411),
    .A1(net1409),
    .A2(net1190),
    .A3(net1199),
    .S1(net210),
    .X(_08587_));
 sg13g2_a21oi_1 _17282_ (.A1(_03067_),
    .A2(_08505_),
    .Y(_08588_),
    .B1(_08488_));
 sg13g2_mux2_1 _17283_ (.A0(_08587_),
    .A1(_08588_),
    .S(net1175),
    .X(_08589_));
 sg13g2_inv_1 _17284_ (.Y(_08590_),
    .A(_08589_));
 sg13g2_nand2_1 _17285_ (.Y(_08591_),
    .A(net1163),
    .B(_08590_));
 sg13g2_o21ai_1 _17286_ (.B1(_08591_),
    .Y(_08592_),
    .A1(net1163),
    .A2(net1133));
 sg13g2_nor2_1 _17287_ (.A(net1139),
    .B(_08592_),
    .Y(_08593_));
 sg13g2_a21oi_1 _17288_ (.A1(net1139),
    .A2(_08585_),
    .Y(_08594_),
    .B1(_08593_));
 sg13g2_nor2_2 _17289_ (.A(net41),
    .B(net1133),
    .Y(_08595_));
 sg13g2_a21oi_1 _17290_ (.A1(net43),
    .A2(_08594_),
    .Y(_08596_),
    .B1(_08595_));
 sg13g2_nand2_1 _17291_ (.Y(_08597_),
    .A(net204),
    .B(_08596_));
 sg13g2_o21ai_1 _17292_ (.B1(_08597_),
    .Y(_08598_),
    .A1(net201),
    .A2(_08576_));
 sg13g2_buf_1 fanout688 (.A(net691),
    .X(net688));
 sg13g2_nand2_1 _17294_ (.Y(_08600_),
    .A(net151),
    .B(net128));
 sg13g2_nand3_1 _17295_ (.B(_02193_),
    .C(net1356),
    .A(net151),
    .Y(_08601_));
 sg13g2_o21ai_1 _17296_ (.B1(_08601_),
    .Y(_08602_),
    .A1(net152),
    .A2(net1356));
 sg13g2_buf_2 fanout687 (.A(net691),
    .X(net687));
 sg13g2_buf_2 fanout686 (.A(rf_wdata_wb_24_),
    .X(net686));
 sg13g2_a221oi_1 _17299_ (.B2(net1422),
    .C1(net1417),
    .B1(_08602_),
    .A1(_02134_),
    .Y(_08605_),
    .A2(_08600_));
 sg13g2_a221oi_1 _17300_ (.B2(net1367),
    .C1(_08605_),
    .B1(_08598_),
    .A1(data_addr_o_10_),
    .Y(_08606_),
    .A2(net1317));
 sg13g2_buf_2 fanout685 (.A(net686),
    .X(net685));
 sg13g2_o21ai_1 _17302_ (.B1(net377),
    .Y(_08608_),
    .A1(net1197),
    .A2(_08606_));
 sg13g2_nor2_2 _17303_ (.A(_04033_),
    .B(net1538),
    .Y(_08609_));
 sg13g2_nor2_2 _17304_ (.A(net1577),
    .B(_08609_),
    .Y(_08610_));
 sg13g2_inv_2 _17305_ (.Y(_08611_),
    .A(_08610_));
 sg13g2_a22oi_1 _17306_ (.Y(_08612_),
    .B1(_08611_),
    .B2(_04918_),
    .A2(net1472),
    .A1(_05012_));
 sg13g2_and3_1 _17307_ (.X(_08613_),
    .A(net397),
    .B(_08608_),
    .C(_08612_));
 sg13g2_a21oi_2 _17308_ (.B1(_08613_),
    .Y(_08614_),
    .A2(net1677),
    .A1(csr_rdata_10_));
 sg13g2_a22oi_1 _17309_ (.Y(_08615_),
    .B1(net1951),
    .B2(data_rdata_i_15_),
    .A2(net1935),
    .A1(data_rdata_i_23_));
 sg13g2_nand2_1 _17310_ (.Y(_08616_),
    .A(data_rdata_i_31_),
    .B(net1944));
 sg13g2_nand2_1 _17311_ (.Y(_08617_),
    .A(_08615_),
    .B(_08616_));
 sg13g2_a21o_1 _17312_ (.A2(net417),
    .A1(data_rdata_i_7_),
    .B1(_08617_),
    .X(_08618_));
 sg13g2_nand2_1 _17313_ (.Y(_08619_),
    .A(\load_store_unit_i.data_sign_ext_q ),
    .B(_08618_));
 sg13g2_nand2_1 _17314_ (.Y(_08620_),
    .A(net1960),
    .B(_08619_));
 sg13g2_buf_2 fanout684 (.A(rf_wdata_wb_24_),
    .X(net684));
 sg13g2_a22oi_1 _17316_ (.Y(_08622_),
    .B1(net414),
    .B2(data_rdata_i_10_),
    .A2(net1947),
    .A1(data_rdata_i_2_));
 sg13g2_buf_2 fanout683 (.A(rf_wdata_wb_24_),
    .X(net683));
 sg13g2_buf_8 fanout682 (.A(\cs_registers_i/_1763_ ),
    .X(net682));
 sg13g2_a22oi_1 _17319_ (.Y(_08625_),
    .B1(net1951),
    .B2(data_rdata_i_18_),
    .A2(net1935),
    .A1(data_rdata_i_26_));
 sg13g2_a21oi_1 _17320_ (.A1(_08622_),
    .A2(_08625_),
    .Y(_08626_),
    .B1(net1959));
 sg13g2_buf_16 fanout681 (.X(net681),
    .A(net682));
 sg13g2_buf_8 fanout680 (.A(\cs_registers_i/_1763_ ),
    .X(net680));
 sg13g2_buf_16 fanout679 (.X(net679),
    .A(net680));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(\cs_registers_i/_2110_ ));
 sg13g2_a221oi_1 _17325_ (.B2(\load_store_unit_i.rdata_q_10_ ),
    .C1(net1931),
    .B1(net1951),
    .A1(\load_store_unit_i.rdata_q_18_ ),
    .Y(_08631_),
    .A2(net1935));
 sg13g2_a21oi_1 _17326_ (.A1(net1931),
    .A2(_08625_),
    .Y(_08632_),
    .B1(_08631_));
 sg13g2_nor2_1 _17327_ (.A(net1960),
    .B(_08632_),
    .Y(_08633_));
 sg13g2_nand4_1 _17328_ (.B(\load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ),
    .C(_01495_),
    .A(net2466),
    .Y(_08634_),
    .D(_01596_));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(net678));
 sg13g2_a21oi_1 _17330_ (.A1(_08622_),
    .A2(_08633_),
    .Y(_08636_),
    .B1(net1646));
 sg13g2_o21ai_1 _17331_ (.B1(_08636_),
    .Y(_08637_),
    .A1(net1602),
    .A2(_08626_));
 sg13g2_o21ai_1 _17332_ (.B1(_08637_),
    .Y(rf_wdata_wb_10_),
    .A1(net1073),
    .A2(_08614_));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net677));
 sg13g2_nand2_2 _17334_ (.Y(_08639_),
    .A(net1538),
    .B(_06016_));
 sg13g2_nor2_1 _17335_ (.A(_05128_),
    .B(_08639_),
    .Y(_08640_));
 sg13g2_buf_1 fanout675 (.A(rf_wdata_wb_21_),
    .X(net675));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674));
 sg13g2_mux2_1 _17338_ (.A0(_08580_),
    .A1(_08587_),
    .S(net1175),
    .X(_08643_));
 sg13g2_a22oi_1 _17339_ (.Y(_08644_),
    .B1(_08423_),
    .B2(_08438_),
    .A2(net1458),
    .A1(net1247));
 sg13g2_nor3_1 _17340_ (.A(net1163),
    .B(_08488_),
    .C(_08644_),
    .Y(_08645_));
 sg13g2_a21oi_2 _17341_ (.B1(_08645_),
    .Y(_08646_),
    .A2(_08643_),
    .A1(net1163));
 sg13g2_nor2_1 _17342_ (.A(net1136),
    .B(_08565_),
    .Y(_08647_));
 sg13g2_a21oi_1 _17343_ (.A1(net1136),
    .A2(_08646_),
    .Y(_08648_),
    .B1(_08647_));
 sg13g2_mux2_1 _17344_ (.A0(_08583_),
    .A1(_08579_),
    .S(net1175),
    .X(_08649_));
 sg13g2_mux4_1 _17345_ (.S0(net1459),
    .A0(net1415),
    .A1(net1413),
    .A2(net1281),
    .A3(net1249),
    .S1(net210),
    .X(_08650_));
 sg13g2_mux2_1 _17346_ (.A0(_08650_),
    .A1(_08582_),
    .S(net1175),
    .X(_08651_));
 sg13g2_mux2_1 _17347_ (.A0(_08649_),
    .A1(_08651_),
    .S(net1162),
    .X(_08652_));
 sg13g2_nor2_1 _17348_ (.A(net1136),
    .B(_08652_),
    .Y(_08653_));
 sg13g2_xnor2_1 _17349_ (.Y(_08654_),
    .A(net1457),
    .B(net203));
 sg13g2_nand2_1 _17350_ (.Y(_08655_),
    .A(_01234_),
    .B(_08654_));
 sg13g2_o21ai_1 _17351_ (.B1(_08655_),
    .Y(_08656_),
    .A1(net1351),
    .A2(_08654_));
 sg13g2_mux4_1 _17352_ (.S0(net1459),
    .A0(net1352),
    .A1(net1283),
    .A2(net1203),
    .A3(net1250),
    .S1(net210),
    .X(_08657_));
 sg13g2_nand2_1 _17353_ (.Y(_08658_),
    .A(net1176),
    .B(_08657_));
 sg13g2_o21ai_1 _17354_ (.B1(_08658_),
    .Y(_08659_),
    .A1(net1176),
    .A2(_08656_));
 sg13g2_mux4_1 _17355_ (.S0(net200),
    .A0(net1413),
    .A1(net1249),
    .A2(net1415),
    .A3(net1282),
    .S1(net1459),
    .X(_08660_));
 sg13g2_mux4_1 _17356_ (.S0(_03067_),
    .A0(net1352),
    .A1(net1283),
    .A2(net1203),
    .A3(net1250),
    .S1(net205),
    .X(_08661_));
 sg13g2_mux2_1 _17357_ (.A0(_08660_),
    .A1(_08661_),
    .S(net1176),
    .X(_08662_));
 sg13g2_mux2_1 _17358_ (.A0(_08659_),
    .A1(_08662_),
    .S(net1162),
    .X(_08663_));
 sg13g2_nor2_1 _17359_ (.A(net1134),
    .B(_08663_),
    .Y(_08664_));
 sg13g2_a22oi_1 _17360_ (.Y(_08665_),
    .B1(_08664_),
    .B2(net1136),
    .A2(_08653_),
    .A1(net41));
 sg13g2_o21ai_1 _17361_ (.B1(_08665_),
    .Y(_08666_),
    .A1(net42),
    .A2(_08648_));
 sg13g2_mux4_1 _17362_ (.S0(net1165),
    .A0(_08496_),
    .A1(_08483_),
    .A2(_08565_),
    .A3(_08493_),
    .S1(net47),
    .X(_08667_));
 sg13g2_nor2_1 _17363_ (.A(net41),
    .B(_08509_),
    .Y(_08668_));
 sg13g2_a21o_1 _17364_ (.A2(_08667_),
    .A1(net44),
    .B1(_08668_),
    .X(_08669_));
 sg13g2_nor2_1 _17365_ (.A(net207),
    .B(_08669_),
    .Y(_08670_));
 sg13g2_a21oi_1 _17366_ (.A1(net209),
    .A2(_08666_),
    .Y(_08671_),
    .B1(_08670_));
 sg13g2_a21oi_1 _17367_ (.A1(_02483_),
    .A2(net130),
    .Y(_08672_),
    .B1(net1414));
 sg13g2_nand3_1 _17368_ (.B(_02483_),
    .C(net1354),
    .A(net1414),
    .Y(_08673_));
 sg13g2_o21ai_1 _17369_ (.B1(_08673_),
    .Y(_08674_),
    .A1(_02483_),
    .A2(net1357));
 sg13g2_a21oi_1 _17370_ (.A1(net1421),
    .A2(_08674_),
    .Y(_08675_),
    .B1(net1416));
 sg13g2_nor2b_1 _17371_ (.A(_08672_),
    .B_N(_08675_),
    .Y(_08676_));
 sg13g2_a221oi_1 _17372_ (.B2(net1366),
    .C1(_08676_),
    .B1(_08671_),
    .A1(data_addr_o_11_),
    .Y(_08677_),
    .A2(net1318));
 sg13g2_o21ai_1 _17373_ (.B1(net375),
    .Y(_08678_),
    .A1(net1196),
    .A2(_08677_));
 sg13g2_o21ai_1 _17374_ (.B1(_08678_),
    .Y(_08679_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .A2(_08610_));
 sg13g2_nor3_2 _17375_ (.A(net1679),
    .B(_08640_),
    .C(_08679_),
    .Y(_08680_));
 sg13g2_a21oi_2 _17376_ (.B1(_08680_),
    .Y(_08681_),
    .A2(net1677),
    .A1(csr_rdata_11_));
 sg13g2_buf_2 fanout673 (.A(net675),
    .X(net673));
 sg13g2_a22oi_1 _17378_ (.Y(_08683_),
    .B1(net414),
    .B2(data_rdata_i_11_),
    .A2(net1950),
    .A1(data_rdata_i_3_));
 sg13g2_a22oi_1 _17379_ (.Y(_08684_),
    .B1(net1955),
    .B2(data_rdata_i_19_),
    .A2(net1939),
    .A1(data_rdata_i_27_));
 sg13g2_a21oi_1 _17380_ (.A1(_08683_),
    .A2(_08684_),
    .Y(_08685_),
    .B1(net1959));
 sg13g2_buf_2 fanout672 (.A(rf_wdata_wb_21_),
    .X(net672));
 sg13g2_a221oi_1 _17382_ (.B2(\load_store_unit_i.rdata_q_11_ ),
    .C1(net1932),
    .B1(net1957),
    .A1(\load_store_unit_i.rdata_q_19_ ),
    .Y(_08687_),
    .A2(net1939));
 sg13g2_a21oi_1 _17383_ (.A1(net1932),
    .A2(_08684_),
    .Y(_08688_),
    .B1(_08687_));
 sg13g2_nor2_1 _17384_ (.A(net1961),
    .B(_08688_),
    .Y(_08689_));
 sg13g2_a21oi_1 _17385_ (.A1(_08683_),
    .A2(_08689_),
    .Y(_08690_),
    .B1(net1646));
 sg13g2_o21ai_1 _17386_ (.B1(_08690_),
    .Y(_08691_),
    .A1(net1602),
    .A2(_08685_));
 sg13g2_o21ai_1 _17387_ (.B1(_08691_),
    .Y(rf_wdata_wb_11_),
    .A1(net1072),
    .A2(_08681_));
 sg13g2_buf_1 fanout671 (.A(net672),
    .X(net671));
 sg13g2_nor2_1 _17389_ (.A(net45),
    .B(_08652_),
    .Y(_08693_));
 sg13g2_a21oi_1 _17390_ (.A1(net46),
    .A2(_08646_),
    .Y(_08694_),
    .B1(_08693_));
 sg13g2_inv_1 _17391_ (.Y(_08695_),
    .A(_08694_));
 sg13g2_a21oi_1 _17392_ (.A1(net44),
    .A2(_08695_),
    .Y(_08696_),
    .B1(_08595_));
 sg13g2_nand2_1 _17393_ (.Y(_08697_),
    .A(net1166),
    .B(net1136));
 sg13g2_mux2_1 _17394_ (.A0(_08493_),
    .A1(_08565_),
    .S(_08697_),
    .X(_08698_));
 sg13g2_mux4_1 _17395_ (.S0(net1164),
    .A0(_08496_),
    .A1(_08483_),
    .A2(_08480_),
    .A3(_08469_),
    .S1(net1137),
    .X(_08699_));
 sg13g2_mux2_1 _17396_ (.A0(_08698_),
    .A1(_08699_),
    .S(net42),
    .X(_08700_));
 sg13g2_mux2_1 _17397_ (.A0(_08696_),
    .A1(_08700_),
    .S(net206),
    .X(_08701_));
 sg13g2_buf_2 fanout670 (.A(net672),
    .X(net670));
 sg13g2_nand2_1 _17399_ (.Y(_08703_),
    .A(net1412),
    .B(net129));
 sg13g2_buf_1 fanout669 (.A(rf_wdata_wb_26_),
    .X(net669));
 sg13g2_nand2_1 _17401_ (.Y(_08705_),
    .A(_02470_),
    .B(net1353));
 sg13g2_o21ai_1 _17402_ (.B1(_08705_),
    .Y(_08706_),
    .A1(net1412),
    .A2(net1353));
 sg13g2_a221oi_1 _17403_ (.B2(net1421),
    .C1(net1416),
    .B1(_08706_),
    .A1(_02469_),
    .Y(_08707_),
    .A2(_08703_));
 sg13g2_a221oi_1 _17404_ (.B2(net1366),
    .C1(_08707_),
    .B1(_08701_),
    .A1(data_addr_o_12_),
    .Y(_08708_),
    .A2(net1317));
 sg13g2_o21ai_1 _17405_ (.B1(net375),
    .Y(_08709_),
    .A1(net1196),
    .A2(_08708_));
 sg13g2_o21ai_1 _17406_ (.B1(_08709_),
    .Y(_08710_),
    .A1(net2114),
    .A2(_08610_));
 sg13g2_a221oi_1 _17407_ (.B2(net1472),
    .C1(_08710_),
    .B1(_05262_),
    .A1(net412),
    .Y(_08711_),
    .A2(net1716));
 sg13g2_a21oi_2 _17408_ (.B1(_08711_),
    .Y(_08712_),
    .A2(net1677),
    .A1(csr_rdata_12_));
 sg13g2_a22oi_1 _17409_ (.Y(_08713_),
    .B1(net414),
    .B2(data_rdata_i_12_),
    .A2(net1948),
    .A1(data_rdata_i_4_));
 sg13g2_a22oi_1 _17410_ (.Y(_08714_),
    .B1(net1957),
    .B2(data_rdata_i_20_),
    .A2(net1939),
    .A1(data_rdata_i_28_));
 sg13g2_a21oi_1 _17411_ (.A1(_08713_),
    .A2(_08714_),
    .Y(_08715_),
    .B1(net1959));
 sg13g2_a221oi_1 _17412_ (.B2(\load_store_unit_i.rdata_q_12_ ),
    .C1(net1934),
    .B1(net1957),
    .A1(\load_store_unit_i.rdata_q_20_ ),
    .Y(_08716_),
    .A2(net1941));
 sg13g2_a21oi_1 _17413_ (.A1(net1932),
    .A2(_08714_),
    .Y(_08717_),
    .B1(_08716_));
 sg13g2_nor2_1 _17414_ (.A(net1961),
    .B(_08717_),
    .Y(_08718_));
 sg13g2_a21oi_1 _17415_ (.A1(_08713_),
    .A2(_08718_),
    .Y(_08719_),
    .B1(net1647));
 sg13g2_o21ai_1 _17416_ (.B1(_08719_),
    .Y(_00490_),
    .A1(net1602),
    .A2(_08715_));
 sg13g2_o21ai_1 _17417_ (.B1(_00490_),
    .Y(rf_wdata_wb_12_),
    .A1(net1073),
    .A2(_08712_));
 sg13g2_mux2_1 _17418_ (.A0(_08657_),
    .A1(_08650_),
    .S(net1176),
    .X(_00491_));
 sg13g2_nor2_1 _17419_ (.A(net1176),
    .B(_08661_),
    .Y(_00492_));
 sg13g2_a21oi_1 _17420_ (.A1(net1176),
    .A2(_08656_),
    .Y(_00493_),
    .B1(_00492_));
 sg13g2_mux2_1 _17421_ (.A0(_00491_),
    .A1(_00493_),
    .S(net1162),
    .X(_00494_));
 sg13g2_nand2_1 _17422_ (.Y(_00495_),
    .A(net1135),
    .B(_08592_));
 sg13g2_o21ai_1 _17423_ (.B1(_00495_),
    .Y(_00496_),
    .A1(net1134),
    .A2(_00494_));
 sg13g2_a21oi_1 _17424_ (.A1(net43),
    .A2(_08585_),
    .Y(_00497_),
    .B1(_08668_));
 sg13g2_mux2_1 _17425_ (.A0(_00496_),
    .A1(_00497_),
    .S(net45),
    .X(_00498_));
 sg13g2_inv_1 _17426_ (.Y(_00499_),
    .A(_08570_));
 sg13g2_nand2_1 _17427_ (.Y(_00500_),
    .A(net46),
    .B(_00499_));
 sg13g2_o21ai_1 _17428_ (.B1(_00500_),
    .Y(_00501_),
    .A1(net45),
    .A2(_08564_));
 sg13g2_nor2_1 _17429_ (.A(net1134),
    .B(_00501_),
    .Y(_00502_));
 sg13g2_nor2_1 _17430_ (.A(_08595_),
    .B(_00502_),
    .Y(_00503_));
 sg13g2_nand2_1 _17431_ (.Y(_00504_),
    .A(net204),
    .B(_00503_));
 sg13g2_o21ai_1 _17432_ (.B1(_00504_),
    .Y(_00505_),
    .A1(net202),
    .A2(_00498_));
 sg13g2_a21oi_1 _17433_ (.A1(_02104_),
    .A2(net130),
    .Y(_00506_),
    .B1(net1352));
 sg13g2_nand3_1 _17434_ (.B(_02104_),
    .C(net1354),
    .A(net1352),
    .Y(_00507_));
 sg13g2_o21ai_1 _17435_ (.B1(_00507_),
    .Y(_00508_),
    .A1(_02104_),
    .A2(net1357));
 sg13g2_a21oi_1 _17436_ (.A1(net1421),
    .A2(_00508_),
    .Y(_00509_),
    .B1(net1416));
 sg13g2_nor2b_1 _17437_ (.A(_00506_),
    .B_N(_00509_),
    .Y(_00510_));
 sg13g2_a221oi_1 _17438_ (.B2(net1367),
    .C1(_00510_),
    .B1(_00505_),
    .A1(data_addr_o_13_),
    .Y(_00511_),
    .A2(net1318));
 sg13g2_o21ai_1 _17439_ (.B1(net375),
    .Y(_00512_),
    .A1(net1196),
    .A2(_00511_));
 sg13g2_o21ai_1 _17440_ (.B1(_00512_),
    .Y(_00513_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .A2(_08610_));
 sg13g2_a221oi_1 _17441_ (.B2(net1472),
    .C1(_00513_),
    .B1(_05356_),
    .A1(net412),
    .Y(_00514_),
    .A2(_01198_));
 sg13g2_a21oi_2 _17442_ (.B1(_00514_),
    .Y(_00515_),
    .A2(net1677),
    .A1(csr_rdata_13_));
 sg13g2_a22oi_1 _17443_ (.Y(_00516_),
    .B1(net414),
    .B2(data_rdata_i_13_),
    .A2(net1949),
    .A1(data_rdata_i_5_));
 sg13g2_a22oi_1 _17444_ (.Y(_00517_),
    .B1(net1956),
    .B2(data_rdata_i_21_),
    .A2(net1940),
    .A1(data_rdata_i_29_));
 sg13g2_a21oi_1 _17445_ (.A1(_00516_),
    .A2(_00517_),
    .Y(_00518_),
    .B1(_08388_));
 sg13g2_a221oi_1 _17446_ (.B2(\load_store_unit_i.rdata_q_13_ ),
    .C1(net1934),
    .B1(net1956),
    .A1(\load_store_unit_i.rdata_q_21_ ),
    .Y(_00519_),
    .A2(net1940));
 sg13g2_a21oi_1 _17447_ (.A1(net1933),
    .A2(_00517_),
    .Y(_00520_),
    .B1(_00519_));
 sg13g2_nor2_1 _17448_ (.A(net1963),
    .B(_00520_),
    .Y(_00521_));
 sg13g2_a21oi_1 _17449_ (.A1(_00516_),
    .A2(_00521_),
    .Y(_00522_),
    .B1(net1647));
 sg13g2_o21ai_1 _17450_ (.B1(_00522_),
    .Y(_00523_),
    .A1(net1602),
    .A2(_00518_));
 sg13g2_o21ai_1 _17451_ (.B1(_00523_),
    .Y(rf_wdata_wb_13_),
    .A1(net1072),
    .A2(_00515_));
 sg13g2_nor2_1 _17452_ (.A(_05470_),
    .B(_08639_),
    .Y(_00524_));
 sg13g2_inv_1 _17453_ (.Y(_00525_),
    .A(_08568_));
 sg13g2_mux2_1 _17454_ (.A0(_00525_),
    .A1(_08562_),
    .S(net1167),
    .X(_00526_));
 sg13g2_nand2_1 _17455_ (.Y(_00527_),
    .A(_08492_),
    .B(_08506_));
 sg13g2_o21ai_1 _17456_ (.B1(_00527_),
    .Y(_00528_),
    .A1(_08509_),
    .A2(_08506_));
 sg13g2_mux2_1 _17457_ (.A0(_08561_),
    .A1(_08572_),
    .S(net1166),
    .X(_00529_));
 sg13g2_mux4_1 _17458_ (.S0(net41),
    .A0(net1133),
    .A1(_00526_),
    .A2(_00528_),
    .A3(_00529_),
    .S1(net1136),
    .X(_00530_));
 sg13g2_mux2_1 _17459_ (.A0(_08584_),
    .A1(_00491_),
    .S(net1162),
    .X(_00531_));
 sg13g2_mux2_1 _17460_ (.A0(_08589_),
    .A1(_08581_),
    .S(net1163),
    .X(_00532_));
 sg13g2_and2_1 _17461_ (.A(net45),
    .B(_00532_),
    .X(_00533_));
 sg13g2_a21oi_1 _17462_ (.A1(net1139),
    .A2(_00531_),
    .Y(_00534_),
    .B1(_00533_));
 sg13g2_a21oi_1 _17463_ (.A1(net43),
    .A2(_00534_),
    .Y(_00535_),
    .B1(_08595_));
 sg13g2_mux2_1 _17464_ (.A0(_00530_),
    .A1(_00535_),
    .S(net202),
    .X(_00536_));
 sg13g2_nand2b_1 _17465_ (.Y(_00537_),
    .B(net129),
    .A_N(net241));
 sg13g2_mux2_1 _17466_ (.A0(net241),
    .A1(_02112_),
    .S(net1353),
    .X(_00538_));
 sg13g2_a221oi_1 _17467_ (.B2(net1421),
    .C1(net1416),
    .B1(_00538_),
    .A1(_01224_),
    .Y(_00539_),
    .A2(_00537_));
 sg13g2_a221oi_1 _17468_ (.B2(net1366),
    .C1(_00539_),
    .B1(_00536_),
    .A1(data_addr_o_14_),
    .Y(_00540_),
    .A2(net1317));
 sg13g2_o21ai_1 _17469_ (.B1(net374),
    .Y(_00541_),
    .A1(net1196),
    .A2(_00540_));
 sg13g2_o21ai_1 _17470_ (.B1(_00541_),
    .Y(_00542_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .A2(_08610_));
 sg13g2_nor3_2 _17471_ (.A(net1679),
    .B(_00524_),
    .C(_00542_),
    .Y(_00543_));
 sg13g2_a21oi_2 _17472_ (.B1(_00543_),
    .Y(_00544_),
    .A2(net1676),
    .A1(csr_rdata_14_));
 sg13g2_o21ai_1 _17473_ (.B1(net1602),
    .Y(_00545_),
    .A1(net1962),
    .A2(_08388_));
 sg13g2_a22oi_1 _17474_ (.Y(_00546_),
    .B1(net1953),
    .B2(data_rdata_i_22_),
    .A2(net1937),
    .A1(data_rdata_i_30_));
 sg13g2_buf_1 fanout668 (.A(net669),
    .X(net668));
 sg13g2_a22oi_1 _17476_ (.Y(_00548_),
    .B1(net1953),
    .B2(\load_store_unit_i.rdata_q_14_ ),
    .A2(net1937),
    .A1(\load_store_unit_i.rdata_q_22_ ));
 sg13g2_a22oi_1 _17477_ (.Y(_00549_),
    .B1(_00548_),
    .B2(net1704),
    .A2(_00546_),
    .A1(_00545_));
 sg13g2_a221oi_1 _17478_ (.B2(data_rdata_i_14_),
    .C1(_00549_),
    .B1(net415),
    .A1(data_rdata_i_6_),
    .Y(_00550_),
    .A2(net1945));
 sg13g2_o21ai_1 _17479_ (.B1(net1648),
    .Y(_00551_),
    .A1(net1931),
    .A2(net1602));
 sg13g2_or2_1 _17480_ (.X(_00552_),
    .B(_00551_),
    .A(_00550_));
 sg13g2_o21ai_1 _17481_ (.B1(_00552_),
    .Y(rf_wdata_wb_14_),
    .A1(net1072),
    .A2(_00544_));
 sg13g2_mux2_1 _17482_ (.A0(_08643_),
    .A1(_08649_),
    .S(net1163),
    .X(_00553_));
 sg13g2_mux2_1 _17483_ (.A0(_08651_),
    .A1(_08659_),
    .S(net1162),
    .X(_00554_));
 sg13g2_mux4_1 _17484_ (.S0(net1139),
    .A0(net1133),
    .A1(_08508_),
    .A2(_00553_),
    .A3(_00554_),
    .S1(_08575_),
    .X(_00555_));
 sg13g2_a21o_1 _17485_ (.A2(net44),
    .A1(_08499_),
    .B1(_08668_),
    .X(_00556_));
 sg13g2_mux2_1 _17486_ (.A0(_00555_),
    .A1(_00556_),
    .S(net200),
    .X(_00557_));
 sg13g2_nand2_1 _17487_ (.Y(_00558_),
    .A(_02526_),
    .B(net129));
 sg13g2_nand3_1 _17488_ (.B(_02526_),
    .C(net1355),
    .A(net1351),
    .Y(_00559_));
 sg13g2_o21ai_1 _17489_ (.B1(_00559_),
    .Y(_00560_),
    .A1(net1343),
    .A2(net1355));
 sg13g2_a221oi_1 _17490_ (.B2(net1422),
    .C1(net1418),
    .B1(_00560_),
    .A1(_01228_),
    .Y(_00561_),
    .A2(_00558_));
 sg13g2_a221oi_1 _17491_ (.B2(net1367),
    .C1(_00561_),
    .B1(_00557_),
    .A1(data_addr_o_15_),
    .Y(_00562_),
    .A2(net1318));
 sg13g2_o21ai_1 _17492_ (.B1(net374),
    .Y(_00563_),
    .A1(net1197),
    .A2(_00562_));
 sg13g2_o21ai_1 _17493_ (.B1(_00563_),
    .Y(_00564_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .A2(_08610_));
 sg13g2_a221oi_1 _17494_ (.B2(net1472),
    .C1(_00564_),
    .B1(_05616_),
    .A1(_01153_),
    .Y(_00565_),
    .A2(_01198_));
 sg13g2_a21oi_2 _17495_ (.B1(_00565_),
    .Y(_00566_),
    .A2(net1677),
    .A1(csr_rdata_15_));
 sg13g2_a22oi_1 _17496_ (.Y(_00567_),
    .B1(net413),
    .B2(data_rdata_i_15_),
    .A2(net1944),
    .A1(data_rdata_i_7_));
 sg13g2_a22oi_1 _17497_ (.Y(_00568_),
    .B1(net1951),
    .B2(data_rdata_i_23_),
    .A2(net1935),
    .A1(data_rdata_i_31_));
 sg13g2_a21oi_1 _17498_ (.A1(_00567_),
    .A2(_00568_),
    .Y(_00569_),
    .B1(net1959));
 sg13g2_a221oi_1 _17499_ (.B2(\load_store_unit_i.rdata_q_15_ ),
    .C1(net1932),
    .B1(net1952),
    .A1(\load_store_unit_i.rdata_q_23_ ),
    .Y(_00570_),
    .A2(net1936));
 sg13g2_a21oi_1 _17500_ (.A1(net1931),
    .A2(_00568_),
    .Y(_00571_),
    .B1(_00570_));
 sg13g2_nor2_1 _17501_ (.A(net1960),
    .B(_00571_),
    .Y(_00572_));
 sg13g2_a21oi_1 _17502_ (.A1(_00567_),
    .A2(_00572_),
    .Y(_00573_),
    .B1(net1646));
 sg13g2_o21ai_1 _17503_ (.B1(_00573_),
    .Y(_00574_),
    .A1(net1602),
    .A2(_00569_));
 sg13g2_o21ai_1 _17504_ (.B1(_00574_),
    .Y(rf_wdata_wb_15_),
    .A1(net1072),
    .A2(_00566_));
 sg13g2_buf_2 fanout667 (.A(net669),
    .X(net667));
 sg13g2_buf_2 fanout666 (.A(rf_wdata_wb_26_),
    .X(net666));
 sg13g2_buf_2 fanout665 (.A(rf_wdata_wb_26_),
    .X(net665));
 sg13g2_buf_8 fanout664 (.A(\cs_registers_i/_0584_ ),
    .X(net664));
 sg13g2_a22oi_1 _17509_ (.Y(_00579_),
    .B1(net1945),
    .B2(data_rdata_i_8_),
    .A2(net1954),
    .A1(\load_store_unit_i.rdata_q_16_ ));
 sg13g2_inv_1 _17510_ (.Y(_00580_),
    .A(_00579_));
 sg13g2_a221oi_1 _17511_ (.B2(data_rdata_i_16_),
    .C1(_00580_),
    .B1(net417),
    .A1(data_rdata_i_0_),
    .Y(_00581_),
    .A2(net1938));
 sg13g2_a21oi_1 _17512_ (.A1(net1960),
    .A2(_08618_),
    .Y(_00582_),
    .B1(_00569_));
 sg13g2_nand2b_1 _17513_ (.Y(_00583_),
    .B(\load_store_unit_i.data_sign_ext_q ),
    .A_N(_00582_));
 sg13g2_buf_16 fanout663 (.X(net663),
    .A(net664));
 sg13g2_o21ai_1 _17515_ (.B1(net1601),
    .Y(_00585_),
    .A1(net1707),
    .A2(_00581_));
 sg13g2_nor2_1 _17516_ (.A(csr_rdata_16_),
    .B(_01199_),
    .Y(_00586_));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662));
 sg13g2_nor3_1 _17518_ (.A(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .B(net1679),
    .C(net341),
    .Y(_00588_));
 sg13g2_mux2_1 _17519_ (.A0(_00555_),
    .A1(_00556_),
    .S(net207),
    .X(_00589_));
 sg13g2_nand2_1 _17520_ (.Y(_00590_),
    .A(_02551_),
    .B(net128));
 sg13g2_buf_1 fanout661 (.A(net663),
    .X(net661));
 sg13g2_nand3_1 _17522_ (.B(_02551_),
    .C(net1356),
    .A(alu_operand_a_ex_16_),
    .Y(_00592_));
 sg13g2_o21ai_1 _17523_ (.B1(_00592_),
    .Y(_00593_),
    .A1(_02551_),
    .A2(net1357));
 sg13g2_a221oi_1 _17524_ (.B2(net1422),
    .C1(net1418),
    .B1(_00593_),
    .A1(_01234_),
    .Y(_00594_),
    .A2(_00590_));
 sg13g2_a221oi_1 _17525_ (.B2(net1367),
    .C1(_00594_),
    .B1(_00589_),
    .A1(data_addr_o_16_),
    .Y(_00595_),
    .A2(net1318));
 sg13g2_nor3_1 _17526_ (.A(_07002_),
    .B(net1196),
    .C(_00595_),
    .Y(_00596_));
 sg13g2_nor3_1 _17527_ (.A(_04033_),
    .B(net299),
    .C(_05748_),
    .Y(_00597_));
 sg13g2_nand2_1 _17528_ (.Y(_00598_),
    .A(_04064_),
    .B(_08609_));
 sg13g2_nor2_1 _17529_ (.A(net1679),
    .B(net1577),
    .Y(_00599_));
 sg13g2_nand2_1 _17530_ (.Y(_00600_),
    .A(_00598_),
    .B(_00599_));
 sg13g2_nor3_1 _17531_ (.A(_00596_),
    .B(_00597_),
    .C(_00600_),
    .Y(_00601_));
 sg13g2_nor4_2 _17532_ (.A(_08551_),
    .B(_00586_),
    .C(_00588_),
    .Y(_00602_),
    .D(_00601_));
 sg13g2_a21o_2 _17533_ (.A2(_00585_),
    .A1(net1648),
    .B1(_00602_),
    .X(rf_wdata_wb_16_));
 sg13g2_nand3b_1 _17534_ (.B(net343),
    .C(_07002_),
    .Y(_00603_),
    .A_N(_05889_));
 sg13g2_o21ai_1 _17535_ (.B1(_00603_),
    .Y(_00604_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .A2(net340));
 sg13g2_nand2_1 _17536_ (.Y(_00605_),
    .A(data_addr_o_17_),
    .B(net1315));
 sg13g2_a21o_1 _17537_ (.A2(net132),
    .A1(_02592_),
    .B1(net1250),
    .X(_00606_));
 sg13g2_nand3_1 _17538_ (.B(_02592_),
    .C(net1361),
    .A(net1250),
    .Y(_00607_));
 sg13g2_o21ai_1 _17539_ (.B1(_00607_),
    .Y(_00608_),
    .A1(_02592_),
    .A2(net1361));
 sg13g2_a21oi_1 _17540_ (.A1(net1425),
    .A2(_00608_),
    .Y(_00609_),
    .B1(net1419));
 sg13g2_buf_16 fanout660 (.X(net660),
    .A(net663));
 sg13g2_mux2_1 _17542_ (.A0(_00530_),
    .A1(_00535_),
    .S(net208),
    .X(_00611_));
 sg13g2_a22oi_1 _17543_ (.Y(_00612_),
    .B1(_00611_),
    .B2(net1364),
    .A2(_00609_),
    .A1(_00606_));
 sg13g2_buf_4 fanout659 (.X(net659),
    .A(net664));
 sg13g2_a21oi_1 _17545_ (.A1(_00605_),
    .A2(_00612_),
    .Y(_00614_),
    .B1(net1194));
 sg13g2_nor2_1 _17546_ (.A(net1680),
    .B(net1075),
    .Y(_00615_));
 sg13g2_o21ai_1 _17547_ (.B1(net1061),
    .Y(_00616_),
    .A1(net355),
    .A2(_00614_));
 sg13g2_a22oi_1 _17548_ (.Y(_00617_),
    .B1(net1956),
    .B2(\load_store_unit_i.rdata_q_17_ ),
    .A2(net1941),
    .A1(data_rdata_i_1_));
 sg13g2_inv_1 _17549_ (.Y(_00618_),
    .A(_00617_));
 sg13g2_a221oi_1 _17550_ (.B2(data_rdata_i_17_),
    .C1(_00618_),
    .B1(net415),
    .A1(data_rdata_i_9_),
    .Y(_00619_),
    .A2(net1950));
 sg13g2_o21ai_1 _17551_ (.B1(net1601),
    .Y(_00620_),
    .A1(net1705),
    .A2(_00619_));
 sg13g2_nor2_2 _17552_ (.A(net396),
    .B(net1075),
    .Y(_00621_));
 sg13g2_a22oi_1 _17553_ (.Y(_00622_),
    .B1(net1060),
    .B2(csr_rdata_17_),
    .A2(_00620_),
    .A1(net1649));
 sg13g2_o21ai_1 _17554_ (.B1(_00622_),
    .Y(rf_wdata_wb_17_),
    .A1(_00604_),
    .A2(_00616_));
 sg13g2_or3_1 _17555_ (.A(net1576),
    .B(_04033_),
    .C(_06000_),
    .X(_00623_));
 sg13g2_o21ai_1 _17556_ (.B1(_00623_),
    .Y(_00624_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_50_ ),
    .A2(net340));
 sg13g2_nand2_1 _17557_ (.Y(_00625_),
    .A(data_addr_o_18_),
    .B(net1315));
 sg13g2_a21o_1 _17558_ (.A2(net132),
    .A1(_02564_),
    .B1(net1203),
    .X(_00626_));
 sg13g2_nand3_1 _17559_ (.B(_02564_),
    .C(net1359),
    .A(net1203),
    .Y(_00627_));
 sg13g2_o21ai_1 _17560_ (.B1(_00627_),
    .Y(_00628_),
    .A1(_02564_),
    .A2(net1359));
 sg13g2_a21oi_1 _17561_ (.A1(net1424),
    .A2(_00628_),
    .Y(_00629_),
    .B1(net1418));
 sg13g2_nand2_1 _17562_ (.Y(_00630_),
    .A(net212),
    .B(_00503_));
 sg13g2_o21ai_1 _17563_ (.B1(_00630_),
    .Y(_00631_),
    .A1(net208),
    .A2(_00498_));
 sg13g2_a22oi_1 _17564_ (.Y(_00632_),
    .B1(_00631_),
    .B2(net1365),
    .A2(_00629_),
    .A1(_00626_));
 sg13g2_a21oi_1 _17565_ (.A1(_00625_),
    .A2(_00632_),
    .Y(_00633_),
    .B1(net1194));
 sg13g2_o21ai_1 _17566_ (.B1(net1061),
    .Y(_00634_),
    .A1(net355),
    .A2(_00633_));
 sg13g2_a22oi_1 _17567_ (.Y(_00635_),
    .B1(net1951),
    .B2(\load_store_unit_i.rdata_q_18_ ),
    .A2(net1935),
    .A1(data_rdata_i_2_));
 sg13g2_inv_1 _17568_ (.Y(_00636_),
    .A(_00635_));
 sg13g2_a221oi_1 _17569_ (.B2(data_rdata_i_18_),
    .C1(_00636_),
    .B1(net416),
    .A1(data_rdata_i_10_),
    .Y(_00637_),
    .A2(net1944));
 sg13g2_o21ai_1 _17570_ (.B1(net1600),
    .Y(_00638_),
    .A1(net1707),
    .A2(_00637_));
 sg13g2_a22oi_1 _17571_ (.Y(_00639_),
    .B1(_00638_),
    .B2(net1650),
    .A2(net1060),
    .A1(csr_rdata_18_));
 sg13g2_o21ai_1 _17572_ (.B1(_00639_),
    .Y(rf_wdata_wb_18_),
    .A1(_00624_),
    .A2(_00634_));
 sg13g2_o21ai_1 _17573_ (.B1(net1061),
    .Y(_00640_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .A2(net340));
 sg13g2_mux2_1 _17574_ (.A0(_08696_),
    .A1(_08700_),
    .S(net202),
    .X(_00641_));
 sg13g2_a21oi_1 _17575_ (.A1(net169),
    .A2(net130),
    .Y(_00642_),
    .B1(net1249));
 sg13g2_nand3_1 _17576_ (.B(net169),
    .C(net1360),
    .A(net1248),
    .Y(_00643_));
 sg13g2_o21ai_1 _17577_ (.B1(_00643_),
    .Y(_00644_),
    .A1(net169),
    .A2(net1360));
 sg13g2_a21oi_1 _17578_ (.A1(net1423),
    .A2(_00644_),
    .Y(_00645_),
    .B1(net1419));
 sg13g2_nor2b_1 _17579_ (.A(_00642_),
    .B_N(_00645_),
    .Y(_00646_));
 sg13g2_a221oi_1 _17580_ (.B2(net1366),
    .C1(_00646_),
    .B1(_00641_),
    .A1(data_addr_o_19_),
    .Y(_00647_),
    .A2(net1317));
 sg13g2_o21ai_1 _17581_ (.B1(net377),
    .Y(_00648_),
    .A1(net1196),
    .A2(_00647_));
 sg13g2_nor2b_1 _17582_ (.A(_00640_),
    .B_N(_00648_),
    .Y(_00649_));
 sg13g2_o21ai_1 _17583_ (.B1(_00649_),
    .Y(_00650_),
    .A1(_07003_),
    .A2(_06132_));
 sg13g2_a22oi_1 _17584_ (.Y(_00651_),
    .B1(net1948),
    .B2(data_rdata_i_11_),
    .A2(net1955),
    .A1(\load_store_unit_i.rdata_q_19_ ));
 sg13g2_inv_1 _17585_ (.Y(_00652_),
    .A(_00651_));
 sg13g2_a221oi_1 _17586_ (.B2(data_rdata_i_19_),
    .C1(_00652_),
    .B1(net416),
    .A1(data_rdata_i_3_),
    .Y(_00653_),
    .A2(net1942));
 sg13g2_o21ai_1 _17587_ (.B1(_00583_),
    .Y(_00654_),
    .A1(net1706),
    .A2(_00653_));
 sg13g2_a22oi_1 _17588_ (.Y(_00655_),
    .B1(_00654_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_19_));
 sg13g2_nand2_2 _17589_ (.Y(rf_wdata_wb_19_),
    .A(_00650_),
    .B(_00655_));
 sg13g2_mux4_1 _17590_ (.S0(net1460),
    .A0(net1202),
    .A1(net88),
    .A2(net1350),
    .A3(net1405),
    .S1(net211),
    .X(_00656_));
 sg13g2_mux4_1 _17591_ (.S0(net1459),
    .A0(net150),
    .A1(alu_operand_a_ex_24_),
    .A2(net1279),
    .A3(alu_operand_a_ex_7_),
    .S1(net210),
    .X(_00657_));
 sg13g2_mux2_1 _17592_ (.A0(_00656_),
    .A1(_00657_),
    .S(net1178),
    .X(_00658_));
 sg13g2_mux4_1 _17593_ (.S0(net206),
    .A0(net1199),
    .A1(net1410),
    .A2(net1190),
    .A3(net1411),
    .S1(net1462),
    .X(_00659_));
 sg13g2_nand2b_1 _17594_ (.Y(_00660_),
    .B(_00659_),
    .A_N(net1178));
 sg13g2_mux4_1 _17595_ (.S0(net1460),
    .A0(net123),
    .A1(net1201),
    .A2(net1407),
    .A3(net1408),
    .S1(net211),
    .X(_00661_));
 sg13g2_nand2_1 _17596_ (.Y(_00662_),
    .A(net1178),
    .B(_00661_));
 sg13g2_nand3_1 _17597_ (.B(_00660_),
    .C(_00662_),
    .A(net1165),
    .Y(_00663_));
 sg13g2_o21ai_1 _17598_ (.B1(_00663_),
    .Y(_00664_),
    .A1(net1165),
    .A2(_00658_));
 sg13g2_nor2_1 _17599_ (.A(net1134),
    .B(_00664_),
    .Y(_00665_));
 sg13g2_a21oi_1 _17600_ (.A1(net1134),
    .A2(_00531_),
    .Y(_00666_),
    .B1(_00665_));
 sg13g2_mux4_1 _17601_ (.S0(net199),
    .A0(net151),
    .A1(net127),
    .A2(net194),
    .A3(net196),
    .S1(net1459),
    .X(_00667_));
 sg13g2_mux2_1 _17602_ (.A0(_00667_),
    .A1(_08660_),
    .S(net1175),
    .X(_00668_));
 sg13g2_nor2b_1 _17603_ (.A(net1169),
    .B_N(_00493_),
    .Y(_00669_));
 sg13g2_a21oi_1 _17604_ (.A1(net1169),
    .A2(_00668_),
    .Y(_00670_),
    .B1(_00669_));
 sg13g2_nor2_1 _17605_ (.A(net41),
    .B(_00532_),
    .Y(_00671_));
 sg13g2_a21oi_1 _17606_ (.A1(net43),
    .A2(_00670_),
    .Y(_00672_),
    .B1(_00671_));
 sg13g2_nor2_1 _17607_ (.A(net1137),
    .B(_00672_),
    .Y(_00673_));
 sg13g2_a21oi_1 _17608_ (.A1(net1137),
    .A2(_00666_),
    .Y(_00674_),
    .B1(_00673_));
 sg13g2_mux2_1 _17609_ (.A0(net1133),
    .A1(_00528_),
    .S(_08503_),
    .X(_00675_));
 sg13g2_mux2_1 _17610_ (.A0(_00674_),
    .A1(_00675_),
    .S(net202),
    .X(_00676_));
 sg13g2_nand2_1 _17611_ (.Y(_00677_),
    .A(net1411),
    .B(net128));
 sg13g2_nand2_1 _17612_ (.Y(_00678_),
    .A(_02347_),
    .B(net1355));
 sg13g2_o21ai_1 _17613_ (.B1(_00678_),
    .Y(_00679_),
    .A1(net1411),
    .A2(net1357));
 sg13g2_a221oi_1 _17614_ (.B2(net1422),
    .C1(net1417),
    .B1(_00679_),
    .A1(net1247),
    .Y(_00680_),
    .A2(_00677_));
 sg13g2_a221oi_1 _17615_ (.B2(net1367),
    .C1(_00680_),
    .B1(_00676_),
    .A1(net1112),
    .Y(_00681_),
    .A2(net1318));
 sg13g2_o21ai_1 _17616_ (.B1(net377),
    .Y(_00682_),
    .A1(net1197),
    .A2(_00681_));
 sg13g2_a22oi_1 _17617_ (.Y(_00683_),
    .B1(_08611_),
    .B2(_04147_),
    .A2(net1472),
    .A1(_04185_));
 sg13g2_and3_2 _17618_ (.X(_00684_),
    .A(net396),
    .B(_00682_),
    .C(_00683_));
 sg13g2_a21oi_2 _17619_ (.B1(_00684_),
    .Y(_00685_),
    .A2(net1676),
    .A1(csr_rdata_1_));
 sg13g2_nand2_1 _17620_ (.Y(_00686_),
    .A(\load_store_unit_i.rdata_q_9_ ),
    .B(net1941));
 sg13g2_a22oi_1 _17621_ (.Y(_00687_),
    .B1(net1949),
    .B2(\load_store_unit_i.rdata_q_17_ ),
    .A2(net1957),
    .A1(\load_store_unit_i.rdata_q_1_ ));
 sg13g2_a21oi_1 _17622_ (.A1(_00686_),
    .A2(_00687_),
    .Y(_00688_),
    .B1(net1706));
 sg13g2_a22oi_1 _17623_ (.Y(_00689_),
    .B1(net1956),
    .B2(data_rdata_i_9_),
    .A2(net1940),
    .A1(data_rdata_i_17_));
 sg13g2_a22oi_1 _17624_ (.Y(_00690_),
    .B1(net1934),
    .B2(\load_store_unit_i.rdata_q_17_ ),
    .A2(net1962),
    .A1(data_rdata_i_25_));
 sg13g2_nand2b_1 _17625_ (.Y(_00691_),
    .B(net1949),
    .A_N(_00690_));
 sg13g2_o21ai_1 _17626_ (.B1(_00691_),
    .Y(_00692_),
    .A1(net1704),
    .A2(_00689_));
 sg13g2_mux2_1 _17627_ (.A0(_00692_),
    .A1(data_rdata_i_1_),
    .S(net413),
    .X(_00693_));
 sg13g2_o21ai_1 _17628_ (.B1(net1651),
    .Y(_00694_),
    .A1(_00688_),
    .A2(_00693_));
 sg13g2_o21ai_1 _17629_ (.B1(_00694_),
    .Y(rf_wdata_wb_1_),
    .A1(net1072),
    .A2(_00685_));
 sg13g2_nor2_2 _17630_ (.A(_06238_),
    .B(_08639_),
    .Y(_00695_));
 sg13g2_nand2_1 _17631_ (.Y(_00696_),
    .A(_07002_),
    .B(net297));
 sg13g2_nor3_1 _17632_ (.A(net1576),
    .B(_04393_),
    .C(_00696_),
    .Y(_00697_));
 sg13g2_a21oi_1 _17633_ (.A1(_06147_),
    .A2(net1577),
    .Y(_00698_),
    .B1(_00697_));
 sg13g2_nor2_1 _17634_ (.A(net201),
    .B(_08669_),
    .Y(_00699_));
 sg13g2_a21oi_1 _17635_ (.A1(net203),
    .A2(_08666_),
    .Y(_00700_),
    .B1(_00699_));
 sg13g2_a21o_1 _17636_ (.A2(_02667_),
    .A1(_01882_),
    .B1(_02653_),
    .X(_00701_));
 sg13g2_a21oi_1 _17637_ (.A1(net129),
    .A2(_00701_),
    .Y(_00702_),
    .B1(net1281));
 sg13g2_nand3_1 _17638_ (.B(net1353),
    .C(_00701_),
    .A(net1281),
    .Y(_00703_));
 sg13g2_o21ai_1 _17639_ (.B1(_00703_),
    .Y(_00704_),
    .A1(net1353),
    .A2(_00701_));
 sg13g2_a21oi_1 _17640_ (.A1(net1421),
    .A2(_00704_),
    .Y(_00705_),
    .B1(net1416));
 sg13g2_nor2b_1 _17641_ (.A(_00702_),
    .B_N(_00705_),
    .Y(_00706_));
 sg13g2_a221oi_1 _17642_ (.B2(net1366),
    .C1(_00706_),
    .B1(_00700_),
    .A1(data_addr_o_20_),
    .Y(_00707_),
    .A2(net1317));
 sg13g2_o21ai_1 _17643_ (.B1(net377),
    .Y(_00708_),
    .A1(net1197),
    .A2(_00707_));
 sg13g2_nand3_1 _17644_ (.B(_00698_),
    .C(_00708_),
    .A(net1061),
    .Y(_00709_));
 sg13g2_a22oi_1 _17645_ (.Y(_00710_),
    .B1(net1955),
    .B2(\load_store_unit_i.rdata_q_20_ ),
    .A2(net1939),
    .A1(data_rdata_i_4_));
 sg13g2_inv_1 _17646_ (.Y(_00711_),
    .A(_00710_));
 sg13g2_a221oi_1 _17647_ (.B2(data_rdata_i_20_),
    .C1(_00711_),
    .B1(net416),
    .A1(data_rdata_i_12_),
    .Y(_00712_),
    .A2(net1948));
 sg13g2_o21ai_1 _17648_ (.B1(net1601),
    .Y(_00713_),
    .A1(net1705),
    .A2(_00712_));
 sg13g2_a22oi_1 _17649_ (.Y(_00714_),
    .B1(_00713_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_20_));
 sg13g2_o21ai_1 _17650_ (.B1(_00714_),
    .Y(rf_wdata_wb_20_),
    .A1(_00695_),
    .A2(_00709_));
 sg13g2_a22oi_1 _17651_ (.Y(_00715_),
    .B1(net1958),
    .B2(\load_store_unit_i.rdata_q_21_ ),
    .A2(net1938),
    .A1(data_rdata_i_5_));
 sg13g2_inv_1 _17652_ (.Y(_00716_),
    .A(_00715_));
 sg13g2_a221oi_1 _17653_ (.B2(data_rdata_i_21_),
    .C1(_00716_),
    .B1(net417),
    .A1(data_rdata_i_13_),
    .Y(_00717_),
    .A2(net1946));
 sg13g2_o21ai_1 _17654_ (.B1(net1601),
    .Y(_00718_),
    .A1(net1705),
    .A2(_00717_));
 sg13g2_nor2_1 _17655_ (.A(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .B(net341),
    .Y(_00719_));
 sg13g2_nand2_1 _17656_ (.Y(_00720_),
    .A(net209),
    .B(_08596_));
 sg13g2_o21ai_1 _17657_ (.B1(_00720_),
    .Y(_00721_),
    .A1(net206),
    .A2(_08576_));
 sg13g2_a21oi_1 _17658_ (.A1(net240),
    .A2(net130),
    .Y(_00722_),
    .B1(net126));
 sg13g2_nand2_1 _17659_ (.Y(_00723_),
    .A(_02736_),
    .B(net1360));
 sg13g2_o21ai_1 _17660_ (.B1(_00723_),
    .Y(_00724_),
    .A1(net240),
    .A2(net1360));
 sg13g2_a21oi_1 _17661_ (.A1(net1423),
    .A2(_00724_),
    .Y(_00725_),
    .B1(net1419));
 sg13g2_nor2b_1 _17662_ (.A(_00722_),
    .B_N(_00725_),
    .Y(_00726_));
 sg13g2_a221oi_1 _17663_ (.B2(net1364),
    .C1(_00726_),
    .B1(_00721_),
    .A1(data_addr_o_21_),
    .Y(_00727_),
    .A2(net1315));
 sg13g2_o21ai_1 _17664_ (.B1(net367),
    .Y(_00728_),
    .A1(net1194),
    .A2(_00727_));
 sg13g2_inv_1 _17665_ (.Y(_00729_),
    .A(_00728_));
 sg13g2_nor3_1 _17666_ (.A(net1576),
    .B(_04479_),
    .C(_00696_),
    .Y(_00730_));
 sg13g2_nor4_1 _17667_ (.A(net1680),
    .B(_00719_),
    .C(_00729_),
    .D(_00730_),
    .Y(_00731_));
 sg13g2_a21oi_1 _17668_ (.A1(csr_rdata_21_),
    .A2(net1681),
    .Y(_00732_),
    .B1(_00731_));
 sg13g2_o21ai_1 _17669_ (.B1(net397),
    .Y(_00733_),
    .A1(_06016_),
    .A2(_00719_));
 sg13g2_nor2_1 _17670_ (.A(_06343_),
    .B(_00733_),
    .Y(_00734_));
 sg13g2_nor3_2 _17671_ (.A(net1075),
    .B(_00732_),
    .C(_00734_),
    .Y(_00735_));
 sg13g2_a21o_2 _17672_ (.A2(_00718_),
    .A1(net1648),
    .B1(_00735_),
    .X(rf_wdata_wb_21_));
 sg13g2_a21oi_1 _17673_ (.A1(net43),
    .A2(_00531_),
    .Y(_00736_),
    .B1(_08668_));
 sg13g2_nand2_1 _17674_ (.Y(_00737_),
    .A(net46),
    .B(_00736_));
 sg13g2_o21ai_1 _17675_ (.B1(_00737_),
    .Y(_00738_),
    .A1(net45),
    .A2(_00672_));
 sg13g2_nand2b_1 _17676_ (.Y(_00739_),
    .B(net45),
    .A_N(_00528_));
 sg13g2_o21ai_1 _17677_ (.B1(_00739_),
    .Y(_00740_),
    .A1(net45),
    .A2(_00526_));
 sg13g2_a21oi_1 _17678_ (.A1(net43),
    .A2(_00740_),
    .Y(_00741_),
    .B1(_08595_));
 sg13g2_nand2_1 _17679_ (.Y(_00742_),
    .A(net209),
    .B(_00741_));
 sg13g2_o21ai_1 _17680_ (.B1(_00742_),
    .Y(_00743_),
    .A1(net207),
    .A2(_00738_));
 sg13g2_a21oi_1 _17681_ (.A1(_02642_),
    .A2(net130),
    .Y(_00744_),
    .B1(net195));
 sg13g2_nand2_1 _17682_ (.Y(_00745_),
    .A(_02766_),
    .B(net1362));
 sg13g2_o21ai_1 _17683_ (.B1(_00745_),
    .Y(_00746_),
    .A1(_02642_),
    .A2(net1360));
 sg13g2_a21oi_1 _17684_ (.A1(net1423),
    .A2(_00746_),
    .Y(_00747_),
    .B1(net1419));
 sg13g2_nor2b_1 _17685_ (.A(_00744_),
    .B_N(_00747_),
    .Y(_00748_));
 sg13g2_a221oi_1 _17686_ (.B2(net1366),
    .C1(_00748_),
    .B1(_00743_),
    .A1(data_addr_o_22_),
    .Y(_00749_),
    .A2(net1317));
 sg13g2_nor3_1 _17687_ (.A(_07002_),
    .B(net1196),
    .C(_00749_),
    .Y(_00750_));
 sg13g2_a21o_1 _17688_ (.A2(_06474_),
    .A1(_07002_),
    .B1(_00750_),
    .X(_00751_));
 sg13g2_and3_1 _17689_ (.X(_00752_),
    .A(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .B(net396),
    .C(net1577));
 sg13g2_a221oi_1 _17690_ (.B2(_00751_),
    .C1(_00752_),
    .B1(_00599_),
    .A1(csr_rdata_22_),
    .Y(_00753_),
    .A2(net1679));
 sg13g2_a22oi_1 _17691_ (.Y(_00754_),
    .B1(net1945),
    .B2(data_rdata_i_14_),
    .A2(net1953),
    .A1(\load_store_unit_i.rdata_q_22_ ));
 sg13g2_inv_1 _17692_ (.Y(_00755_),
    .A(_00754_));
 sg13g2_a221oi_1 _17693_ (.B2(data_rdata_i_22_),
    .C1(_00755_),
    .B1(net416),
    .A1(data_rdata_i_6_),
    .Y(_00756_),
    .A2(net1937));
 sg13g2_o21ai_1 _17694_ (.B1(net1600),
    .Y(_00757_),
    .A1(net1705),
    .A2(_00756_));
 sg13g2_nand2_1 _17695_ (.Y(_00758_),
    .A(net1648),
    .B(_00757_));
 sg13g2_o21ai_1 _17696_ (.B1(_00758_),
    .Y(rf_wdata_wb_22_),
    .A1(net1072),
    .A2(_00753_));
 sg13g2_nor2_2 _17697_ (.A(_06563_),
    .B(_08639_),
    .Y(_00759_));
 sg13g2_or2_1 _17698_ (.X(_00760_),
    .B(net340),
    .A(\ex_block_i.alu_i.imd_val_q_i_55_ ));
 sg13g2_nand3_1 _17699_ (.B(_04656_),
    .C(_08609_),
    .A(net342),
    .Y(_00761_));
 sg13g2_mux2_1 _17700_ (.A0(_08508_),
    .A1(_00553_),
    .S(net1139),
    .X(_00762_));
 sg13g2_inv_1 _17701_ (.Y(_00763_),
    .A(_08595_));
 sg13g2_o21ai_1 _17702_ (.B1(_00763_),
    .Y(_00764_),
    .A1(net1135),
    .A2(_00762_));
 sg13g2_inv_1 _17703_ (.Y(_00765_),
    .A(_08497_));
 sg13g2_mux4_1 _17704_ (.S0(net1134),
    .A0(_08471_),
    .A1(_00765_),
    .A2(_08485_),
    .A3(_08509_),
    .S1(net47),
    .X(_00766_));
 sg13g2_or2_1 _17705_ (.X(_00767_),
    .B(_00766_),
    .A(net207));
 sg13g2_o21ai_1 _17706_ (.B1(_00767_),
    .Y(_00768_),
    .A1(net201),
    .A2(_00764_));
 sg13g2_a21oi_1 _17707_ (.A1(net1344),
    .A2(net131),
    .Y(_00769_),
    .B1(net149));
 sg13g2_nand3_1 _17708_ (.B(net1344),
    .C(net1353),
    .A(net150),
    .Y(_00770_));
 sg13g2_o21ai_1 _17709_ (.B1(_00770_),
    .Y(_00771_),
    .A1(_02039_),
    .A2(net1353));
 sg13g2_a21oi_1 _17710_ (.A1(net1422),
    .A2(_00771_),
    .Y(_00772_),
    .B1(net1417));
 sg13g2_nor2b_1 _17711_ (.A(_00769_),
    .B_N(_00772_),
    .Y(_00773_));
 sg13g2_a221oi_1 _17712_ (.B2(net1368),
    .C1(_00773_),
    .B1(_00768_),
    .A1(data_addr_o_23_),
    .Y(_00774_),
    .A2(net1319));
 sg13g2_o21ai_1 _17713_ (.B1(net377),
    .Y(_00775_),
    .A1(net1195),
    .A2(_00774_));
 sg13g2_nand4_1 _17714_ (.B(_00760_),
    .C(_00761_),
    .A(net1061),
    .Y(_00776_),
    .D(_00775_));
 sg13g2_a22oi_1 _17715_ (.Y(_00777_),
    .B1(net1944),
    .B2(data_rdata_i_15_),
    .A2(net1952),
    .A1(\load_store_unit_i.rdata_q_23_ ));
 sg13g2_inv_1 _17716_ (.Y(_00778_),
    .A(_00777_));
 sg13g2_a221oi_1 _17717_ (.B2(data_rdata_i_23_),
    .C1(_00778_),
    .B1(net416),
    .A1(data_rdata_i_7_),
    .Y(_00779_),
    .A2(net1936));
 sg13g2_o21ai_1 _17718_ (.B1(net1600),
    .Y(_00780_),
    .A1(net1707),
    .A2(_00779_));
 sg13g2_a22oi_1 _17719_ (.Y(_00781_),
    .B1(_00780_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_23_));
 sg13g2_o21ai_1 _17720_ (.B1(_00781_),
    .Y(rf_wdata_wb_23_),
    .A1(_00759_),
    .A2(_00776_));
 sg13g2_a22oi_1 _17721_ (.Y(_00782_),
    .B1(net1946),
    .B2(data_rdata_i_16_),
    .A2(net1938),
    .A1(data_rdata_i_8_));
 sg13g2_inv_1 _17722_ (.Y(_00783_),
    .A(_00782_));
 sg13g2_a221oi_1 _17723_ (.B2(data_rdata_i_24_),
    .C1(_00783_),
    .B1(net415),
    .A1(data_rdata_i_0_),
    .Y(_00784_),
    .A2(net1954));
 sg13g2_o21ai_1 _17724_ (.B1(net1600),
    .Y(_00785_),
    .A1(net1707),
    .A2(_00784_));
 sg13g2_nor2_1 _17725_ (.A(csr_rdata_24_),
    .B(net397),
    .Y(_00786_));
 sg13g2_nand2b_1 _17726_ (.Y(_00787_),
    .B(_08662_),
    .A_N(net1162));
 sg13g2_mux2_1 _17727_ (.A0(_00657_),
    .A1(_00667_),
    .S(net1175),
    .X(_00788_));
 sg13g2_nand2_1 _17728_ (.Y(_00789_),
    .A(net1162),
    .B(_00788_));
 sg13g2_nand3_1 _17729_ (.B(_00787_),
    .C(_00789_),
    .A(net1137),
    .Y(_00790_));
 sg13g2_o21ai_1 _17730_ (.B1(_00790_),
    .Y(_00791_),
    .A1(net1139),
    .A2(_00554_));
 sg13g2_nor2_1 _17731_ (.A(net1135),
    .B(_00791_),
    .Y(_00792_));
 sg13g2_a21oi_1 _17732_ (.A1(net1135),
    .A2(_00762_),
    .Y(_00793_),
    .B1(_00792_));
 sg13g2_a21oi_1 _17733_ (.A1(_08497_),
    .A2(net1120),
    .Y(_00794_),
    .B1(_08510_));
 sg13g2_and2_1 _17734_ (.A(net206),
    .B(_00794_),
    .X(_00795_));
 sg13g2_a21oi_1 _17735_ (.A1(net203),
    .A2(_00793_),
    .Y(_00796_),
    .B1(_00795_));
 sg13g2_a21oi_1 _17736_ (.A1(_02060_),
    .A2(net132),
    .Y(_00797_),
    .B1(net125));
 sg13g2_nand3_1 _17737_ (.B(_02060_),
    .C(net1361),
    .A(net125),
    .Y(_00798_));
 sg13g2_o21ai_1 _17738_ (.B1(_00798_),
    .Y(_00799_),
    .A1(_02060_),
    .A2(net1361));
 sg13g2_a21oi_1 _17739_ (.A1(net1423),
    .A2(_00799_),
    .Y(_00800_),
    .B1(net1419));
 sg13g2_nor2b_1 _17740_ (.A(_00797_),
    .B_N(_00800_),
    .Y(_00801_));
 sg13g2_a221oi_1 _17741_ (.B2(net1364),
    .C1(_00801_),
    .B1(_00796_),
    .A1(data_addr_o_24_),
    .Y(_00802_),
    .A2(net1315));
 sg13g2_o21ai_1 _17742_ (.B1(net374),
    .Y(_00803_),
    .A1(net1194),
    .A2(_00802_));
 sg13g2_nor2_1 _17743_ (.A(net1677),
    .B(_00803_),
    .Y(_00804_));
 sg13g2_nor4_1 _17744_ (.A(_04030_),
    .B(net1075),
    .C(_00786_),
    .D(_00804_),
    .Y(_00805_));
 sg13g2_nand2_1 _17745_ (.Y(_00806_),
    .A(csr_rdata_24_),
    .B(net1677));
 sg13g2_or2_1 _17746_ (.X(_00807_),
    .B(net339),
    .A(net556));
 sg13g2_nand4_1 _17747_ (.B(_07003_),
    .C(_00803_),
    .A(net397),
    .Y(_00808_),
    .D(_00807_));
 sg13g2_a21oi_1 _17748_ (.A1(_00806_),
    .A2(_00808_),
    .Y(_00809_),
    .B1(net1075));
 sg13g2_a221oi_1 _17749_ (.B2(_06653_),
    .C1(_00809_),
    .B1(_00805_),
    .A1(net1650),
    .Y(_00810_),
    .A2(_00785_));
 sg13g2_inv_2 _17750_ (.Y(rf_wdata_wb_24_),
    .A(_00810_));
 sg13g2_nand2b_1 _17751_ (.Y(_00811_),
    .B(_08571_),
    .A_N(net1166));
 sg13g2_mux2_1 _17752_ (.A0(_08452_),
    .A1(_08462_),
    .S(net1177),
    .X(_00812_));
 sg13g2_nand2_1 _17753_ (.Y(_00813_),
    .A(net1166),
    .B(_00812_));
 sg13g2_nand3_1 _17754_ (.B(_00811_),
    .C(_00813_),
    .A(net1138),
    .Y(_00814_));
 sg13g2_o21ai_1 _17755_ (.B1(_00814_),
    .Y(_00815_),
    .A1(net1136),
    .A2(_00529_));
 sg13g2_mux2_1 _17756_ (.A0(_00740_),
    .A1(_00815_),
    .S(net42),
    .X(_00816_));
 sg13g2_a21oi_1 _17757_ (.A1(net1120),
    .A2(_00532_),
    .Y(_00817_),
    .B1(_08510_));
 sg13g2_and2_1 _17758_ (.A(net206),
    .B(_00817_),
    .X(_00818_));
 sg13g2_a21oi_1 _17759_ (.A1(net203),
    .A2(_00816_),
    .Y(_00819_),
    .B1(_00818_));
 sg13g2_nand3_1 _17760_ (.B(_01993_),
    .C(net1362),
    .A(net1202),
    .Y(_00820_));
 sg13g2_o21ai_1 _17761_ (.B1(_00820_),
    .Y(_00821_),
    .A1(_01993_),
    .A2(net1361));
 sg13g2_a21oi_1 _17762_ (.A1(_01993_),
    .A2(net130),
    .Y(_00822_),
    .B1(net1202));
 sg13g2_nand2b_1 _17763_ (.Y(_00823_),
    .B(_08545_),
    .A_N(_00822_));
 sg13g2_a21oi_1 _17764_ (.A1(net1425),
    .A2(_00821_),
    .Y(_00824_),
    .B1(_00823_));
 sg13g2_a221oi_1 _17765_ (.B2(net1364),
    .C1(_00824_),
    .B1(_00819_),
    .A1(data_addr_o_25_),
    .Y(_00825_),
    .A2(net1315));
 sg13g2_or2_1 _17766_ (.X(_00826_),
    .B(_00825_),
    .A(net1195));
 sg13g2_nand2_1 _17767_ (.Y(_00827_),
    .A(net1540),
    .B(_06738_));
 sg13g2_o21ai_1 _17768_ (.B1(_00827_),
    .Y(_00828_),
    .A1(net1540),
    .A2(_04901_));
 sg13g2_o21ai_1 _17769_ (.B1(net1061),
    .Y(_00829_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .A2(net340));
 sg13g2_a221oi_1 _17770_ (.B2(_06016_),
    .C1(_00829_),
    .B1(_00828_),
    .A1(net381),
    .Y(_00830_),
    .A2(_00826_));
 sg13g2_a22oi_1 _17771_ (.Y(_00831_),
    .B1(net1949),
    .B2(data_rdata_i_17_),
    .A2(net1940),
    .A1(data_rdata_i_9_));
 sg13g2_inv_1 _17772_ (.Y(_00832_),
    .A(_00831_));
 sg13g2_a221oi_1 _17773_ (.B2(data_rdata_i_25_),
    .C1(_00832_),
    .B1(net416),
    .A1(data_rdata_i_1_),
    .Y(_00833_),
    .A2(net1956));
 sg13g2_o21ai_1 _17774_ (.B1(net1601),
    .Y(_00834_),
    .A1(net1705),
    .A2(_00833_));
 sg13g2_a22oi_1 _17775_ (.Y(_00835_),
    .B1(_00834_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_25_));
 sg13g2_nand2b_2 _17776_ (.Y(rf_wdata_wb_25_),
    .B(_00835_),
    .A_N(_00830_));
 sg13g2_nor2_1 _17777_ (.A(_06800_),
    .B(_08639_),
    .Y(_00836_));
 sg13g2_or2_1 _17778_ (.X(_00837_),
    .B(net340),
    .A(\ex_block_i.alu_i.imd_val_q_i_58_ ));
 sg13g2_nand3_1 _17779_ (.B(_05012_),
    .C(_08609_),
    .A(net342),
    .Y(_00838_));
 sg13g2_a21oi_1 _17780_ (.A1(net1120),
    .A2(_00499_),
    .Y(_00839_),
    .B1(_08510_));
 sg13g2_mux2_1 _17781_ (.A0(_00668_),
    .A1(_00658_),
    .S(net1162),
    .X(_00840_));
 sg13g2_mux2_1 _17782_ (.A0(_08585_),
    .A1(_00840_),
    .S(net41),
    .X(_00841_));
 sg13g2_nand2_1 _17783_ (.Y(_00842_),
    .A(net1139),
    .B(_00841_));
 sg13g2_o21ai_1 _17784_ (.B1(_00842_),
    .Y(_00843_),
    .A1(net1139),
    .A2(_00496_));
 sg13g2_nor2_1 _17785_ (.A(net208),
    .B(_00843_),
    .Y(_00844_));
 sg13g2_a21oi_1 _17786_ (.A1(net212),
    .A2(_00839_),
    .Y(_00845_),
    .B1(_00844_));
 sg13g2_nand2_1 _17787_ (.Y(_00846_),
    .A(_02800_),
    .B(net1360));
 sg13g2_o21ai_1 _17788_ (.B1(_00846_),
    .Y(_00847_),
    .A1(net1278),
    .A2(net1361));
 sg13g2_a21oi_1 _17789_ (.A1(net1278),
    .A2(net130),
    .Y(_00848_),
    .B1(net87));
 sg13g2_nand2b_1 _17790_ (.Y(_00849_),
    .B(_08545_),
    .A_N(_00848_));
 sg13g2_a21oi_1 _17791_ (.A1(net1423),
    .A2(_00847_),
    .Y(_00850_),
    .B1(_00849_));
 sg13g2_a221oi_1 _17792_ (.B2(net1365),
    .C1(_00850_),
    .B1(_00845_),
    .A1(data_addr_o_26_),
    .Y(_00851_),
    .A2(net1316));
 sg13g2_o21ai_1 _17793_ (.B1(net376),
    .Y(_00852_),
    .A1(net1195),
    .A2(_00851_));
 sg13g2_nand4_1 _17794_ (.B(_00837_),
    .C(_00838_),
    .A(net1061),
    .Y(_00853_),
    .D(_00852_));
 sg13g2_a22oi_1 _17795_ (.Y(_00854_),
    .B1(net1944),
    .B2(data_rdata_i_18_),
    .A2(net1935),
    .A1(data_rdata_i_10_));
 sg13g2_inv_1 _17796_ (.Y(_00855_),
    .A(_00854_));
 sg13g2_a221oi_1 _17797_ (.B2(data_rdata_i_26_),
    .C1(_00855_),
    .B1(net416),
    .A1(data_rdata_i_2_),
    .Y(_00856_),
    .A2(net1952));
 sg13g2_o21ai_1 _17798_ (.B1(net1600),
    .Y(_00857_),
    .A1(net1707),
    .A2(_00856_));
 sg13g2_a22oi_1 _17799_ (.Y(_00858_),
    .B1(_00857_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_26_));
 sg13g2_o21ai_1 _17800_ (.B1(_00858_),
    .Y(rf_wdata_wb_26_),
    .A1(_00836_),
    .A2(_00853_));
 sg13g2_nor2_1 _17801_ (.A(_06880_),
    .B(_08639_),
    .Y(_00859_));
 sg13g2_mux4_1 _17802_ (.S0(net1164),
    .A0(_08464_),
    .A1(_08455_),
    .A2(_08480_),
    .A3(_08469_),
    .S1(net47),
    .X(_00860_));
 sg13g2_mux2_1 _17803_ (.A0(_08667_),
    .A1(_00860_),
    .S(net41),
    .X(_00861_));
 sg13g2_nor2_1 _17804_ (.A(net1133),
    .B(net1120),
    .Y(_00862_));
 sg13g2_a21oi_1 _17805_ (.A1(net1120),
    .A2(_08646_),
    .Y(_00863_),
    .B1(_00862_));
 sg13g2_mux2_1 _17806_ (.A0(_00861_),
    .A1(_00863_),
    .S(net208),
    .X(_00864_));
 sg13g2_a21oi_1 _17807_ (.A1(_01896_),
    .A2(net131),
    .Y(_00865_),
    .B1(net122));
 sg13g2_nand3_1 _17808_ (.B(_01896_),
    .C(net1358),
    .A(net123),
    .Y(_00866_));
 sg13g2_o21ai_1 _17809_ (.B1(_00866_),
    .Y(_00867_),
    .A1(_01896_),
    .A2(net1358));
 sg13g2_a21oi_1 _17810_ (.A1(net1424),
    .A2(_00867_),
    .Y(_00868_),
    .B1(net1418));
 sg13g2_nor2b_1 _17811_ (.A(_00865_),
    .B_N(_00868_),
    .Y(_00869_));
 sg13g2_a221oi_1 _17812_ (.B2(net1365),
    .C1(_00869_),
    .B1(_00864_),
    .A1(data_addr_o_27_),
    .Y(_00870_),
    .A2(net1316));
 sg13g2_o21ai_1 _17813_ (.B1(net375),
    .Y(_00871_),
    .A1(net1195),
    .A2(_00870_));
 sg13g2_nor3_1 _17814_ (.A(net1576),
    .B(_05128_),
    .C(_00696_),
    .Y(_00872_));
 sg13g2_a21oi_1 _17815_ (.A1(_01899_),
    .A2(net1576),
    .Y(_00873_),
    .B1(_00872_));
 sg13g2_nand3_1 _17816_ (.B(_00871_),
    .C(_00873_),
    .A(_00615_),
    .Y(_00874_));
 sg13g2_a22oi_1 _17817_ (.Y(_00875_),
    .B1(net1948),
    .B2(data_rdata_i_19_),
    .A2(net1939),
    .A1(data_rdata_i_11_));
 sg13g2_inv_1 _17818_ (.Y(_00876_),
    .A(_00875_));
 sg13g2_a221oi_1 _17819_ (.B2(data_rdata_i_27_),
    .C1(_00876_),
    .B1(net415),
    .A1(data_rdata_i_3_),
    .Y(_00877_),
    .A2(net1955));
 sg13g2_o21ai_1 _17820_ (.B1(net1601),
    .Y(_00878_),
    .A1(net1705),
    .A2(_00877_));
 sg13g2_a22oi_1 _17821_ (.Y(_00879_),
    .B1(_00878_),
    .B2(net1649),
    .A2(net1060),
    .A1(csr_rdata_27_));
 sg13g2_o21ai_1 _17822_ (.B1(_00879_),
    .Y(rf_wdata_wb_27_),
    .A1(_00859_),
    .A2(_00874_));
 sg13g2_nand2_1 _17823_ (.Y(_00880_),
    .A(net1178),
    .B(_00656_));
 sg13g2_nand2b_1 _17824_ (.Y(_00881_),
    .B(_00661_),
    .A_N(net1178));
 sg13g2_nand3_1 _17825_ (.B(_00880_),
    .C(_00881_),
    .A(net1165),
    .Y(_00882_));
 sg13g2_o21ai_1 _17826_ (.B1(_00882_),
    .Y(_00883_),
    .A1(net1165),
    .A2(_00788_));
 sg13g2_nor2_1 _17827_ (.A(net42),
    .B(_08694_),
    .Y(_00884_));
 sg13g2_a221oi_1 _17828_ (.B2(_08503_),
    .C1(_00884_),
    .B1(_00883_),
    .A1(net46),
    .Y(_00885_),
    .A2(_08664_));
 sg13g2_nand2_1 _17829_ (.Y(_00886_),
    .A(net1168),
    .B(_08503_));
 sg13g2_mux2_1 _17830_ (.A0(_08493_),
    .A1(net1133),
    .S(_00886_),
    .X(_00887_));
 sg13g2_mux2_1 _17831_ (.A0(_00885_),
    .A1(_00887_),
    .S(net207),
    .X(_00888_));
 sg13g2_a21oi_1 _17832_ (.A1(net1346),
    .A2(net131),
    .Y(_00889_),
    .B1(net1200));
 sg13g2_nand3_1 _17833_ (.B(net1346),
    .C(net1358),
    .A(net1200),
    .Y(_00890_));
 sg13g2_o21ai_1 _17834_ (.B1(_00890_),
    .Y(_00891_),
    .A1(_01936_),
    .A2(net1358));
 sg13g2_a21oi_1 _17835_ (.A1(net1423),
    .A2(_00891_),
    .Y(_00892_),
    .B1(net1419));
 sg13g2_nor2b_1 _17836_ (.A(_00889_),
    .B_N(_00892_),
    .Y(_00893_));
 sg13g2_a221oi_1 _17837_ (.B2(net1364),
    .C1(_00893_),
    .B1(_00888_),
    .A1(data_addr_o_28_),
    .Y(_00894_),
    .A2(net1315));
 sg13g2_o21ai_1 _17838_ (.B1(net375),
    .Y(_00895_),
    .A1(net1194),
    .A2(_00894_));
 sg13g2_o21ai_1 _17839_ (.B1(_07002_),
    .Y(_00896_),
    .A1(net1540),
    .A2(_05262_));
 sg13g2_nand2_1 _17840_ (.Y(_00897_),
    .A(_06894_),
    .B(net1578));
 sg13g2_o21ai_1 _17841_ (.B1(_00897_),
    .Y(_00898_),
    .A1(net1576),
    .A2(_00896_));
 sg13g2_o21ai_1 _17842_ (.B1(_00898_),
    .Y(_00899_),
    .A1(_04044_),
    .A2(_06985_));
 sg13g2_nand3_1 _17843_ (.B(_00895_),
    .C(_00899_),
    .A(net1061),
    .Y(_00900_));
 sg13g2_a22oi_1 _17844_ (.Y(_00901_),
    .B1(net1948),
    .B2(data_rdata_i_20_),
    .A2(net1939),
    .A1(data_rdata_i_12_));
 sg13g2_inv_1 _17845_ (.Y(_00902_),
    .A(_00901_));
 sg13g2_a221oi_1 _17846_ (.B2(data_rdata_i_28_),
    .C1(_00902_),
    .B1(net415),
    .A1(data_rdata_i_4_),
    .Y(_00903_),
    .A2(net1955));
 sg13g2_o21ai_1 _17847_ (.B1(net1601),
    .Y(_00904_),
    .A1(net1705),
    .A2(_00903_));
 sg13g2_a22oi_1 _17848_ (.Y(_00905_),
    .B1(_00904_),
    .B2(net1649),
    .A2(_00621_),
    .A1(csr_rdata_28_));
 sg13g2_nand2_2 _17849_ (.Y(rf_wdata_wb_28_),
    .A(_00900_),
    .B(_00905_));
 sg13g2_nor2b_1 _17850_ (.A(net1179),
    .B_N(_08442_),
    .Y(_00906_));
 sg13g2_a21oi_1 _17851_ (.A1(net1179),
    .A2(_08451_),
    .Y(_00907_),
    .B1(_00906_));
 sg13g2_nor2_1 _17852_ (.A(net1167),
    .B(_00812_),
    .Y(_00908_));
 sg13g2_a21oi_1 _17853_ (.A1(net1166),
    .A2(_00907_),
    .Y(_00909_),
    .B1(_00908_));
 sg13g2_nand2_1 _17854_ (.Y(_00910_),
    .A(net1138),
    .B(_00909_));
 sg13g2_o21ai_1 _17855_ (.B1(_00910_),
    .Y(_00911_),
    .A1(net1136),
    .A2(_08574_));
 sg13g2_mux2_1 _17856_ (.A0(_00501_),
    .A1(_00911_),
    .S(net42),
    .X(_00912_));
 sg13g2_inv_1 _17857_ (.Y(_00913_),
    .A(_08592_));
 sg13g2_a21o_1 _17858_ (.A2(_00913_),
    .A1(net1120),
    .B1(_08510_),
    .X(_00914_));
 sg13g2_mux2_1 _17859_ (.A0(_00912_),
    .A1(_00914_),
    .S(net207),
    .X(_00915_));
 sg13g2_a21oi_1 _17860_ (.A1(_01964_),
    .A2(net131),
    .Y(_00916_),
    .B1(net1198));
 sg13g2_nand3_1 _17861_ (.B(_01964_),
    .C(net1360),
    .A(net1198),
    .Y(_00917_));
 sg13g2_o21ai_1 _17862_ (.B1(_00917_),
    .Y(_00918_),
    .A1(net1345),
    .A2(net1360));
 sg13g2_a21oi_1 _17863_ (.A1(net1423),
    .A2(_00918_),
    .Y(_00919_),
    .B1(net1419));
 sg13g2_nor2b_1 _17864_ (.A(_00916_),
    .B_N(_00919_),
    .Y(_00920_));
 sg13g2_a221oi_1 _17865_ (.B2(net1364),
    .C1(_00920_),
    .B1(_00915_),
    .A1(data_addr_o_29_),
    .Y(_00921_),
    .A2(net1315));
 sg13g2_a21oi_1 _17866_ (.A1(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .A2(_04030_),
    .Y(_00922_),
    .B1(net1680));
 sg13g2_o21ai_1 _17867_ (.B1(_00922_),
    .Y(_00923_),
    .A1(_08548_),
    .A2(_00921_));
 sg13g2_nor2_2 _17868_ (.A(_07050_),
    .B(_00923_),
    .Y(_00924_));
 sg13g2_o21ai_1 _17869_ (.B1(_08552_),
    .Y(_00925_),
    .A1(csr_rdata_29_),
    .A2(net396));
 sg13g2_a22oi_1 _17870_ (.Y(_00926_),
    .B1(net1946),
    .B2(data_rdata_i_21_),
    .A2(net1938),
    .A1(data_rdata_i_13_));
 sg13g2_inv_1 _17871_ (.Y(_00927_),
    .A(_00926_));
 sg13g2_a221oi_1 _17872_ (.B2(data_rdata_i_29_),
    .C1(_00927_),
    .B1(net416),
    .A1(data_rdata_i_5_),
    .Y(_00928_),
    .A2(net1956));
 sg13g2_o21ai_1 _17873_ (.B1(net1600),
    .Y(_00929_),
    .A1(net1705),
    .A2(_00928_));
 sg13g2_nand2_2 _17874_ (.Y(_00930_),
    .A(net1648),
    .B(_00929_));
 sg13g2_o21ai_1 _17875_ (.B1(_00930_),
    .Y(rf_wdata_wb_29_),
    .A1(_00924_),
    .A2(_00925_));
 sg13g2_mux2_1 _17876_ (.A0(_00912_),
    .A1(_00914_),
    .S(net202),
    .X(_00931_));
 sg13g2_a21oi_1 _17877_ (.A1(net1398),
    .A2(net130),
    .Y(_00932_),
    .B1(net1409));
 sg13g2_nand3_1 _17878_ (.B(net1398),
    .C(net1356),
    .A(net1409),
    .Y(_00933_));
 sg13g2_o21ai_1 _17879_ (.B1(_00933_),
    .Y(_00934_),
    .A1(net1398),
    .A2(net1356));
 sg13g2_a21oi_1 _17880_ (.A1(net1422),
    .A2(_00934_),
    .Y(_00935_),
    .B1(net1417));
 sg13g2_nor2b_1 _17881_ (.A(_00932_),
    .B_N(_00935_),
    .Y(_00936_));
 sg13g2_a221oi_1 _17882_ (.B2(net1364),
    .C1(_00936_),
    .B1(_00931_),
    .A1(data_addr_o_2_),
    .Y(_00937_),
    .A2(net1316));
 sg13g2_o21ai_1 _17883_ (.B1(net376),
    .Y(_00938_),
    .A1(net1194),
    .A2(_00937_));
 sg13g2_a22oi_1 _17884_ (.Y(_00939_),
    .B1(_08611_),
    .B2(_04190_),
    .A2(_07195_),
    .A1(_04264_));
 sg13g2_and3_1 _17885_ (.X(_00940_),
    .A(net396),
    .B(_00938_),
    .C(_00939_));
 sg13g2_a21oi_2 _17886_ (.B1(_00940_),
    .Y(_00941_),
    .A2(net1676),
    .A1(csr_rdata_2_));
 sg13g2_nand2_1 _17887_ (.Y(_00942_),
    .A(\load_store_unit_i.rdata_q_2_ ),
    .B(net1951));
 sg13g2_a22oi_1 _17888_ (.Y(_00943_),
    .B1(net1944),
    .B2(\load_store_unit_i.rdata_q_18_ ),
    .A2(net1935),
    .A1(\load_store_unit_i.rdata_q_10_ ));
 sg13g2_a21oi_1 _17889_ (.A1(_00942_),
    .A2(_00943_),
    .Y(_00944_),
    .B1(net1707));
 sg13g2_a22oi_1 _17890_ (.Y(_00945_),
    .B1(net1951),
    .B2(data_rdata_i_10_),
    .A2(net1935),
    .A1(data_rdata_i_18_));
 sg13g2_a22oi_1 _17891_ (.Y(_00946_),
    .B1(net1931),
    .B2(\load_store_unit_i.rdata_q_18_ ),
    .A2(net1960),
    .A1(data_rdata_i_26_));
 sg13g2_nand2b_1 _17892_ (.Y(_00947_),
    .B(net1944),
    .A_N(_00946_));
 sg13g2_o21ai_1 _17893_ (.B1(_00947_),
    .Y(_00948_),
    .A1(net1704),
    .A2(_00945_));
 sg13g2_mux2_1 _17894_ (.A0(_00948_),
    .A1(data_rdata_i_2_),
    .S(net413),
    .X(_00949_));
 sg13g2_o21ai_1 _17895_ (.B1(net1651),
    .Y(_00950_),
    .A1(_00944_),
    .A2(_00949_));
 sg13g2_o21ai_1 _17896_ (.B1(_00950_),
    .Y(rf_wdata_wb_2_),
    .A1(net1074),
    .A2(_00941_));
 sg13g2_a22oi_1 _17897_ (.Y(_00951_),
    .B1(net1945),
    .B2(data_rdata_i_22_),
    .A2(net1937),
    .A1(data_rdata_i_14_));
 sg13g2_inv_1 _17898_ (.Y(_00952_),
    .A(_00951_));
 sg13g2_a221oi_1 _17899_ (.B2(data_rdata_i_30_),
    .C1(_00952_),
    .B1(net415),
    .A1(data_rdata_i_6_),
    .Y(_00953_),
    .A2(net1953));
 sg13g2_nand2b_1 _17900_ (.Y(_00954_),
    .B(net1704),
    .A_N(_00953_));
 sg13g2_a21o_2 _17901_ (.A2(_00954_),
    .A1(net1600),
    .B1(net1646),
    .X(_00955_));
 sg13g2_o21ai_1 _17902_ (.B1(_08552_),
    .Y(_00956_),
    .A1(csr_rdata_30_),
    .A2(net396));
 sg13g2_mux2_1 _17903_ (.A0(_00674_),
    .A1(_00675_),
    .S(net207),
    .X(_00957_));
 sg13g2_nand3_1 _17904_ (.B(_01867_),
    .C(net1361),
    .A(net1190),
    .Y(_00958_));
 sg13g2_o21ai_1 _17905_ (.B1(_00958_),
    .Y(_00959_),
    .A1(_01867_),
    .A2(net1361));
 sg13g2_a21oi_1 _17906_ (.A1(_01867_),
    .A2(net132),
    .Y(_00960_),
    .B1(net1190));
 sg13g2_nand2b_1 _17907_ (.Y(_00961_),
    .B(_08545_),
    .A_N(_00960_));
 sg13g2_a21oi_1 _17908_ (.A1(net1423),
    .A2(_00959_),
    .Y(_00962_),
    .B1(_00961_));
 sg13g2_a221oi_1 _17909_ (.B2(net1366),
    .C1(_00962_),
    .B1(_00957_),
    .A1(data_addr_o_30_),
    .Y(_00963_),
    .A2(net1317));
 sg13g2_or2_1 _17910_ (.X(_00964_),
    .B(_00963_),
    .A(_08548_));
 sg13g2_a21oi_2 _17911_ (.B1(net1680),
    .Y(_00965_),
    .A2(net1577),
    .A1(\ex_block_i.alu_i.imd_val_q_i_62_ ));
 sg13g2_and3_1 _17912_ (.X(_00966_),
    .A(_00955_),
    .B(_00964_),
    .C(_00965_));
 sg13g2_a22oi_1 _17913_ (.Y(rf_wdata_wb_30_),
    .B1(_00966_),
    .B2(_07103_),
    .A2(_00956_),
    .A1(_00955_));
 sg13g2_a22oi_1 _17914_ (.Y(_00967_),
    .B1(net1944),
    .B2(data_rdata_i_23_),
    .A2(net1936),
    .A1(data_rdata_i_15_));
 sg13g2_inv_1 _17915_ (.Y(_00968_),
    .A(_00967_));
 sg13g2_a221oi_1 _17916_ (.B2(data_rdata_i_31_),
    .C1(_00968_),
    .B1(net415),
    .A1(data_rdata_i_7_),
    .Y(_00969_),
    .A2(net1952));
 sg13g2_nand2b_1 _17917_ (.Y(_00970_),
    .B(net1704),
    .A_N(_00969_));
 sg13g2_a21oi_2 _17918_ (.B1(net1646),
    .Y(_00971_),
    .A2(_00970_),
    .A1(net1600));
 sg13g2_nor3_2 _17919_ (.A(_01846_),
    .B(net376),
    .C(net342),
    .Y(_00972_));
 sg13g2_mux2_1 _17920_ (.A0(_08501_),
    .A1(_08511_),
    .S(net207),
    .X(_00973_));
 sg13g2_nand2_1 _17921_ (.Y(_00974_),
    .A(net81),
    .B(net128));
 sg13g2_nand3_1 _17922_ (.B(_01813_),
    .C(net1354),
    .A(net81),
    .Y(_00975_));
 sg13g2_o21ai_1 _17923_ (.B1(_00975_),
    .Y(_00976_),
    .A1(net81),
    .A2(net1354));
 sg13g2_a221oi_1 _17924_ (.B2(net1421),
    .C1(net1416),
    .B1(_00976_),
    .A1(_01808_),
    .Y(_00977_),
    .A2(_00974_));
 sg13g2_a221oi_1 _17925_ (.B2(net1368),
    .C1(_00977_),
    .B1(_00973_),
    .A1(net37),
    .Y(_00978_),
    .A2(net1319));
 sg13g2_nor2_1 _17926_ (.A(_08548_),
    .B(_00978_),
    .Y(_00979_));
 sg13g2_nor4_1 _17927_ (.A(net1677),
    .B(_00971_),
    .C(_00972_),
    .D(_00979_),
    .Y(_00980_));
 sg13g2_nand2b_1 _17928_ (.Y(_00981_),
    .B(net1678),
    .A_N(csr_rdata_31_));
 sg13g2_a21oi_1 _17929_ (.A1(_08552_),
    .A2(_00981_),
    .Y(_00982_),
    .B1(_00971_));
 sg13g2_a21oi_2 _17930_ (.B1(_00982_),
    .Y(rf_wdata_wb_31_),
    .A2(_00980_),
    .A1(_07153_));
 sg13g2_mux2_1 _17931_ (.A0(_00885_),
    .A1(_00887_),
    .S(net201),
    .X(_00983_));
 sg13g2_a21oi_1 _17932_ (.A1(_02287_),
    .A2(net131),
    .Y(_00984_),
    .B1(net1408));
 sg13g2_nand3_1 _17933_ (.B(_02287_),
    .C(net1356),
    .A(net1408),
    .Y(_00985_));
 sg13g2_o21ai_1 _17934_ (.B1(_00985_),
    .Y(_00986_),
    .A1(_02287_),
    .A2(net1359));
 sg13g2_a21oi_1 _17935_ (.A1(net1424),
    .A2(_00986_),
    .Y(_00987_),
    .B1(net1418));
 sg13g2_nor2b_1 _17936_ (.A(_00984_),
    .B_N(_00987_),
    .Y(_00988_));
 sg13g2_a221oi_1 _17937_ (.B2(net1367),
    .C1(_00988_),
    .B1(_00983_),
    .A1(data_addr_o_3_),
    .Y(_00989_),
    .A2(net1318));
 sg13g2_nor4_1 _17938_ (.A(net1577),
    .B(_07002_),
    .C(net1197),
    .D(_00989_),
    .Y(_00990_));
 sg13g2_a221oi_1 _17939_ (.B2(\ex_block_i.alu_i.imd_val_q_i_35_ ),
    .C1(net1679),
    .B1(_08611_),
    .A1(_04326_),
    .Y(_00991_),
    .A2(net1472));
 sg13g2_nor2b_2 _17940_ (.A(_00990_),
    .B_N(_00991_),
    .Y(_00992_));
 sg13g2_o21ai_1 _17941_ (.B1(_08552_),
    .Y(_00993_),
    .A1(csr_rdata_3_),
    .A2(net396));
 sg13g2_nand2_1 _17942_ (.Y(_00994_),
    .A(\load_store_unit_i.rdata_q_3_ ),
    .B(net1955));
 sg13g2_a22oi_1 _17943_ (.Y(_00995_),
    .B1(net1948),
    .B2(\load_store_unit_i.rdata_q_19_ ),
    .A2(net1939),
    .A1(\load_store_unit_i.rdata_q_11_ ));
 sg13g2_a21oi_1 _17944_ (.A1(_00994_),
    .A2(_00995_),
    .Y(_00996_),
    .B1(net1706));
 sg13g2_a22oi_1 _17945_ (.Y(_00997_),
    .B1(net1955),
    .B2(data_rdata_i_11_),
    .A2(net1939),
    .A1(data_rdata_i_19_));
 sg13g2_a22oi_1 _17946_ (.Y(_00998_),
    .B1(net1932),
    .B2(\load_store_unit_i.rdata_q_19_ ),
    .A2(net1961),
    .A1(data_rdata_i_27_));
 sg13g2_nand2b_1 _17947_ (.Y(_00999_),
    .B(net1948),
    .A_N(_00998_));
 sg13g2_o21ai_1 _17948_ (.B1(_00999_),
    .Y(_01000_),
    .A1(net1704),
    .A2(_00997_));
 sg13g2_mux2_1 _17949_ (.A0(_01000_),
    .A1(data_rdata_i_3_),
    .S(net413),
    .X(_01001_));
 sg13g2_o21ai_1 _17950_ (.B1(net1648),
    .Y(_01002_),
    .A1(_00996_),
    .A2(_01001_));
 sg13g2_o21ai_1 _17951_ (.B1(_01002_),
    .Y(rf_wdata_wb_3_),
    .A1(_00992_),
    .A2(_00993_));
 sg13g2_mux2_1 _17952_ (.A0(_00861_),
    .A1(_00863_),
    .S(net200),
    .X(_01003_));
 sg13g2_a21oi_1 _17953_ (.A1(net1399),
    .A2(net131),
    .Y(_01004_),
    .B1(net1406));
 sg13g2_nand3_1 _17954_ (.B(net1399),
    .C(net1358),
    .A(net1406),
    .Y(_01005_));
 sg13g2_o21ai_1 _17955_ (.B1(_01005_),
    .Y(_01006_),
    .A1(_02259_),
    .A2(net1359));
 sg13g2_a21oi_1 _17956_ (.A1(net1424),
    .A2(_01006_),
    .Y(_01007_),
    .B1(net1418));
 sg13g2_nor2b_1 _17957_ (.A(_01004_),
    .B_N(_01007_),
    .Y(_01008_));
 sg13g2_a221oi_1 _17958_ (.B2(net1365),
    .C1(_01008_),
    .B1(_01003_),
    .A1(data_addr_o_4_),
    .Y(_01009_),
    .A2(net1316));
 sg13g2_or2_1 _17959_ (.X(_01010_),
    .B(_01009_),
    .A(net1195));
 sg13g2_o21ai_1 _17960_ (.B1(_07003_),
    .Y(_01011_),
    .A1(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .A2(net340));
 sg13g2_a221oi_1 _17961_ (.B2(_04396_),
    .C1(net1680),
    .B1(_01011_),
    .A1(net381),
    .Y(_01012_),
    .A2(_01010_));
 sg13g2_a21oi_2 _17962_ (.B1(_01012_),
    .Y(_01013_),
    .A2(net1676),
    .A1(csr_rdata_4_));
 sg13g2_nand2_1 _17963_ (.Y(_01014_),
    .A(\load_store_unit_i.rdata_q_4_ ),
    .B(net1955));
 sg13g2_a22oi_1 _17964_ (.Y(_01015_),
    .B1(net1948),
    .B2(\load_store_unit_i.rdata_q_20_ ),
    .A2(net1941),
    .A1(\load_store_unit_i.rdata_q_12_ ));
 sg13g2_a21oi_1 _17965_ (.A1(_01014_),
    .A2(_01015_),
    .Y(_01016_),
    .B1(net1706));
 sg13g2_a22oi_1 _17966_ (.Y(_01017_),
    .B1(net1956),
    .B2(data_rdata_i_12_),
    .A2(net1940),
    .A1(data_rdata_i_20_));
 sg13g2_a22oi_1 _17967_ (.Y(_01018_),
    .B1(net1933),
    .B2(\load_store_unit_i.rdata_q_20_ ),
    .A2(net1962),
    .A1(data_rdata_i_28_));
 sg13g2_nand2b_1 _17968_ (.Y(_01019_),
    .B(net1949),
    .A_N(_01018_));
 sg13g2_o21ai_1 _17969_ (.B1(_01019_),
    .Y(_01020_),
    .A1(net1704),
    .A2(_01017_));
 sg13g2_mux2_1 _17970_ (.A0(_01020_),
    .A1(data_rdata_i_4_),
    .S(net413),
    .X(_01021_));
 sg13g2_o21ai_1 _17971_ (.B1(net1648),
    .Y(_01022_),
    .A1(_01016_),
    .A2(_01021_));
 sg13g2_o21ai_1 _17972_ (.B1(_01022_),
    .Y(rf_wdata_wb_4_),
    .A1(net1074),
    .A2(_01013_));
 sg13g2_and2_1 _17973_ (.A(\load_store_unit_i.rdata_q_5_ ),
    .B(net1954),
    .X(_01023_));
 sg13g2_a221oi_1 _17974_ (.B2(\load_store_unit_i.rdata_q_21_ ),
    .C1(_01023_),
    .B1(net1949),
    .A1(\load_store_unit_i.rdata_q_13_ ),
    .Y(_01024_),
    .A2(net1940));
 sg13g2_a22oi_1 _17975_ (.Y(_01025_),
    .B1(net1954),
    .B2(data_rdata_i_13_),
    .A2(net1940),
    .A1(data_rdata_i_21_));
 sg13g2_a22oi_1 _17976_ (.Y(_01026_),
    .B1(net1933),
    .B2(\load_store_unit_i.rdata_q_21_ ),
    .A2(net1962),
    .A1(data_rdata_i_29_));
 sg13g2_nand2b_1 _17977_ (.Y(_01027_),
    .B(net1949),
    .A_N(_01026_));
 sg13g2_o21ai_1 _17978_ (.B1(_01027_),
    .Y(_01028_),
    .A1(_08404_),
    .A2(_01025_));
 sg13g2_nand2b_1 _17979_ (.Y(_01029_),
    .B(net414),
    .A_N(data_rdata_i_5_));
 sg13g2_o21ai_1 _17980_ (.B1(_01029_),
    .Y(_01030_),
    .A1(net413),
    .A2(_01028_));
 sg13g2_o21ai_1 _17981_ (.B1(_01030_),
    .Y(_01031_),
    .A1(net1706),
    .A2(_01024_));
 sg13g2_nor2_1 _17982_ (.A(net201),
    .B(_00843_),
    .Y(_01032_));
 sg13g2_a21oi_1 _17983_ (.A1(net203),
    .A2(_00839_),
    .Y(_01033_),
    .B1(_01032_));
 sg13g2_a21oi_1 _17984_ (.A1(_02435_),
    .A2(net131),
    .Y(_01034_),
    .B1(net1404));
 sg13g2_nand3_1 _17985_ (.B(_02435_),
    .C(net1358),
    .A(net1404),
    .Y(_01035_));
 sg13g2_o21ai_1 _17986_ (.B1(_01035_),
    .Y(_01036_),
    .A1(_02435_),
    .A2(net1358));
 sg13g2_a21oi_1 _17987_ (.A1(net1424),
    .A2(_01036_),
    .Y(_01037_),
    .B1(net1418));
 sg13g2_nor2b_1 _17988_ (.A(_01034_),
    .B_N(_01037_),
    .Y(_01038_));
 sg13g2_a221oi_1 _17989_ (.B2(net1365),
    .C1(_01038_),
    .B1(_01033_),
    .A1(data_addr_o_5_),
    .Y(_01039_),
    .A2(net1316));
 sg13g2_mux2_1 _17990_ (.A0(\ex_block_i.alu_i.imd_val_q_i_37_ ),
    .A1(_04479_),
    .S(_04144_),
    .X(_01040_));
 sg13g2_a21oi_1 _17991_ (.A1(net360),
    .A2(_01040_),
    .Y(_01041_),
    .B1(net1680));
 sg13g2_o21ai_1 _17992_ (.B1(_01041_),
    .Y(_01042_),
    .A1(_08548_),
    .A2(_01039_));
 sg13g2_inv_1 _17993_ (.Y(_01043_),
    .A(csr_rdata_5_));
 sg13g2_a21oi_1 _17994_ (.A1(_01043_),
    .A2(net1678),
    .Y(_01044_),
    .B1(net1075));
 sg13g2_a22oi_1 _17995_ (.Y(_01045_),
    .B1(_01042_),
    .B2(_01044_),
    .A2(_01031_),
    .A1(net1650));
 sg13g2_inv_2 _17996_ (.Y(rf_wdata_wb_5_),
    .A(_01045_));
 sg13g2_nor2_1 _17997_ (.A(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .B(net341),
    .Y(_01046_));
 sg13g2_nor3_1 _17998_ (.A(net1577),
    .B(_04033_),
    .C(_04560_),
    .Y(_01047_));
 sg13g2_and2_1 _17999_ (.A(net199),
    .B(_00817_),
    .X(_01048_));
 sg13g2_a21oi_1 _18000_ (.A1(net209),
    .A2(_00816_),
    .Y(_01049_),
    .B1(_01048_));
 sg13g2_nand2_1 _18001_ (.Y(_01050_),
    .A(net1349),
    .B(net128));
 sg13g2_nand3_1 _18002_ (.B(_02388_),
    .C(net1355),
    .A(net1349),
    .Y(_01051_));
 sg13g2_o21ai_1 _18003_ (.B1(_01051_),
    .Y(_01052_),
    .A1(net1349),
    .A2(net1356));
 sg13g2_a221oi_1 _18004_ (.B2(net1424),
    .C1(net1418),
    .B1(_01052_),
    .A1(_02387_),
    .Y(_01053_),
    .A2(_01050_));
 sg13g2_a221oi_1 _18005_ (.B2(net1365),
    .C1(_01053_),
    .B1(_01049_),
    .A1(data_addr_o_6_),
    .Y(_01054_),
    .A2(net1316));
 sg13g2_o21ai_1 _18006_ (.B1(net374),
    .Y(_01055_),
    .A1(net1195),
    .A2(_01054_));
 sg13g2_inv_1 _18007_ (.Y(_01056_),
    .A(_01055_));
 sg13g2_nor4_2 _18008_ (.A(net1680),
    .B(_01046_),
    .C(_01047_),
    .Y(_01057_),
    .D(_01056_));
 sg13g2_a21oi_2 _18009_ (.B1(_01057_),
    .Y(_01058_),
    .A2(net1676),
    .A1(csr_rdata_6_));
 sg13g2_nand2_1 _18010_ (.Y(_01059_),
    .A(\load_store_unit_i.rdata_q_6_ ),
    .B(net1953));
 sg13g2_a22oi_1 _18011_ (.Y(_01060_),
    .B1(net1945),
    .B2(\load_store_unit_i.rdata_q_22_ ),
    .A2(net1937),
    .A1(\load_store_unit_i.rdata_q_14_ ));
 sg13g2_a21oi_1 _18012_ (.A1(_01059_),
    .A2(_01060_),
    .Y(_01061_),
    .B1(net1707));
 sg13g2_a22oi_1 _18013_ (.Y(_01062_),
    .B1(net1953),
    .B2(data_rdata_i_14_),
    .A2(net1937),
    .A1(data_rdata_i_22_));
 sg13g2_a22oi_1 _18014_ (.Y(_01063_),
    .B1(net1933),
    .B2(\load_store_unit_i.rdata_q_22_ ),
    .A2(net1962),
    .A1(data_rdata_i_30_));
 sg13g2_nand2b_1 _18015_ (.Y(_01064_),
    .B(net1945),
    .A_N(_01063_));
 sg13g2_o21ai_1 _18016_ (.B1(_01064_),
    .Y(_01065_),
    .A1(_08404_),
    .A2(_01062_));
 sg13g2_mux2_1 _18017_ (.A0(_01065_),
    .A1(data_rdata_i_6_),
    .S(net413),
    .X(_01066_));
 sg13g2_o21ai_1 _18018_ (.B1(net1648),
    .Y(_01067_),
    .A1(_01061_),
    .A2(_01066_));
 sg13g2_o21ai_1 _18019_ (.B1(_01067_),
    .Y(rf_wdata_wb_6_),
    .A1(net1073),
    .A2(_01058_));
 sg13g2_nor2b_1 _18020_ (.A(net415),
    .B_N(net1960),
    .Y(_01068_));
 sg13g2_a221oi_1 _18021_ (.B2(\load_store_unit_i.rdata_q_7_ ),
    .C1(net1931),
    .B1(net1951),
    .A1(\load_store_unit_i.rdata_q_15_ ),
    .Y(_01069_),
    .A2(net1936));
 sg13g2_a21oi_1 _18022_ (.A1(net1931),
    .A2(_08615_),
    .Y(_01070_),
    .B1(_01069_));
 sg13g2_a21oi_1 _18023_ (.A1(\load_store_unit_i.rdata_q_23_ ),
    .A2(net1947),
    .Y(_01071_),
    .B1(_01070_));
 sg13g2_a21oi_1 _18024_ (.A1(net1960),
    .A2(net1959),
    .Y(_01072_),
    .B1(_01071_));
 sg13g2_a221oi_1 _18025_ (.B2(_01068_),
    .C1(_01072_),
    .B1(_08617_),
    .A1(data_rdata_i_7_),
    .Y(_01073_),
    .A2(net417));
 sg13g2_nand2_1 _18026_ (.Y(_01074_),
    .A(csr_rdata_7_),
    .B(net1678));
 sg13g2_and2_1 _18027_ (.A(net199),
    .B(_00794_),
    .X(_01075_));
 sg13g2_a21oi_1 _18028_ (.A1(net209),
    .A2(_00793_),
    .Y(_01076_),
    .B1(_01075_));
 sg13g2_nand2_1 _18029_ (.Y(_01077_),
    .A(net148),
    .B(net128));
 sg13g2_nand2_1 _18030_ (.Y(_01078_),
    .A(_02166_),
    .B(net1355));
 sg13g2_o21ai_1 _18031_ (.B1(_01078_),
    .Y(_01079_),
    .A1(net148),
    .A2(net1355));
 sg13g2_a221oi_1 _18032_ (.B2(net1422),
    .C1(net1417),
    .B1(_01079_),
    .A1(_02164_),
    .Y(_01080_),
    .A2(_01077_));
 sg13g2_a221oi_1 _18033_ (.B2(net1365),
    .C1(_01080_),
    .B1(_01076_),
    .A1(data_addr_o_7_),
    .Y(_01081_),
    .A2(net1316));
 sg13g2_o21ai_1 _18034_ (.B1(net376),
    .Y(_01082_),
    .A1(net1194),
    .A2(_01081_));
 sg13g2_a22oi_1 _18035_ (.Y(_01083_),
    .B1(_08611_),
    .B2(_02204_),
    .A2(net1472),
    .A1(_04656_));
 sg13g2_nand3_1 _18036_ (.B(_01082_),
    .C(_01083_),
    .A(_01199_),
    .Y(_01084_));
 sg13g2_a21o_2 _18037_ (.A2(_01084_),
    .A1(_01074_),
    .B1(net1075),
    .X(_01085_));
 sg13g2_o21ai_1 _18038_ (.B1(_01085_),
    .Y(rf_wdata_wb_7_),
    .A1(net1646),
    .A2(_01073_));
 sg13g2_nand2b_1 _18039_ (.Y(_01086_),
    .B(net206),
    .A_N(_00766_));
 sg13g2_o21ai_1 _18040_ (.B1(_01086_),
    .Y(_01087_),
    .A1(net206),
    .A2(_00764_));
 sg13g2_nand2_1 _18041_ (.Y(_01088_),
    .A(net1279),
    .B(net128));
 sg13g2_nand2_1 _18042_ (.Y(_01089_),
    .A(_02167_),
    .B(net1355));
 sg13g2_o21ai_1 _18043_ (.B1(_01089_),
    .Y(_01090_),
    .A1(net1279),
    .A2(net1355));
 sg13g2_a221oi_1 _18044_ (.B2(net1422),
    .C1(net1416),
    .B1(_01090_),
    .A1(net1401),
    .Y(_01091_),
    .A2(_01088_));
 sg13g2_a221oi_1 _18045_ (.B2(net1368),
    .C1(_01091_),
    .B1(_01087_),
    .A1(data_addr_o_8_),
    .Y(_01092_),
    .A2(net1319));
 sg13g2_o21ai_1 _18046_ (.B1(net374),
    .Y(_01093_),
    .A1(net1195),
    .A2(_01092_));
 sg13g2_inv_1 _18047_ (.Y(_01094_),
    .A(_01093_));
 sg13g2_nor2_1 _18048_ (.A(_04756_),
    .B(_08639_),
    .Y(_01095_));
 sg13g2_nor2_1 _18049_ (.A(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .B(_08610_),
    .Y(_01096_));
 sg13g2_nor4_2 _18050_ (.A(net1679),
    .B(_01094_),
    .C(_01095_),
    .Y(_01097_),
    .D(_01096_));
 sg13g2_a21oi_2 _18051_ (.B1(_01097_),
    .Y(_01098_),
    .A2(net1678),
    .A1(csr_rdata_8_));
 sg13g2_a22oi_1 _18052_ (.Y(_01099_),
    .B1(net414),
    .B2(data_rdata_i_8_),
    .A2(net1946),
    .A1(data_rdata_i_0_));
 sg13g2_a22oi_1 _18053_ (.Y(_01100_),
    .B1(net1954),
    .B2(data_rdata_i_16_),
    .A2(net1938),
    .A1(data_rdata_i_24_));
 sg13g2_a21oi_1 _18054_ (.A1(_01099_),
    .A2(_01100_),
    .Y(_01101_),
    .B1(net1959));
 sg13g2_a221oi_1 _18055_ (.B2(\load_store_unit_i.rdata_q_8_ ),
    .C1(net1933),
    .B1(net1954),
    .A1(\load_store_unit_i.rdata_q_16_ ),
    .Y(_01102_),
    .A2(net1938));
 sg13g2_a21oi_1 _18056_ (.A1(net1933),
    .A2(_01100_),
    .Y(_01103_),
    .B1(_01102_));
 sg13g2_nor2_1 _18057_ (.A(net1962),
    .B(_01103_),
    .Y(_01104_));
 sg13g2_a21oi_1 _18058_ (.A1(_01099_),
    .A2(_01104_),
    .Y(_01105_),
    .B1(net1646));
 sg13g2_o21ai_1 _18059_ (.B1(_01105_),
    .Y(_01106_),
    .A1(net1602),
    .A2(_01101_));
 sg13g2_o21ai_1 _18060_ (.B1(_01106_),
    .Y(rf_wdata_wb_8_),
    .A1(net1072),
    .A2(_01098_));
 sg13g2_nor2_1 _18061_ (.A(net2115),
    .B(_08610_),
    .Y(_01107_));
 sg13g2_nor2_1 _18062_ (.A(_04901_),
    .B(_08639_),
    .Y(_01108_));
 sg13g2_nand2_1 _18063_ (.Y(_01109_),
    .A(net203),
    .B(_00741_));
 sg13g2_o21ai_1 _18064_ (.B1(_01109_),
    .Y(_01110_),
    .A1(net201),
    .A2(_00738_));
 sg13g2_nand2_1 _18065_ (.Y(_01111_),
    .A(net193),
    .B(net128));
 sg13g2_nand3_1 _18066_ (.B(_02194_),
    .C(net1353),
    .A(net193),
    .Y(_01112_));
 sg13g2_o21ai_1 _18067_ (.B1(_01112_),
    .Y(_01113_),
    .A1(net192),
    .A2(net1354));
 sg13g2_a221oi_1 _18068_ (.B2(net1421),
    .C1(net1416),
    .B1(_01113_),
    .A1(_02148_),
    .Y(_01114_),
    .A2(_01111_));
 sg13g2_a221oi_1 _18069_ (.B2(net1366),
    .C1(_01114_),
    .B1(_01110_),
    .A1(data_addr_o_9_),
    .Y(_01115_),
    .A2(net1317));
 sg13g2_o21ai_1 _18070_ (.B1(net374),
    .Y(_01116_),
    .A1(net1196),
    .A2(_01115_));
 sg13g2_inv_1 _18071_ (.Y(_01117_),
    .A(_01116_));
 sg13g2_nor4_2 _18072_ (.A(net1679),
    .B(_01107_),
    .C(_01108_),
    .Y(_01118_),
    .D(_01117_));
 sg13g2_a21oi_2 _18073_ (.B1(_01118_),
    .Y(_01119_),
    .A2(net1676),
    .A1(csr_rdata_9_));
 sg13g2_a22oi_1 _18074_ (.Y(_01120_),
    .B1(net414),
    .B2(data_rdata_i_9_),
    .A2(net1949),
    .A1(data_rdata_i_1_));
 sg13g2_a22oi_1 _18075_ (.Y(_01121_),
    .B1(net1956),
    .B2(data_rdata_i_17_),
    .A2(net1941),
    .A1(data_rdata_i_25_));
 sg13g2_a21oi_1 _18076_ (.A1(_01120_),
    .A2(_01121_),
    .Y(_01122_),
    .B1(net1959));
 sg13g2_a221oi_1 _18077_ (.B2(\load_store_unit_i.rdata_q_9_ ),
    .C1(net1934),
    .B1(net1957),
    .A1(\load_store_unit_i.rdata_q_17_ ),
    .Y(_01123_),
    .A2(net1940));
 sg13g2_a21oi_1 _18078_ (.A1(net1933),
    .A2(_01121_),
    .Y(_01124_),
    .B1(_01123_));
 sg13g2_nor2_1 _18079_ (.A(net1962),
    .B(_01124_),
    .Y(_01125_));
 sg13g2_a21oi_1 _18080_ (.A1(_01120_),
    .A2(_01125_),
    .Y(_01126_),
    .B1(net1646));
 sg13g2_o21ai_1 _18081_ (.B1(_01126_),
    .Y(_01127_),
    .A1(_08620_),
    .A2(_01122_));
 sg13g2_o21ai_1 _18082_ (.B1(_01127_),
    .Y(rf_wdata_wb_9_),
    .A1(net1072),
    .A2(_01119_));
 sg13g2_nand2_2 _18083_ (.Y(rf_we_wb),
    .A(net1647),
    .B(net1074));
 sg13g2_tielo _09591__7 (.L_LO(net7));
 sg13g2_dfrbp_2 \crash_dump_o[100]_reg  (.RESET_B(net2331),
    .D(_00000_),
    .Q(crash_dump_o_100_),
    .Q_N(_09094_),
    .CLK(clknet_leaf_251_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[101]_reg  (.RESET_B(net2333),
    .D(_00001_),
    .Q(crash_dump_o_101_),
    .Q_N(_09093_),
    .CLK(clknet_leaf_251_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[102]_reg  (.RESET_B(net2331),
    .D(_00002_),
    .Q(crash_dump_o_102_),
    .Q_N(_09092_),
    .CLK(clknet_leaf_251_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[103]_reg  (.RESET_B(net2331),
    .D(_00003_),
    .Q(crash_dump_o_103_),
    .Q_N(_09091_),
    .CLK(clknet_leaf_251_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[104]_reg  (.RESET_B(net2338),
    .D(_00004_),
    .Q(crash_dump_o_104_),
    .Q_N(_09090_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[105]_reg  (.RESET_B(net2332),
    .D(_00005_),
    .Q(crash_dump_o_105_),
    .Q_N(_09089_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[106]_reg  (.RESET_B(net2332),
    .D(_00006_),
    .Q(crash_dump_o_106_),
    .Q_N(_09088_),
    .CLK(clknet_leaf_250_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[107]_reg  (.RESET_B(net2322),
    .D(_00007_),
    .Q(crash_dump_o_107_),
    .Q_N(_09087_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[108]_reg  (.RESET_B(net2333),
    .D(_00008_),
    .Q(crash_dump_o_108_),
    .Q_N(_09086_),
    .CLK(clknet_leaf_252_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[109]_reg  (.RESET_B(net2332),
    .D(_00009_),
    .Q(crash_dump_o_109_),
    .Q_N(_09085_),
    .CLK(clknet_leaf_250_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[110]_reg  (.RESET_B(net2338),
    .D(_00010_),
    .Q(crash_dump_o_110_),
    .Q_N(_09084_),
    .CLK(clknet_leaf_250_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[111]_reg  (.RESET_B(net2320),
    .D(_00011_),
    .Q(crash_dump_o_111_),
    .Q_N(_09083_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[112]_reg  (.RESET_B(net2333),
    .D(_00012_),
    .Q(crash_dump_o_112_),
    .Q_N(_09082_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[113]_reg  (.RESET_B(net2333),
    .D(_00013_),
    .Q(crash_dump_o_113_),
    .Q_N(_09081_),
    .CLK(clknet_leaf_252_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[114]_reg  (.RESET_B(net2342),
    .D(_00014_),
    .Q(crash_dump_o_114_),
    .Q_N(_09080_),
    .CLK(clknet_leaf_250_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[115]_reg  (.RESET_B(net2333),
    .D(_00015_),
    .Q(crash_dump_o_115_),
    .Q_N(_09079_),
    .CLK(clknet_leaf_252_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[116]_reg  (.RESET_B(net2340),
    .D(_00016_),
    .Q(crash_dump_o_116_),
    .Q_N(_09078_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[117]_reg  (.RESET_B(net2324),
    .D(_00017_),
    .Q(crash_dump_o_117_),
    .Q_N(_09077_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[118]_reg  (.RESET_B(net2334),
    .D(_00018_),
    .Q(crash_dump_o_118_),
    .Q_N(_09076_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[119]_reg  (.RESET_B(net2334),
    .D(_00019_),
    .Q(crash_dump_o_119_),
    .Q_N(_09075_),
    .CLK(clknet_leaf_251_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[120]_reg  (.RESET_B(net2334),
    .D(_00020_),
    .Q(crash_dump_o_120_),
    .Q_N(_09074_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[121]_reg  (.RESET_B(net2341),
    .D(_00021_),
    .Q(crash_dump_o_121_),
    .Q_N(_09073_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[122]_reg  (.RESET_B(net2333),
    .D(_00022_),
    .Q(crash_dump_o_122_),
    .Q_N(_09072_),
    .CLK(clknet_leaf_252_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[123]_reg  (.RESET_B(net2341),
    .D(_00023_),
    .Q(crash_dump_o_123_),
    .Q_N(_09071_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[124]_reg  (.RESET_B(net2339),
    .D(_00024_),
    .Q(crash_dump_o_124_),
    .Q_N(_09070_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[125]_reg  (.RESET_B(net2341),
    .D(_00025_),
    .Q(crash_dump_o_125_),
    .Q_N(_09069_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[126]_reg  (.RESET_B(net2341),
    .D(_00026_),
    .Q(crash_dump_o_126_),
    .Q_N(_09068_),
    .CLK(clknet_leaf_241_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[127]_reg  (.RESET_B(net2340),
    .D(_00027_),
    .Q(crash_dump_o_127_),
    .Q_N(_09067_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[32]_reg  (.RESET_B(net2321),
    .D(_00028_),
    .Q(crash_dump_o_32_),
    .Q_N(_09066_),
    .CLK(clknet_leaf_226_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[33]_reg  (.RESET_B(net2321),
    .D(_00029_),
    .Q(crash_dump_o_33_),
    .Q_N(_09065_),
    .CLK(clknet_leaf_287_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[34]_reg  (.RESET_B(net2314),
    .D(_00030_),
    .Q(crash_dump_o_34_),
    .Q_N(_09064_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[35]_reg  (.RESET_B(net2313),
    .D(_00031_),
    .Q(crash_dump_o_35_),
    .Q_N(_09063_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[36]_reg  (.RESET_B(net2311),
    .D(_00032_),
    .Q(crash_dump_o_36_),
    .Q_N(_09062_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[37]_reg  (.RESET_B(net2313),
    .D(_00033_),
    .Q(crash_dump_o_37_),
    .Q_N(_09061_),
    .CLK(clknet_leaf_242_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[38]_reg  (.RESET_B(net2311),
    .D(_00034_),
    .Q(crash_dump_o_38_),
    .Q_N(_09060_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[39]_reg  (.RESET_B(net2313),
    .D(_00035_),
    .Q(crash_dump_o_39_),
    .Q_N(_09059_),
    .CLK(clknet_leaf_242_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[40]_reg  (.RESET_B(net2315),
    .D(_00036_),
    .Q(crash_dump_o_40_),
    .Q_N(_09058_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[41]_reg  (.RESET_B(net2315),
    .D(_00037_),
    .Q(crash_dump_o_41_),
    .Q_N(_09057_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[42]_reg  (.RESET_B(net2328),
    .D(_00038_),
    .Q(crash_dump_o_42_),
    .Q_N(_09056_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[43]_reg  (.RESET_B(net2315),
    .D(_00039_),
    .Q(crash_dump_o_43_),
    .Q_N(_09055_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[44]_reg  (.RESET_B(net2314),
    .D(_00040_),
    .Q(crash_dump_o_44_),
    .Q_N(_09054_),
    .CLK(clknet_leaf_243_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[45]_reg  (.RESET_B(net2314),
    .D(_00041_),
    .Q(crash_dump_o_45_),
    .Q_N(_09053_),
    .CLK(clknet_leaf_244_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[46]_reg  (.RESET_B(net2333),
    .D(_00042_),
    .Q(crash_dump_o_46_),
    .Q_N(_09052_),
    .CLK(clknet_leaf_242_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[47]_reg  (.RESET_B(net2314),
    .D(_00043_),
    .Q(crash_dump_o_47_),
    .Q_N(_09051_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[48]_reg  (.RESET_B(net2315),
    .D(_00044_),
    .Q(crash_dump_o_48_),
    .Q_N(_09050_),
    .CLK(clknet_leaf_237_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[49]_reg  (.RESET_B(net2327),
    .D(_00045_),
    .Q(crash_dump_o_49_),
    .Q_N(_09049_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[50]_reg  (.RESET_B(net2327),
    .D(_00046_),
    .Q(crash_dump_o_50_),
    .Q_N(_09048_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[51]_reg  (.RESET_B(net2327),
    .D(_00047_),
    .Q(crash_dump_o_51_),
    .Q_N(_09047_),
    .CLK(clknet_leaf_238_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[52]_reg  (.RESET_B(net2329),
    .D(_00048_),
    .Q(crash_dump_o_52_),
    .Q_N(_09046_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[53]_reg  (.RESET_B(net2329),
    .D(_00049_),
    .Q(crash_dump_o_53_),
    .Q_N(_09045_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[54]_reg  (.RESET_B(net2331),
    .D(_00050_),
    .Q(crash_dump_o_54_),
    .Q_N(_09044_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[55]_reg  (.RESET_B(net2329),
    .D(_00051_),
    .Q(crash_dump_o_55_),
    .Q_N(_09043_),
    .CLK(clknet_leaf_238_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[56]_reg  (.RESET_B(net2328),
    .D(_00052_),
    .Q(crash_dump_o_56_),
    .Q_N(_09042_),
    .CLK(clknet_leaf_238_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[57]_reg  (.RESET_B(net2328),
    .D(_00053_),
    .Q(crash_dump_o_57_),
    .Q_N(_09041_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[58]_reg  (.RESET_B(net2328),
    .D(_00054_),
    .Q(crash_dump_o_58_),
    .Q_N(_09040_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[59]_reg  (.RESET_B(net2329),
    .D(_00055_),
    .Q(crash_dump_o_59_),
    .Q_N(_09039_),
    .CLK(clknet_leaf_237_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[60]_reg  (.RESET_B(net2329),
    .D(_00056_),
    .Q(crash_dump_o_60_),
    .Q_N(_09038_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[61]_reg  (.RESET_B(net2332),
    .D(_00057_),
    .Q(crash_dump_o_61_),
    .Q_N(_09037_),
    .CLK(clknet_leaf_245_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[62]_reg  (.RESET_B(net2329),
    .D(_00058_),
    .Q(crash_dump_o_62_),
    .Q_N(_09036_),
    .CLK(clknet_leaf_238_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[63]_reg  (.RESET_B(net2331),
    .D(_00059_),
    .Q(crash_dump_o_63_),
    .Q_N(_09035_),
    .CLK(clknet_leaf_237_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[65]_reg  (.RESET_B(net2362),
    .D(_00060_),
    .Q(crash_dump_o_65_),
    .Q_N(_09034_),
    .CLK(clknet_leaf_56_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[66]_reg  (.RESET_B(net2346),
    .D(_00061_),
    .Q(crash_dump_o_66_),
    .Q_N(_09033_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[67]_reg  (.RESET_B(net2344),
    .D(_00062_),
    .Q(crash_dump_o_67_),
    .Q_N(_09032_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[68]_reg  (.RESET_B(net2345),
    .D(_00063_),
    .Q(crash_dump_o_68_),
    .Q_N(_09031_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[69]_reg  (.RESET_B(net2344),
    .D(_00064_),
    .Q(crash_dump_o_69_),
    .Q_N(_09030_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[70]_reg  (.RESET_B(net2345),
    .D(_00065_),
    .Q(crash_dump_o_70_),
    .Q_N(_09029_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[71]_reg  (.RESET_B(net2344),
    .D(_00066_),
    .Q(crash_dump_o_71_),
    .Q_N(_09028_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[72]_reg  (.RESET_B(net2344),
    .D(_00067_),
    .Q(crash_dump_o_72_),
    .Q_N(_09027_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[73]_reg  (.RESET_B(net2344),
    .D(_00068_),
    .Q(crash_dump_o_73_),
    .Q_N(_09026_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[74]_reg  (.RESET_B(net2345),
    .D(_00069_),
    .Q(crash_dump_o_74_),
    .Q_N(_09025_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[75]_reg  (.RESET_B(net2345),
    .D(_00070_),
    .Q(crash_dump_o_75_),
    .Q_N(_09024_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[76]_reg  (.RESET_B(net2345),
    .D(_00071_),
    .Q(crash_dump_o_76_),
    .Q_N(_09023_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[77]_reg  (.RESET_B(net2345),
    .D(_00072_),
    .Q(crash_dump_o_77_),
    .Q_N(_09022_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[78]_reg  (.RESET_B(net2345),
    .D(_00073_),
    .Q(crash_dump_o_78_),
    .Q_N(_09021_),
    .CLK(clknet_leaf_235_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[79]_reg  (.RESET_B(net2345),
    .D(_00074_),
    .Q(crash_dump_o_79_),
    .Q_N(_09020_),
    .CLK(clknet_leaf_235_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[80]_reg  (.RESET_B(net2342),
    .D(_00075_),
    .Q(crash_dump_o_80_),
    .Q_N(_09019_),
    .CLK(clknet_leaf_231_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[81]_reg  (.RESET_B(net2346),
    .D(_00076_),
    .Q(crash_dump_o_81_),
    .Q_N(_09018_),
    .CLK(clknet_leaf_233_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[82]_reg  (.RESET_B(net2346),
    .D(_00077_),
    .Q(crash_dump_o_82_),
    .Q_N(_09017_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[83]_reg  (.RESET_B(net2340),
    .D(_00078_),
    .Q(crash_dump_o_83_),
    .Q_N(_09016_),
    .CLK(clknet_leaf_237_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[84]_reg  (.RESET_B(net2340),
    .D(_00079_),
    .Q(crash_dump_o_84_),
    .Q_N(_09015_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[85]_reg  (.RESET_B(net2340),
    .D(_00080_),
    .Q(crash_dump_o_85_),
    .Q_N(_09014_),
    .CLK(clknet_leaf_236_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[86]_reg  (.RESET_B(net2341),
    .D(_00081_),
    .Q(crash_dump_o_86_),
    .Q_N(_09013_),
    .CLK(clknet_leaf_235_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[87]_reg  (.RESET_B(net2341),
    .D(_00082_),
    .Q(crash_dump_o_87_),
    .Q_N(_09012_),
    .CLK(clknet_leaf_235_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[88]_reg  (.RESET_B(net2341),
    .D(_00083_),
    .Q(crash_dump_o_88_),
    .Q_N(_09011_),
    .CLK(clknet_leaf_235_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[89]_reg  (.RESET_B(net2342),
    .D(_00084_),
    .Q(crash_dump_o_89_),
    .Q_N(_09010_),
    .CLK(clknet_leaf_236_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[90]_reg  (.RESET_B(net2343),
    .D(_00085_),
    .Q(crash_dump_o_90_),
    .Q_N(_09009_),
    .CLK(clknet_leaf_239_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[91]_reg  (.RESET_B(net2340),
    .D(_00086_),
    .Q(crash_dump_o_91_),
    .Q_N(_09008_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[92]_reg  (.RESET_B(net2341),
    .D(_00087_),
    .Q(crash_dump_o_92_),
    .Q_N(_09007_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[93]_reg  (.RESET_B(net2342),
    .D(_00088_),
    .Q(crash_dump_o_93_),
    .Q_N(_09006_),
    .CLK(clknet_leaf_236_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[94]_reg  (.RESET_B(net2340),
    .D(_00089_),
    .Q(crash_dump_o_94_),
    .Q_N(_09005_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[95]_reg  (.RESET_B(net2340),
    .D(_00090_),
    .Q(crash_dump_o_95_),
    .Q_N(_09004_),
    .CLK(clknet_leaf_234_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[96]_reg  (.RESET_B(net2343),
    .D(_00091_),
    .Q(crash_dump_o_96_),
    .Q_N(_09003_),
    .CLK(clknet_leaf_240_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[97]_reg  (.RESET_B(net2362),
    .D(_00092_),
    .Q(crash_dump_o_97_),
    .Q_N(\csr_mtval_1__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_MUX__Y_B ),
    .CLK(clknet_leaf_56_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[98]_reg  (.RESET_B(net2333),
    .D(_00093_),
    .Q(crash_dump_o_98_),
    .Q_N(_09002_),
    .CLK(clknet_leaf_242_clk_i));
 sg13g2_dfrbp_2 \crash_dump_o[99]_reg  (.RESET_B(net2334),
    .D(_00094_),
    .Q(crash_dump_o_99_),
    .Q_N(_09001_),
    .CLK(clknet_leaf_242_clk_i));
 sg13g2_or2_1 \cs_registers_i/_2923_  (.X(\cs_registers_i/_0472_ ),
    .B(net99),
    .A(net1276));
 sg13g2_buf_8 fanout658 (.A(\cs_registers_i/_0656_ ),
    .X(net658));
 sg13g2_buf_16 fanout657 (.X(net657),
    .A(net658));
 sg13g2_buf_16 fanout656 (.X(net656),
    .A(net657));
 sg13g2_nand2b_2 \cs_registers_i/_2927_  (.Y(\cs_registers_i/_0476_ ),
    .B(net1235),
    .A_N(net61));
 sg13g2_nor2_2 \cs_registers_i/_2928_  (.A(net1192),
    .B(\cs_registers_i/_0476_ ),
    .Y(\cs_registers_i/_0477_ ));
 sg13g2_buf_16 fanout655 (.X(net655),
    .A(net657));
 sg13g2_buf_16 fanout654 (.X(net654),
    .A(net658));
 sg13g2_buf_8 fanout653 (.A(\cs_registers_i/_1591_ ),
    .X(net653));
 sg13g2_nand2b_1 \cs_registers_i/_2932_  (.Y(\cs_registers_i/_0481_ ),
    .B(net1270),
    .A_N(net1267));
 sg13g2_buf_16 fanout652 (.X(net652),
    .A(net653));
 sg13g2_buf_16 fanout651 (.X(net651),
    .A(net652));
 sg13g2_nand2_1 \cs_registers_i/_2935_  (.Y(\cs_registers_i/_0484_ ),
    .A(net1273),
    .B(net144));
 sg13g2_nand3_1 \cs_registers_i/_2936_  (.B(csr_addr_8_),
    .C(csr_addr_10_),
    .A(csr_addr_9_),
    .Y(\cs_registers_i/_0485_ ));
 sg13g2_nor4_1 \cs_registers_i/_2937_  (.A(csr_addr_11_),
    .B(\cs_registers_i/_0481_ ),
    .C(\cs_registers_i/_0484_ ),
    .D(\cs_registers_i/_0485_ ),
    .Y(\cs_registers_i/_0486_ ));
 sg13g2_buf_16 fanout650 (.X(net650),
    .A(net653));
 sg13g2_buf_16 fanout649 (.X(net649),
    .A(net653));
 sg13g2_buf_8 fanout648 (.A(\cs_registers_i/_1591_ ),
    .X(net648));
 sg13g2_or3_2 \cs_registers_i/_2941_  (.A(net1271),
    .B(net1269),
    .C(net144),
    .X(\cs_registers_i/_0490_ ));
 sg13g2_buf_8 fanout647 (.A(net648),
    .X(net647));
 sg13g2_nor2b_1 \cs_registers_i/_2943_  (.A(net101),
    .B_N(net1238),
    .Y(\cs_registers_i/_0492_ ));
 sg13g2_nor4_1 \cs_registers_i/_2944_  (.A(csr_addr_4_),
    .B(net61),
    .C(\cs_registers_i/_0490_ ),
    .D(net1174),
    .Y(\cs_registers_i/_0493_ ));
 sg13g2_buf_16 fanout646 (.X(net646),
    .A(net648));
 sg13g2_buf_8 fanout645 (.A(\cs_registers_i/_1690_ ),
    .X(net645));
 sg13g2_buf_16 fanout644 (.X(net644),
    .A(net645));
 sg13g2_nand2b_1 \cs_registers_i/_2948_  (.Y(\cs_registers_i/_0497_ ),
    .B(net1267),
    .A_N(net1271));
 sg13g2_nor4_1 \cs_registers_i/_2949_  (.A(net1273),
    .B(net100),
    .C(net146),
    .D(\cs_registers_i/_0497_ ),
    .Y(\cs_registers_i/_0498_ ));
 sg13g2_buf_4 fanout643 (.X(net643),
    .A(\cs_registers_i/_1690_ ));
 sg13g2_nand2_2 \cs_registers_i/_2951_  (.Y(\cs_registers_i/_0500_ ),
    .A(csr_addr_9_),
    .B(csr_addr_8_));
 sg13g2_or2_1 \cs_registers_i/_2952_  (.X(\cs_registers_i/_0501_ ),
    .B(csr_addr_11_),
    .A(csr_addr_10_));
 sg13g2_nor3_1 \cs_registers_i/_2953_  (.A(net1276),
    .B(\cs_registers_i/_0500_ ),
    .C(\cs_registers_i/_0501_ ),
    .Y(\cs_registers_i/_0502_ ));
 sg13g2_o21ai_1 \cs_registers_i/_2954_  (.B1(\cs_registers_i/_0502_ ),
    .Y(\cs_registers_i/_0503_ ),
    .A1(\cs_registers_i/_0493_ ),
    .A2(\cs_registers_i/_0498_ ));
 sg13g2_inv_1 \cs_registers_i/_2955_  (.Y(\cs_registers_i/_0504_ ),
    .A(net1270));
 sg13g2_or2_2 \cs_registers_i/_2956_  (.X(\cs_registers_i/_0505_ ),
    .B(net144),
    .A(net1267));
 sg13g2_or4_2 \cs_registers_i/_2957_  (.A(net1276),
    .B(net101),
    .C(net61),
    .D(net1238),
    .X(\cs_registers_i/_0506_ ));
 sg13g2_nor4_1 \cs_registers_i/_2958_  (.A(net1273),
    .B(\cs_registers_i/_0504_ ),
    .C(\cs_registers_i/_0505_ ),
    .D(\cs_registers_i/_0506_ ),
    .Y(\cs_registers_i/_0507_ ));
 sg13g2_or4_2 \cs_registers_i/_2959_  (.A(net1273),
    .B(net1270),
    .C(net1267),
    .D(net144),
    .X(\cs_registers_i/_0508_ ));
 sg13g2_nor3_1 \cs_registers_i/_2960_  (.A(net1192),
    .B(\cs_registers_i/_0476_ ),
    .C(\cs_registers_i/_0508_ ),
    .Y(\cs_registers_i/_0509_ ));
 sg13g2_nor2_1 \cs_registers_i/_2961_  (.A(\cs_registers_i/_0500_ ),
    .B(\cs_registers_i/_0501_ ),
    .Y(\cs_registers_i/_0510_ ));
 sg13g2_o21ai_1 \cs_registers_i/_2962_  (.B1(net56),
    .Y(\cs_registers_i/_0511_ ),
    .A1(net1118),
    .A2(\cs_registers_i/_0509_ ));
 sg13g2_nor2_1 \cs_registers_i/_2963_  (.A(csr_addr_10_),
    .B(net1277),
    .Y(\cs_registers_i/_0512_ ));
 sg13g2_nor2b_1 \cs_registers_i/_2964_  (.A(net1274),
    .B_N(net1268),
    .Y(\cs_registers_i/_0513_ ));
 sg13g2_buf_8 fanout642 (.A(net643),
    .X(net642));
 sg13g2_nor2b_1 \cs_registers_i/_2966_  (.A(net1268),
    .B_N(net1274),
    .Y(\cs_registers_i/_0515_ ));
 sg13g2_and2_1 \cs_registers_i/_2967_  (.A(csr_addr_10_),
    .B(net1277),
    .X(\cs_registers_i/_0516_ ));
 sg13g2_a22oi_1 \cs_registers_i/_2968_  (.Y(\cs_registers_i/_0517_ ),
    .B1(\cs_registers_i/_0515_ ),
    .B2(\cs_registers_i/_0516_ ),
    .A2(\cs_registers_i/_0513_ ),
    .A1(\cs_registers_i/_0512_ ));
 sg13g2_nand2b_2 \cs_registers_i/_2969_  (.Y(\cs_registers_i/_0518_ ),
    .B(net101),
    .A_N(net1276));
 sg13g2_nor3_2 \cs_registers_i/_2970_  (.A(net61),
    .B(net1242),
    .C(\cs_registers_i/_0518_ ),
    .Y(\cs_registers_i/_0519_ ));
 sg13g2_nor3_1 \cs_registers_i/_2971_  (.A(net1271),
    .B(net145),
    .C(\cs_registers_i/_0500_ ),
    .Y(\cs_registers_i/_0520_ ));
 sg13g2_nand3b_1 \cs_registers_i/_2972_  (.B(net40),
    .C(\cs_registers_i/_0520_ ),
    .Y(\cs_registers_i/_0521_ ),
    .A_N(\cs_registers_i/_0517_ ));
 sg13g2_nand3_1 \cs_registers_i/_2973_  (.B(\cs_registers_i/_0511_ ),
    .C(\cs_registers_i/_0521_ ),
    .A(\cs_registers_i/_0503_ ),
    .Y(\cs_registers_i/_0522_ ));
 sg13g2_buf_8 fanout641 (.A(\cs_registers_i/_1703_ ),
    .X(net641));
 sg13g2_nor2_2 \cs_registers_i/_2975_  (.A(net1274),
    .B(net1275),
    .Y(\cs_registers_i/_0524_ ));
 sg13g2_nor2_1 \cs_registers_i/_2976_  (.A(net99),
    .B(net74),
    .Y(\cs_registers_i/_0525_ ));
 sg13g2_nand3_1 \cs_registers_i/_2977_  (.B(\cs_registers_i/_0524_ ),
    .C(\cs_registers_i/_0525_ ),
    .A(net1235),
    .Y(\cs_registers_i/_0526_ ));
 sg13g2_nand2b_1 \cs_registers_i/_2978_  (.Y(\cs_registers_i/_0527_ ),
    .B(net1277),
    .A_N(csr_addr_10_));
 sg13g2_nor3_1 \cs_registers_i/_2979_  (.A(net1271),
    .B(\cs_registers_i/_0500_ ),
    .C(\cs_registers_i/_0527_ ),
    .Y(\cs_registers_i/_0528_ ));
 sg13g2_nand2_2 \cs_registers_i/_2980_  (.Y(\cs_registers_i/_0529_ ),
    .A(net74),
    .B(net1238));
 sg13g2_nand3b_1 \cs_registers_i/_2981_  (.B(\cs_registers_i/_0524_ ),
    .C(\cs_registers_i/_0529_ ),
    .Y(\cs_registers_i/_0530_ ),
    .A_N(net100));
 sg13g2_nor4_1 \cs_registers_i/_2982_  (.A(\cs_registers_i/_0504_ ),
    .B(net145),
    .C(\cs_registers_i/_0500_ ),
    .D(\cs_registers_i/_0501_ ),
    .Y(\cs_registers_i/_0531_ ));
 sg13g2_a22oi_1 \cs_registers_i/_2983_  (.Y(\cs_registers_i/_0532_ ),
    .B1(\cs_registers_i/_0530_ ),
    .B2(\cs_registers_i/_0531_ ),
    .A2(\cs_registers_i/_0528_ ),
    .A1(\cs_registers_i/_0526_ ));
 sg13g2_nor3_1 \cs_registers_i/_2984_  (.A(net1277),
    .B(\cs_registers_i/_0481_ ),
    .C(\cs_registers_i/_0484_ ),
    .Y(\cs_registers_i/_0533_ ));
 sg13g2_inv_1 \cs_registers_i/_2985_  (.Y(\cs_registers_i/_0534_ ),
    .A(net1277));
 sg13g2_nand2b_2 \cs_registers_i/_2986_  (.Y(\cs_registers_i/_0535_ ),
    .B(net1274),
    .A_N(net1272));
 sg13g2_xnor2_1 \cs_registers_i/_2987_  (.Y(\cs_registers_i/_0536_ ),
    .A(net74),
    .B(net1231));
 sg13g2_nor4_1 \cs_registers_i/_2988_  (.A(\cs_registers_i/_0534_ ),
    .B(\cs_registers_i/_0505_ ),
    .C(\cs_registers_i/_0535_ ),
    .D(\cs_registers_i/_0536_ ),
    .Y(\cs_registers_i/_0537_ ));
 sg13g2_nor2_1 \cs_registers_i/_2989_  (.A(net1192),
    .B(\cs_registers_i/_0485_ ),
    .Y(\cs_registers_i/_0538_ ));
 sg13g2_o21ai_1 \cs_registers_i/_2990_  (.B1(\cs_registers_i/_0538_ ),
    .Y(\cs_registers_i/_0539_ ),
    .A1(\cs_registers_i/_0533_ ),
    .A2(\cs_registers_i/_0537_ ));
 sg13g2_o21ai_1 \cs_registers_i/_2991_  (.B1(\cs_registers_i/_0539_ ),
    .Y(\cs_registers_i/_0540_ ),
    .A1(net1267),
    .A2(\cs_registers_i/_0532_ ));
 sg13g2_and2_1 \cs_registers_i/_2992_  (.A(csr_addr_9_),
    .B(csr_addr_8_),
    .X(\cs_registers_i/_0541_ ));
 sg13g2_nand2_1 \cs_registers_i/_2993_  (.Y(\cs_registers_i/_0542_ ),
    .A(\cs_registers_i/_0541_ ),
    .B(\cs_registers_i/_0512_ ));
 sg13g2_nor2_1 \cs_registers_i/_2994_  (.A(\cs_registers_i/_0505_ ),
    .B(\cs_registers_i/_0535_ ),
    .Y(\cs_registers_i/_0543_ ));
 sg13g2_nor2_2 \cs_registers_i/_2995_  (.A(net1276),
    .B(net101),
    .Y(\cs_registers_i/_0544_ ));
 sg13g2_nor2_1 \cs_registers_i/_2996_  (.A(net61),
    .B(net1238),
    .Y(\cs_registers_i/_0545_ ));
 sg13g2_and2_1 \cs_registers_i/_2997_  (.A(\cs_registers_i/_0544_ ),
    .B(net1131),
    .X(\cs_registers_i/_0546_ ));
 sg13g2_buf_16 fanout640 (.X(net640),
    .A(net641));
 sg13g2_mux2_1 \cs_registers_i/_2999_  (.A0(net1276),
    .A1(\cs_registers_i/_0524_ ),
    .S(net99),
    .X(\cs_registers_i/_0548_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3000_  (.A(net1235),
    .B_N(net61),
    .Y(\cs_registers_i/_0549_ ));
 sg13g2_nor3_2 \cs_registers_i/_3001_  (.A(net1270),
    .B(net1267),
    .C(net146),
    .Y(\cs_registers_i/_0550_ ));
 sg13g2_and2_1 \cs_registers_i/_3002_  (.A(\cs_registers_i/_0549_ ),
    .B(net1191),
    .X(\cs_registers_i/_0551_ ));
 sg13g2_inv_1 \cs_registers_i/_3003_  (.Y(\cs_registers_i/_0552_ ),
    .A(net1274));
 sg13g2_nand3b_1 \cs_registers_i/_3004_  (.B(net146),
    .C(net1270),
    .Y(\cs_registers_i/_0553_ ),
    .A_N(net1267));
 sg13g2_a21oi_1 \cs_registers_i/_3005_  (.A1(\cs_registers_i/_0552_ ),
    .A2(net1192),
    .Y(\cs_registers_i/_0554_ ),
    .B1(\cs_registers_i/_0553_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3006_  (.B2(\cs_registers_i/_0551_ ),
    .C1(\cs_registers_i/_0554_ ),
    .B1(\cs_registers_i/_0548_ ),
    .A1(\cs_registers_i/_0543_ ),
    .Y(\cs_registers_i/_0555_ ),
    .A2(net1117));
 sg13g2_nor2_1 \cs_registers_i/_3007_  (.A(net1277),
    .B(\cs_registers_i/_0485_ ),
    .Y(\cs_registers_i/_0556_ ));
 sg13g2_or2_2 \cs_registers_i/_3008_  (.X(\cs_registers_i/_0557_ ),
    .B(net1272),
    .A(net1274));
 sg13g2_nand2_1 \cs_registers_i/_3009_  (.Y(\cs_registers_i/_0558_ ),
    .A(net1269),
    .B(net145));
 sg13g2_nor4_1 \cs_registers_i/_3010_  (.A(net1192),
    .B(\cs_registers_i/_0476_ ),
    .C(\cs_registers_i/_0557_ ),
    .D(\cs_registers_i/_0558_ ),
    .Y(\cs_registers_i/_0559_ ));
 sg13g2_nand4_1 \cs_registers_i/_3011_  (.B(csr_addr_8_),
    .C(csr_addr_10_),
    .A(csr_addr_9_),
    .Y(\cs_registers_i/_0560_ ),
    .D(net1277));
 sg13g2_nor3_2 \cs_registers_i/_3012_  (.A(\cs_registers_i/_0505_ ),
    .B(\cs_registers_i/_0535_ ),
    .C(\cs_registers_i/_0560_ ),
    .Y(\cs_registers_i/_0561_ ));
 sg13g2_inv_1 \cs_registers_i/_3013_  (.Y(\cs_registers_i/_0562_ ),
    .A(net1239));
 sg13g2_xnor2_1 \cs_registers_i/_3014_  (.Y(\cs_registers_i/_0563_ ),
    .A(net101),
    .B(net74));
 sg13g2_nor3_1 \cs_registers_i/_3015_  (.A(csr_addr_3_),
    .B(net53),
    .C(\cs_registers_i/_0563_ ),
    .Y(\cs_registers_i/_0564_ ));
 sg13g2_inv_1 \cs_registers_i/_3016_  (.Y(\cs_registers_i/_0565_ ),
    .A(csr_access));
 sg13g2_a221oi_1 \cs_registers_i/_3017_  (.B2(\cs_registers_i/_0564_ ),
    .C1(\cs_registers_i/_0565_ ),
    .B1(\cs_registers_i/_0561_ ),
    .A1(\cs_registers_i/_0556_ ),
    .Y(\cs_registers_i/_0566_ ),
    .A2(\cs_registers_i/_0559_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3018_  (.B1(\cs_registers_i/_0566_ ),
    .Y(\cs_registers_i/_0567_ ),
    .A1(net1172),
    .A2(\cs_registers_i/_0555_ ));
 sg13g2_nor3_2 \cs_registers_i/_3019_  (.A(\cs_registers_i/_0522_ ),
    .B(\cs_registers_i/_0540_ ),
    .C(\cs_registers_i/_0567_ ),
    .Y(\cs_registers_i/_0568_ ));
 sg13g2_buf_16 fanout639 (.X(net639),
    .A(net641));
 sg13g2_or2_1 \cs_registers_i/_3021_  (.X(\cs_registers_i/_0570_ ),
    .B(csr_op_0_),
    .A(csr_op_1_));
 sg13g2_nand2_2 \cs_registers_i/_3022_  (.Y(\cs_registers_i/_0571_ ),
    .A(csr_op_en),
    .B(\cs_registers_i/_0570_ ));
 sg13g2_nand3b_1 \cs_registers_i/_3023_  (.B(\cs_registers_i/_0544_ ),
    .C(net60),
    .Y(\cs_registers_i/_0572_ ),
    .A_N(debug_mode));
 sg13g2_nand2b_1 \cs_registers_i/_3024_  (.Y(\cs_registers_i/_0573_ ),
    .B(csr_addr_8_),
    .A_N(\id_stage_i.controller_i.priv_mode_i_0_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3025_  (.Y(\cs_registers_i/_0574_ ),
    .B(csr_addr_9_),
    .A_N(net2116));
 sg13g2_nor2b_1 \cs_registers_i/_3026_  (.A(csr_addr_9_),
    .B_N(net2116),
    .Y(\cs_registers_i/_0575_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3027_  (.A1(\cs_registers_i/_0573_ ),
    .A2(\cs_registers_i/_0574_ ),
    .Y(\cs_registers_i/_0576_ ),
    .B1(\cs_registers_i/_0575_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3028_  (.B2(\cs_registers_i/_0554_ ),
    .C1(\cs_registers_i/_0576_ ),
    .B1(net57),
    .A1(\cs_registers_i/_0570_ ),
    .Y(\cs_registers_i/_0577_ ),
    .A2(\cs_registers_i/_0516_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3029_  (.B1(\cs_registers_i/_0565_ ),
    .Y(\cs_registers_i/_0578_ ),
    .A2(\cs_registers_i/_0577_ ),
    .A1(\cs_registers_i/_0572_ ));
 sg13g2_nor2_2 \cs_registers_i/_3030_  (.A(\cs_registers_i/_0571_ ),
    .B(\cs_registers_i/_0578_ ),
    .Y(\cs_registers_i/_0579_ ));
 sg13g2_nor2b_2 \cs_registers_i/_3031_  (.A(\cs_registers_i/_0568_ ),
    .B_N(\cs_registers_i/_0579_ ),
    .Y(\cs_registers_i/_0580_ ));
 sg13g2_and2_2 \cs_registers_i/_3032_  (.A(net60),
    .B(net722),
    .X(\cs_registers_i/_0581_ ));
 sg13g2_buf_8 fanout638 (.A(\cs_registers_i/_1703_ ),
    .X(net638));
 sg13g2_and2_1 \cs_registers_i/_3034_  (.A(net255),
    .B(debug_csr_save),
    .X(\cs_registers_i/_0583_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3035_  (.B1(net1313),
    .Y(\cs_registers_i/_0584_ ),
    .A2(\cs_registers_i/_0581_ ),
    .A1(\cs_registers_i/_0477_ ));
 sg13g2_buf_16 fanout637 (.X(net637),
    .A(net638));
 sg13g2_buf_8 fanout636 (.A(\cs_registers_i/_1707_ ),
    .X(net636));
 sg13g2_buf_16 fanout635 (.X(net635),
    .A(net636));
 sg13g2_mux2_2 \cs_registers_i/_3039_  (.A0(crash_dump_o_96_),
    .A1(net6),
    .S(net1483),
    .X(\cs_registers_i/_0588_ ));
 sg13g2_buf_16 fanout634 (.X(net634),
    .A(net635));
 sg13g2_a22oi_1 \cs_registers_i/_3041_  (.Y(\cs_registers_i/_0590_ ),
    .B1(\cs_registers_i/_0588_ ),
    .B2(net1308),
    .A2(net664),
    .A1(csr_depc_0_));
 sg13g2_inv_1 \cs_registers_i/_3042_  (.Y(\cs_registers_i/_0010_ ),
    .A(\cs_registers_i/_0590_ ));
 sg13g2_buf_16 fanout633 (.X(net633),
    .A(net634));
 sg13g2_nand2_1 \cs_registers_i/_3044_  (.Y(\cs_registers_i/_0592_ ),
    .A(csr_depc_10_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3045_  (.A0(crash_dump_o_106_),
    .A1(crash_dump_o_74_),
    .S(net1480),
    .X(\cs_registers_i/_0593_ ));
 sg13g2_nand2_1 \cs_registers_i/_3046_  (.Y(\cs_registers_i/_0594_ ),
    .A(csr_op_1_),
    .B(csr_op_0_));
 sg13g2_buf_16 fanout632 (.X(net632),
    .A(net636));
 sg13g2_o21ai_1 \cs_registers_i/_3048_  (.B1(csr_op_1_),
    .Y(\cs_registers_i/_0596_ ),
    .A1(\cs_registers_i/_0522_ ),
    .A2(\cs_registers_i/_0540_ ));
 sg13g2_buf_16 fanout631 (.X(net631),
    .A(net636));
 sg13g2_nor2_2 \cs_registers_i/_3050_  (.A(\cs_registers_i/_0476_ ),
    .B(\cs_registers_i/_0518_ ),
    .Y(\cs_registers_i/_0598_ ));
 sg13g2_nor3_2 \cs_registers_i/_3051_  (.A(\cs_registers_i/_0500_ ),
    .B(\cs_registers_i/_0501_ ),
    .C(\cs_registers_i/_0508_ ),
    .Y(\cs_registers_i/_0599_ ));
 sg13g2_and2_2 \cs_registers_i/_3052_  (.A(\cs_registers_i/_0598_ ),
    .B(\cs_registers_i/_0599_ ),
    .X(\cs_registers_i/_0600_ ));
 sg13g2_or2_2 \cs_registers_i/_3053_  (.X(\cs_registers_i/_0601_ ),
    .B(net1275),
    .A(net1274));
 sg13g2_buf_8 fanout630 (.A(\cs_registers_i/_1825_ ),
    .X(net630));
 sg13g2_nand2b_2 \cs_registers_i/_3055_  (.Y(\cs_registers_i/_0603_ ),
    .B(net1267),
    .A_N(net144));
 sg13g2_nor4_1 \cs_registers_i/_3056_  (.A(net100),
    .B(net1270),
    .C(\cs_registers_i/_0601_ ),
    .D(\cs_registers_i/_0603_ ),
    .Y(\cs_registers_i/_0604_ ));
 sg13g2_and2_2 \cs_registers_i/_3057_  (.A(net56),
    .B(net1160),
    .X(\cs_registers_i/_0605_ ));
 sg13g2_buf_16 fanout629 (.X(net629),
    .A(net630));
 sg13g2_buf_16 fanout628 (.X(net628),
    .A(net629));
 sg13g2_buf_16 fanout627 (.X(net627),
    .A(net629));
 sg13g2_buf_16 fanout626 (.X(net626),
    .A(net630));
 sg13g2_buf_2 fanout625 (.A(\cs_registers_i/_2188_ ),
    .X(net625));
 sg13g2_buf_2 fanout624 (.A(\cs_registers_i/_2330_ ),
    .X(net624));
 sg13g2_and2_1 \cs_registers_i/_3064_  (.A(crash_dump_o_10_),
    .B(net1234),
    .X(\cs_registers_i/_0612_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3065_  (.A1(net54),
    .A2(\cs_registers_i/mscratch_q_10_ ),
    .Y(\cs_registers_i/_0613_ ),
    .B1(\cs_registers_i/_0612_ ));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_16 fanout621 (.X(net621),
    .A(net623));
 sg13g2_buf_8 fanout620 (.A(\cs_registers_i/_2333_ ),
    .X(net620));
 sg13g2_buf_16 fanout619 (.X(net619),
    .A(net620));
 sg13g2_nand3_1 \cs_registers_i/_3071_  (.B(net1233),
    .C(\cs_registers_i/mtval_q_10_ ),
    .A(net76),
    .Y(\cs_registers_i/_0619_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3072_  (.B1(\cs_registers_i/_0619_ ),
    .Y(\cs_registers_i/_0620_ ),
    .A1(net64),
    .A2(\cs_registers_i/_0613_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3073_  (.Y(\cs_registers_i/_0621_ ),
    .B1(\cs_registers_i/_0605_ ),
    .B2(\cs_registers_i/_0620_ ),
    .A2(\cs_registers_i/_0600_ ),
    .A1(csr_mtvec_10_));
 sg13g2_buf_16 fanout618 (.X(net618),
    .A(net619));
 sg13g2_buf_16 fanout617 (.X(net617),
    .A(net620));
 sg13g2_mux2_1 \cs_registers_i/_3076_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .A1(\cs_registers_i/mhpmcounter_1866_ ),
    .S(net68),
    .X(\cs_registers_i/_0624_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3077_  (.A(csr_addr_10_),
    .B_N(net1277),
    .Y(\cs_registers_i/_0625_ ));
 sg13g2_nor2_2 \cs_registers_i/_3078_  (.A(net99),
    .B(net1235),
    .Y(\cs_registers_i/_0626_ ));
 sg13g2_nand4_1 \cs_registers_i/_3079_  (.B(\cs_registers_i/_0524_ ),
    .C(\cs_registers_i/_0625_ ),
    .A(\cs_registers_i/_0541_ ),
    .Y(\cs_registers_i/_0627_ ),
    .D(\cs_registers_i/_0626_ ));
 sg13g2_nor2_2 \cs_registers_i/_3080_  (.A(\cs_registers_i/_0490_ ),
    .B(net1158),
    .Y(\cs_registers_i/_0628_ ));
 sg13g2_nor2_1 \cs_registers_i/_3081_  (.A(net1272),
    .B(net1268),
    .Y(\cs_registers_i/_0629_ ));
 sg13g2_and2_1 \cs_registers_i/_3082_  (.A(net144),
    .B(\cs_registers_i/_0629_ ),
    .X(\cs_registers_i/_0630_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3083_  (.A(net1158),
    .B_N(net1156),
    .Y(\cs_registers_i/_0631_ ));
 sg13g2_buf_16 fanout616 (.X(net616),
    .A(net620));
 sg13g2_buf_8 fanout615 (.A(\cs_registers_i/_2361_ ),
    .X(net615));
 sg13g2_mux2_1 \cs_registers_i/_3086_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_42_ ),
    .A1(\cs_registers_i/mhpmcounter_1898_ ),
    .S(net69),
    .X(\cs_registers_i/_0634_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3087_  (.Y(\cs_registers_i/_0635_ ),
    .B1(net1130),
    .B2(\cs_registers_i/_0634_ ),
    .A2(\cs_registers_i/_0628_ ),
    .A1(\cs_registers_i/_0624_ ));
 sg13g2_nor2b_2 \cs_registers_i/_3088_  (.A(net1235),
    .B_N(net99),
    .Y(\cs_registers_i/_0636_ ));
 sg13g2_buf_16 fanout614 (.X(net614),
    .A(net615));
 sg13g2_buf_16 fanout613 (.X(net613),
    .A(net614));
 sg13g2_a21oi_1 \cs_registers_i/_3091_  (.A1(hart_id_i_10_),
    .A2(net1155),
    .Y(\cs_registers_i/_0639_ ),
    .B1(net1174));
 sg13g2_or2_1 \cs_registers_i/_3092_  (.X(\cs_registers_i/_0640_ ),
    .B(net64),
    .A(net1275));
 sg13g2_buf_16 fanout612 (.X(net612),
    .A(net614));
 sg13g2_nor2_1 \cs_registers_i/_3094_  (.A(\cs_registers_i/_0639_ ),
    .B(net1100),
    .Y(\cs_registers_i/_0642_ ));
 sg13g2_buf_16 fanout611 (.X(net611),
    .A(net615));
 sg13g2_mux4_1 \cs_registers_i/_3096_  (.S0(net70),
    .A0(\cs_registers_i/dcsr_q_10_ ),
    .A1(\cs_registers_i/dscratch0_q_10_ ),
    .A2(csr_depc_10_),
    .A3(\cs_registers_i/dscratch1_q_10_ ),
    .S1(net1232),
    .X(\cs_registers_i/_0644_ ));
 sg13g2_and2_1 \cs_registers_i/_3097_  (.A(\cs_registers_i/_0544_ ),
    .B(net59),
    .X(\cs_registers_i/_0645_ ));
 sg13g2_buf_16 fanout610 (.X(net610),
    .A(net611));
 sg13g2_buf_16 fanout609 (.X(net609),
    .A(net615));
 sg13g2_or4_2 \cs_registers_i/_3100_  (.A(net1273),
    .B(\cs_registers_i/_0504_ ),
    .C(net1172),
    .D(\cs_registers_i/_0505_ ),
    .X(\cs_registers_i/_0648_ ));
 sg13g2_nor2_2 \cs_registers_i/_3101_  (.A(\cs_registers_i/_0506_ ),
    .B(\cs_registers_i/_0648_ ),
    .Y(\cs_registers_i/_0649_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3102_  (.B2(net1150),
    .C1(\cs_registers_i/_0649_ ),
    .B1(\cs_registers_i/_0644_ ),
    .A1(\cs_registers_i/_0561_ ),
    .Y(\cs_registers_i/_0650_ ),
    .A2(\cs_registers_i/_0642_ ));
 sg13g2_and3_2 \cs_registers_i/_3103_  (.X(\cs_registers_i/_0651_ ),
    .A(\cs_registers_i/_0621_ ),
    .B(\cs_registers_i/_0635_ ),
    .C(\cs_registers_i/_0650_ ));
 sg13g2_nor3_1 \cs_registers_i/_3104_  (.A(net152),
    .B(net1089),
    .C(\cs_registers_i/_0651_ ),
    .Y(\cs_registers_i/_0652_ ));
 sg13g2_a21o_2 \cs_registers_i/_3105_  (.A2(net260),
    .A1(net151),
    .B1(\cs_registers_i/_0652_ ),
    .X(\cs_registers_i/_0653_ ));
 sg13g2_buf_16 fanout608 (.X(net608),
    .A(net609));
 sg13g2_nand2_2 \cs_registers_i/_3107_  (.Y(\cs_registers_i/_0655_ ),
    .A(net257),
    .B(debug_csr_save));
 sg13g2_and3_1 \cs_registers_i/_3108_  (.X(\cs_registers_i/_0656_ ),
    .A(\cs_registers_i/_0655_ ),
    .B(\cs_registers_i/_0477_ ),
    .C(\cs_registers_i/_0581_ ));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_16 fanout606 (.X(net606),
    .A(net608));
 sg13g2_a22oi_1 \cs_registers_i/_3111_  (.Y(\cs_registers_i/_0659_ ),
    .B1(\cs_registers_i/_0653_ ),
    .B2(net656),
    .A2(\cs_registers_i/_0593_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3112_  (.Y(\cs_registers_i/_0011_ ),
    .A(\cs_registers_i/_0592_ ),
    .B(\cs_registers_i/_0659_ ));
 sg13g2_nand2_1 \cs_registers_i/_3113_  (.Y(\cs_registers_i/_0660_ ),
    .A(csr_depc_11_),
    .B(net660));
 sg13g2_mux2_1 \cs_registers_i/_3114_  (.A0(crash_dump_o_107_),
    .A1(crash_dump_o_75_),
    .S(net1483),
    .X(\cs_registers_i/_0661_ ));
 sg13g2_buf_8 fanout605 (.A(net615),
    .X(net605));
 sg13g2_buf_16 fanout604 (.X(net604),
    .A(net615));
 sg13g2_and2_1 \cs_registers_i/_3117_  (.A(net100),
    .B(net1231),
    .X(\cs_registers_i/_0664_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3118_  (.Y(\cs_registers_i/_0665_ ),
    .B1(\cs_registers_i/_0664_ ),
    .B2(csr_mtvec_11_),
    .A2(\cs_registers_i/_0626_ ),
    .A1(\cs_registers_i/mstatus_q_2_ ));
 sg13g2_buf_2 fanout603 (.A(rf_wdata_wb_25_),
    .X(net603));
 sg13g2_nor4_2 \cs_registers_i/_3120_  (.A(net71),
    .B(net1270),
    .C(\cs_registers_i/_0601_ ),
    .Y(\cs_registers_i/_0667_ ),
    .D(\cs_registers_i/_0505_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3121_  (.Y(\cs_registers_i/_0668_ ),
    .B(\cs_registers_i/_0667_ ),
    .A_N(\cs_registers_i/_0665_ ));
 sg13g2_nor2b_2 \cs_registers_i/_3122_  (.A(net1272),
    .B_N(net1268),
    .Y(\cs_registers_i/_0669_ ));
 sg13g2_nor2b_2 \cs_registers_i/_3123_  (.A(net1268),
    .B_N(net1272),
    .Y(\cs_registers_i/_0670_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3124_  (.A1(\cs_registers_i/mscratch_q_11_ ),
    .A2(\cs_registers_i/_0669_ ),
    .Y(\cs_registers_i/_0671_ ),
    .B1(\cs_registers_i/_0670_ ));
 sg13g2_or2_1 \cs_registers_i/_3125_  (.X(\cs_registers_i/_0672_ ),
    .B(net64),
    .A(net100));
 sg13g2_nor4_2 \cs_registers_i/_3126_  (.A(net1236),
    .B(net145),
    .C(\cs_registers_i/_0601_ ),
    .Y(\cs_registers_i/_0673_ ),
    .D(\cs_registers_i/_0672_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3127_  (.Y(\cs_registers_i/_0674_ ),
    .B(\cs_registers_i/_0673_ ),
    .A_N(\cs_registers_i/_0671_ ));
 sg13g2_or4_2 \cs_registers_i/_3128_  (.A(net80),
    .B(net1270),
    .C(\cs_registers_i/_0601_ ),
    .D(\cs_registers_i/_0603_ ),
    .X(\cs_registers_i/_0675_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3129_  (.Y(\cs_registers_i/_0676_ ),
    .B1(net1155),
    .B2(irq_external_i),
    .A2(net1174),
    .A1(crash_dump_o_11_));
 sg13g2_or2_1 \cs_registers_i/_3130_  (.X(\cs_registers_i/_0677_ ),
    .B(\cs_registers_i/_0676_ ),
    .A(\cs_registers_i/_0675_ ));
 sg13g2_nor4_2 \cs_registers_i/_3131_  (.A(net1192),
    .B(\cs_registers_i/_0529_ ),
    .C(\cs_registers_i/_0557_ ),
    .Y(\cs_registers_i/_0678_ ),
    .D(\cs_registers_i/_0603_ ));
 sg13g2_nand2_1 \cs_registers_i/_3132_  (.Y(\cs_registers_i/_0679_ ),
    .A(\cs_registers_i/mtval_q_11_ ),
    .B(\cs_registers_i/_0678_ ));
 sg13g2_nand4_1 \cs_registers_i/_3133_  (.B(\cs_registers_i/_0674_ ),
    .C(\cs_registers_i/_0677_ ),
    .A(\cs_registers_i/_0668_ ),
    .Y(\cs_registers_i/_0680_ ),
    .D(\cs_registers_i/_0679_ ));
 sg13g2_buf_2 fanout602 (.A(rf_wdata_wb_25_),
    .X(net602));
 sg13g2_buf_2 fanout601 (.A(rf_wdata_wb_25_),
    .X(net601));
 sg13g2_mux4_1 \cs_registers_i/_3136_  (.S0(net68),
    .A0(\cs_registers_i/dcsr_q_11_ ),
    .A1(\cs_registers_i/dscratch0_q_11_ ),
    .A2(csr_depc_11_),
    .A3(\cs_registers_i/dscratch1_q_11_ ),
    .S1(net1243),
    .X(\cs_registers_i/_0683_ ));
 sg13g2_buf_1 fanout600 (.A(net601),
    .X(net600));
 sg13g2_mux2_1 \cs_registers_i/_3138_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_11_ ),
    .A1(\cs_registers_i/mhpmcounter_1867_ ),
    .S(net62),
    .X(\cs_registers_i/_0685_ ));
 sg13g2_nand2_1 \cs_registers_i/_3139_  (.Y(\cs_registers_i/_0686_ ),
    .A(\cs_registers_i/_0550_ ),
    .B(\cs_registers_i/_0685_ ));
 sg13g2_buf_2 fanout599 (.A(net600),
    .X(net599));
 sg13g2_mux2_1 \cs_registers_i/_3141_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ),
    .A1(\cs_registers_i/mhpmcounter_1899_ ),
    .S(net62),
    .X(\cs_registers_i/_0688_ ));
 sg13g2_nand3_1 \cs_registers_i/_3142_  (.B(\cs_registers_i/_0629_ ),
    .C(\cs_registers_i/_0688_ ),
    .A(net146),
    .Y(\cs_registers_i/_0689_ ));
 sg13g2_buf_8 fanout598 (.A(\cs_registers_i/_1412_ ),
    .X(net598));
 sg13g2_a21o_1 \cs_registers_i/_3144_  (.A2(\cs_registers_i/_0689_ ),
    .A1(\cs_registers_i/_0686_ ),
    .B1(net1159),
    .X(\cs_registers_i/_0691_ ));
 sg13g2_buf_16 fanout597 (.X(net597),
    .A(net598));
 sg13g2_nand3_1 \cs_registers_i/_3146_  (.B(net40),
    .C(\cs_registers_i/_0599_ ),
    .A(\cs_registers_i/mie_q_16_ ),
    .Y(\cs_registers_i/_0693_ ));
 sg13g2_nand3_1 \cs_registers_i/_3147_  (.B(net40),
    .C(\cs_registers_i/_0561_ ),
    .A(hart_id_i_11_),
    .Y(\cs_registers_i/_0694_ ));
 sg13g2_nand3_1 \cs_registers_i/_3148_  (.B(\cs_registers_i/_0693_ ),
    .C(\cs_registers_i/_0694_ ),
    .A(\cs_registers_i/_0691_ ),
    .Y(\cs_registers_i/_0695_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3149_  (.B2(net1152),
    .C1(\cs_registers_i/_0695_ ),
    .B1(\cs_registers_i/_0683_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0696_ ),
    .A2(\cs_registers_i/_0680_ ));
 sg13g2_nor3_1 \cs_registers_i/_3150_  (.A(net1415),
    .B(net1088),
    .C(\cs_registers_i/_0696_ ),
    .Y(\cs_registers_i/_0697_ ));
 sg13g2_a21o_2 \cs_registers_i/_3151_  (.A2(net261),
    .A1(net1414),
    .B1(\cs_registers_i/_0697_ ),
    .X(\cs_registers_i/_0698_ ));
 sg13g2_buf_16 fanout596 (.X(net596),
    .A(net597));
 sg13g2_a22oi_1 \cs_registers_i/_3153_  (.Y(\cs_registers_i/_0700_ ),
    .B1(net1070),
    .B2(net658),
    .A2(\cs_registers_i/_0661_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3154_  (.Y(\cs_registers_i/_0012_ ),
    .A(\cs_registers_i/_0660_ ),
    .B(\cs_registers_i/_0700_ ));
 sg13g2_nand2_1 \cs_registers_i/_3155_  (.Y(\cs_registers_i/_0701_ ),
    .A(csr_depc_12_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3156_  (.A0(crash_dump_o_108_),
    .A1(crash_dump_o_76_),
    .S(net1480),
    .X(\cs_registers_i/_0702_ ));
 sg13g2_buf_16 fanout595 (.X(net595),
    .A(net596));
 sg13g2_buf_16 fanout594 (.X(net594),
    .A(net598));
 sg13g2_buf_16 fanout593 (.X(net593),
    .A(net594));
 sg13g2_buf_16 fanout592 (.X(net592),
    .A(net593));
 sg13g2_and2_1 \cs_registers_i/_3161_  (.A(crash_dump_o_12_),
    .B(net1240),
    .X(\cs_registers_i/_0707_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3162_  (.A1(net55),
    .A2(\cs_registers_i/mscratch_q_12_ ),
    .Y(\cs_registers_i/_0708_ ),
    .B1(\cs_registers_i/_0707_ ));
 sg13g2_nand3_1 \cs_registers_i/_3163_  (.B(net1238),
    .C(\cs_registers_i/mtval_q_12_ ),
    .A(net75),
    .Y(\cs_registers_i/_0709_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3164_  (.B1(\cs_registers_i/_0709_ ),
    .Y(\cs_registers_i/_0710_ ),
    .A1(net73),
    .A2(\cs_registers_i/_0708_ ));
 sg13g2_inv_1 \cs_registers_i/_3165_  (.Y(\cs_registers_i/_0711_ ),
    .A(net1174));
 sg13g2_o21ai_1 \cs_registers_i/_3166_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_44_ ),
    .Y(\cs_registers_i/_0712_ ),
    .A1(\cs_registers_i/_0601_ ),
    .A2(\cs_registers_i/_0711_ ));
 sg13g2_nand2_1 \cs_registers_i/_3167_  (.Y(\cs_registers_i/_0713_ ),
    .A(net77),
    .B(\cs_registers_i/mhpmcounter_1900_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3168_  (.B1(\cs_registers_i/_0713_ ),
    .Y(\cs_registers_i/_0714_ ),
    .A1(net73),
    .A2(\cs_registers_i/_0712_ ));
 sg13g2_and2_1 \cs_registers_i/_3169_  (.A(net40),
    .B(\cs_registers_i/_0561_ ),
    .X(\cs_registers_i/_0715_ ));
 sg13g2_buf_16 fanout591 (.X(net591),
    .A(net598));
 sg13g2_nor2b_2 \cs_registers_i/_3171_  (.A(net74),
    .B_N(net1238),
    .Y(\cs_registers_i/_0717_ ));
 sg13g2_nand2_1 \cs_registers_i/_3172_  (.Y(\cs_registers_i/_0718_ ),
    .A(net1275),
    .B(net99));
 sg13g2_or3_1 \cs_registers_i/_3173_  (.A(\cs_registers_i/_0490_ ),
    .B(net1131),
    .C(\cs_registers_i/_0718_ ),
    .X(\cs_registers_i/_0719_ ));
 sg13g2_nor4_2 \cs_registers_i/_3174_  (.A(net1274),
    .B(net1272),
    .C(net1268),
    .Y(\cs_registers_i/_0720_ ),
    .D(net147));
 sg13g2_o21ai_1 \cs_registers_i/_3175_  (.B1(\cs_registers_i/_0720_ ),
    .Y(\cs_registers_i/_0721_ ),
    .A1(net1131),
    .A2(\cs_registers_i/_0718_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3176_  (.B2(\cs_registers_i/_0721_ ),
    .C1(net1158),
    .B1(\cs_registers_i/_0719_ ),
    .A1(\cs_registers_i/_0544_ ),
    .Y(\cs_registers_i/_0722_ ),
    .A2(\cs_registers_i/_0717_ ));
 sg13g2_inv_1 \cs_registers_i/_3177_  (.Y(\cs_registers_i/_0723_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_12_ ));
 sg13g2_nand2_1 \cs_registers_i/_3178_  (.Y(\cs_registers_i/_0724_ ),
    .A(net76),
    .B(\cs_registers_i/mhpmcounter_1868_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3179_  (.B1(\cs_registers_i/_0724_ ),
    .Y(\cs_registers_i/_0725_ ),
    .A1(net66),
    .A2(\cs_registers_i/_0723_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3180_  (.Y(\cs_registers_i/_0726_ ),
    .B1(\cs_registers_i/_0722_ ),
    .B2(\cs_registers_i/_0725_ ),
    .A2(net1098),
    .A1(hart_id_i_12_));
 sg13g2_buf_16 fanout590 (.X(net590),
    .A(net591));
 sg13g2_mux4_1 \cs_registers_i/_3182_  (.S0(net67),
    .A0(debug_ebreaku),
    .A1(\cs_registers_i/dscratch0_q_12_ ),
    .A2(csr_depc_12_),
    .A3(\cs_registers_i/dscratch1_q_12_ ),
    .S1(net1240),
    .X(\cs_registers_i/_0728_ ));
 sg13g2_buf_16 fanout589 (.X(net589),
    .A(net590));
 sg13g2_nor2_1 \cs_registers_i/_3184_  (.A(net1231),
    .B(\cs_registers_i/mstatus_q_3_ ),
    .Y(\cs_registers_i/_0730_ ));
 sg13g2_nand2_1 \cs_registers_i/_3185_  (.Y(\cs_registers_i/_0731_ ),
    .A(csr_mtvec_12_),
    .B(net1234));
 sg13g2_o21ai_1 \cs_registers_i/_3186_  (.B1(\cs_registers_i/_0731_ ),
    .Y(\cs_registers_i/_0732_ ),
    .A1(net101),
    .A2(\cs_registers_i/_0730_ ));
 sg13g2_a21o_1 \cs_registers_i/_3187_  (.A2(\cs_registers_i/_0732_ ),
    .A1(\cs_registers_i/_0667_ ),
    .B1(net1118),
    .X(\cs_registers_i/_0733_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3188_  (.Y(\cs_registers_i/_0734_ ),
    .B1(\cs_registers_i/_0733_ ),
    .B2(net58),
    .A2(\cs_registers_i/_0728_ ),
    .A1(net1150));
 sg13g2_nand2_1 \cs_registers_i/_3189_  (.Y(\cs_registers_i/_0735_ ),
    .A(\cs_registers_i/_0726_ ),
    .B(\cs_registers_i/_0734_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3190_  (.B2(net1130),
    .C1(\cs_registers_i/_0735_ ),
    .B1(\cs_registers_i/_0714_ ),
    .A1(\cs_registers_i/_0605_ ),
    .Y(\cs_registers_i/_0736_ ),
    .A2(\cs_registers_i/_0710_ ));
 sg13g2_nor3_1 \cs_registers_i/_3191_  (.A(net1412),
    .B(net1090),
    .C(\cs_registers_i/_0736_ ),
    .Y(\cs_registers_i/_0737_ ));
 sg13g2_a21o_2 \cs_registers_i/_3192_  (.A2(net261),
    .A1(net1412),
    .B1(\cs_registers_i/_0737_ ),
    .X(\cs_registers_i/_0738_ ));
 sg13g2_buf_16 fanout588 (.X(net588),
    .A(net590));
 sg13g2_a22oi_1 \cs_registers_i/_3194_  (.Y(\cs_registers_i/_0740_ ),
    .B1(net1029),
    .B2(net656),
    .A2(\cs_registers_i/_0702_ ),
    .A1(net1313));
 sg13g2_nand2_1 \cs_registers_i/_3195_  (.Y(\cs_registers_i/_0013_ ),
    .A(\cs_registers_i/_0701_ ),
    .B(\cs_registers_i/_0740_ ));
 sg13g2_nand2_1 \cs_registers_i/_3196_  (.Y(\cs_registers_i/_0741_ ),
    .A(csr_depc_13_),
    .B(net659));
 sg13g2_mux2_2 \cs_registers_i/_3197_  (.A0(crash_dump_o_109_),
    .A1(crash_dump_o_77_),
    .S(net1480),
    .X(\cs_registers_i/_0742_ ));
 sg13g2_buf_2 fanout587 (.A(\cs_registers_i/_1727_ ),
    .X(net587));
 sg13g2_buf_4 fanout586 (.X(net586),
    .A(\cs_registers_i/_1727_ ));
 sg13g2_buf_2 fanout585 (.A(rf_wdata_wb_27_),
    .X(net585));
 sg13g2_buf_2 fanout584 (.A(rf_wdata_wb_27_),
    .X(net584));
 sg13g2_mux2_1 \cs_registers_i/_3202_  (.A0(crash_dump_o_13_),
    .A1(\cs_registers_i/mtval_q_13_ ),
    .S(net65),
    .X(\cs_registers_i/_0747_ ));
 sg13g2_nand3_1 \cs_registers_i/_3203_  (.B(net1161),
    .C(\cs_registers_i/_0747_ ),
    .A(net1234),
    .Y(\cs_registers_i/_0748_ ));
 sg13g2_nor3_2 \cs_registers_i/_3204_  (.A(\cs_registers_i/_0476_ ),
    .B(\cs_registers_i/_0508_ ),
    .C(\cs_registers_i/_0518_ ),
    .Y(\cs_registers_i/_0749_ ));
 sg13g2_nand2_1 \cs_registers_i/_3205_  (.Y(\cs_registers_i/_0750_ ),
    .A(csr_mtvec_13_),
    .B(\cs_registers_i/_0749_ ));
 sg13g2_nand2_1 \cs_registers_i/_3206_  (.Y(\cs_registers_i/_0751_ ),
    .A(\cs_registers_i/_0748_ ),
    .B(\cs_registers_i/_0750_ ));
 sg13g2_mux4_1 \cs_registers_i/_3207_  (.S0(net69),
    .A0(\cs_registers_i/dcsr_q_13_ ),
    .A1(\cs_registers_i/dscratch0_q_13_ ),
    .A2(csr_depc_13_),
    .A3(\cs_registers_i/dscratch1_q_13_ ),
    .S1(net1237),
    .X(\cs_registers_i/_0752_ ));
 sg13g2_buf_2 fanout583 (.A(rf_wdata_wb_27_),
    .X(net583));
 sg13g2_mux2_1 \cs_registers_i/_3209_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_13_ ),
    .A1(\cs_registers_i/mhpmcounter_1869_ ),
    .S(net70),
    .X(\cs_registers_i/_0754_ ));
 sg13g2_mux2_1 \cs_registers_i/_3210_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_45_ ),
    .A1(\cs_registers_i/mhpmcounter_1901_ ),
    .S(net70),
    .X(\cs_registers_i/_0755_ ));
 sg13g2_buf_1 fanout582 (.A(net583),
    .X(net582));
 sg13g2_a22oi_1 \cs_registers_i/_3212_  (.Y(\cs_registers_i/_0757_ ),
    .B1(\cs_registers_i/_0755_ ),
    .B2(net1157),
    .A2(\cs_registers_i/_0754_ ),
    .A1(\cs_registers_i/_0550_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3213_  (.A1(\cs_registers_i/mscratch_q_13_ ),
    .A2(\cs_registers_i/_0669_ ),
    .Y(\cs_registers_i/_0758_ ),
    .B1(\cs_registers_i/_0670_ ));
 sg13g2_nor2_1 \cs_registers_i/_3214_  (.A(net1172),
    .B(\cs_registers_i/_0758_ ),
    .Y(\cs_registers_i/_0759_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3215_  (.Y(\cs_registers_i/_0760_ ),
    .B1(\cs_registers_i/_0759_ ),
    .B2(\cs_registers_i/_0673_ ),
    .A2(net1096),
    .A1(hart_id_i_13_));
 sg13g2_o21ai_1 \cs_registers_i/_3216_  (.B1(\cs_registers_i/_0760_ ),
    .Y(\cs_registers_i/_0761_ ),
    .A1(net1158),
    .A2(\cs_registers_i/_0757_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3217_  (.B2(net1151),
    .C1(\cs_registers_i/_0761_ ),
    .B1(\cs_registers_i/_0752_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0762_ ),
    .A2(\cs_registers_i/_0751_ ));
 sg13g2_nor3_1 \cs_registers_i/_3218_  (.A(alu_operand_a_ex_13_),
    .B(net1089),
    .C(\cs_registers_i/_0762_ ),
    .Y(\cs_registers_i/_0763_ ));
 sg13g2_a21o_2 \cs_registers_i/_3219_  (.A2(net262),
    .A1(alu_operand_a_ex_13_),
    .B1(\cs_registers_i/_0763_ ),
    .X(\cs_registers_i/_0764_ ));
 sg13g2_buf_2 fanout581 (.A(net583),
    .X(net581));
 sg13g2_a22oi_1 \cs_registers_i/_3221_  (.Y(\cs_registers_i/_0766_ ),
    .B1(net1057),
    .B2(net654),
    .A2(\cs_registers_i/_0742_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3222_  (.Y(\cs_registers_i/_0014_ ),
    .A(\cs_registers_i/_0741_ ),
    .B(\cs_registers_i/_0766_ ));
 sg13g2_nand2_1 \cs_registers_i/_3223_  (.Y(\cs_registers_i/_0767_ ),
    .A(csr_depc_14_),
    .B(net659));
 sg13g2_mux2_1 \cs_registers_i/_3224_  (.A0(crash_dump_o_110_),
    .A1(crash_dump_o_78_),
    .S(net1483),
    .X(\cs_registers_i/_0768_ ));
 sg13g2_buf_2 fanout580 (.A(rf_wdata_wb_28_),
    .X(net580));
 sg13g2_and2_1 \cs_registers_i/_3226_  (.A(net61),
    .B(net1238),
    .X(\cs_registers_i/_0770_ ));
 sg13g2_buf_2 fanout579 (.A(net580),
    .X(net579));
 sg13g2_mux2_1 \cs_registers_i/_3228_  (.A0(\cs_registers_i/mscratch_q_14_ ),
    .A1(crash_dump_o_14_),
    .S(net1231),
    .X(\cs_registers_i/_0772_ ));
 sg13g2_inv_1 \cs_registers_i/_3229_  (.Y(\cs_registers_i/_0773_ ),
    .A(net61));
 sg13g2_buf_2 fanout578 (.A(rf_wdata_wb_28_),
    .X(net578));
 sg13g2_a22oi_1 \cs_registers_i/_3231_  (.Y(\cs_registers_i/_0775_ ),
    .B1(\cs_registers_i/_0772_ ),
    .B2(net1114),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_14_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3232_  (.A(\cs_registers_i/_0775_ ),
    .B_N(net1160),
    .Y(\cs_registers_i/_0776_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3233_  (.B1(net56),
    .Y(\cs_registers_i/_0777_ ),
    .A1(net1119),
    .A2(\cs_registers_i/_0776_ ));
 sg13g2_buf_2 fanout577 (.A(rf_wdata_wb_28_),
    .X(net577));
 sg13g2_nand2_1 \cs_registers_i/_3235_  (.Y(\cs_registers_i/_0779_ ),
    .A(hart_id_i_14_),
    .B(net1098));
 sg13g2_mux2_2 \cs_registers_i/_3236_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .A1(\cs_registers_i/mhpmcounter_1902_ ),
    .S(net72),
    .X(\cs_registers_i/_0780_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3237_  (.Y(\cs_registers_i/_0781_ ),
    .B1(\cs_registers_i/_0780_ ),
    .B2(net1130),
    .A2(\cs_registers_i/_0600_ ),
    .A1(csr_mtvec_14_));
 sg13g2_mux4_1 \cs_registers_i/_3238_  (.S0(net67),
    .A0(\cs_registers_i/dcsr_q_14_ ),
    .A1(\cs_registers_i/dscratch0_q_14_ ),
    .A2(csr_depc_14_),
    .A3(\cs_registers_i/dscratch1_q_14_ ),
    .S1(net1237),
    .X(\cs_registers_i/_0782_ ));
 sg13g2_inv_1 \cs_registers_i/_3239_  (.Y(\cs_registers_i/_0783_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ));
 sg13g2_buf_4 fanout576 (.X(net576),
    .A(rf_wdata_wb_30_));
 sg13g2_nand2_1 \cs_registers_i/_3241_  (.Y(\cs_registers_i/_0785_ ),
    .A(net80),
    .B(\cs_registers_i/mhpmcounter_1870_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3242_  (.B1(\cs_registers_i/_0785_ ),
    .Y(\cs_registers_i/_0786_ ),
    .A1(net69),
    .A2(\cs_registers_i/_0783_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3243_  (.Y(\cs_registers_i/_0787_ ),
    .B1(\cs_registers_i/_0786_ ),
    .B2(\cs_registers_i/_0722_ ),
    .A2(\cs_registers_i/_0782_ ),
    .A1(net1152));
 sg13g2_and4_2 \cs_registers_i/_3244_  (.A(\cs_registers_i/_0777_ ),
    .B(\cs_registers_i/_0779_ ),
    .C(\cs_registers_i/_0781_ ),
    .D(\cs_registers_i/_0787_ ),
    .X(\cs_registers_i/_0788_ ));
 sg13g2_nor3_1 \cs_registers_i/_3245_  (.A(net1283),
    .B(net1088),
    .C(\cs_registers_i/_0788_ ),
    .Y(\cs_registers_i/_0789_ ));
 sg13g2_a21o_2 \cs_registers_i/_3246_  (.A2(net261),
    .A1(net1283),
    .B1(\cs_registers_i/_0789_ ),
    .X(\cs_registers_i/_0790_ ));
 sg13g2_buf_4 fanout575 (.X(net575),
    .A(net576));
 sg13g2_a22oi_1 \cs_registers_i/_3248_  (.Y(\cs_registers_i/_0792_ ),
    .B1(net1056),
    .B2(net654),
    .A2(\cs_registers_i/_0768_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3249_  (.Y(\cs_registers_i/_0015_ ),
    .A(\cs_registers_i/_0767_ ),
    .B(\cs_registers_i/_0792_ ));
 sg13g2_nand2_1 \cs_registers_i/_3250_  (.Y(\cs_registers_i/_0793_ ),
    .A(csr_depc_15_),
    .B(net659));
 sg13g2_mux2_1 \cs_registers_i/_3251_  (.A0(crash_dump_o_111_),
    .A1(crash_dump_o_79_),
    .S(net1483),
    .X(\cs_registers_i/_0794_ ));
 sg13g2_mux2_1 \cs_registers_i/_3252_  (.A0(\cs_registers_i/mscratch_q_15_ ),
    .A1(crash_dump_o_15_),
    .S(net1234),
    .X(\cs_registers_i/_0795_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3253_  (.Y(\cs_registers_i/_0796_ ),
    .B1(\cs_registers_i/_0795_ ),
    .B2(net1114),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_15_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3254_  (.A(\cs_registers_i/_0796_ ),
    .B_N(net1161),
    .Y(\cs_registers_i/_0797_ ));
 sg13g2_a21o_1 \cs_registers_i/_3255_  (.A2(\cs_registers_i/_0749_ ),
    .A1(csr_mtvec_15_),
    .B1(net1118),
    .X(\cs_registers_i/_0798_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3256_  (.B1(net56),
    .Y(\cs_registers_i/_0799_ ),
    .A1(\cs_registers_i/_0797_ ),
    .A2(\cs_registers_i/_0798_ ));
 sg13g2_mux2_1 \cs_registers_i/_3257_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_15_ ),
    .A1(\cs_registers_i/mhpmcounter_1871_ ),
    .S(net73),
    .X(\cs_registers_i/_0800_ ));
 sg13g2_nand2_1 \cs_registers_i/_3258_  (.Y(\cs_registers_i/_0801_ ),
    .A(\cs_registers_i/_0722_ ),
    .B(\cs_registers_i/_0800_ ));
 sg13g2_mux4_1 \cs_registers_i/_3259_  (.S0(net65),
    .A0(debug_ebreakm),
    .A1(\cs_registers_i/dscratch0_q_15_ ),
    .A2(csr_depc_15_),
    .A3(\cs_registers_i/dscratch1_q_15_ ),
    .S1(net1232),
    .X(\cs_registers_i/_0802_ ));
 sg13g2_nand2_1 \cs_registers_i/_3260_  (.Y(\cs_registers_i/_0803_ ),
    .A(net1150),
    .B(\cs_registers_i/_0802_ ));
 sg13g2_mux2_1 \cs_registers_i/_3261_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_47_ ),
    .A1(\cs_registers_i/mhpmcounter_1903_ ),
    .S(net63),
    .X(\cs_registers_i/_0804_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3262_  (.Y(\cs_registers_i/_0805_ ),
    .B1(\cs_registers_i/_0804_ ),
    .B2(net1129),
    .A2(net1095),
    .A1(hart_id_i_15_));
 sg13g2_and4_2 \cs_registers_i/_3263_  (.A(\cs_registers_i/_0799_ ),
    .B(\cs_registers_i/_0801_ ),
    .C(\cs_registers_i/_0803_ ),
    .D(\cs_registers_i/_0805_ ),
    .X(\cs_registers_i/_0806_ ));
 sg13g2_nor3_1 \cs_registers_i/_3264_  (.A(net1351),
    .B(net1090),
    .C(\cs_registers_i/_0806_ ),
    .Y(\cs_registers_i/_0807_ ));
 sg13g2_a21o_2 \cs_registers_i/_3265_  (.A2(net260),
    .A1(net1351),
    .B1(\cs_registers_i/_0807_ ),
    .X(\cs_registers_i/_0808_ ));
 sg13g2_buf_2 fanout574 (.A(net575),
    .X(net574));
 sg13g2_a22oi_1 \cs_registers_i/_3267_  (.Y(\cs_registers_i/_0810_ ),
    .B1(net1068),
    .B2(net654),
    .A2(\cs_registers_i/_0794_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3268_  (.Y(\cs_registers_i/_0016_ ),
    .A(\cs_registers_i/_0793_ ),
    .B(\cs_registers_i/_0810_ ));
 sg13g2_nand2_1 \cs_registers_i/_3269_  (.Y(\cs_registers_i/_0811_ ),
    .A(csr_depc_16_),
    .B(net660));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_mux2_2 \cs_registers_i/_3271_  (.A0(crash_dump_o_112_),
    .A1(crash_dump_o_80_),
    .S(net1481),
    .X(\cs_registers_i/_0813_ ));
 sg13g2_nor4_2 \cs_registers_i/_3272_  (.A(net1273),
    .B(net80),
    .C(\cs_registers_i/_0490_ ),
    .Y(\cs_registers_i/_0814_ ),
    .D(\cs_registers_i/_0518_ ));
 sg13g2_mux2_1 \cs_registers_i/_3273_  (.A0(\cs_registers_i/mie_q_0_ ),
    .A1(csr_mtvec_16_),
    .S(net1242),
    .X(\cs_registers_i/_0815_ ));
 sg13g2_nand2_1 \cs_registers_i/_3274_  (.Y(\cs_registers_i/_0816_ ),
    .A(net1094),
    .B(\cs_registers_i/_0815_ ));
 sg13g2_mux2_1 \cs_registers_i/_3275_  (.A0(crash_dump_o_16_),
    .A1(\cs_registers_i/mtval_q_16_ ),
    .S(net62),
    .X(\cs_registers_i/_0817_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3276_  (.A(net75),
    .B_N(net100),
    .Y(\cs_registers_i/_0818_ ));
 sg13g2_and2_2 \cs_registers_i/_3277_  (.A(net53),
    .B(\cs_registers_i/_0818_ ),
    .X(\cs_registers_i/_0819_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3278_  (.Y(\cs_registers_i/_0820_ ),
    .B1(\cs_registers_i/_0819_ ),
    .B2(irq_fast_i_0_),
    .A2(\cs_registers_i/_0817_ ),
    .A1(net1174));
 sg13g2_nor3_2 \cs_registers_i/_3279_  (.A(net144),
    .B(\cs_registers_i/_0601_ ),
    .C(\cs_registers_i/_0497_ ),
    .Y(\cs_registers_i/_0821_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3280_  (.Y(\cs_registers_i/_0822_ ),
    .B(\cs_registers_i/_0821_ ),
    .A_N(\cs_registers_i/_0820_ ));
 sg13g2_nand3b_1 \cs_registers_i/_3281_  (.B(\cs_registers_i/_0816_ ),
    .C(\cs_registers_i/_0822_ ),
    .Y(\cs_registers_i/_0823_ ),
    .A_N(net1119));
 sg13g2_mux4_1 \cs_registers_i/_3282_  (.S0(net69),
    .A0(\cs_registers_i/dcsr_q_16_ ),
    .A1(\cs_registers_i/dscratch0_q_16_ ),
    .A2(csr_depc_16_),
    .A3(\cs_registers_i/dscratch1_q_16_ ),
    .S1(net1237),
    .X(\cs_registers_i/_0824_ ));
 sg13g2_mux2_1 \cs_registers_i/_3283_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .A1(\cs_registers_i/mhpmcounter_1872_ ),
    .S(net72),
    .X(\cs_registers_i/_0825_ ));
 sg13g2_nand2_1 \cs_registers_i/_3284_  (.Y(\cs_registers_i/_0826_ ),
    .A(\cs_registers_i/_0628_ ),
    .B(\cs_registers_i/_0825_ ));
 sg13g2_nor3_2 \cs_registers_i/_3285_  (.A(net1172),
    .B(\cs_registers_i/_0557_ ),
    .C(\cs_registers_i/_0603_ ),
    .Y(\cs_registers_i/_0827_ ));
 sg13g2_nand3_1 \cs_registers_i/_3286_  (.B(\cs_registers_i/_0546_ ),
    .C(net1149),
    .A(\cs_registers_i/mscratch_q_16_ ),
    .Y(\cs_registers_i/_0828_ ));
 sg13g2_mux2_1 \cs_registers_i/_3287_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .A1(\cs_registers_i/mhpmcounter_1904_ ),
    .S(net70),
    .X(\cs_registers_i/_0829_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3288_  (.Y(\cs_registers_i/_0830_ ),
    .B1(\cs_registers_i/_0829_ ),
    .B2(net1129),
    .A2(net1095),
    .A1(hart_id_i_16_));
 sg13g2_nand3_1 \cs_registers_i/_3289_  (.B(\cs_registers_i/_0828_ ),
    .C(\cs_registers_i/_0830_ ),
    .A(\cs_registers_i/_0826_ ),
    .Y(\cs_registers_i/_0831_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3290_  (.B2(net1152),
    .C1(\cs_registers_i/_0831_ ),
    .B1(\cs_registers_i/_0824_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0832_ ),
    .A2(\cs_registers_i/_0823_ ));
 sg13g2_nor3_1 \cs_registers_i/_3291_  (.A(alu_operand_a_ex_16_),
    .B(net1090),
    .C(\cs_registers_i/_0832_ ),
    .Y(\cs_registers_i/_0833_ ));
 sg13g2_a21o_2 \cs_registers_i/_3292_  (.A2(net260),
    .A1(alu_operand_a_ex_16_),
    .B1(\cs_registers_i/_0833_ ),
    .X(\cs_registers_i/_0834_ ));
 sg13g2_buf_1 fanout572 (.A(rf_wdata_wb_29_),
    .X(net572));
 sg13g2_a22oi_1 \cs_registers_i/_3294_  (.Y(\cs_registers_i/_0836_ ),
    .B1(net1055),
    .B2(net655),
    .A2(\cs_registers_i/_0813_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3295_  (.Y(\cs_registers_i/_0017_ ),
    .A(\cs_registers_i/_0811_ ),
    .B(\cs_registers_i/_0836_ ));
 sg13g2_nand2_1 \cs_registers_i/_3296_  (.Y(\cs_registers_i/_0837_ ),
    .A(csr_depc_17_),
    .B(net660));
 sg13g2_buf_2 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout570 (.A(net571),
    .X(net570));
 sg13g2_mux2_2 \cs_registers_i/_3299_  (.A0(crash_dump_o_113_),
    .A1(crash_dump_o_81_),
    .S(net1482),
    .X(\cs_registers_i/_0840_ ));
 sg13g2_buf_2 fanout569 (.A(rf_wdata_wb_29_),
    .X(net569));
 sg13g2_nor2_2 \cs_registers_i/_3301_  (.A(net101),
    .B(\cs_registers_i/_0529_ ),
    .Y(\cs_registers_i/_0842_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3302_  (.Y(\cs_registers_i/_0843_ ),
    .B1(\cs_registers_i/_0842_ ),
    .B2(\cs_registers_i/mtval_q_17_ ),
    .A2(\cs_registers_i/_0819_ ),
    .A1(irq_fast_i_1_));
 sg13g2_nand2b_1 \cs_registers_i/_3303_  (.Y(\cs_registers_i/_0844_ ),
    .B(\cs_registers_i/_0821_ ),
    .A_N(\cs_registers_i/_0843_ ));
 sg13g2_mux2_1 \cs_registers_i/_3304_  (.A0(\cs_registers_i/mscratch_q_17_ ),
    .A1(crash_dump_o_17_),
    .S(net1241),
    .X(\cs_registers_i/_0845_ ));
 sg13g2_nand3_1 \cs_registers_i/_3305_  (.B(net1161),
    .C(\cs_registers_i/_0845_ ),
    .A(\cs_registers_i/_0773_ ),
    .Y(\cs_registers_i/_0846_ ));
 sg13g2_inv_1 \cs_registers_i/_3306_  (.Y(\cs_registers_i/_0847_ ),
    .A(\cs_registers_i/mstatus_q_1_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3307_  (.A1(\cs_registers_i/_0847_ ),
    .A2(\cs_registers_i/_0504_ ),
    .Y(\cs_registers_i/_0848_ ),
    .B1(net1269));
 sg13g2_mux2_1 \cs_registers_i/_3308_  (.A0(\cs_registers_i/mie_q_1_ ),
    .A1(csr_mtvec_17_),
    .S(net1241),
    .X(\cs_registers_i/_0849_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3309_  (.Y(\cs_registers_i/_0850_ ),
    .B1(\cs_registers_i/_0849_ ),
    .B2(net1094),
    .A2(\cs_registers_i/_0848_ ),
    .A1(\cs_registers_i/_0673_ ));
 sg13g2_nand3_1 \cs_registers_i/_3310_  (.B(\cs_registers_i/_0846_ ),
    .C(\cs_registers_i/_0850_ ),
    .A(\cs_registers_i/_0844_ ),
    .Y(\cs_registers_i/_0851_ ));
 sg13g2_mux4_1 \cs_registers_i/_3311_  (.S0(net66),
    .A0(\cs_registers_i/dcsr_q_17_ ),
    .A1(\cs_registers_i/dscratch0_q_17_ ),
    .A2(csr_depc_17_),
    .A3(\cs_registers_i/dscratch1_q_17_ ),
    .S1(net1244),
    .X(\cs_registers_i/_0852_ ));
 sg13g2_mux2_1 \cs_registers_i/_3312_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .A1(\cs_registers_i/mhpmcounter_1905_ ),
    .S(net70),
    .X(\cs_registers_i/_0853_ ));
 sg13g2_mux2_1 \cs_registers_i/_3313_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_17_ ),
    .A1(\cs_registers_i/mhpmcounter_1873_ ),
    .S(net72),
    .X(\cs_registers_i/_0854_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3314_  (.Y(\cs_registers_i/_0855_ ),
    .B1(\cs_registers_i/_0854_ ),
    .B2(\cs_registers_i/_0550_ ),
    .A2(\cs_registers_i/_0853_ ),
    .A1(net1157));
 sg13g2_nand2_1 \cs_registers_i/_3315_  (.Y(\cs_registers_i/_0856_ ),
    .A(hart_id_i_17_),
    .B(net1095));
 sg13g2_o21ai_1 \cs_registers_i/_3316_  (.B1(\cs_registers_i/_0856_ ),
    .Y(\cs_registers_i/_0857_ ),
    .A1(net1158),
    .A2(\cs_registers_i/_0855_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3317_  (.B2(net1152),
    .C1(\cs_registers_i/_0857_ ),
    .B1(\cs_registers_i/_0852_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0858_ ),
    .A2(\cs_registers_i/_0851_ ));
 sg13g2_nor3_1 \cs_registers_i/_3318_  (.A(net1251),
    .B(net1091),
    .C(\cs_registers_i/_0858_ ),
    .Y(\cs_registers_i/_0859_ ));
 sg13g2_a21o_2 \cs_registers_i/_3319_  (.A2(net260),
    .A1(net1251),
    .B1(\cs_registers_i/_0859_ ),
    .X(\cs_registers_i/_0860_ ));
 sg13g2_buf_1 fanout568 (.A(net569),
    .X(net568));
 sg13g2_a22oi_1 \cs_registers_i/_3321_  (.Y(\cs_registers_i/_0862_ ),
    .B1(net1053),
    .B2(net655),
    .A2(\cs_registers_i/_0840_ ),
    .A1(net1310));
 sg13g2_nand2_1 \cs_registers_i/_3322_  (.Y(\cs_registers_i/_0018_ ),
    .A(\cs_registers_i/_0837_ ),
    .B(\cs_registers_i/_0862_ ));
 sg13g2_nand2_1 \cs_registers_i/_3323_  (.Y(\cs_registers_i/_0863_ ),
    .A(csr_depc_18_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3324_  (.A0(crash_dump_o_114_),
    .A1(crash_dump_o_82_),
    .S(net1480),
    .X(\cs_registers_i/_0864_ ));
 sg13g2_mux2_1 \cs_registers_i/_3325_  (.A0(\cs_registers_i/mie_q_2_ ),
    .A1(csr_mtvec_18_),
    .S(net1239),
    .X(\cs_registers_i/_0865_ ));
 sg13g2_a21o_1 \cs_registers_i/_3326_  (.A2(\cs_registers_i/_0865_ ),
    .A1(net1094),
    .B1(net1118),
    .X(\cs_registers_i/_0866_ ));
 sg13g2_buf_2 fanout567 (.A(net569),
    .X(net567));
 sg13g2_buf_4 fanout566 (.X(net566),
    .A(rf_wdata_wb_31_));
 sg13g2_a22oi_1 \cs_registers_i/_3329_  (.Y(\cs_registers_i/_0869_ ),
    .B1(net1132),
    .B2(\cs_registers_i/mscratch_q_18_ ),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_18_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3330_  (.Y(\cs_registers_i/_0870_ ),
    .B1(\cs_registers_i/_0636_ ),
    .B2(irq_fast_i_2_),
    .A2(net1173),
    .A1(crash_dump_o_18_));
 sg13g2_or2_1 \cs_registers_i/_3331_  (.X(\cs_registers_i/_0871_ ),
    .B(\cs_registers_i/_0870_ ),
    .A(net1101));
 sg13g2_o21ai_1 \cs_registers_i/_3332_  (.B1(\cs_registers_i/_0871_ ),
    .Y(\cs_registers_i/_0872_ ),
    .A1(net1193),
    .A2(\cs_registers_i/_0869_ ));
 sg13g2_buf_2 fanout565 (.A(net566),
    .X(net565));
 sg13g2_mux4_1 \cs_registers_i/_3334_  (.S0(net69),
    .A0(\cs_registers_i/dcsr_q_18_ ),
    .A1(\cs_registers_i/dscratch0_q_18_ ),
    .A2(csr_depc_18_),
    .A3(\cs_registers_i/dscratch1_q_18_ ),
    .S1(net1237),
    .X(\cs_registers_i/_0874_ ));
 sg13g2_nand2_1 \cs_registers_i/_3335_  (.Y(\cs_registers_i/_0875_ ),
    .A(net1150),
    .B(\cs_registers_i/_0874_ ));
 sg13g2_nand3_1 \cs_registers_i/_3336_  (.B(\cs_registers_i/_0625_ ),
    .C(\cs_registers_i/_0629_ ),
    .A(\cs_registers_i/_0541_ ),
    .Y(\cs_registers_i/_0876_ ));
 sg13g2_nor4_2 \cs_registers_i/_3337_  (.A(net99),
    .B(net1235),
    .C(\cs_registers_i/_0601_ ),
    .Y(\cs_registers_i/_0877_ ),
    .D(\cs_registers_i/_0876_ ));
 sg13g2_mux4_1 \cs_registers_i/_3338_  (.S0(net65),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_18_ ),
    .A1(\cs_registers_i/mhpmcounter_1874_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_50_ ),
    .A3(\cs_registers_i/mhpmcounter_1906_ ),
    .S1(net147),
    .X(\cs_registers_i/_0878_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3339_  (.Y(\cs_registers_i/_0879_ ),
    .B1(\cs_registers_i/_0877_ ),
    .B2(\cs_registers_i/_0878_ ),
    .A2(net1096),
    .A1(hart_id_i_18_));
 sg13g2_nand2_1 \cs_registers_i/_3340_  (.Y(\cs_registers_i/_0880_ ),
    .A(\cs_registers_i/_0875_ ),
    .B(\cs_registers_i/_0879_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3341_  (.B2(net1148),
    .C1(\cs_registers_i/_0880_ ),
    .B1(\cs_registers_i/_0872_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0881_ ),
    .A2(\cs_registers_i/_0866_ ));
 sg13g2_nor3_1 \cs_registers_i/_3342_  (.A(alu_operand_a_ex_18_),
    .B(net1091),
    .C(\cs_registers_i/_0881_ ),
    .Y(\cs_registers_i/_0882_ ));
 sg13g2_a21o_2 \cs_registers_i/_3343_  (.A2(net262),
    .A1(alu_operand_a_ex_18_),
    .B1(\cs_registers_i/_0882_ ),
    .X(\cs_registers_i/_0883_ ));
 sg13g2_buf_2 fanout564 (.A(net566),
    .X(net564));
 sg13g2_a22oi_1 \cs_registers_i/_3345_  (.Y(\cs_registers_i/_0885_ ),
    .B1(net1051),
    .B2(net656),
    .A2(\cs_registers_i/_0864_ ),
    .A1(net1314));
 sg13g2_nand2_1 \cs_registers_i/_3346_  (.Y(\cs_registers_i/_0019_ ),
    .A(\cs_registers_i/_0863_ ),
    .B(\cs_registers_i/_0885_ ));
 sg13g2_nand2_1 \cs_registers_i/_3347_  (.Y(\cs_registers_i/_0886_ ),
    .A(csr_depc_19_),
    .B(net660));
 sg13g2_mux2_2 \cs_registers_i/_3348_  (.A0(crash_dump_o_115_),
    .A1(crash_dump_o_83_),
    .S(net1480),
    .X(\cs_registers_i/_0887_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3349_  (.Y(\cs_registers_i/_0888_ ),
    .B1(\cs_registers_i/_0636_ ),
    .B2(irq_fast_i_3_),
    .A2(net1173),
    .A1(crash_dump_o_19_));
 sg13g2_a22oi_1 \cs_registers_i/_3350_  (.Y(\cs_registers_i/_0889_ ),
    .B1(net1132),
    .B2(\cs_registers_i/mscratch_q_19_ ),
    .A2(net1116),
    .A1(\cs_registers_i/mtval_q_19_ ));
 sg13g2_inv_1 \cs_registers_i/_3351_  (.Y(\cs_registers_i/_0890_ ),
    .A(\cs_registers_i/_0889_ ));
 sg13g2_mux2_1 \cs_registers_i/_3352_  (.A0(\cs_registers_i/mie_q_3_ ),
    .A1(csr_mtvec_19_),
    .S(net1240),
    .X(\cs_registers_i/_0891_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3353_  (.B2(net1094),
    .C1(net1118),
    .B1(\cs_registers_i/_0891_ ),
    .A1(net1161),
    .Y(\cs_registers_i/_0892_ ),
    .A2(\cs_registers_i/_0890_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3354_  (.B1(\cs_registers_i/_0892_ ),
    .Y(\cs_registers_i/_0893_ ),
    .A1(\cs_registers_i/_0675_ ),
    .A2(\cs_registers_i/_0888_ ));
 sg13g2_mux4_1 \cs_registers_i/_3355_  (.S0(net68),
    .A0(\cs_registers_i/dcsr_q_19_ ),
    .A1(\cs_registers_i/dscratch0_q_19_ ),
    .A2(csr_depc_19_),
    .A3(\cs_registers_i/dscratch1_q_19_ ),
    .S1(net1243),
    .X(\cs_registers_i/_0894_ ));
 sg13g2_or2_1 \cs_registers_i/_3356_  (.X(\cs_registers_i/_0895_ ),
    .B(net1159),
    .A(\cs_registers_i/_0490_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3357_  (.A(net76),
    .B_N(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .Y(\cs_registers_i/_0896_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3358_  (.B1(\cs_registers_i/_0896_ ),
    .Y(\cs_registers_i/_0897_ ),
    .A2(\cs_registers_i/mhpmcounter_1875_ ),
    .A1(net75));
 sg13g2_mux2_1 \cs_registers_i/_3359_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_51_ ),
    .A1(\cs_registers_i/mhpmcounter_1907_ ),
    .S(net63),
    .X(\cs_registers_i/_0898_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3360_  (.Y(\cs_registers_i/_0899_ ),
    .B1(\cs_registers_i/_0898_ ),
    .B2(net1130),
    .A2(net1096),
    .A1(hart_id_i_19_));
 sg13g2_o21ai_1 \cs_registers_i/_3361_  (.B1(\cs_registers_i/_0899_ ),
    .Y(\cs_registers_i/_0900_ ),
    .A1(\cs_registers_i/_0895_ ),
    .A2(\cs_registers_i/_0897_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3362_  (.B2(net1151),
    .C1(\cs_registers_i/_0900_ ),
    .B1(\cs_registers_i/_0894_ ),
    .A1(net57),
    .Y(\cs_registers_i/_0901_ ),
    .A2(\cs_registers_i/_0893_ ));
 sg13g2_nor3_1 \cs_registers_i/_3363_  (.A(net1249),
    .B(net1089),
    .C(\cs_registers_i/_0901_ ),
    .Y(\cs_registers_i/_0902_ ));
 sg13g2_a21o_2 \cs_registers_i/_3364_  (.A2(net260),
    .A1(net1249),
    .B1(\cs_registers_i/_0902_ ),
    .X(\cs_registers_i/_0903_ ));
 sg13g2_buf_2 fanout563 (.A(net566),
    .X(net563));
 sg13g2_a22oi_1 \cs_registers_i/_3366_  (.Y(\cs_registers_i/_0905_ ),
    .B1(net1050),
    .B2(net655),
    .A2(\cs_registers_i/_0887_ ),
    .A1(net1310));
 sg13g2_nand2_1 \cs_registers_i/_3367_  (.Y(\cs_registers_i/_0020_ ),
    .A(\cs_registers_i/_0886_ ),
    .B(\cs_registers_i/_0905_ ));
 sg13g2_buf_2 fanout562 (.A(net566),
    .X(net562));
 sg13g2_nand2_1 \cs_registers_i/_3369_  (.Y(\cs_registers_i/_0907_ ),
    .A(csr_depc_1_),
    .B(net659));
 sg13g2_mux2_1 \cs_registers_i/_3370_  (.A0(crash_dump_o_97_),
    .A1(net560),
    .S(net1483),
    .X(\cs_registers_i/_0908_ ));
 sg13g2_mux2_1 \cs_registers_i/_3371_  (.A0(\cs_registers_i/dscratch0_q_1_ ),
    .A1(\cs_registers_i/dscratch1_q_1_ ),
    .S(net1245),
    .X(\cs_registers_i/_0909_ ));
 sg13g2_nand2_1 \cs_registers_i/_3372_  (.Y(\cs_registers_i/_0910_ ),
    .A(net80),
    .B(\cs_registers_i/_0909_ ));
 sg13g2_nand3_1 \cs_registers_i/_3373_  (.B(net54),
    .C(\cs_registers_i/dcsr_q_1_ ),
    .A(net1114),
    .Y(\cs_registers_i/_0911_ ));
 sg13g2_nand2_2 \cs_registers_i/_3374_  (.Y(\cs_registers_i/_0912_ ),
    .A(\cs_registers_i/_0544_ ),
    .B(net59));
 sg13g2_a21o_1 \cs_registers_i/_3375_  (.A2(\cs_registers_i/_0911_ ),
    .A1(\cs_registers_i/_0910_ ),
    .B1(\cs_registers_i/_0912_ ),
    .X(\cs_registers_i/_0913_ ));
 sg13g2_mux2_1 \cs_registers_i/_3376_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .A1(\cs_registers_i/mhpmcounter_1889_ ),
    .S(net64),
    .X(\cs_registers_i/_0914_ ));
 sg13g2_inv_1 \cs_registers_i/_3377_  (.Y(\cs_registers_i/_0915_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_1_ ));
 sg13g2_nand2_1 \cs_registers_i/_3378_  (.Y(\cs_registers_i/_0916_ ),
    .A(net74),
    .B(\cs_registers_i/mhpmcounter_1857_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3379_  (.B1(\cs_registers_i/_0916_ ),
    .Y(\cs_registers_i/_0917_ ),
    .A1(net71),
    .A2(\cs_registers_i/_0915_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3380_  (.Y(\cs_registers_i/_0918_ ),
    .B1(\cs_registers_i/_0917_ ),
    .B2(net1191),
    .A2(\cs_registers_i/_0914_ ),
    .A1(net1156));
 sg13g2_or2_1 \cs_registers_i/_3381_  (.X(\cs_registers_i/_0919_ ),
    .B(\cs_registers_i/_0918_ ),
    .A(net1159));
 sg13g2_mux4_1 \cs_registers_i/_3382_  (.S0(net67),
    .A0(\cs_registers_i/mscratch_q_1_ ),
    .A1(\cs_registers_i/mcause_q_1_ ),
    .A2(crash_dump_o_1_),
    .A3(\cs_registers_i/mtval_q_1_ ),
    .S1(net1231),
    .X(\cs_registers_i/_0920_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3383_  (.Y(\cs_registers_i/_0921_ ),
    .B1(\cs_registers_i/_0605_ ),
    .B2(\cs_registers_i/_0920_ ),
    .A2(\cs_registers_i/_0600_ ),
    .A1(csr_mtvec_1_));
 sg13g2_or3_1 \cs_registers_i/_3384_  (.A(\cs_registers_i/_0505_ ),
    .B(\cs_registers_i/_0535_ ),
    .C(\cs_registers_i/_0560_ ),
    .X(\cs_registers_i/_0922_ ));
 sg13g2_nor2_1 \cs_registers_i/_3385_  (.A(net1275),
    .B(\cs_registers_i/_0922_ ),
    .Y(\cs_registers_i/_0923_ ));
 sg13g2_nand3_1 \cs_registers_i/_3386_  (.B(hart_id_i_1_),
    .C(net1131),
    .A(net102),
    .Y(\cs_registers_i/_0924_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3387_  (.B1(\cs_registers_i/_0924_ ),
    .Y(\cs_registers_i/_0925_ ),
    .A1(net100),
    .A2(\cs_registers_i/_0536_ ));
 sg13g2_inv_1 \cs_registers_i/_3388_  (.Y(\cs_registers_i/_0926_ ),
    .A(csr_depc_1_));
 sg13g2_nand2_1 \cs_registers_i/_3389_  (.Y(\cs_registers_i/_0927_ ),
    .A(net1235),
    .B(\cs_registers_i/_0525_ ));
 sg13g2_nor3_1 \cs_registers_i/_3390_  (.A(\cs_registers_i/_0926_ ),
    .B(net1275),
    .C(\cs_registers_i/_0927_ ),
    .Y(\cs_registers_i/_0928_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3391_  (.Y(\cs_registers_i/_0929_ ),
    .B1(\cs_registers_i/_0928_ ),
    .B2(net60),
    .A2(\cs_registers_i/_0925_ ),
    .A1(\cs_registers_i/_0923_ ));
 sg13g2_and4_2 \cs_registers_i/_3392_  (.A(\cs_registers_i/_0913_ ),
    .B(\cs_registers_i/_0919_ ),
    .C(\cs_registers_i/_0921_ ),
    .D(\cs_registers_i/_0929_ ),
    .X(\cs_registers_i/_0930_ ));
 sg13g2_nor3_1 \cs_registers_i/_3393_  (.A(net1411),
    .B(net1088),
    .C(\cs_registers_i/_0930_ ),
    .Y(\cs_registers_i/_0931_ ));
 sg13g2_a21o_2 \cs_registers_i/_3394_  (.A2(net260),
    .A1(alu_operand_a_ex_1_),
    .B1(\cs_registers_i/_0931_ ),
    .X(\cs_registers_i/_0932_ ));
 sg13g2_buf_2 fanout561 (.A(crash_dump_o_65_),
    .X(net561));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_a22oi_1 \cs_registers_i/_3397_  (.Y(\cs_registers_i/_0935_ ),
    .B1(net1067),
    .B2(net654),
    .A2(\cs_registers_i/_0908_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3398_  (.Y(\cs_registers_i/_0021_ ),
    .A(\cs_registers_i/_0907_ ),
    .B(\cs_registers_i/_0935_ ));
 sg13g2_nand2_1 \cs_registers_i/_3399_  (.Y(\cs_registers_i/_0936_ ),
    .A(csr_depc_20_),
    .B(net661));
 sg13g2_mux2_2 \cs_registers_i/_3400_  (.A0(crash_dump_o_116_),
    .A1(crash_dump_o_84_),
    .S(net1480),
    .X(\cs_registers_i/_0937_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3401_  (.A(net102),
    .B_N(\cs_registers_i/mscratch_q_20_ ),
    .Y(\cs_registers_i/_0938_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3402_  (.A1(net102),
    .A2(irq_fast_i_4_),
    .Y(\cs_registers_i/_0939_ ),
    .B1(\cs_registers_i/_0938_ ));
 sg13g2_nor3_1 \cs_registers_i/_3403_  (.A(net1236),
    .B(net1100),
    .C(\cs_registers_i/_0939_ ),
    .Y(\cs_registers_i/_0940_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3404_  (.A(net74),
    .B_N(crash_dump_o_20_),
    .Y(\cs_registers_i/_0941_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3405_  (.A1(net76),
    .A2(\cs_registers_i/mtval_q_20_ ),
    .Y(\cs_registers_i/_0942_ ),
    .B1(\cs_registers_i/_0941_ ));
 sg13g2_nor3_1 \cs_registers_i/_3406_  (.A(net53),
    .B(net1193),
    .C(\cs_registers_i/_0942_ ),
    .Y(\cs_registers_i/_0943_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3407_  (.B1(net1149),
    .Y(\cs_registers_i/_0944_ ),
    .A1(\cs_registers_i/_0940_ ),
    .A2(\cs_registers_i/_0943_ ));
 sg13g2_mux2_1 \cs_registers_i/_3408_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_20_ ),
    .A1(\cs_registers_i/mhpmcounter_1876_ ),
    .S(net73),
    .X(\cs_registers_i/_0945_ ));
 sg13g2_nand2_2 \cs_registers_i/_3409_  (.Y(\cs_registers_i/_0946_ ),
    .A(net57),
    .B(\cs_registers_i/_0720_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3410_  (.Y(\cs_registers_i/_0947_ ),
    .B1(\cs_registers_i/_0598_ ),
    .B2(csr_mtvec_20_),
    .A2(\cs_registers_i/_0519_ ),
    .A1(\cs_registers_i/mie_q_4_ ));
 sg13g2_nor2_2 \cs_registers_i/_3411_  (.A(net1192),
    .B(\cs_registers_i/_0529_ ),
    .Y(\cs_registers_i/_0948_ ));
 sg13g2_nand3_1 \cs_registers_i/_3412_  (.B(net59),
    .C(\cs_registers_i/_0948_ ),
    .A(\cs_registers_i/dscratch1_q_20_ ),
    .Y(\cs_registers_i/_0949_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3413_  (.B1(\cs_registers_i/_0949_ ),
    .Y(\cs_registers_i/_0950_ ),
    .A1(\cs_registers_i/_0946_ ),
    .A2(\cs_registers_i/_0947_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3414_  (.B2(\cs_registers_i/_0628_ ),
    .C1(\cs_registers_i/_0950_ ),
    .B1(\cs_registers_i/_0945_ ),
    .A1(hart_id_i_20_),
    .Y(\cs_registers_i/_0951_ ),
    .A2(net1098));
 sg13g2_mux2_2 \cs_registers_i/_3415_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_52_ ),
    .A1(\cs_registers_i/mhpmcounter_1908_ ),
    .S(net63),
    .X(\cs_registers_i/_0952_ ));
 sg13g2_and2_1 \cs_registers_i/_3416_  (.A(csr_depc_20_),
    .B(net1243),
    .X(\cs_registers_i/_0953_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3417_  (.A1(net54),
    .A2(\cs_registers_i/dcsr_q_20_ ),
    .Y(\cs_registers_i/_0954_ ),
    .B1(\cs_registers_i/_0953_ ));
 sg13g2_nand3_1 \cs_registers_i/_3418_  (.B(net54),
    .C(\cs_registers_i/dscratch0_q_20_ ),
    .A(net77),
    .Y(\cs_registers_i/_0955_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3419_  (.B1(\cs_registers_i/_0955_ ),
    .Y(\cs_registers_i/_0956_ ),
    .A1(net66),
    .A2(\cs_registers_i/_0954_ ));
 sg13g2_inv_1 \cs_registers_i/_3420_  (.Y(\cs_registers_i/_0957_ ),
    .A(\cs_registers_i/_0511_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3421_  (.B2(net1153),
    .C1(\cs_registers_i/_0957_ ),
    .B1(\cs_registers_i/_0956_ ),
    .A1(net1130),
    .Y(\cs_registers_i/_0958_ ),
    .A2(\cs_registers_i/_0952_ ));
 sg13g2_and3_2 \cs_registers_i/_3422_  (.X(\cs_registers_i/_0959_ ),
    .A(\cs_registers_i/_0944_ ),
    .B(\cs_registers_i/_0951_ ),
    .C(\cs_registers_i/_0958_ ));
 sg13g2_nor3_1 \cs_registers_i/_3423_  (.A(net1282),
    .B(net1089),
    .C(\cs_registers_i/_0959_ ),
    .Y(\cs_registers_i/_0960_ ));
 sg13g2_a21o_2 \cs_registers_i/_3424_  (.A2(net262),
    .A1(net1282),
    .B1(\cs_registers_i/_0960_ ),
    .X(\cs_registers_i/_0961_ ));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net561));
 sg13g2_a22oi_1 \cs_registers_i/_3426_  (.Y(\cs_registers_i/_0963_ ),
    .B1(net1049),
    .B2(net657),
    .A2(\cs_registers_i/_0937_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3427_  (.Y(\cs_registers_i/_0022_ ),
    .A(\cs_registers_i/_0936_ ),
    .B(\cs_registers_i/_0963_ ));
 sg13g2_nand2_1 \cs_registers_i/_3428_  (.Y(\cs_registers_i/_0964_ ),
    .A(csr_depc_21_),
    .B(net661));
 sg13g2_mux2_2 \cs_registers_i/_3429_  (.A0(crash_dump_o_117_),
    .A1(crash_dump_o_85_),
    .S(net1482),
    .X(\cs_registers_i/_0965_ ));
 sg13g2_mux2_1 \cs_registers_i/_3430_  (.A0(\cs_registers_i/mscratch_q_21_ ),
    .A1(crash_dump_o_21_),
    .S(net1240),
    .X(\cs_registers_i/_0966_ ));
 sg13g2_nand3_1 \cs_registers_i/_3431_  (.B(net1161),
    .C(\cs_registers_i/_0966_ ),
    .A(\cs_registers_i/_0773_ ),
    .Y(\cs_registers_i/_0967_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3432_  (.Y(\cs_registers_i/_0968_ ),
    .B1(\cs_registers_i/_0842_ ),
    .B2(\cs_registers_i/mtval_q_21_ ),
    .A2(\cs_registers_i/_0819_ ),
    .A1(irq_fast_i_5_));
 sg13g2_nand2b_1 \cs_registers_i/_3433_  (.Y(\cs_registers_i/_0969_ ),
    .B(\cs_registers_i/_0821_ ),
    .A_N(\cs_registers_i/_0968_ ));
 sg13g2_mux2_1 \cs_registers_i/_3434_  (.A0(\cs_registers_i/mie_q_5_ ),
    .A1(csr_mtvec_21_),
    .S(net1239),
    .X(\cs_registers_i/_0970_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3435_  (.Y(\cs_registers_i/_0971_ ),
    .B1(\cs_registers_i/_0970_ ),
    .B2(net102),
    .A2(\cs_registers_i/_0626_ ),
    .A1(csr_mstatus_tw));
 sg13g2_inv_1 \cs_registers_i/_3436_  (.Y(\cs_registers_i/_0972_ ),
    .A(\cs_registers_i/_0971_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3437_  (.A1(\cs_registers_i/_0667_ ),
    .A2(\cs_registers_i/_0972_ ),
    .Y(\cs_registers_i/_0973_ ),
    .B1(net1118));
 sg13g2_nand3_1 \cs_registers_i/_3438_  (.B(\cs_registers_i/_0969_ ),
    .C(\cs_registers_i/_0973_ ),
    .A(\cs_registers_i/_0967_ ),
    .Y(\cs_registers_i/_0974_ ));
 sg13g2_mux4_1 \cs_registers_i/_3439_  (.S0(net66),
    .A0(\cs_registers_i/dcsr_q_21_ ),
    .A1(\cs_registers_i/dscratch0_q_21_ ),
    .A2(csr_depc_21_),
    .A3(\cs_registers_i/dscratch1_q_21_ ),
    .S1(net1244),
    .X(\cs_registers_i/_0975_ ));
 sg13g2_mux2_1 \cs_registers_i/_3440_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_53_ ),
    .A1(\cs_registers_i/mhpmcounter_1909_ ),
    .S(net63),
    .X(\cs_registers_i/_0976_ ));
 sg13g2_mux2_1 \cs_registers_i/_3441_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_21_ ),
    .A1(\cs_registers_i/mhpmcounter_1877_ ),
    .S(net71),
    .X(\cs_registers_i/_0977_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3442_  (.Y(\cs_registers_i/_0978_ ),
    .B1(\cs_registers_i/_0977_ ),
    .B2(net1191),
    .A2(\cs_registers_i/_0976_ ),
    .A1(net1157));
 sg13g2_nand2_1 \cs_registers_i/_3443_  (.Y(\cs_registers_i/_0979_ ),
    .A(hart_id_i_21_),
    .B(net1095));
 sg13g2_o21ai_1 \cs_registers_i/_3444_  (.B1(\cs_registers_i/_0979_ ),
    .Y(\cs_registers_i/_0980_ ),
    .A1(net1158),
    .A2(\cs_registers_i/_0978_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3445_  (.B2(net1152),
    .C1(\cs_registers_i/_0980_ ),
    .B1(\cs_registers_i/_0975_ ),
    .A1(net58),
    .Y(\cs_registers_i/_0981_ ),
    .A2(\cs_registers_i/_0974_ ));
 sg13g2_nor3_1 \cs_registers_i/_3446_  (.A(net126),
    .B(net1091),
    .C(\cs_registers_i/_0981_ ),
    .Y(\cs_registers_i/_0982_ ));
 sg13g2_a21o_2 \cs_registers_i/_3447_  (.A2(net259),
    .A1(net127),
    .B1(\cs_registers_i/_0982_ ),
    .X(\cs_registers_i/_0983_ ));
 sg13g2_buf_4 fanout558 (.X(net558),
    .A(net561));
 sg13g2_a22oi_1 \cs_registers_i/_3449_  (.Y(\cs_registers_i/_0985_ ),
    .B1(net1047),
    .B2(net657),
    .A2(\cs_registers_i/_0965_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3450_  (.Y(\cs_registers_i/_0023_ ),
    .A(\cs_registers_i/_0964_ ),
    .B(\cs_registers_i/_0985_ ));
 sg13g2_nand2_1 \cs_registers_i/_3451_  (.Y(\cs_registers_i/_0986_ ),
    .A(csr_depc_22_),
    .B(net661));
 sg13g2_mux2_2 \cs_registers_i/_3452_  (.A0(crash_dump_o_118_),
    .A1(crash_dump_o_86_),
    .S(net1480),
    .X(\cs_registers_i/_0987_ ));
 sg13g2_nand2_1 \cs_registers_i/_3453_  (.Y(\cs_registers_i/_0988_ ),
    .A(\cs_registers_i/dcsr_q_22_ ),
    .B(net60));
 sg13g2_a21oi_1 \cs_registers_i/_3454_  (.A1(\cs_registers_i/_0648_ ),
    .A2(\cs_registers_i/_0988_ ),
    .Y(\cs_registers_i/_0989_ ),
    .B1(\cs_registers_i/_0506_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3455_  (.Y(\cs_registers_i/_0990_ ),
    .B1(\cs_registers_i/_0598_ ),
    .B2(csr_mtvec_22_),
    .A2(\cs_registers_i/_0519_ ),
    .A1(\cs_registers_i/mie_q_6_ ));
 sg13g2_inv_1 \cs_registers_i/_3456_  (.Y(\cs_registers_i/_0991_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_22_ ));
 sg13g2_nand2_1 \cs_registers_i/_3457_  (.Y(\cs_registers_i/_0992_ ),
    .A(net77),
    .B(\cs_registers_i/mhpmcounter_1878_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3458_  (.B1(\cs_registers_i/_0992_ ),
    .Y(\cs_registers_i/_0993_ ),
    .A1(net68),
    .A2(\cs_registers_i/_0991_ ));
 sg13g2_nand2_1 \cs_registers_i/_3459_  (.Y(\cs_registers_i/_0994_ ),
    .A(\cs_registers_i/_0628_ ),
    .B(\cs_registers_i/_0993_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3460_  (.B1(\cs_registers_i/_0994_ ),
    .Y(\cs_registers_i/_0995_ ),
    .A1(\cs_registers_i/_0946_ ),
    .A2(\cs_registers_i/_0990_ ));
 sg13g2_mux2_1 \cs_registers_i/_3461_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_54_ ),
    .A1(\cs_registers_i/mhpmcounter_1910_ ),
    .S(net63),
    .X(\cs_registers_i/_0996_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3462_  (.Y(\cs_registers_i/_0997_ ),
    .B1(\cs_registers_i/_0996_ ),
    .B2(net1129),
    .A2(net1095),
    .A1(hart_id_i_22_));
 sg13g2_inv_1 \cs_registers_i/_3463_  (.Y(\cs_registers_i/_0998_ ),
    .A(\cs_registers_i/_0997_ ));
 sg13g2_mux2_1 \cs_registers_i/_3464_  (.A0(\cs_registers_i/dscratch0_q_22_ ),
    .A1(\cs_registers_i/dscratch1_q_22_ ),
    .S(net1243),
    .X(\cs_registers_i/_0999_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3465_  (.Y(\cs_registers_i/_1000_ ),
    .B1(\cs_registers_i/_0999_ ),
    .B2(net77),
    .A2(\cs_registers_i/_0717_ ),
    .A1(csr_depc_22_));
 sg13g2_a22oi_1 \cs_registers_i/_3466_  (.Y(\cs_registers_i/_1001_ ),
    .B1(\cs_registers_i/_0636_ ),
    .B2(irq_fast_i_6_),
    .A2(net1173),
    .A1(crash_dump_o_22_));
 sg13g2_nor2_1 \cs_registers_i/_3467_  (.A(net1101),
    .B(\cs_registers_i/_1001_ ),
    .Y(\cs_registers_i/_1002_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3468_  (.Y(\cs_registers_i/_1003_ ),
    .B1(net1132),
    .B2(\cs_registers_i/mscratch_q_22_ ),
    .A2(net1116),
    .A1(\cs_registers_i/mtval_q_22_ ));
 sg13g2_nor2_1 \cs_registers_i/_3469_  (.A(net1193),
    .B(\cs_registers_i/_1003_ ),
    .Y(\cs_registers_i/_1004_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3470_  (.B1(net1148),
    .Y(\cs_registers_i/_1005_ ),
    .A1(\cs_registers_i/_1002_ ),
    .A2(\cs_registers_i/_1004_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3471_  (.B1(\cs_registers_i/_1005_ ),
    .Y(\cs_registers_i/_1006_ ),
    .A1(\cs_registers_i/_0912_ ),
    .A2(\cs_registers_i/_1000_ ));
 sg13g2_nor4_2 \cs_registers_i/_3472_  (.A(\cs_registers_i/_0989_ ),
    .B(\cs_registers_i/_0995_ ),
    .C(\cs_registers_i/_0998_ ),
    .Y(\cs_registers_i/_1007_ ),
    .D(\cs_registers_i/_1006_ ));
 sg13g2_nor3_1 \cs_registers_i/_3473_  (.A(net195),
    .B(net1089),
    .C(\cs_registers_i/_1007_ ),
    .Y(\cs_registers_i/_1008_ ));
 sg13g2_a21o_2 \cs_registers_i/_3474_  (.A2(net262),
    .A1(net196),
    .B1(\cs_registers_i/_1008_ ),
    .X(\cs_registers_i/_1009_ ));
 sg13g2_buf_2 fanout557 (.A(net561),
    .X(net557));
 sg13g2_a22oi_1 \cs_registers_i/_3476_  (.Y(\cs_registers_i/_1011_ ),
    .B1(net1027),
    .B2(net655),
    .A2(\cs_registers_i/_0987_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3477_  (.Y(\cs_registers_i/_0024_ ),
    .A(\cs_registers_i/_0986_ ),
    .B(\cs_registers_i/_1011_ ));
 sg13g2_nand2_1 \cs_registers_i/_3478_  (.Y(\cs_registers_i/_1012_ ),
    .A(csr_depc_23_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3479_  (.A0(crash_dump_o_119_),
    .A1(crash_dump_o_87_),
    .S(net1479),
    .X(\cs_registers_i/_1013_ ));
 sg13g2_mux4_1 \cs_registers_i/_3480_  (.S0(net65),
    .A0(\cs_registers_i/dcsr_q_23_ ),
    .A1(\cs_registers_i/dscratch0_q_23_ ),
    .A2(csr_depc_23_),
    .A3(\cs_registers_i/dscratch1_q_23_ ),
    .S1(net1237),
    .X(\cs_registers_i/_1014_ ));
 sg13g2_nor3_1 \cs_registers_i/_3481_  (.A(net1273),
    .B(net145),
    .C(\cs_registers_i/_0497_ ),
    .Y(\cs_registers_i/_1015_ ));
 sg13g2_nand3_1 \cs_registers_i/_3482_  (.B(\cs_registers_i/_0477_ ),
    .C(\cs_registers_i/_1015_ ),
    .A(crash_dump_o_23_),
    .Y(\cs_registers_i/_1016_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3483_  (.Y(\cs_registers_i/_1017_ ),
    .B1(\cs_registers_i/_0842_ ),
    .B2(\cs_registers_i/mtval_q_23_ ),
    .A2(\cs_registers_i/_0819_ ),
    .A1(irq_fast_i_7_));
 sg13g2_nand2b_1 \cs_registers_i/_3484_  (.Y(\cs_registers_i/_1018_ ),
    .B(\cs_registers_i/_0821_ ),
    .A_N(\cs_registers_i/_1017_ ));
 sg13g2_mux2_1 \cs_registers_i/_3485_  (.A0(\cs_registers_i/mie_q_7_ ),
    .A1(csr_mtvec_23_),
    .S(net1242),
    .X(\cs_registers_i/_1019_ ));
 sg13g2_nand2_1 \cs_registers_i/_3486_  (.Y(\cs_registers_i/_1020_ ),
    .A(net1094),
    .B(\cs_registers_i/_1019_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3487_  (.A1(\cs_registers_i/mscratch_q_23_ ),
    .A2(\cs_registers_i/_0669_ ),
    .Y(\cs_registers_i/_1021_ ),
    .B1(\cs_registers_i/_0670_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3488_  (.Y(\cs_registers_i/_1022_ ),
    .B(\cs_registers_i/_0673_ ),
    .A_N(\cs_registers_i/_1021_ ));
 sg13g2_nand4_1 \cs_registers_i/_3489_  (.B(\cs_registers_i/_1018_ ),
    .C(\cs_registers_i/_1020_ ),
    .A(\cs_registers_i/_1016_ ),
    .Y(\cs_registers_i/_1023_ ),
    .D(\cs_registers_i/_1022_ ));
 sg13g2_mux2_1 \cs_registers_i/_3490_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_55_ ),
    .A1(\cs_registers_i/mhpmcounter_1911_ ),
    .S(net73),
    .X(\cs_registers_i/_1024_ ));
 sg13g2_mux2_1 \cs_registers_i/_3491_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_23_ ),
    .A1(\cs_registers_i/mhpmcounter_1879_ ),
    .S(net67),
    .X(\cs_registers_i/_1025_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3492_  (.Y(\cs_registers_i/_1026_ ),
    .B1(\cs_registers_i/_1025_ ),
    .B2(net1191),
    .A2(\cs_registers_i/_1024_ ),
    .A1(net1157));
 sg13g2_nand2_1 \cs_registers_i/_3493_  (.Y(\cs_registers_i/_1027_ ),
    .A(hart_id_i_23_),
    .B(net1095));
 sg13g2_o21ai_1 \cs_registers_i/_3494_  (.B1(\cs_registers_i/_1027_ ),
    .Y(\cs_registers_i/_1028_ ),
    .A1(net1158),
    .A2(\cs_registers_i/_1026_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3495_  (.B2(net57),
    .C1(\cs_registers_i/_1028_ ),
    .B1(\cs_registers_i/_1023_ ),
    .A1(net1154),
    .Y(\cs_registers_i/_1029_ ),
    .A2(\cs_registers_i/_1014_ ));
 sg13g2_nor2_2 \cs_registers_i/_3496_  (.A(net1093),
    .B(\cs_registers_i/_1029_ ),
    .Y(\cs_registers_i/_1030_ ));
 sg13g2_mux2_2 \cs_registers_i/_3497_  (.A0(\cs_registers_i/_1030_ ),
    .A1(net259),
    .S(net149),
    .X(\cs_registers_i/_1031_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3498_  (.Y(\cs_registers_i/_1032_ ),
    .B1(net1046),
    .B2(net656),
    .A2(\cs_registers_i/_1013_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3499_  (.Y(\cs_registers_i/_0025_ ),
    .A(\cs_registers_i/_1012_ ),
    .B(\cs_registers_i/_1032_ ));
 sg13g2_nand2_1 \cs_registers_i/_3500_  (.Y(\cs_registers_i/_1033_ ),
    .A(csr_depc_24_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3501_  (.A0(crash_dump_o_120_),
    .A1(crash_dump_o_88_),
    .S(net1479),
    .X(\cs_registers_i/_1034_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3502_  (.A1(\cs_registers_i/mscratch_q_24_ ),
    .A2(\cs_registers_i/_0669_ ),
    .Y(\cs_registers_i/_1035_ ),
    .B1(\cs_registers_i/_0670_ ));
 sg13g2_or4_1 \cs_registers_i/_3503_  (.A(net1273),
    .B(net146),
    .C(\cs_registers_i/_0506_ ),
    .D(\cs_registers_i/_1035_ ),
    .X(\cs_registers_i/_1036_ ));
 sg13g2_mux2_1 \cs_registers_i/_3504_  (.A0(\cs_registers_i/mie_q_8_ ),
    .A1(csr_mtvec_24_),
    .S(net1241),
    .X(\cs_registers_i/_1037_ ));
 sg13g2_nand2_1 \cs_registers_i/_3505_  (.Y(\cs_registers_i/_1038_ ),
    .A(\cs_registers_i/_0814_ ),
    .B(\cs_registers_i/_1037_ ));
 sg13g2_mux2_1 \cs_registers_i/_3506_  (.A0(crash_dump_o_24_),
    .A1(\cs_registers_i/mtval_q_24_ ),
    .S(net62),
    .X(\cs_registers_i/_1039_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3507_  (.Y(\cs_registers_i/_1040_ ),
    .B1(\cs_registers_i/_1039_ ),
    .B2(net1174),
    .A2(\cs_registers_i/_0819_ ),
    .A1(irq_fast_i_8_));
 sg13g2_nand2b_1 \cs_registers_i/_3508_  (.Y(\cs_registers_i/_1041_ ),
    .B(\cs_registers_i/_0821_ ),
    .A_N(\cs_registers_i/_1040_ ));
 sg13g2_nand3_1 \cs_registers_i/_3509_  (.B(\cs_registers_i/_1038_ ),
    .C(\cs_registers_i/_1041_ ),
    .A(\cs_registers_i/_1036_ ),
    .Y(\cs_registers_i/_1042_ ));
 sg13g2_mux4_1 \cs_registers_i/_3510_  (.S0(net68),
    .A0(\cs_registers_i/dcsr_q_24_ ),
    .A1(\cs_registers_i/dscratch0_q_24_ ),
    .A2(csr_depc_24_),
    .A3(\cs_registers_i/dscratch1_q_24_ ),
    .S1(net1243),
    .X(\cs_registers_i/_1043_ ));
 sg13g2_inv_1 \cs_registers_i/_3511_  (.Y(\cs_registers_i/_1044_ ),
    .A(net1130));
 sg13g2_nor2b_1 \cs_registers_i/_3512_  (.A(net76),
    .B_N(\cs_registers_i/mcycle_counter_i.counter_val_o_56_ ),
    .Y(\cs_registers_i/_1045_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3513_  (.B1(\cs_registers_i/_1045_ ),
    .Y(\cs_registers_i/_1046_ ),
    .A2(\cs_registers_i/mhpmcounter_1912_ ),
    .A1(net77));
 sg13g2_mux2_1 \cs_registers_i/_3514_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .A1(\cs_registers_i/mhpmcounter_1880_ ),
    .S(net71),
    .X(\cs_registers_i/_1047_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3515_  (.Y(\cs_registers_i/_1048_ ),
    .B1(\cs_registers_i/_1047_ ),
    .B2(\cs_registers_i/_0628_ ),
    .A2(net1097),
    .A1(hart_id_i_24_));
 sg13g2_o21ai_1 \cs_registers_i/_3516_  (.B1(\cs_registers_i/_1048_ ),
    .Y(\cs_registers_i/_1049_ ),
    .A1(\cs_registers_i/_1044_ ),
    .A2(\cs_registers_i/_1046_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3517_  (.B2(net1152),
    .C1(\cs_registers_i/_1049_ ),
    .B1(\cs_registers_i/_1043_ ),
    .A1(net58),
    .Y(\cs_registers_i/_1050_ ),
    .A2(\cs_registers_i/_1042_ ));
 sg13g2_nor3_1 \cs_registers_i/_3518_  (.A(net125),
    .B(net1089),
    .C(\cs_registers_i/_1050_ ),
    .Y(\cs_registers_i/_1051_ ));
 sg13g2_a21o_2 \cs_registers_i/_3519_  (.A2(net262),
    .A1(alu_operand_a_ex_24_),
    .B1(\cs_registers_i/_1051_ ),
    .X(\cs_registers_i/_1052_ ));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(\ex_block_i.alu_i.imd_val_q_i_56_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3521_  (.Y(\cs_registers_i/_1054_ ),
    .B1(net1044),
    .B2(net656),
    .A2(\cs_registers_i/_1034_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3522_  (.Y(\cs_registers_i/_0026_ ),
    .A(\cs_registers_i/_1033_ ),
    .B(\cs_registers_i/_1054_ ));
 sg13g2_nand2_1 \cs_registers_i/_3523_  (.Y(\cs_registers_i/_1055_ ),
    .A(csr_depc_25_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3524_  (.A0(crash_dump_o_121_),
    .A1(crash_dump_o_89_),
    .S(net1479),
    .X(\cs_registers_i/_1056_ ));
 sg13g2_and2_1 \cs_registers_i/_3525_  (.A(csr_depc_25_),
    .B(net1246),
    .X(\cs_registers_i/_1057_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3526_  (.A1(net55),
    .A2(\cs_registers_i/dcsr_q_25_ ),
    .Y(\cs_registers_i/_1058_ ),
    .B1(\cs_registers_i/_1057_ ));
 sg13g2_nor3_1 \cs_registers_i/_3527_  (.A(net72),
    .B(\cs_registers_i/_0912_ ),
    .C(\cs_registers_i/_1058_ ),
    .Y(\cs_registers_i/_1059_ ));
 sg13g2_or2_1 \cs_registers_i/_3528_  (.X(\cs_registers_i/_1060_ ),
    .B(\cs_registers_i/_0648_ ),
    .A(\cs_registers_i/_0506_ ));
 sg13g2_and2_2 \cs_registers_i/_3529_  (.A(\cs_registers_i/_0544_ ),
    .B(\cs_registers_i/_0549_ ),
    .X(\cs_registers_i/_1061_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3530_  (.Y(\cs_registers_i/_1062_ ),
    .B1(\cs_registers_i/_1061_ ),
    .B2(\cs_registers_i/dscratch0_q_25_ ),
    .A2(\cs_registers_i/_0948_ ),
    .A1(\cs_registers_i/dscratch1_q_25_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3531_  (.Y(\cs_registers_i/_1063_ ),
    .B(net59),
    .A_N(\cs_registers_i/_1062_ ));
 sg13g2_nand2_1 \cs_registers_i/_3532_  (.Y(\cs_registers_i/_1064_ ),
    .A(hart_id_i_25_),
    .B(net1097));
 sg13g2_mux4_1 \cs_registers_i/_3533_  (.S0(net144),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_25_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_57_ ),
    .A2(\cs_registers_i/mhpmcounter_1881_ ),
    .A3(\cs_registers_i/mhpmcounter_1913_ ),
    .S1(csr_addr_1_),
    .X(\cs_registers_i/_1065_ ));
 sg13g2_nand2_1 \cs_registers_i/_3534_  (.Y(\cs_registers_i/_1066_ ),
    .A(\cs_registers_i/_0877_ ),
    .B(\cs_registers_i/_1065_ ));
 sg13g2_nand4_1 \cs_registers_i/_3535_  (.B(\cs_registers_i/_1063_ ),
    .C(\cs_registers_i/_1064_ ),
    .A(\cs_registers_i/_1060_ ),
    .Y(\cs_registers_i/_1067_ ),
    .D(\cs_registers_i/_1066_ ));
 sg13g2_nand2_1 \cs_registers_i/_3536_  (.Y(\cs_registers_i/_1068_ ),
    .A(net57),
    .B(net1094));
 sg13g2_and2_1 \cs_registers_i/_3537_  (.A(csr_mtvec_25_),
    .B(net1239),
    .X(\cs_registers_i/_1069_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3538_  (.A1(net55),
    .A2(\cs_registers_i/mie_q_9_ ),
    .Y(\cs_registers_i/_1070_ ),
    .B1(\cs_registers_i/_1069_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3539_  (.Y(\cs_registers_i/_1071_ ),
    .B1(net1155),
    .B2(irq_fast_i_9_),
    .A2(net1173),
    .A1(crash_dump_o_25_));
 sg13g2_nor2_1 \cs_registers_i/_3540_  (.A(net1101),
    .B(\cs_registers_i/_1071_ ),
    .Y(\cs_registers_i/_1072_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3541_  (.Y(\cs_registers_i/_1073_ ),
    .B1(net1132),
    .B2(\cs_registers_i/mscratch_q_25_ ),
    .A2(net1116),
    .A1(\cs_registers_i/mtval_q_25_ ));
 sg13g2_nor2_1 \cs_registers_i/_3542_  (.A(net1193),
    .B(\cs_registers_i/_1073_ ),
    .Y(\cs_registers_i/_1074_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3543_  (.B1(net1148),
    .Y(\cs_registers_i/_1075_ ),
    .A1(\cs_registers_i/_1072_ ),
    .A2(\cs_registers_i/_1074_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3544_  (.B1(\cs_registers_i/_1075_ ),
    .Y(\cs_registers_i/_1076_ ),
    .A1(\cs_registers_i/_1068_ ),
    .A2(\cs_registers_i/_1070_ ));
 sg13g2_nor3_2 \cs_registers_i/_3545_  (.A(\cs_registers_i/_1059_ ),
    .B(\cs_registers_i/_1067_ ),
    .C(\cs_registers_i/_1076_ ),
    .Y(\cs_registers_i/_1077_ ));
 sg13g2_nor3_1 \cs_registers_i/_3546_  (.A(net1202),
    .B(net1093),
    .C(\cs_registers_i/_1077_ ),
    .Y(\cs_registers_i/_1078_ ));
 sg13g2_a21o_2 \cs_registers_i/_3547_  (.A2(net259),
    .A1(alu_operand_a_ex_25_),
    .B1(\cs_registers_i/_1078_ ),
    .X(\cs_registers_i/_1079_ ));
 sg13g2_buf_2 fanout555 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0_ ),
    .X(net555));
 sg13g2_a22oi_1 \cs_registers_i/_3549_  (.Y(\cs_registers_i/_1081_ ),
    .B1(net1043),
    .B2(net656),
    .A2(\cs_registers_i/_1056_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3550_  (.Y(\cs_registers_i/_0027_ ),
    .A(\cs_registers_i/_1055_ ),
    .B(\cs_registers_i/_1081_ ));
 sg13g2_nand2_1 \cs_registers_i/_3551_  (.Y(\cs_registers_i/_1082_ ),
    .A(csr_depc_26_),
    .B(net662));
 sg13g2_buf_4 fanout554 (.X(net554),
    .A(net555));
 sg13g2_mux2_2 \cs_registers_i/_3553_  (.A0(crash_dump_o_122_),
    .A1(crash_dump_o_90_),
    .S(net1479),
    .X(\cs_registers_i/_1084_ ));
 sg13g2_mux2_1 \cs_registers_i/_3554_  (.A0(\cs_registers_i/mie_q_10_ ),
    .A1(csr_mtvec_26_),
    .S(net1239),
    .X(\cs_registers_i/_1085_ ));
 sg13g2_nand3_1 \cs_registers_i/_3555_  (.B(net1094),
    .C(\cs_registers_i/_1085_ ),
    .A(net57),
    .Y(\cs_registers_i/_1086_ ));
 sg13g2_mux2_1 \cs_registers_i/_3556_  (.A0(\cs_registers_i/dcsr_q_26_ ),
    .A1(csr_depc_26_),
    .S(net1240),
    .X(\cs_registers_i/_1087_ ));
 sg13g2_nand3_1 \cs_registers_i/_3557_  (.B(net1151),
    .C(\cs_registers_i/_1087_ ),
    .A(\cs_registers_i/_0773_ ),
    .Y(\cs_registers_i/_1088_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3558_  (.Y(\cs_registers_i/_1089_ ),
    .B1(\cs_registers_i/_1061_ ),
    .B2(\cs_registers_i/dscratch0_q_26_ ),
    .A2(\cs_registers_i/_0948_ ),
    .A1(\cs_registers_i/dscratch1_q_26_ ));
 sg13g2_inv_1 \cs_registers_i/_3559_  (.Y(\cs_registers_i/_1090_ ),
    .A(\cs_registers_i/_1089_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3560_  (.Y(\cs_registers_i/_1091_ ),
    .B1(\cs_registers_i/_1090_ ),
    .B2(net60),
    .A2(net1097),
    .A1(hart_id_i_26_));
 sg13g2_a22oi_1 \cs_registers_i/_3561_  (.Y(\cs_registers_i/_1092_ ),
    .B1(net1132),
    .B2(\cs_registers_i/mscratch_q_26_ ),
    .A2(net1116),
    .A1(\cs_registers_i/mtval_q_26_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3562_  (.Y(\cs_registers_i/_1093_ ),
    .B1(net1155),
    .B2(irq_fast_i_10_),
    .A2(net1173),
    .A1(crash_dump_o_26_));
 sg13g2_or2_1 \cs_registers_i/_3563_  (.X(\cs_registers_i/_1094_ ),
    .B(\cs_registers_i/_1093_ ),
    .A(net1100));
 sg13g2_o21ai_1 \cs_registers_i/_3564_  (.B1(\cs_registers_i/_1094_ ),
    .Y(\cs_registers_i/_1095_ ),
    .A1(net1193),
    .A2(\cs_registers_i/_1092_ ));
 sg13g2_mux4_1 \cs_registers_i/_3565_  (.S0(net66),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_26_ ),
    .A1(\cs_registers_i/mhpmcounter_1882_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_58_ ),
    .A3(\cs_registers_i/mhpmcounter_1914_ ),
    .S1(net147),
    .X(\cs_registers_i/_1096_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3566_  (.B2(\cs_registers_i/_0877_ ),
    .C1(\cs_registers_i/_0649_ ),
    .B1(\cs_registers_i/_1096_ ),
    .A1(net1148),
    .Y(\cs_registers_i/_1097_ ),
    .A2(\cs_registers_i/_1095_ ));
 sg13g2_and4_2 \cs_registers_i/_3567_  (.A(\cs_registers_i/_1086_ ),
    .B(\cs_registers_i/_1088_ ),
    .C(\cs_registers_i/_1091_ ),
    .D(\cs_registers_i/_1097_ ),
    .X(\cs_registers_i/_1098_ ));
 sg13g2_nor3_1 \cs_registers_i/_3568_  (.A(net87),
    .B(net1089),
    .C(\cs_registers_i/_1098_ ),
    .Y(\cs_registers_i/_1099_ ));
 sg13g2_a21o_2 \cs_registers_i/_3569_  (.A2(net259),
    .A1(net88),
    .B1(\cs_registers_i/_1099_ ),
    .X(\cs_registers_i/_1100_ ));
 sg13g2_buf_4 fanout553 (.X(net553),
    .A(\id_stage_i.controller_i.instr_i_11_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3571_  (.Y(\cs_registers_i/_1102_ ),
    .B1(net1066),
    .B2(net656),
    .A2(\cs_registers_i/_1084_ ),
    .A1(net1312));
 sg13g2_nand2_1 \cs_registers_i/_3572_  (.Y(\cs_registers_i/_0028_ ),
    .A(\cs_registers_i/_1082_ ),
    .B(\cs_registers_i/_1102_ ));
 sg13g2_nand2_1 \cs_registers_i/_3573_  (.Y(\cs_registers_i/_1103_ ),
    .A(csr_depc_27_),
    .B(net660));
 sg13g2_mux2_2 \cs_registers_i/_3574_  (.A0(crash_dump_o_123_),
    .A1(crash_dump_o_91_),
    .S(net1479),
    .X(\cs_registers_i/_1104_ ));
 sg13g2_nand2_1 \cs_registers_i/_3575_  (.Y(\cs_registers_i/_1105_ ),
    .A(\cs_registers_i/dcsr_q_27_ ),
    .B(net59));
 sg13g2_a21oi_1 \cs_registers_i/_3576_  (.A1(\cs_registers_i/_0648_ ),
    .A2(\cs_registers_i/_1105_ ),
    .Y(\cs_registers_i/_1106_ ),
    .B1(\cs_registers_i/_0506_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3577_  (.Y(\cs_registers_i/_1107_ ),
    .B1(\cs_registers_i/_0598_ ),
    .B2(csr_mtvec_27_),
    .A2(\cs_registers_i/_0519_ ),
    .A1(\cs_registers_i/mie_q_11_ ));
 sg13g2_inv_1 \cs_registers_i/_3578_  (.Y(\cs_registers_i/_1108_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_27_ ));
 sg13g2_nand2_1 \cs_registers_i/_3579_  (.Y(\cs_registers_i/_1109_ ),
    .A(net77),
    .B(\cs_registers_i/mhpmcounter_1883_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3580_  (.B1(\cs_registers_i/_1109_ ),
    .Y(\cs_registers_i/_1110_ ),
    .A1(net73),
    .A2(\cs_registers_i/_1108_ ));
 sg13g2_nand2_1 \cs_registers_i/_3581_  (.Y(\cs_registers_i/_1111_ ),
    .A(\cs_registers_i/_0628_ ),
    .B(\cs_registers_i/_1110_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3582_  (.B1(\cs_registers_i/_1111_ ),
    .Y(\cs_registers_i/_1112_ ),
    .A1(\cs_registers_i/_0946_ ),
    .A2(\cs_registers_i/_1107_ ));
 sg13g2_inv_1 \cs_registers_i/_3583_  (.Y(\cs_registers_i/_1113_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_59_ ));
 sg13g2_nand2_1 \cs_registers_i/_3584_  (.Y(\cs_registers_i/_1114_ ),
    .A(net77),
    .B(\cs_registers_i/mhpmcounter_1915_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3585_  (.B1(\cs_registers_i/_1114_ ),
    .Y(\cs_registers_i/_1115_ ),
    .A1(net67),
    .A2(\cs_registers_i/_1113_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3586_  (.Y(\cs_registers_i/_1116_ ),
    .B1(\cs_registers_i/_1115_ ),
    .B2(net1130),
    .A2(net1098),
    .A1(hart_id_i_27_));
 sg13g2_inv_1 \cs_registers_i/_3587_  (.Y(\cs_registers_i/_1117_ ),
    .A(\cs_registers_i/_1116_ ));
 sg13g2_mux2_1 \cs_registers_i/_3588_  (.A0(\cs_registers_i/dscratch0_q_27_ ),
    .A1(\cs_registers_i/dscratch1_q_27_ ),
    .S(net1243),
    .X(\cs_registers_i/_1118_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3589_  (.Y(\cs_registers_i/_1119_ ),
    .B1(\cs_registers_i/_1118_ ),
    .B2(net75),
    .A2(\cs_registers_i/_0717_ ),
    .A1(csr_depc_27_));
 sg13g2_a22oi_1 \cs_registers_i/_3590_  (.Y(\cs_registers_i/_1120_ ),
    .B1(net1155),
    .B2(irq_fast_i_11_),
    .A2(net1173),
    .A1(crash_dump_o_27_));
 sg13g2_nor2_1 \cs_registers_i/_3591_  (.A(net1101),
    .B(\cs_registers_i/_1120_ ),
    .Y(\cs_registers_i/_1121_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3592_  (.Y(\cs_registers_i/_1122_ ),
    .B1(net1131),
    .B2(\cs_registers_i/mscratch_q_27_ ),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_27_ ));
 sg13g2_nor2_1 \cs_registers_i/_3593_  (.A(net1193),
    .B(\cs_registers_i/_1122_ ),
    .Y(\cs_registers_i/_1123_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3594_  (.B1(net1148),
    .Y(\cs_registers_i/_1124_ ),
    .A1(\cs_registers_i/_1121_ ),
    .A2(\cs_registers_i/_1123_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3595_  (.B1(\cs_registers_i/_1124_ ),
    .Y(\cs_registers_i/_1125_ ),
    .A1(\cs_registers_i/_0912_ ),
    .A2(\cs_registers_i/_1119_ ));
 sg13g2_nor4_2 \cs_registers_i/_3596_  (.A(\cs_registers_i/_1106_ ),
    .B(\cs_registers_i/_1112_ ),
    .C(\cs_registers_i/_1117_ ),
    .Y(\cs_registers_i/_1126_ ),
    .D(\cs_registers_i/_1125_ ));
 sg13g2_nor3_1 \cs_registers_i/_3597_  (.A(net122),
    .B(net1090),
    .C(\cs_registers_i/_1126_ ),
    .Y(\cs_registers_i/_1127_ ));
 sg13g2_a21o_2 \cs_registers_i/_3598_  (.A2(net261),
    .A1(net124),
    .B1(\cs_registers_i/_1127_ ),
    .X(\cs_registers_i/_1128_ ));
 sg13g2_buf_1 fanout552 (.A(\id_stage_i.controller_i.instr_i_13_ ),
    .X(net552));
 sg13g2_a22oi_1 \cs_registers_i/_3600_  (.Y(\cs_registers_i/_1130_ ),
    .B1(net1026),
    .B2(net655),
    .A2(\cs_registers_i/_1104_ ),
    .A1(net1310));
 sg13g2_nand2_1 \cs_registers_i/_3601_  (.Y(\cs_registers_i/_0029_ ),
    .A(\cs_registers_i/_1103_ ),
    .B(\cs_registers_i/_1130_ ));
 sg13g2_nand2_1 \cs_registers_i/_3602_  (.Y(\cs_registers_i/_1131_ ),
    .A(csr_depc_28_),
    .B(net660));
 sg13g2_mux2_2 \cs_registers_i/_3603_  (.A0(crash_dump_o_124_),
    .A1(crash_dump_o_92_),
    .S(net1482),
    .X(\cs_registers_i/_1132_ ));
 sg13g2_and2_1 \cs_registers_i/_3604_  (.A(csr_depc_28_),
    .B(net1234),
    .X(\cs_registers_i/_1133_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3605_  (.A1(net55),
    .A2(\cs_registers_i/dcsr_q_28_ ),
    .Y(\cs_registers_i/_1134_ ),
    .B1(\cs_registers_i/_1133_ ));
 sg13g2_nor3_1 \cs_registers_i/_3606_  (.A(net72),
    .B(\cs_registers_i/_0912_ ),
    .C(\cs_registers_i/_1134_ ),
    .Y(\cs_registers_i/_1135_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3607_  (.Y(\cs_registers_i/_1136_ ),
    .B1(\cs_registers_i/_1061_ ),
    .B2(\cs_registers_i/dscratch0_q_28_ ),
    .A2(\cs_registers_i/_0948_ ),
    .A1(\cs_registers_i/dscratch1_q_28_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3608_  (.Y(\cs_registers_i/_1137_ ),
    .B(net59),
    .A_N(\cs_registers_i/_1136_ ));
 sg13g2_nand2_1 \cs_registers_i/_3609_  (.Y(\cs_registers_i/_1138_ ),
    .A(hart_id_i_28_),
    .B(net1097));
 sg13g2_mux4_1 \cs_registers_i/_3610_  (.S0(net66),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .A1(\cs_registers_i/mhpmcounter_1884_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_60_ ),
    .A3(\cs_registers_i/mhpmcounter_1916_ ),
    .S1(net147),
    .X(\cs_registers_i/_1139_ ));
 sg13g2_nand2_1 \cs_registers_i/_3611_  (.Y(\cs_registers_i/_1140_ ),
    .A(\cs_registers_i/_0877_ ),
    .B(\cs_registers_i/_1139_ ));
 sg13g2_nand4_1 \cs_registers_i/_3612_  (.B(\cs_registers_i/_1137_ ),
    .C(\cs_registers_i/_1138_ ),
    .A(\cs_registers_i/_1060_ ),
    .Y(\cs_registers_i/_1141_ ),
    .D(\cs_registers_i/_1140_ ));
 sg13g2_and2_1 \cs_registers_i/_3613_  (.A(csr_mtvec_28_),
    .B(net1239),
    .X(\cs_registers_i/_1142_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3614_  (.A1(net55),
    .A2(\cs_registers_i/mie_q_12_ ),
    .Y(\cs_registers_i/_1143_ ),
    .B1(\cs_registers_i/_1142_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3615_  (.Y(\cs_registers_i/_1144_ ),
    .B1(net1155),
    .B2(irq_fast_i_12_),
    .A2(net1173),
    .A1(crash_dump_o_28_));
 sg13g2_nor2_1 \cs_registers_i/_3616_  (.A(net1100),
    .B(\cs_registers_i/_1144_ ),
    .Y(\cs_registers_i/_1145_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3617_  (.Y(\cs_registers_i/_1146_ ),
    .B1(net1131),
    .B2(\cs_registers_i/mscratch_q_28_ ),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_28_ ));
 sg13g2_nor2_1 \cs_registers_i/_3618_  (.A(net1193),
    .B(\cs_registers_i/_1146_ ),
    .Y(\cs_registers_i/_1147_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3619_  (.B1(net1148),
    .Y(\cs_registers_i/_1148_ ),
    .A1(\cs_registers_i/_1145_ ),
    .A2(\cs_registers_i/_1147_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3620_  (.B1(\cs_registers_i/_1148_ ),
    .Y(\cs_registers_i/_1149_ ),
    .A1(\cs_registers_i/_1068_ ),
    .A2(\cs_registers_i/_1143_ ));
 sg13g2_nor3_2 \cs_registers_i/_3621_  (.A(\cs_registers_i/_1135_ ),
    .B(\cs_registers_i/_1141_ ),
    .C(\cs_registers_i/_1149_ ),
    .Y(\cs_registers_i/_1150_ ));
 sg13g2_nor3_1 \cs_registers_i/_3622_  (.A(net1201),
    .B(net1090),
    .C(\cs_registers_i/_1150_ ),
    .Y(\cs_registers_i/_1151_ ));
 sg13g2_a21o_2 \cs_registers_i/_3623_  (.A2(net261),
    .A1(net1201),
    .B1(\cs_registers_i/_1151_ ),
    .X(\cs_registers_i/_1152_ ));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_a22oi_1 \cs_registers_i/_3625_  (.Y(\cs_registers_i/_1154_ ),
    .B1(net1042),
    .B2(net655),
    .A2(\cs_registers_i/_1132_ ),
    .A1(net1310));
 sg13g2_nand2_1 \cs_registers_i/_3626_  (.Y(\cs_registers_i/_0030_ ),
    .A(\cs_registers_i/_1131_ ),
    .B(\cs_registers_i/_1154_ ));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_nand2_1 \cs_registers_i/_3628_  (.Y(\cs_registers_i/_1156_ ),
    .A(csr_depc_29_),
    .B(net663));
 sg13g2_mux2_2 \cs_registers_i/_3629_  (.A0(crash_dump_o_125_),
    .A1(crash_dump_o_93_),
    .S(net1479),
    .X(\cs_registers_i/_1157_ ));
 sg13g2_mux2_1 \cs_registers_i/_3630_  (.A0(\cs_registers_i/mie_q_13_ ),
    .A1(csr_mtvec_29_),
    .S(net1239),
    .X(\cs_registers_i/_1158_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3631_  (.A1(net1094),
    .A2(\cs_registers_i/_1158_ ),
    .Y(\cs_registers_i/_1159_ ),
    .B1(net1118));
 sg13g2_nand2b_1 \cs_registers_i/_3632_  (.Y(\cs_registers_i/_1160_ ),
    .B(net57),
    .A_N(\cs_registers_i/_1159_ ));
 sg13g2_nand3_1 \cs_registers_i/_3633_  (.B(net59),
    .C(\cs_registers_i/_1061_ ),
    .A(\cs_registers_i/dscratch0_q_29_ ),
    .Y(\cs_registers_i/_1161_ ));
 sg13g2_nand2_1 \cs_registers_i/_3634_  (.Y(\cs_registers_i/_1162_ ),
    .A(hart_id_i_29_),
    .B(net1098));
 sg13g2_mux2_1 \cs_registers_i/_3635_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_29_ ),
    .A1(\cs_registers_i/mhpmcounter_1885_ ),
    .S(net64),
    .X(\cs_registers_i/_1163_ ));
 sg13g2_mux2_1 \cs_registers_i/_3636_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_61_ ),
    .A1(\cs_registers_i/mhpmcounter_1917_ ),
    .S(net64),
    .X(\cs_registers_i/_1164_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3637_  (.Y(\cs_registers_i/_1165_ ),
    .B1(\cs_registers_i/_1164_ ),
    .B2(net1156),
    .A2(\cs_registers_i/_1163_ ),
    .A1(net1191));
 sg13g2_or2_1 \cs_registers_i/_3638_  (.X(\cs_registers_i/_1166_ ),
    .B(\cs_registers_i/_1165_ ),
    .A(net1159));
 sg13g2_and2_1 \cs_registers_i/_3639_  (.A(csr_depc_29_),
    .B(net1240),
    .X(\cs_registers_i/_1167_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3640_  (.B1(\cs_registers_i/_1167_ ),
    .Y(\cs_registers_i/_1168_ ),
    .A2(\cs_registers_i/dcsr_q_29_ ),
    .A1(net53));
 sg13g2_nand3_1 \cs_registers_i/_3641_  (.B(net1235),
    .C(\cs_registers_i/dscratch1_q_29_ ),
    .A(net75),
    .Y(\cs_registers_i/_1169_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3642_  (.B1(\cs_registers_i/_1169_ ),
    .Y(\cs_registers_i/_1170_ ),
    .A1(net69),
    .A2(\cs_registers_i/_1168_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3643_  (.Y(\cs_registers_i/_1171_ ),
    .B1(net1131),
    .B2(\cs_registers_i/mscratch_q_29_ ),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_29_ ));
 sg13g2_nand3b_1 \cs_registers_i/_3644_  (.B(irq_fast_i_13_),
    .C(net101),
    .Y(\cs_registers_i/_1172_ ),
    .A_N(net1242));
 sg13g2_nand3b_1 \cs_registers_i/_3645_  (.B(net1238),
    .C(crash_dump_o_29_),
    .Y(\cs_registers_i/_1173_ ),
    .A_N(net99));
 sg13g2_a21o_1 \cs_registers_i/_3646_  (.A2(\cs_registers_i/_1173_ ),
    .A1(\cs_registers_i/_1172_ ),
    .B1(net1100),
    .X(\cs_registers_i/_1174_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3647_  (.B1(\cs_registers_i/_1174_ ),
    .Y(\cs_registers_i/_1175_ ),
    .A1(net1192),
    .A2(\cs_registers_i/_1171_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3648_  (.Y(\cs_registers_i/_1176_ ),
    .B1(\cs_registers_i/_1175_ ),
    .B2(net1149),
    .A2(\cs_registers_i/_1170_ ),
    .A1(net1152));
 sg13g2_and4_1 \cs_registers_i/_3649_  (.A(\cs_registers_i/_1161_ ),
    .B(\cs_registers_i/_1162_ ),
    .C(\cs_registers_i/_1166_ ),
    .D(\cs_registers_i/_1176_ ),
    .X(\cs_registers_i/_1177_ ));
 sg13g2_nor2_2 \cs_registers_i/_3650_  (.A(\cs_registers_i/_0522_ ),
    .B(\cs_registers_i/_0540_ ),
    .Y(\cs_registers_i/_1178_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3651_  (.B1(\cs_registers_i/_1178_ ),
    .Y(csr_rdata_29_),
    .A2(\cs_registers_i/_1177_ ),
    .A1(\cs_registers_i/_1160_ ));
 sg13g2_nand2_1 \cs_registers_i/_3652_  (.Y(\cs_registers_i/_1179_ ),
    .A(csr_op_1_),
    .B(csr_rdata_29_));
 sg13g2_nand2_1 \cs_registers_i/_3653_  (.Y(\cs_registers_i/_1180_ ),
    .A(net1198),
    .B(net263));
 sg13g2_o21ai_1 \cs_registers_i/_3654_  (.B1(\cs_registers_i/_1180_ ),
    .Y(\cs_registers_i/_1181_ ),
    .A1(net1198),
    .A2(\cs_registers_i/_1179_ ));
 sg13g2_buf_4 fanout549 (.X(net549),
    .A(net552));
 sg13g2_buf_2 fanout548 (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .X(net548));
 sg13g2_a22oi_1 \cs_registers_i/_3657_  (.Y(\cs_registers_i/_1184_ ),
    .B1(net1040),
    .B2(net657),
    .A2(\cs_registers_i/_1157_ ),
    .A1(net1314));
 sg13g2_nand2_1 \cs_registers_i/_3658_  (.Y(\cs_registers_i/_0031_ ),
    .A(\cs_registers_i/_1156_ ),
    .B(\cs_registers_i/_1184_ ));
 sg13g2_nand2_1 \cs_registers_i/_3659_  (.Y(\cs_registers_i/_1185_ ),
    .A(csr_depc_2_),
    .B(net662));
 sg13g2_mux2_2 \cs_registers_i/_3660_  (.A0(crash_dump_o_98_),
    .A1(crash_dump_o_66_),
    .S(net1481),
    .X(\cs_registers_i/_1186_ ));
 sg13g2_inv_1 \cs_registers_i/_3661_  (.Y(\cs_registers_i/_1187_ ),
    .A(\cs_registers_i/_0673_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3662_  (.Y(\cs_registers_i/_1188_ ),
    .B1(\cs_registers_i/_0669_ ),
    .B2(\cs_registers_i/mscratch_q_2_ ),
    .A2(\cs_registers_i/_0670_ ),
    .A1(\cs_registers_i/mcountinhibit_2_ ));
 sg13g2_a21o_1 \cs_registers_i/_3663_  (.A2(\cs_registers_i/_0598_ ),
    .A1(csr_mtvec_2_),
    .B1(\cs_registers_i/_0477_ ),
    .X(\cs_registers_i/_1189_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3664_  (.Y(\cs_registers_i/_1190_ ),
    .B1(\cs_registers_i/_0549_ ),
    .B2(\cs_registers_i/mcause_q_2_ ),
    .A2(\cs_registers_i/_0717_ ),
    .A1(crash_dump_o_2_));
 sg13g2_nor2b_1 \cs_registers_i/_3665_  (.A(\cs_registers_i/_1190_ ),
    .B_N(net1160),
    .Y(\cs_registers_i/_1191_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3666_  (.B2(\cs_registers_i/_0720_ ),
    .C1(\cs_registers_i/_1191_ ),
    .B1(\cs_registers_i/_1189_ ),
    .A1(\cs_registers_i/mtval_q_2_ ),
    .Y(\cs_registers_i/_1192_ ),
    .A2(\cs_registers_i/_0678_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3667_  (.B1(\cs_registers_i/_1192_ ),
    .Y(\cs_registers_i/_1193_ ),
    .A1(\cs_registers_i/_1187_ ),
    .A2(\cs_registers_i/_1188_ ));
 sg13g2_mux4_1 \cs_registers_i/_3668_  (.S0(net67),
    .A0(debug_single_step),
    .A1(\cs_registers_i/dscratch0_q_2_ ),
    .A2(csr_depc_2_),
    .A3(\cs_registers_i/dscratch1_q_2_ ),
    .S1(net1241),
    .X(\cs_registers_i/_1194_ ));
 sg13g2_inv_1 \cs_registers_i/_3669_  (.Y(\cs_registers_i/_1195_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_2_ ));
 sg13g2_nor2_1 \cs_registers_i/_3670_  (.A(net68),
    .B(\cs_registers_i/_1195_ ),
    .Y(\cs_registers_i/_1196_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3671_  (.A1(net75),
    .A2(\cs_registers_i/mhpmcounter_1858_ ),
    .Y(\cs_registers_i/_1197_ ),
    .B1(\cs_registers_i/_1196_ ));
 sg13g2_mux2_1 \cs_registers_i/_3672_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .A1(\cs_registers_i/mhpmcounter_1890_ ),
    .S(net63),
    .X(\cs_registers_i/_1198_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3673_  (.Y(\cs_registers_i/_1199_ ),
    .B1(\cs_registers_i/_1198_ ),
    .B2(net1129),
    .A2(net1095),
    .A1(hart_id_i_2_));
 sg13g2_o21ai_1 \cs_registers_i/_3674_  (.B1(\cs_registers_i/_1199_ ),
    .Y(\cs_registers_i/_1200_ ),
    .A1(\cs_registers_i/_0895_ ),
    .A2(\cs_registers_i/_1197_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3675_  (.B2(net1154),
    .C1(\cs_registers_i/_1200_ ),
    .B1(\cs_registers_i/_1194_ ),
    .A1(net57),
    .Y(\cs_registers_i/_1201_ ),
    .A2(\cs_registers_i/_1193_ ));
 sg13g2_nor3_1 \cs_registers_i/_3676_  (.A(net1410),
    .B(net1093),
    .C(\cs_registers_i/_1201_ ),
    .Y(\cs_registers_i/_1202_ ));
 sg13g2_a21o_1 \cs_registers_i/_3677_  (.A2(net261),
    .A1(net1410),
    .B1(\cs_registers_i/_1202_ ),
    .X(\cs_registers_i/_1203_ ));
 sg13g2_buf_2 fanout547 (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .X(net547));
 sg13g2_a22oi_1 \cs_registers_i/_3679_  (.Y(\cs_registers_i/_1205_ ),
    .B1(net1039),
    .B2(net656),
    .A2(\cs_registers_i/_1186_ ),
    .A1(net1312));
 sg13g2_nand2_1 \cs_registers_i/_3680_  (.Y(\cs_registers_i/_0032_ ),
    .A(\cs_registers_i/_1185_ ),
    .B(\cs_registers_i/_1205_ ));
 sg13g2_nand2_1 \cs_registers_i/_3681_  (.Y(\cs_registers_i/_1206_ ),
    .A(csr_depc_30_),
    .B(net661));
 sg13g2_mux2_2 \cs_registers_i/_3682_  (.A0(crash_dump_o_126_),
    .A1(crash_dump_o_94_),
    .S(net1479),
    .X(\cs_registers_i/_1207_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3683_  (.A(net1086),
    .B_N(csr_op_1_),
    .Y(\cs_registers_i/_1208_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3684_  (.Y(\cs_registers_i/_1209_ ),
    .B1(\cs_registers_i/_0842_ ),
    .B2(\cs_registers_i/mtval_q_30_ ),
    .A2(\cs_registers_i/_0819_ ),
    .A1(irq_fast_i_14_));
 sg13g2_nor2_1 \cs_registers_i/_3685_  (.A(net1276),
    .B(\cs_registers_i/_1209_ ),
    .Y(\cs_registers_i/_1210_ ));
 sg13g2_and2_1 \cs_registers_i/_3686_  (.A(crash_dump_o_30_),
    .B(net1241),
    .X(\cs_registers_i/_1211_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3687_  (.A1(net54),
    .A2(\cs_registers_i/mscratch_q_30_ ),
    .Y(\cs_registers_i/_1212_ ),
    .B1(\cs_registers_i/_1211_ ));
 sg13g2_nor3_1 \cs_registers_i/_3688_  (.A(net72),
    .B(net1193),
    .C(\cs_registers_i/_1212_ ),
    .Y(\cs_registers_i/_1213_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3689_  (.B1(net1149),
    .Y(\cs_registers_i/_1214_ ),
    .A1(\cs_registers_i/_1210_ ),
    .A2(\cs_registers_i/_1213_ ));
 sg13g2_mux4_1 \cs_registers_i/_3690_  (.S0(net68),
    .A0(\cs_registers_i/dcsr_q_30_ ),
    .A1(\cs_registers_i/dscratch0_q_30_ ),
    .A2(csr_depc_30_),
    .A3(\cs_registers_i/dscratch1_q_30_ ),
    .S1(net1243),
    .X(\cs_registers_i/_1215_ ));
 sg13g2_nand2_1 \cs_registers_i/_3691_  (.Y(\cs_registers_i/_1216_ ),
    .A(net1153),
    .B(\cs_registers_i/_1215_ ));
 sg13g2_mux4_1 \cs_registers_i/_3692_  (.S0(net71),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_30_ ),
    .A1(\cs_registers_i/mhpmcounter_1886_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_62_ ),
    .A3(\cs_registers_i/mhpmcounter_1918_ ),
    .S1(net147),
    .X(\cs_registers_i/_1217_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3693_  (.Y(\cs_registers_i/_1218_ ),
    .B1(\cs_registers_i/_0598_ ),
    .B2(csr_mtvec_30_),
    .A2(net40),
    .A1(\cs_registers_i/mie_q_14_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3694_  (.B1(\cs_registers_i/_0511_ ),
    .Y(\cs_registers_i/_1219_ ),
    .A1(\cs_registers_i/_0946_ ),
    .A2(\cs_registers_i/_1218_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3695_  (.B2(\cs_registers_i/_1217_ ),
    .C1(\cs_registers_i/_1219_ ),
    .B1(\cs_registers_i/_0877_ ),
    .A1(hart_id_i_30_),
    .Y(\cs_registers_i/_1220_ ),
    .A2(net1097));
 sg13g2_nand3_1 \cs_registers_i/_3696_  (.B(\cs_registers_i/_1216_ ),
    .C(\cs_registers_i/_1220_ ),
    .A(\cs_registers_i/_1214_ ),
    .Y(\cs_registers_i/_1221_ ));
 sg13g2_nand2_1 \cs_registers_i/_3697_  (.Y(\cs_registers_i/_1222_ ),
    .A(\cs_registers_i/_1208_ ),
    .B(\cs_registers_i/_1221_ ));
 sg13g2_nand2_1 \cs_registers_i/_3698_  (.Y(\cs_registers_i/_1223_ ),
    .A(net1190),
    .B(net263));
 sg13g2_o21ai_1 \cs_registers_i/_3699_  (.B1(\cs_registers_i/_1223_ ),
    .Y(\cs_registers_i/_1224_ ),
    .A1(alu_operand_a_ex_30_),
    .A2(\cs_registers_i/_1222_ ));
 sg13g2_buf_4 fanout546 (.X(net546),
    .A(\id_stage_i.controller_i.instr_i_16_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3701_  (.Y(\cs_registers_i/_1226_ ),
    .B1(net1037),
    .B2(net657),
    .A2(\cs_registers_i/_1207_ ),
    .A1(net1310));
 sg13g2_nand2_1 \cs_registers_i/_3702_  (.Y(\cs_registers_i/_0033_ ),
    .A(\cs_registers_i/_1206_ ),
    .B(\cs_registers_i/_1226_ ));
 sg13g2_nand2_1 \cs_registers_i/_3703_  (.Y(\cs_registers_i/_1227_ ),
    .A(csr_depc_31_),
    .B(net663));
 sg13g2_mux2_2 \cs_registers_i/_3704_  (.A0(crash_dump_o_127_),
    .A1(crash_dump_o_95_),
    .S(net1479),
    .X(\cs_registers_i/_1228_ ));
 sg13g2_mux4_1 \cs_registers_i/_3705_  (.S0(net67),
    .A0(\cs_registers_i/dcsr_q_31_ ),
    .A1(\cs_registers_i/dscratch0_q_31_ ),
    .A2(csr_depc_31_),
    .A3(\cs_registers_i/dscratch1_q_31_ ),
    .S1(net1241),
    .X(\cs_registers_i/_1229_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3706_  (.Y(\cs_registers_i/_1230_ ),
    .B1(net1155),
    .B2(irq_fast_i_15_),
    .A2(net1173),
    .A1(crash_dump_o_31_));
 sg13g2_nor2b_1 \cs_registers_i/_3707_  (.A(net1231),
    .B_N(\cs_registers_i/mcause_q_6_ ),
    .Y(\cs_registers_i/_1231_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3708_  (.A1(net1234),
    .A2(\cs_registers_i/mtval_q_31_ ),
    .Y(\cs_registers_i/_1232_ ),
    .B1(\cs_registers_i/_1231_ ));
 sg13g2_nand3_1 \cs_registers_i/_3709_  (.B(net53),
    .C(\cs_registers_i/mscratch_q_31_ ),
    .A(net1114),
    .Y(\cs_registers_i/_1233_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3710_  (.B1(\cs_registers_i/_1233_ ),
    .Y(\cs_registers_i/_1234_ ),
    .A1(net1114),
    .A2(\cs_registers_i/_1232_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3711_  (.A1(net1160),
    .A2(\cs_registers_i/_1234_ ),
    .Y(\cs_registers_i/_1235_ ),
    .B1(net1118));
 sg13g2_o21ai_1 \cs_registers_i/_3712_  (.B1(\cs_registers_i/_1235_ ),
    .Y(\cs_registers_i/_1236_ ),
    .A1(\cs_registers_i/_0675_ ),
    .A2(\cs_registers_i/_1230_ ));
 sg13g2_and2_1 \cs_registers_i/_3713_  (.A(csr_mtvec_31_),
    .B(net1239),
    .X(\cs_registers_i/_1237_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3714_  (.A1(net54),
    .A2(\cs_registers_i/mie_q_15_ ),
    .Y(\cs_registers_i/_1238_ ),
    .B1(\cs_registers_i/_1237_ ));
 sg13g2_mux4_1 \cs_registers_i/_3715_  (.S0(net145),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_31_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_63_ ),
    .A2(\cs_registers_i/mhpmcounter_1887_ ),
    .A3(\cs_registers_i/mhpmcounter_1919_ ),
    .S1(csr_addr_1_),
    .X(\cs_registers_i/_1239_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3716_  (.Y(\cs_registers_i/_1240_ ),
    .B1(\cs_registers_i/_0877_ ),
    .B2(\cs_registers_i/_1239_ ),
    .A2(net1097),
    .A1(hart_id_i_31_));
 sg13g2_o21ai_1 \cs_registers_i/_3717_  (.B1(\cs_registers_i/_1240_ ),
    .Y(\cs_registers_i/_1241_ ),
    .A1(\cs_registers_i/_1068_ ),
    .A2(\cs_registers_i/_1238_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3718_  (.B2(net56),
    .C1(\cs_registers_i/_1241_ ),
    .B1(\cs_registers_i/_1236_ ),
    .A1(net1151),
    .Y(\cs_registers_i/_1242_ ),
    .A2(\cs_registers_i/_1229_ ));
 sg13g2_nor3_1 \cs_registers_i/_3719_  (.A(net81),
    .B(net1089),
    .C(\cs_registers_i/_1242_ ),
    .Y(\cs_registers_i/_1243_ ));
 sg13g2_a21o_2 \cs_registers_i/_3720_  (.A2(net260),
    .A1(net81),
    .B1(\cs_registers_i/_1243_ ),
    .X(\cs_registers_i/_1244_ ));
 sg13g2_buf_4 fanout545 (.X(net545),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3722_  (.Y(\cs_registers_i/_1246_ ),
    .B1(net1035),
    .B2(net657),
    .A2(\cs_registers_i/_1228_ ),
    .A1(net1311));
 sg13g2_nand2_1 \cs_registers_i/_3723_  (.Y(\cs_registers_i/_0034_ ),
    .A(\cs_registers_i/_1227_ ),
    .B(\cs_registers_i/_1246_ ));
 sg13g2_nand2_1 \cs_registers_i/_3724_  (.Y(\cs_registers_i/_1247_ ),
    .A(csr_depc_3_),
    .B(net659));
 sg13g2_mux2_2 \cs_registers_i/_3725_  (.A0(crash_dump_o_99_),
    .A1(crash_dump_o_67_),
    .S(net1481),
    .X(\cs_registers_i/_1248_ ));
 sg13g2_mux4_1 \cs_registers_i/_3726_  (.S0(net71),
    .A0(\cs_registers_i/mscratch_q_3_ ),
    .A1(\cs_registers_i/mcause_q_3_ ),
    .A2(crash_dump_o_3_),
    .A3(\cs_registers_i/mtval_q_3_ ),
    .S1(net1233),
    .X(\cs_registers_i/_1249_ ));
 sg13g2_nand2_1 \cs_registers_i/_3727_  (.Y(\cs_registers_i/_1250_ ),
    .A(net1160),
    .B(\cs_registers_i/_1249_ ));
 sg13g2_nand3_1 \cs_registers_i/_3728_  (.B(net1117),
    .C(\cs_registers_i/_0720_ ),
    .A(csr_mstatus_mie),
    .Y(\cs_registers_i/_1251_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3729_  (.A1(\cs_registers_i/_1250_ ),
    .A2(\cs_registers_i/_1251_ ),
    .Y(\cs_registers_i/_1252_ ),
    .B1(net1172));
 sg13g2_mux2_2 \cs_registers_i/_3730_  (.A0(\cs_registers_i/dscratch0_q_3_ ),
    .A1(\cs_registers_i/dscratch1_q_3_ ),
    .S(net1244),
    .X(\cs_registers_i/_1253_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3731_  (.Y(\cs_registers_i/_1254_ ),
    .B1(\cs_registers_i/_1253_ ),
    .B2(net75),
    .A2(\cs_registers_i/_0717_ ),
    .A1(csr_depc_3_));
 sg13g2_nor2_1 \cs_registers_i/_3732_  (.A(\cs_registers_i/_0912_ ),
    .B(\cs_registers_i/_1254_ ),
    .Y(\cs_registers_i/_1255_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3733_  (.A(net1268),
    .B_N(\cs_registers_i/mie_q_18_ ),
    .Y(\cs_registers_i/_1256_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3734_  (.A1(net1268),
    .A2(irq_software_i),
    .Y(\cs_registers_i/_1257_ ),
    .B1(\cs_registers_i/_1256_ ));
 sg13g2_nor4_1 \cs_registers_i/_3735_  (.A(net145),
    .B(\cs_registers_i/_0542_ ),
    .C(\cs_registers_i/_0557_ ),
    .D(\cs_registers_i/_1257_ ),
    .Y(\cs_registers_i/_1258_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3736_  (.A1(hart_id_i_3_),
    .A2(\cs_registers_i/_0561_ ),
    .Y(\cs_registers_i/_1259_ ),
    .B1(\cs_registers_i/_1258_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3737_  (.A(\cs_registers_i/_1259_ ),
    .B_N(net40),
    .Y(\cs_registers_i/_1260_ ));
 sg13g2_nand3_1 \cs_registers_i/_3738_  (.B(net56),
    .C(\cs_registers_i/_0749_ ),
    .A(csr_mtvec_3_),
    .Y(\cs_registers_i/_1261_ ));
 sg13g2_mux2_1 \cs_registers_i/_3739_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_35_ ),
    .A1(\cs_registers_i/mhpmcounter_1891_ ),
    .S(net65),
    .X(\cs_registers_i/_1262_ ));
 sg13g2_nand2_1 \cs_registers_i/_3740_  (.Y(\cs_registers_i/_1263_ ),
    .A(net1129),
    .B(\cs_registers_i/_1262_ ));
 sg13g2_and2_1 \cs_registers_i/_3741_  (.A(\cs_registers_i/dcsr_q_3_ ),
    .B(net1117),
    .X(\cs_registers_i/_1264_ ));
 sg13g2_inv_1 \cs_registers_i/_3742_  (.Y(\cs_registers_i/_1265_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_3_ ));
 sg13g2_nand2_1 \cs_registers_i/_3743_  (.Y(\cs_registers_i/_1266_ ),
    .A(net76),
    .B(\cs_registers_i/mhpmcounter_1859_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3744_  (.B1(\cs_registers_i/_1266_ ),
    .Y(\cs_registers_i/_1267_ ),
    .A1(net71),
    .A2(\cs_registers_i/_1265_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3745_  (.Y(\cs_registers_i/_1268_ ),
    .B1(\cs_registers_i/_1267_ ),
    .B2(\cs_registers_i/_0628_ ),
    .A2(\cs_registers_i/_1264_ ),
    .A1(net59));
 sg13g2_nand4_1 \cs_registers_i/_3746_  (.B(\cs_registers_i/_1261_ ),
    .C(\cs_registers_i/_1263_ ),
    .A(\cs_registers_i/_1060_ ),
    .Y(\cs_registers_i/_1269_ ),
    .D(\cs_registers_i/_1268_ ));
 sg13g2_nor4_2 \cs_registers_i/_3747_  (.A(\cs_registers_i/_1252_ ),
    .B(\cs_registers_i/_1255_ ),
    .C(\cs_registers_i/_1260_ ),
    .Y(\cs_registers_i/_1270_ ),
    .D(\cs_registers_i/_1269_ ));
 sg13g2_nor3_1 \cs_registers_i/_3748_  (.A(net1408),
    .B(net1088),
    .C(\cs_registers_i/_1270_ ),
    .Y(\cs_registers_i/_1271_ ));
 sg13g2_a21o_2 \cs_registers_i/_3749_  (.A2(net261),
    .A1(alu_operand_a_ex_3_),
    .B1(\cs_registers_i/_1271_ ),
    .X(\cs_registers_i/_1272_ ));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3751_  (.Y(\cs_registers_i/_1274_ ),
    .B1(net1033),
    .B2(net654),
    .A2(\cs_registers_i/_1248_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3752_  (.Y(\cs_registers_i/_0035_ ),
    .A(\cs_registers_i/_1247_ ),
    .B(\cs_registers_i/_1274_ ));
 sg13g2_nand2_1 \cs_registers_i/_3753_  (.Y(\cs_registers_i/_1275_ ),
    .A(csr_depc_4_),
    .B(net659));
 sg13g2_mux2_2 \cs_registers_i/_3754_  (.A0(crash_dump_o_100_),
    .A1(crash_dump_o_68_),
    .S(net1482),
    .X(\cs_registers_i/_1276_ ));
 sg13g2_mux4_1 \cs_registers_i/_3755_  (.S0(net64),
    .A0(\cs_registers_i/dcsr_q_4_ ),
    .A1(\cs_registers_i/dscratch0_q_4_ ),
    .A2(csr_depc_4_),
    .A3(\cs_registers_i/dscratch1_q_4_ ),
    .S1(net1237),
    .X(\cs_registers_i/_1277_ ));
 sg13g2_a21o_1 \cs_registers_i/_3756_  (.A2(\cs_registers_i/_0749_ ),
    .A1(csr_mtvec_4_),
    .B1(net1119),
    .X(\cs_registers_i/_1278_ ));
 sg13g2_nand2_1 \cs_registers_i/_3757_  (.Y(\cs_registers_i/_1279_ ),
    .A(hart_id_i_4_),
    .B(net1096));
 sg13g2_mux4_1 \cs_registers_i/_3758_  (.S0(net62),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .A1(\cs_registers_i/mhpmcounter_1860_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_36_ ),
    .A3(\cs_registers_i/mhpmcounter_1892_ ),
    .S1(net147),
    .X(\cs_registers_i/_1280_ ));
 sg13g2_mux4_1 \cs_registers_i/_3759_  (.S0(net73),
    .A0(\cs_registers_i/mscratch_q_4_ ),
    .A1(\cs_registers_i/mcause_q_4_ ),
    .A2(crash_dump_o_4_),
    .A3(\cs_registers_i/mtval_q_4_ ),
    .S1(net1233),
    .X(\cs_registers_i/_1281_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3760_  (.Y(\cs_registers_i/_1282_ ),
    .B1(\cs_registers_i/_1281_ ),
    .B2(\cs_registers_i/_0605_ ),
    .A2(\cs_registers_i/_1280_ ),
    .A1(\cs_registers_i/_0877_ ));
 sg13g2_nand2_1 \cs_registers_i/_3761_  (.Y(\cs_registers_i/_1283_ ),
    .A(\cs_registers_i/_1279_ ),
    .B(\cs_registers_i/_1282_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3762_  (.B2(net56),
    .C1(\cs_registers_i/_1283_ ),
    .B1(\cs_registers_i/_1278_ ),
    .A1(net1150),
    .Y(\cs_registers_i/_1284_ ),
    .A2(\cs_registers_i/_1277_ ));
 sg13g2_nor3_1 \cs_registers_i/_3763_  (.A(net1407),
    .B(net1088),
    .C(\cs_registers_i/_1284_ ),
    .Y(\cs_registers_i/_1285_ ));
 sg13g2_a21o_2 \cs_registers_i/_3764_  (.A2(net259),
    .A1(net1407),
    .B1(\cs_registers_i/_1285_ ),
    .X(\cs_registers_i/_1286_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3765_  (.Y(\cs_registers_i/_1287_ ),
    .B1(net1032),
    .B2(net654),
    .A2(\cs_registers_i/_1276_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3766_  (.Y(\cs_registers_i/_0036_ ),
    .A(\cs_registers_i/_1275_ ),
    .B(\cs_registers_i/_1287_ ));
 sg13g2_nand2_1 \cs_registers_i/_3767_  (.Y(\cs_registers_i/_1288_ ),
    .A(csr_depc_5_),
    .B(net659));
 sg13g2_mux2_2 \cs_registers_i/_3768_  (.A0(crash_dump_o_101_),
    .A1(crash_dump_o_69_),
    .S(net1481),
    .X(\cs_registers_i/_1289_ ));
 sg13g2_nor2_2 \cs_registers_i/_3769_  (.A(net100),
    .B(net1114),
    .Y(\cs_registers_i/_1290_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3770_  (.A1(hart_id_i_5_),
    .A2(\cs_registers_i/_0818_ ),
    .Y(\cs_registers_i/_1291_ ),
    .B1(\cs_registers_i/_1290_ ));
 sg13g2_nor4_1 \cs_registers_i/_3771_  (.A(net1275),
    .B(net1232),
    .C(\cs_registers_i/_0922_ ),
    .D(\cs_registers_i/_1291_ ),
    .Y(\cs_registers_i/_1292_ ));
 sg13g2_mux4_1 \cs_registers_i/_3772_  (.S0(net71),
    .A0(\cs_registers_i/mscratch_q_5_ ),
    .A1(\cs_registers_i/mcause_q_5_ ),
    .A2(crash_dump_o_5_),
    .A3(\cs_registers_i/mtval_q_5_ ),
    .S1(net1233),
    .X(\cs_registers_i/_1293_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3773_  (.B2(net1160),
    .C1(net1119),
    .B1(\cs_registers_i/_1293_ ),
    .A1(csr_mtvec_5_),
    .Y(\cs_registers_i/_1294_ ),
    .A2(\cs_registers_i/_0749_ ));
 sg13g2_nor2_1 \cs_registers_i/_3774_  (.A(net1172),
    .B(\cs_registers_i/_1294_ ),
    .Y(\cs_registers_i/_1295_ ));
 sg13g2_mux2_1 \cs_registers_i/_3775_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_37_ ),
    .A1(\cs_registers_i/mhpmcounter_1893_ ),
    .S(net65),
    .X(\cs_registers_i/_1296_ ));
 sg13g2_mux2_1 \cs_registers_i/_3776_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_5_ ),
    .A1(\cs_registers_i/mhpmcounter_1861_ ),
    .S(net69),
    .X(\cs_registers_i/_1297_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3777_  (.Y(\cs_registers_i/_1298_ ),
    .B1(\cs_registers_i/_1297_ ),
    .B2(net1191),
    .A2(\cs_registers_i/_1296_ ),
    .A1(net1156));
 sg13g2_mux4_1 \cs_registers_i/_3778_  (.S0(net65),
    .A0(\cs_registers_i/dcsr_q_5_ ),
    .A1(\cs_registers_i/dscratch0_q_5_ ),
    .A2(csr_depc_5_),
    .A3(\cs_registers_i/dscratch1_q_5_ ),
    .S1(net1232),
    .X(\cs_registers_i/_1299_ ));
 sg13g2_nand2_1 \cs_registers_i/_3779_  (.Y(\cs_registers_i/_1300_ ),
    .A(net1150),
    .B(\cs_registers_i/_1299_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3780_  (.B1(\cs_registers_i/_1300_ ),
    .Y(\cs_registers_i/_1301_ ),
    .A1(net1158),
    .A2(\cs_registers_i/_1298_ ));
 sg13g2_nor3_2 \cs_registers_i/_3781_  (.A(\cs_registers_i/_1292_ ),
    .B(\cs_registers_i/_1295_ ),
    .C(\cs_registers_i/_1301_ ),
    .Y(\cs_registers_i/_1302_ ));
 sg13g2_nor3_1 \cs_registers_i/_3782_  (.A(net1405),
    .B(net1088),
    .C(\cs_registers_i/_1302_ ),
    .Y(\cs_registers_i/_1303_ ));
 sg13g2_a21o_2 \cs_registers_i/_3783_  (.A2(net260),
    .A1(net1405),
    .B1(\cs_registers_i/_1303_ ),
    .X(\cs_registers_i/_1304_ ));
 sg13g2_buf_4 fanout543 (.X(net543),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3785_  (.Y(\cs_registers_i/_1306_ ),
    .B1(net1065),
    .B2(net654),
    .A2(\cs_registers_i/_1289_ ),
    .A1(net1308));
 sg13g2_nand2_1 \cs_registers_i/_3786_  (.Y(\cs_registers_i/_0037_ ),
    .A(\cs_registers_i/_1288_ ),
    .B(\cs_registers_i/_1306_ ));
 sg13g2_nand2_1 \cs_registers_i/_3787_  (.Y(\cs_registers_i/_1307_ ),
    .A(csr_depc_6_),
    .B(net660));
 sg13g2_mux2_2 \cs_registers_i/_3788_  (.A0(crash_dump_o_102_),
    .A1(crash_dump_o_70_),
    .S(net1481),
    .X(\cs_registers_i/_1308_ ));
 sg13g2_mux2_1 \cs_registers_i/_3789_  (.A0(\cs_registers_i/mscratch_q_6_ ),
    .A1(crash_dump_o_6_),
    .S(net1231),
    .X(\cs_registers_i/_1309_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3790_  (.Y(\cs_registers_i/_1310_ ),
    .B1(\cs_registers_i/_1309_ ),
    .B2(net1114),
    .A2(net1115),
    .A1(\cs_registers_i/mtval_q_6_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3791_  (.A(\cs_registers_i/_1310_ ),
    .B_N(net1160),
    .Y(\cs_registers_i/_1311_ ));
 sg13g2_a21o_1 \cs_registers_i/_3792_  (.A2(\cs_registers_i/_0749_ ),
    .A1(csr_mtvec_6_),
    .B1(net1119),
    .X(\cs_registers_i/_1312_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3793_  (.B1(net56),
    .Y(\cs_registers_i/_1313_ ),
    .A1(\cs_registers_i/_1311_ ),
    .A2(\cs_registers_i/_1312_ ));
 sg13g2_mux2_1 \cs_registers_i/_3794_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_6_ ),
    .A1(\cs_registers_i/mhpmcounter_1862_ ),
    .S(net66),
    .X(\cs_registers_i/_1314_ ));
 sg13g2_nand2_1 \cs_registers_i/_3795_  (.Y(\cs_registers_i/_1315_ ),
    .A(\cs_registers_i/_0722_ ),
    .B(\cs_registers_i/_1314_ ));
 sg13g2_mux4_1 \cs_registers_i/_3796_  (.S0(net62),
    .A0(\cs_registers_i/dcsr_q_6_ ),
    .A1(\cs_registers_i/dscratch0_q_6_ ),
    .A2(csr_depc_6_),
    .A3(\cs_registers_i/dscratch1_q_6_ ),
    .S1(net1244),
    .X(\cs_registers_i/_1316_ ));
 sg13g2_nand2_1 \cs_registers_i/_3797_  (.Y(\cs_registers_i/_1317_ ),
    .A(net1152),
    .B(\cs_registers_i/_1316_ ));
 sg13g2_mux2_1 \cs_registers_i/_3798_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_38_ ),
    .A1(\cs_registers_i/mhpmcounter_1894_ ),
    .S(net70),
    .X(\cs_registers_i/_1318_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3799_  (.Y(\cs_registers_i/_1319_ ),
    .B1(\cs_registers_i/_1318_ ),
    .B2(net1129),
    .A2(net1095),
    .A1(hart_id_i_6_));
 sg13g2_and4_2 \cs_registers_i/_3800_  (.A(\cs_registers_i/_1313_ ),
    .B(\cs_registers_i/_1315_ ),
    .C(\cs_registers_i/_1317_ ),
    .D(\cs_registers_i/_1319_ ),
    .X(\cs_registers_i/_1320_ ));
 sg13g2_nor3_1 \cs_registers_i/_3801_  (.A(net1350),
    .B(net1090),
    .C(\cs_registers_i/_1320_ ),
    .Y(\cs_registers_i/_1321_ ));
 sg13g2_a21o_2 \cs_registers_i/_3802_  (.A2(net259),
    .A1(net1350),
    .B1(\cs_registers_i/_1321_ ),
    .X(\cs_registers_i/_1322_ ));
 sg13g2_buf_4 fanout542 (.X(net542),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3804_  (.Y(\cs_registers_i/_1324_ ),
    .B1(net1064),
    .B2(net655),
    .A2(\cs_registers_i/_1308_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3805_  (.Y(\cs_registers_i/_0038_ ),
    .A(\cs_registers_i/_1307_ ),
    .B(\cs_registers_i/_1324_ ));
 sg13g2_nand2_1 \cs_registers_i/_3806_  (.Y(\cs_registers_i/_1325_ ),
    .A(csr_depc_7_),
    .B(net660));
 sg13g2_mux2_2 \cs_registers_i/_3807_  (.A0(crash_dump_o_103_),
    .A1(crash_dump_o_71_),
    .S(net1481),
    .X(\cs_registers_i/_1326_ ));
 sg13g2_and2_1 \cs_registers_i/_3808_  (.A(net148),
    .B(net263),
    .X(\cs_registers_i/_1327_ ));
 sg13g2_mux2_1 \cs_registers_i/_3809_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .A1(\cs_registers_i/mhpmcounter_1895_ ),
    .S(net63),
    .X(\cs_registers_i/_1328_ ));
 sg13g2_nand2_1 \cs_registers_i/_3810_  (.Y(\cs_registers_i/_1329_ ),
    .A(net1129),
    .B(\cs_registers_i/_1328_ ));
 sg13g2_mux4_1 \cs_registers_i/_3811_  (.S0(net68),
    .A0(\cs_registers_i/dcsr_q_7_ ),
    .A1(\cs_registers_i/dscratch0_q_7_ ),
    .A2(csr_depc_7_),
    .A3(\cs_registers_i/dscratch1_q_7_ ),
    .S1(net1243),
    .X(\cs_registers_i/_1330_ ));
 sg13g2_nand2_1 \cs_registers_i/_3812_  (.Y(\cs_registers_i/_1331_ ),
    .A(net1153),
    .B(\cs_registers_i/_1330_ ));
 sg13g2_inv_1 \cs_registers_i/_3813_  (.Y(\cs_registers_i/_1332_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_7_ ));
 sg13g2_nand2_1 \cs_registers_i/_3814_  (.Y(\cs_registers_i/_1333_ ),
    .A(net74),
    .B(\cs_registers_i/mhpmcounter_1863_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3815_  (.B1(\cs_registers_i/_1333_ ),
    .Y(\cs_registers_i/_1334_ ),
    .A1(net72),
    .A2(\cs_registers_i/_1332_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3816_  (.Y(\cs_registers_i/_1335_ ),
    .B1(\cs_registers_i/_1334_ ),
    .B2(\cs_registers_i/_0628_ ),
    .A2(net1097),
    .A1(hart_id_i_7_));
 sg13g2_nor2b_1 \cs_registers_i/_3817_  (.A(net102),
    .B_N(\cs_registers_i/mscratch_q_7_ ),
    .Y(\cs_registers_i/_1336_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3818_  (.A1(net102),
    .A2(irq_timer_i),
    .Y(\cs_registers_i/_1337_ ),
    .B1(\cs_registers_i/_1336_ ));
 sg13g2_nor3_1 \cs_registers_i/_3819_  (.A(net1236),
    .B(net1100),
    .C(\cs_registers_i/_1337_ ),
    .Y(\cs_registers_i/_1338_ ));
 sg13g2_mux2_1 \cs_registers_i/_3820_  (.A0(crash_dump_o_7_),
    .A1(\cs_registers_i/mtval_q_7_ ),
    .S(net70),
    .X(\cs_registers_i/_1339_ ));
 sg13g2_nand3_1 \cs_registers_i/_3821_  (.B(\cs_registers_i/_0544_ ),
    .C(\cs_registers_i/_1339_ ),
    .A(net1236),
    .Y(\cs_registers_i/_1340_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3822_  (.Y(\cs_registers_i/_1341_ ),
    .B(\cs_registers_i/_1340_ ),
    .A_N(\cs_registers_i/_1338_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3823_  (.Y(\cs_registers_i/_1342_ ),
    .B1(\cs_registers_i/_0664_ ),
    .B2(csr_mtvec_7_),
    .A2(\cs_registers_i/_0626_ ),
    .A1(\cs_registers_i/mstatus_q_4_ ));
 sg13g2_nand2_1 \cs_registers_i/_3824_  (.Y(\cs_registers_i/_1343_ ),
    .A(\cs_registers_i/mie_q_17_ ),
    .B(net40));
 sg13g2_o21ai_1 \cs_registers_i/_3825_  (.B1(\cs_registers_i/_1343_ ),
    .Y(\cs_registers_i/_1344_ ),
    .A1(net1100),
    .A2(\cs_registers_i/_1342_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3826_  (.B2(\cs_registers_i/_0599_ ),
    .C1(\cs_registers_i/_0649_ ),
    .B1(\cs_registers_i/_1344_ ),
    .A1(net1149),
    .Y(\cs_registers_i/_1345_ ),
    .A2(\cs_registers_i/_1341_ ));
 sg13g2_nand4_1 \cs_registers_i/_3827_  (.B(\cs_registers_i/_1331_ ),
    .C(\cs_registers_i/_1335_ ),
    .A(\cs_registers_i/_1329_ ),
    .Y(\cs_registers_i/_1346_ ),
    .D(\cs_registers_i/_1345_ ));
 sg13g2_nand3b_1 \cs_registers_i/_3828_  (.B(\cs_registers_i/_1208_ ),
    .C(\cs_registers_i/_1346_ ),
    .Y(\cs_registers_i/_1347_ ),
    .A_N(net148));
 sg13g2_nand2b_2 \cs_registers_i/_3829_  (.Y(\cs_registers_i/_1348_ ),
    .B(\cs_registers_i/_1347_ ),
    .A_N(\cs_registers_i/_1327_ ));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3831_  (.Y(\cs_registers_i/_1350_ ),
    .B1(net1031),
    .B2(net655),
    .A2(\cs_registers_i/_1326_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3832_  (.Y(\cs_registers_i/_0039_ ),
    .A(\cs_registers_i/_1325_ ),
    .B(\cs_registers_i/_1350_ ));
 sg13g2_nand2_1 \cs_registers_i/_3833_  (.Y(\cs_registers_i/_1351_ ),
    .A(csr_depc_8_),
    .B(net664));
 sg13g2_mux2_2 \cs_registers_i/_3834_  (.A0(crash_dump_o_104_),
    .A1(crash_dump_o_72_),
    .S(net1482),
    .X(\cs_registers_i/_1352_ ));
 sg13g2_and2_1 \cs_registers_i/_3835_  (.A(crash_dump_o_8_),
    .B(net1234),
    .X(\cs_registers_i/_1353_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3836_  (.A1(net53),
    .A2(\cs_registers_i/mscratch_q_8_ ),
    .Y(\cs_registers_i/_1354_ ),
    .B1(\cs_registers_i/_1353_ ));
 sg13g2_nand2_1 \cs_registers_i/_3837_  (.Y(\cs_registers_i/_1355_ ),
    .A(\cs_registers_i/mtval_q_8_ ),
    .B(net1115));
 sg13g2_o21ai_1 \cs_registers_i/_3838_  (.B1(\cs_registers_i/_1355_ ),
    .Y(\cs_registers_i/_1356_ ),
    .A1(net65),
    .A2(\cs_registers_i/_1354_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3839_  (.Y(\cs_registers_i/_1357_ ),
    .B1(\cs_registers_i/_1356_ ),
    .B2(net1160),
    .A2(\cs_registers_i/_0749_ ),
    .A1(csr_mtvec_8_));
 sg13g2_nor2_1 \cs_registers_i/_3840_  (.A(net1172),
    .B(\cs_registers_i/_1357_ ),
    .Y(\cs_registers_i/_1358_ ));
 sg13g2_mux4_1 \cs_registers_i/_3841_  (.S0(net69),
    .A0(\cs_registers_i/dcsr_q_8_ ),
    .A1(\cs_registers_i/dscratch0_q_8_ ),
    .A2(csr_depc_8_),
    .A3(\cs_registers_i/dscratch1_q_8_ ),
    .S1(net1244),
    .X(\cs_registers_i/_1359_ ));
 sg13g2_inv_1 \cs_registers_i/_3842_  (.Y(\cs_registers_i/_1360_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_8_ ));
 sg13g2_nand2_1 \cs_registers_i/_3843_  (.Y(\cs_registers_i/_1361_ ),
    .A(net77),
    .B(\cs_registers_i/mhpmcounter_1864_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3844_  (.B1(\cs_registers_i/_1361_ ),
    .Y(\cs_registers_i/_1362_ ),
    .A1(net66),
    .A2(\cs_registers_i/_1360_ ));
 sg13g2_mux2_1 \cs_registers_i/_3845_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .A1(\cs_registers_i/mhpmcounter_1896_ ),
    .S(net70),
    .X(\cs_registers_i/_1363_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3846_  (.Y(\cs_registers_i/_1364_ ),
    .B1(\cs_registers_i/_1363_ ),
    .B2(net1156),
    .A2(\cs_registers_i/_1362_ ),
    .A1(net1191));
 sg13g2_o21ai_1 \cs_registers_i/_3847_  (.B1(\cs_registers_i/_0511_ ),
    .Y(\cs_registers_i/_1365_ ),
    .A1(net1159),
    .A2(\cs_registers_i/_1364_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3848_  (.B2(net1153),
    .C1(\cs_registers_i/_1365_ ),
    .B1(\cs_registers_i/_1359_ ),
    .A1(hart_id_i_8_),
    .Y(\cs_registers_i/_1366_ ),
    .A2(net1097));
 sg13g2_nor2b_2 \cs_registers_i/_3849_  (.A(\cs_registers_i/_1358_ ),
    .B_N(\cs_registers_i/_1366_ ),
    .Y(\cs_registers_i/_1367_ ));
 sg13g2_nor3_1 \cs_registers_i/_3850_  (.A(net1280),
    .B(net1093),
    .C(\cs_registers_i/_1367_ ),
    .Y(\cs_registers_i/_1368_ ));
 sg13g2_a21o_2 \cs_registers_i/_3851_  (.A2(net261),
    .A1(net1280),
    .B1(\cs_registers_i/_1368_ ),
    .X(\cs_registers_i/_1369_ ));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3853_  (.Y(\cs_registers_i/_1371_ ),
    .B1(net1025),
    .B2(net658),
    .A2(\cs_registers_i/_1352_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3854_  (.Y(\cs_registers_i/_0040_ ),
    .A(\cs_registers_i/_1351_ ),
    .B(\cs_registers_i/_1371_ ));
 sg13g2_nand2_1 \cs_registers_i/_3855_  (.Y(\cs_registers_i/_1372_ ),
    .A(csr_depc_9_),
    .B(net659));
 sg13g2_mux2_2 \cs_registers_i/_3856_  (.A0(crash_dump_o_105_),
    .A1(crash_dump_o_73_),
    .S(net1481),
    .X(\cs_registers_i/_1373_ ));
 sg13g2_mux2_1 \cs_registers_i/_3857_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ),
    .A1(\cs_registers_i/mhpmcounter_1897_ ),
    .S(net63),
    .X(\cs_registers_i/_1374_ ));
 sg13g2_nand2_1 \cs_registers_i/_3858_  (.Y(\cs_registers_i/_1375_ ),
    .A(net1129),
    .B(\cs_registers_i/_1374_ ));
 sg13g2_mux4_1 \cs_registers_i/_3859_  (.S0(net67),
    .A0(\cs_registers_i/dcsr_q_9_ ),
    .A1(\cs_registers_i/dscratch0_q_9_ ),
    .A2(csr_depc_9_),
    .A3(\cs_registers_i/dscratch1_q_9_ ),
    .S1(net1232),
    .X(\cs_registers_i/_1376_ ));
 sg13g2_nand2_1 \cs_registers_i/_3860_  (.Y(\cs_registers_i/_1377_ ),
    .A(net1150),
    .B(\cs_registers_i/_1376_ ));
 sg13g2_and2_1 \cs_registers_i/_3861_  (.A(crash_dump_o_9_),
    .B(net1234),
    .X(\cs_registers_i/_1378_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3862_  (.A1(net54),
    .A2(\cs_registers_i/mscratch_q_9_ ),
    .Y(\cs_registers_i/_1379_ ),
    .B1(\cs_registers_i/_1378_ ));
 sg13g2_nand3_1 \cs_registers_i/_3863_  (.B(net1232),
    .C(\cs_registers_i/mtval_q_9_ ),
    .A(net75),
    .Y(\cs_registers_i/_1380_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3864_  (.B1(\cs_registers_i/_1380_ ),
    .Y(\cs_registers_i/_1381_ ),
    .A1(net72),
    .A2(\cs_registers_i/_1379_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3865_  (.Y(\cs_registers_i/_1382_ ),
    .B1(\cs_registers_i/_0605_ ),
    .B2(\cs_registers_i/_1381_ ),
    .A2(\cs_registers_i/_0600_ ),
    .A1(csr_mtvec_9_));
 sg13g2_a21oi_1 \cs_registers_i/_3866_  (.A1(hart_id_i_9_),
    .A2(net1155),
    .Y(\cs_registers_i/_1383_ ),
    .B1(net1174));
 sg13g2_nor3_1 \cs_registers_i/_3867_  (.A(\cs_registers_i/_0922_ ),
    .B(net1100),
    .C(\cs_registers_i/_1383_ ),
    .Y(\cs_registers_i/_1384_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3868_  (.B1(\cs_registers_i/_0552_ ),
    .Y(\cs_registers_i/_1385_ ),
    .A1(net1131),
    .A2(\cs_registers_i/_0718_ ));
 sg13g2_nand2_1 \cs_registers_i/_3869_  (.Y(\cs_registers_i/_1386_ ),
    .A(net1191),
    .B(\cs_registers_i/_1385_ ));
 sg13g2_nand2_1 \cs_registers_i/_3870_  (.Y(\cs_registers_i/_1387_ ),
    .A(net1275),
    .B(\cs_registers_i/_0672_ ));
 sg13g2_nand3_1 \cs_registers_i/_3871_  (.B(\cs_registers_i/_0720_ ),
    .C(\cs_registers_i/_1387_ ),
    .A(\cs_registers_i/_0927_ ),
    .Y(\cs_registers_i/_1388_ ));
 sg13g2_nand2_1 \cs_registers_i/_3872_  (.Y(\cs_registers_i/_1389_ ),
    .A(net1114),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ));
 sg13g2_nand2_1 \cs_registers_i/_3873_  (.Y(\cs_registers_i/_1390_ ),
    .A(net76),
    .B(\cs_registers_i/mhpmcounter_1865_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3874_  (.B2(\cs_registers_i/_1390_ ),
    .C1(net1159),
    .B1(\cs_registers_i/_1389_ ),
    .A1(\cs_registers_i/_1386_ ),
    .Y(\cs_registers_i/_1391_ ),
    .A2(\cs_registers_i/_1388_ ));
 sg13g2_nor3_1 \cs_registers_i/_3875_  (.A(\cs_registers_i/_0649_ ),
    .B(\cs_registers_i/_1384_ ),
    .C(\cs_registers_i/_1391_ ),
    .Y(\cs_registers_i/_1392_ ));
 sg13g2_nand4_1 \cs_registers_i/_3876_  (.B(\cs_registers_i/_1377_ ),
    .C(\cs_registers_i/_1382_ ),
    .A(\cs_registers_i/_1375_ ),
    .Y(\cs_registers_i/_1393_ ),
    .D(\cs_registers_i/_1392_ ));
 sg13g2_nand2_1 \cs_registers_i/_3877_  (.Y(\cs_registers_i/_1394_ ),
    .A(\cs_registers_i/_1208_ ),
    .B(\cs_registers_i/_1393_ ));
 sg13g2_nand2_1 \cs_registers_i/_3878_  (.Y(\cs_registers_i/_1395_ ),
    .A(net192),
    .B(net263));
 sg13g2_o21ai_1 \cs_registers_i/_3879_  (.B1(\cs_registers_i/_1395_ ),
    .Y(\cs_registers_i/_1396_ ),
    .A1(net192),
    .A2(\cs_registers_i/_1394_ ));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(net546));
 sg13g2_a22oi_1 \cs_registers_i/_3881_  (.Y(\cs_registers_i/_1398_ ),
    .B1(net1030),
    .B2(net654),
    .A2(\cs_registers_i/_1373_ ),
    .A1(net1309));
 sg13g2_nand2_1 \cs_registers_i/_3882_  (.Y(\cs_registers_i/_0041_ ),
    .A(\cs_registers_i/_1372_ ),
    .B(\cs_registers_i/_1398_ ));
 sg13g2_nor2_2 \cs_registers_i/_3883_  (.A(debug_csr_save),
    .B(debug_mode),
    .Y(\cs_registers_i/_1399_ ));
 sg13g2_and2_2 \cs_registers_i/_3884_  (.A(net255),
    .B(\cs_registers_i/_1399_ ),
    .X(\cs_registers_i/_1400_ ));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net546));
 sg13g2_buf_1 fanout537 (.A(\id_stage_i.controller_i.instr_i_16_ ),
    .X(net537));
 sg13g2_buf_8 fanout536 (.A(\id_stage_i.controller_i.instr_i_16_ ),
    .X(net536));
 sg13g2_and2_1 \cs_registers_i/_3888_  (.A(net344),
    .B(\id_stage_i.controller_i.nmi_mode_o ),
    .X(\cs_registers_i/_1404_ ));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(net536));
 sg13g2_buf_4 fanout534 (.X(net534),
    .A(net536));
 sg13g2_a22oi_1 \cs_registers_i/_3891_  (.Y(\cs_registers_i/_1407_ ),
    .B1(net290),
    .B2(\cs_registers_i/mstack_epc_q_0_ ),
    .A2(net1293),
    .A1(\cs_registers_i/_0588_ ));
 sg13g2_nand2_1 \cs_registers_i/_3892_  (.Y(\cs_registers_i/_1408_ ),
    .A(\cs_registers_i/_0544_ ),
    .B(\cs_registers_i/_0717_ ));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(net536));
 sg13g2_nand2_2 \cs_registers_i/_3894_  (.Y(\cs_registers_i/_1410_ ),
    .A(net722),
    .B(net1148));
 sg13g2_nor2_1 \cs_registers_i/_3895_  (.A(net1298),
    .B(net290),
    .Y(\cs_registers_i/_1411_ ));
 sg13g2_o21ai_1 \cs_registers_i/_3896_  (.B1(\cs_registers_i/_1411_ ),
    .Y(\cs_registers_i/_1412_ ),
    .A1(\cs_registers_i/_1408_ ),
    .A2(\cs_registers_i/_1410_ ));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(net536));
 sg13g2_buf_2 fanout531 (.A(net536),
    .X(net531));
 sg13g2_nor2_2 \cs_registers_i/_3899_  (.A(crash_dump_o_0_),
    .B(net588),
    .Y(\cs_registers_i/_1415_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3900_  (.B1(\cs_registers_i/_1415_ ),
    .Y(\cs_registers_i/_0042_ ),
    .A2(net588),
    .A1(\cs_registers_i/_1407_ ));
 sg13g2_buf_2 fanout530 (.A(\id_stage_i.controller_i.instr_i_17_ ),
    .X(net530));
 sg13g2_or2_2 \cs_registers_i/_3902_  (.X(\cs_registers_i/_1417_ ),
    .B(debug_mode),
    .A(debug_csr_save));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(\id_stage_i.controller_i.instr_i_17_ ));
 sg13g2_nand2b_1 \cs_registers_i/_3904_  (.Y(\cs_registers_i/_1419_ ),
    .B(net345),
    .A_N(\id_stage_i.controller_i.nmi_mode_o ));
 sg13g2_o21ai_1 \cs_registers_i/_3905_  (.B1(\cs_registers_i/_1419_ ),
    .Y(\cs_registers_i/_1420_ ),
    .A1(net344),
    .A2(net255));
 sg13g2_a21o_1 \cs_registers_i/_3906_  (.A2(\cs_registers_i/_1417_ ),
    .A1(net256),
    .B1(\cs_registers_i/_1420_ ),
    .X(\cs_registers_i/_1421_ ));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(\id_stage_i.controller_i.instr_i_17_ ));
 sg13g2_buf_4 fanout527 (.X(net527),
    .A(\id_stage_i.controller_i.instr_i_17_ ));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(\id_stage_i.controller_i.instr_i_17_ ));
 sg13g2_and2_1 \cs_registers_i/_3910_  (.A(\cs_registers_i/mstack_epc_q_10_ ),
    .B(net291),
    .X(\cs_registers_i/_1425_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3911_  (.B2(net1059),
    .C1(\cs_registers_i/_1425_ ),
    .B1(net154),
    .A1(\cs_registers_i/_0593_ ),
    .Y(\cs_registers_i/_1426_ ),
    .A2(net1307));
 sg13g2_nor2_2 \cs_registers_i/_3912_  (.A(crash_dump_o_10_),
    .B(net595),
    .Y(\cs_registers_i/_1427_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3913_  (.A1(net595),
    .A2(\cs_registers_i/_1426_ ),
    .Y(\cs_registers_i/_0043_ ),
    .B1(\cs_registers_i/_1427_ ));
 sg13g2_mux2_1 \cs_registers_i/_3914_  (.A0(\cs_registers_i/_0661_ ),
    .A1(net1070),
    .S(\cs_registers_i/_1417_ ),
    .X(\cs_registers_i/_1428_ ));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(\id_stage_i.controller_i.instr_i_17_ ));
 sg13g2_mux2_2 \cs_registers_i/_3916_  (.A0(net256),
    .A1(\id_stage_i.controller_i.nmi_mode_o ),
    .S(net344),
    .X(\cs_registers_i/_1430_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3917_  (.A(\cs_registers_i/_1430_ ),
    .B_N(net263),
    .Y(\cs_registers_i/_1431_ ));
 sg13g2_nor4_1 \cs_registers_i/_3918_  (.A(net1414),
    .B(net1092),
    .C(\cs_registers_i/_0696_ ),
    .D(\cs_registers_i/_1430_ ),
    .Y(\cs_registers_i/_1432_ ));
 sg13g2_a21o_1 \cs_registers_i/_3919_  (.A2(\cs_registers_i/_1431_ ),
    .A1(net1414),
    .B1(\cs_registers_i/_1432_ ),
    .X(\cs_registers_i/_1433_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3920_  (.B2(net256),
    .C1(\cs_registers_i/_1433_ ),
    .B1(\cs_registers_i/_1428_ ),
    .A1(\cs_registers_i/mstack_epc_q_11_ ),
    .Y(\cs_registers_i/_1434_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_3921_  (.A(crash_dump_o_11_),
    .B(net591),
    .Y(\cs_registers_i/_1435_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3922_  (.A1(net591),
    .A2(\cs_registers_i/_1434_ ),
    .Y(\cs_registers_i/_0044_ ),
    .B1(\cs_registers_i/_1435_ ));
 sg13g2_and2_1 \cs_registers_i/_3923_  (.A(\cs_registers_i/mstack_epc_q_12_ ),
    .B(net291),
    .X(\cs_registers_i/_1436_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3924_  (.B2(net1028),
    .C1(\cs_registers_i/_1436_ ),
    .B1(net154),
    .A1(\cs_registers_i/_0702_ ),
    .Y(\cs_registers_i/_1437_ ),
    .A2(net1307));
 sg13g2_nor2_2 \cs_registers_i/_3925_  (.A(crash_dump_o_12_),
    .B(net595),
    .Y(\cs_registers_i/_1438_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3926_  (.B1(\cs_registers_i/_1438_ ),
    .Y(\cs_registers_i/_0045_ ),
    .A2(\cs_registers_i/_1437_ ),
    .A1(net595));
 sg13g2_and2_1 \cs_registers_i/_3927_  (.A(\cs_registers_i/mstack_epc_q_13_ ),
    .B(net291),
    .X(\cs_registers_i/_1439_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3928_  (.B2(net1057),
    .C1(\cs_registers_i/_1439_ ),
    .B1(net154),
    .A1(\cs_registers_i/_0742_ ),
    .Y(\cs_registers_i/_1440_ ),
    .A2(net1306));
 sg13g2_nor2_2 \cs_registers_i/_3929_  (.A(crash_dump_o_13_),
    .B(net597),
    .Y(\cs_registers_i/_1441_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3930_  (.B1(\cs_registers_i/_1441_ ),
    .Y(\cs_registers_i/_0046_ ),
    .A2(\cs_registers_i/_1440_ ),
    .A1(net597));
 sg13g2_mux2_1 \cs_registers_i/_3931_  (.A0(\cs_registers_i/_0768_ ),
    .A1(net1056),
    .S(\cs_registers_i/_1417_ ),
    .X(\cs_registers_i/_1442_ ));
 sg13g2_nor4_1 \cs_registers_i/_3932_  (.A(alu_operand_a_ex_14_),
    .B(net1092),
    .C(\cs_registers_i/_0788_ ),
    .D(\cs_registers_i/_1430_ ),
    .Y(\cs_registers_i/_1443_ ));
 sg13g2_a21o_1 \cs_registers_i/_3933_  (.A2(\cs_registers_i/_1431_ ),
    .A1(alu_operand_a_ex_14_),
    .B1(\cs_registers_i/_1443_ ),
    .X(\cs_registers_i/_1444_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3934_  (.B2(net256),
    .C1(\cs_registers_i/_1444_ ),
    .B1(\cs_registers_i/_1442_ ),
    .A1(\cs_registers_i/mstack_epc_q_14_ ),
    .Y(\cs_registers_i/_1445_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_3935_  (.A(crash_dump_o_14_),
    .B(net589),
    .Y(\cs_registers_i/_1446_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3936_  (.B1(\cs_registers_i/_1446_ ),
    .Y(\cs_registers_i/_0047_ ),
    .A2(\cs_registers_i/_1445_ ),
    .A1(net589));
 sg13g2_mux2_1 \cs_registers_i/_3937_  (.A0(\cs_registers_i/_0794_ ),
    .A1(net1068),
    .S(\cs_registers_i/_1417_ ),
    .X(\cs_registers_i/_1447_ ));
 sg13g2_nor4_1 \cs_registers_i/_3938_  (.A(alu_operand_a_ex_15_),
    .B(net1090),
    .C(\cs_registers_i/_0806_ ),
    .D(\cs_registers_i/_1430_ ),
    .Y(\cs_registers_i/_1448_ ));
 sg13g2_a21o_1 \cs_registers_i/_3939_  (.A2(\cs_registers_i/_1431_ ),
    .A1(alu_operand_a_ex_15_),
    .B1(\cs_registers_i/_1448_ ),
    .X(\cs_registers_i/_1449_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3940_  (.B2(net256),
    .C1(\cs_registers_i/_1449_ ),
    .B1(\cs_registers_i/_1447_ ),
    .A1(\cs_registers_i/mstack_epc_q_15_ ),
    .Y(\cs_registers_i/_1450_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_3941_  (.A(crash_dump_o_15_),
    .B(net590),
    .Y(\cs_registers_i/_1451_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3942_  (.A1(net590),
    .A2(\cs_registers_i/_1450_ ),
    .Y(\cs_registers_i/_0048_ ),
    .B1(\cs_registers_i/_1451_ ));
 sg13g2_and2_1 \cs_registers_i/_3943_  (.A(net263),
    .B(net153),
    .X(\cs_registers_i/_1452_ ));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_nor2b_1 \cs_registers_i/_3946_  (.A(net1088),
    .B_N(net153),
    .Y(\cs_registers_i/_1455_ ));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_nor2_1 \cs_registers_i/_3948_  (.A(alu_operand_a_ex_16_),
    .B(\cs_registers_i/_0832_ ),
    .Y(\cs_registers_i/_1457_ ));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3951_  (.Y(\cs_registers_i/_1460_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_epc_q_16_ ),
    .A2(net1303),
    .A1(\cs_registers_i/_0813_ ));
 sg13g2_inv_1 \cs_registers_i/_3952_  (.Y(\cs_registers_i/_1461_ ),
    .A(\cs_registers_i/_1460_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3953_  (.B2(\cs_registers_i/_1457_ ),
    .C1(\cs_registers_i/_1461_ ),
    .B1(net1078),
    .A1(alu_operand_a_ex_16_),
    .Y(\cs_registers_i/_1462_ ),
    .A2(net1205));
 sg13g2_nor2_2 \cs_registers_i/_3954_  (.A(crash_dump_o_16_),
    .B(net592),
    .Y(\cs_registers_i/_1463_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3955_  (.A1(net594),
    .A2(\cs_registers_i/_1462_ ),
    .Y(\cs_registers_i/_0049_ ),
    .B1(\cs_registers_i/_1463_ ));
 sg13g2_nor2_1 \cs_registers_i/_3956_  (.A(net1251),
    .B(\cs_registers_i/_0858_ ),
    .Y(\cs_registers_i/_1464_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3957_  (.Y(\cs_registers_i/_1465_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_17_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_0840_ ));
 sg13g2_inv_1 \cs_registers_i/_3958_  (.Y(\cs_registers_i/_1466_ ),
    .A(\cs_registers_i/_1465_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3959_  (.B2(\cs_registers_i/_1464_ ),
    .C1(\cs_registers_i/_1466_ ),
    .B1(net1077),
    .A1(net1251),
    .Y(\cs_registers_i/_1467_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_3960_  (.A(crash_dump_o_17_),
    .B(net592),
    .Y(\cs_registers_i/_1468_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3961_  (.A1(net592),
    .A2(\cs_registers_i/_1467_ ),
    .Y(\cs_registers_i/_0050_ ),
    .B1(\cs_registers_i/_1468_ ));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_and2_1 \cs_registers_i/_3963_  (.A(\cs_registers_i/mstack_epc_q_18_ ),
    .B(net291),
    .X(\cs_registers_i/_1470_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3964_  (.B2(net1051),
    .C1(\cs_registers_i/_1470_ ),
    .B1(net154),
    .A1(\cs_registers_i/_0864_ ),
    .Y(\cs_registers_i/_1471_ ),
    .A2(net1307));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_nor2_2 \cs_registers_i/_3966_  (.A(crash_dump_o_18_),
    .B(net595),
    .Y(\cs_registers_i/_1473_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3967_  (.A1(net595),
    .A2(\cs_registers_i/_1471_ ),
    .Y(\cs_registers_i/_0051_ ),
    .B1(\cs_registers_i/_1473_ ));
 sg13g2_nor2_1 \cs_registers_i/_3968_  (.A(net1249),
    .B(\cs_registers_i/_0901_ ),
    .Y(\cs_registers_i/_1474_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3969_  (.Y(\cs_registers_i/_1475_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_19_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_0887_ ));
 sg13g2_inv_1 \cs_registers_i/_3970_  (.Y(\cs_registers_i/_1476_ ),
    .A(\cs_registers_i/_1475_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3971_  (.B2(\cs_registers_i/_1474_ ),
    .C1(\cs_registers_i/_1476_ ),
    .B1(net1077),
    .A1(net1249),
    .Y(\cs_registers_i/_1477_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_3972_  (.A(crash_dump_o_19_),
    .B(net593),
    .Y(\cs_registers_i/_1478_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3973_  (.B1(\cs_registers_i/_1478_ ),
    .Y(\cs_registers_i/_0052_ ),
    .A2(\cs_registers_i/_1477_ ),
    .A1(net592));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net524));
 sg13g2_and2_1 \cs_registers_i/_3975_  (.A(\cs_registers_i/mstack_epc_q_1_ ),
    .B(net291),
    .X(\cs_registers_i/_1480_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3976_  (.B2(net1067),
    .C1(\cs_registers_i/_1480_ ),
    .B1(net154),
    .A1(\cs_registers_i/_0908_ ),
    .Y(\cs_registers_i/_1481_ ),
    .A2(net1296));
 sg13g2_nor2_2 \cs_registers_i/_3977_  (.A(crash_dump_o_1_),
    .B(net597),
    .Y(\cs_registers_i/_1482_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3978_  (.A1(net597),
    .A2(\cs_registers_i/_1481_ ),
    .Y(\cs_registers_i/_0053_ ),
    .B1(\cs_registers_i/_1482_ ));
 sg13g2_nor2_1 \cs_registers_i/_3979_  (.A(net1282),
    .B(\cs_registers_i/_0959_ ),
    .Y(\cs_registers_i/_1483_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3980_  (.Y(\cs_registers_i/_1484_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_20_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_0937_ ));
 sg13g2_inv_1 \cs_registers_i/_3981_  (.Y(\cs_registers_i/_1485_ ),
    .A(\cs_registers_i/_1484_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3982_  (.B2(\cs_registers_i/_1483_ ),
    .C1(\cs_registers_i/_1485_ ),
    .B1(net1077),
    .A1(net1282),
    .Y(\cs_registers_i/_1486_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_3983_  (.A(crash_dump_o_20_),
    .B(net593),
    .Y(\cs_registers_i/_1487_ ));
 sg13g2_a21oi_2 \cs_registers_i/_3984_  (.B1(\cs_registers_i/_1487_ ),
    .Y(\cs_registers_i/_0054_ ),
    .A2(\cs_registers_i/_1486_ ),
    .A1(net593));
 sg13g2_nor2_1 \cs_registers_i/_3985_  (.A(net126),
    .B(\cs_registers_i/_0981_ ),
    .Y(\cs_registers_i/_1488_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3986_  (.Y(\cs_registers_i/_1489_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_21_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_0965_ ));
 sg13g2_inv_1 \cs_registers_i/_3987_  (.Y(\cs_registers_i/_1490_ ),
    .A(\cs_registers_i/_1489_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3988_  (.B2(\cs_registers_i/_1488_ ),
    .C1(\cs_registers_i/_1490_ ),
    .B1(net1077),
    .A1(net127),
    .Y(\cs_registers_i/_1491_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_3989_  (.A(crash_dump_o_21_),
    .B(net593),
    .Y(\cs_registers_i/_1492_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3990_  (.A1(net593),
    .A2(\cs_registers_i/_1491_ ),
    .Y(\cs_registers_i/_0055_ ),
    .B1(\cs_registers_i/_1492_ ));
 sg13g2_nor2_1 \cs_registers_i/_3991_  (.A(net195),
    .B(\cs_registers_i/_1007_ ),
    .Y(\cs_registers_i/_1493_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3992_  (.Y(\cs_registers_i/_1494_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_22_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_0987_ ));
 sg13g2_inv_1 \cs_registers_i/_3993_  (.Y(\cs_registers_i/_1495_ ),
    .A(\cs_registers_i/_1494_ ));
 sg13g2_a221oi_1 \cs_registers_i/_3994_  (.B2(\cs_registers_i/_1493_ ),
    .C1(\cs_registers_i/_1495_ ),
    .B1(net1077),
    .A1(net196),
    .Y(\cs_registers_i/_1496_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_3995_  (.A(crash_dump_o_22_),
    .B(net593),
    .Y(\cs_registers_i/_1497_ ));
 sg13g2_a21oi_1 \cs_registers_i/_3996_  (.A1(net593),
    .A2(\cs_registers_i/_1496_ ),
    .Y(\cs_registers_i/_0056_ ),
    .B1(\cs_registers_i/_1497_ ));
 sg13g2_nor2_1 \cs_registers_i/_3997_  (.A(net149),
    .B(\cs_registers_i/_1029_ ),
    .Y(\cs_registers_i/_1498_ ));
 sg13g2_a22oi_1 \cs_registers_i/_3998_  (.Y(\cs_registers_i/_1499_ ),
    .B1(net292),
    .B2(\cs_registers_i/mstack_epc_q_23_ ),
    .A2(net1294),
    .A1(\cs_registers_i/_1013_ ));
 sg13g2_inv_1 \cs_registers_i/_3999_  (.Y(\cs_registers_i/_1500_ ),
    .A(\cs_registers_i/_1499_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4000_  (.B2(\cs_registers_i/_1498_ ),
    .C1(\cs_registers_i/_1500_ ),
    .B1(net1079),
    .A1(net150),
    .Y(\cs_registers_i/_1501_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4001_  (.A(crash_dump_o_23_),
    .B(net588),
    .Y(\cs_registers_i/_1502_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4002_  (.B1(\cs_registers_i/_1502_ ),
    .Y(\cs_registers_i/_0057_ ),
    .A2(\cs_registers_i/_1501_ ),
    .A1(net588));
 sg13g2_and2_1 \cs_registers_i/_4003_  (.A(\cs_registers_i/mstack_epc_q_24_ ),
    .B(net291),
    .X(\cs_registers_i/_1503_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4004_  (.B2(net1044),
    .C1(\cs_registers_i/_1503_ ),
    .B1(net154),
    .A1(\cs_registers_i/_1034_ ),
    .Y(\cs_registers_i/_1504_ ),
    .A2(net1307));
 sg13g2_nor2_2 \cs_registers_i/_4005_  (.A(crash_dump_o_24_),
    .B(net595),
    .Y(\cs_registers_i/_1505_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4006_  (.A1(net595),
    .A2(\cs_registers_i/_1504_ ),
    .Y(\cs_registers_i/_0058_ ),
    .B1(\cs_registers_i/_1505_ ));
 sg13g2_nor2_1 \cs_registers_i/_4007_  (.A(alu_operand_a_ex_25_),
    .B(\cs_registers_i/_1077_ ),
    .Y(\cs_registers_i/_1506_ ));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net524));
 sg13g2_a22oi_1 \cs_registers_i/_4009_  (.Y(\cs_registers_i/_1508_ ),
    .B1(net294),
    .B2(\cs_registers_i/mstack_epc_q_25_ ),
    .A2(net1303),
    .A1(\cs_registers_i/_1056_ ));
 sg13g2_inv_1 \cs_registers_i/_4010_  (.Y(\cs_registers_i/_1509_ ),
    .A(\cs_registers_i/_1508_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4011_  (.B2(\cs_registers_i/_1506_ ),
    .C1(\cs_registers_i/_1509_ ),
    .B1(net1078),
    .A1(alu_operand_a_ex_25_),
    .Y(\cs_registers_i/_1510_ ),
    .A2(net1205));
 sg13g2_nor2_2 \cs_registers_i/_4012_  (.A(crash_dump_o_25_),
    .B(net594),
    .Y(\cs_registers_i/_1511_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4013_  (.B1(\cs_registers_i/_1511_ ),
    .Y(\cs_registers_i/_0059_ ),
    .A2(\cs_registers_i/_1510_ ),
    .A1(net594));
 sg13g2_nor2_1 \cs_registers_i/_4014_  (.A(net87),
    .B(\cs_registers_i/_1098_ ),
    .Y(\cs_registers_i/_1512_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4015_  (.Y(\cs_registers_i/_1513_ ),
    .B1(net294),
    .B2(\cs_registers_i/mstack_epc_q_26_ ),
    .A2(net1303),
    .A1(\cs_registers_i/_1084_ ));
 sg13g2_inv_1 \cs_registers_i/_4016_  (.Y(\cs_registers_i/_1514_ ),
    .A(\cs_registers_i/_1513_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4017_  (.B2(\cs_registers_i/_1512_ ),
    .C1(\cs_registers_i/_1514_ ),
    .B1(net1077),
    .A1(net88),
    .Y(\cs_registers_i/_1515_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_4018_  (.A(crash_dump_o_26_),
    .B(net592),
    .Y(\cs_registers_i/_1516_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4019_  (.B1(\cs_registers_i/_1516_ ),
    .Y(\cs_registers_i/_0060_ ),
    .A2(\cs_registers_i/_1515_ ),
    .A1(net592));
 sg13g2_nor2_1 \cs_registers_i/_4020_  (.A(net122),
    .B(\cs_registers_i/_1126_ ),
    .Y(\cs_registers_i/_1517_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4021_  (.Y(\cs_registers_i/_1518_ ),
    .B1(net294),
    .B2(\cs_registers_i/mstack_epc_q_27_ ),
    .A2(net1303),
    .A1(\cs_registers_i/_1104_ ));
 sg13g2_inv_1 \cs_registers_i/_4022_  (.Y(\cs_registers_i/_1519_ ),
    .A(\cs_registers_i/_1518_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4023_  (.B2(\cs_registers_i/_1517_ ),
    .C1(\cs_registers_i/_1519_ ),
    .B1(net1078),
    .A1(net124),
    .Y(\cs_registers_i/_1520_ ),
    .A2(net1205));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(net524));
 sg13g2_nor2_2 \cs_registers_i/_4025_  (.A(crash_dump_o_27_),
    .B(net594),
    .Y(\cs_registers_i/_1522_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4026_  (.A1(net594),
    .A2(\cs_registers_i/_1520_ ),
    .Y(\cs_registers_i/_0061_ ),
    .B1(\cs_registers_i/_1522_ ));
 sg13g2_nor2_1 \cs_registers_i/_4027_  (.A(net1201),
    .B(\cs_registers_i/_1150_ ),
    .Y(\cs_registers_i/_1523_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4028_  (.Y(\cs_registers_i/_1524_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_epc_q_28_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_1132_ ));
 sg13g2_inv_1 \cs_registers_i/_4029_  (.Y(\cs_registers_i/_1525_ ),
    .A(\cs_registers_i/_1524_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4030_  (.B2(\cs_registers_i/_1523_ ),
    .C1(\cs_registers_i/_1525_ ),
    .B1(net1077),
    .A1(net1200),
    .Y(\cs_registers_i/_1526_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_4031_  (.A(crash_dump_o_28_),
    .B(net592),
    .Y(\cs_registers_i/_1527_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4032_  (.A1(net592),
    .A2(\cs_registers_i/_1526_ ),
    .Y(\cs_registers_i/_0062_ ),
    .B1(\cs_registers_i/_1527_ ));
 sg13g2_buf_4 fanout514 (.X(net514),
    .A(net524));
 sg13g2_and2_1 \cs_registers_i/_4034_  (.A(\cs_registers_i/mstack_epc_q_29_ ),
    .B(net291),
    .X(\cs_registers_i/_1529_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4035_  (.B2(net1040),
    .C1(\cs_registers_i/_1529_ ),
    .B1(net154),
    .A1(\cs_registers_i/_1157_ ),
    .Y(\cs_registers_i/_1530_ ),
    .A2(net1307));
 sg13g2_nor2_2 \cs_registers_i/_4036_  (.A(crash_dump_o_29_),
    .B(net596),
    .Y(\cs_registers_i/_1531_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4037_  (.B1(\cs_registers_i/_1531_ ),
    .Y(\cs_registers_i/_0063_ ),
    .A2(\cs_registers_i/_1530_ ),
    .A1(net596));
 sg13g2_and2_1 \cs_registers_i/_4038_  (.A(\cs_registers_i/mstack_epc_q_2_ ),
    .B(net290),
    .X(\cs_registers_i/_1532_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4039_  (.B2(net1039),
    .C1(\cs_registers_i/_1532_ ),
    .B1(net153),
    .A1(\cs_registers_i/_1186_ ),
    .Y(\cs_registers_i/_1533_ ),
    .A2(net1307));
 sg13g2_nor2_2 \cs_registers_i/_4040_  (.A(crash_dump_o_2_),
    .B(net596),
    .Y(\cs_registers_i/_1534_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4041_  (.A1(net596),
    .A2(\cs_registers_i/_1533_ ),
    .Y(\cs_registers_i/_0064_ ),
    .B1(\cs_registers_i/_1534_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4042_  (.A(alu_operand_a_ex_30_),
    .B_N(\cs_registers_i/_1221_ ),
    .Y(\cs_registers_i/_1535_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4043_  (.Y(\cs_registers_i/_1536_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_epc_q_30_ ),
    .A2(net1302),
    .A1(\cs_registers_i/_1207_ ));
 sg13g2_inv_1 \cs_registers_i/_4044_  (.Y(\cs_registers_i/_1537_ ),
    .A(\cs_registers_i/_1536_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4045_  (.B2(\cs_registers_i/_1535_ ),
    .C1(\cs_registers_i/_1537_ ),
    .B1(net1077),
    .A1(alu_operand_a_ex_30_),
    .Y(\cs_registers_i/_1538_ ),
    .A2(net1204));
 sg13g2_nor2_2 \cs_registers_i/_4046_  (.A(crash_dump_o_30_),
    .B(net594),
    .Y(\cs_registers_i/_1539_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4047_  (.A1(net598),
    .A2(\cs_registers_i/_1538_ ),
    .Y(\cs_registers_i/_0065_ ),
    .B1(\cs_registers_i/_1539_ ));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(\id_stage_i.controller_i.instr_i_20_ ));
 sg13g2_and2_1 \cs_registers_i/_4049_  (.A(\cs_registers_i/_1228_ ),
    .B(net1307),
    .X(\cs_registers_i/_1541_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4050_  (.B2(net1035),
    .C1(\cs_registers_i/_1541_ ),
    .B1(net153),
    .A1(\cs_registers_i/mstack_epc_q_31_ ),
    .Y(\cs_registers_i/_1542_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_4051_  (.A(crash_dump_o_31_),
    .B(net596),
    .Y(\cs_registers_i/_1543_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4052_  (.A1(net596),
    .A2(\cs_registers_i/_1542_ ),
    .Y(\cs_registers_i/_0066_ ),
    .B1(\cs_registers_i/_1543_ ));
 sg13g2_and2_1 \cs_registers_i/_4053_  (.A(\cs_registers_i/mstack_epc_q_3_ ),
    .B(net290),
    .X(\cs_registers_i/_1544_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4054_  (.B2(net1033),
    .C1(\cs_registers_i/_1544_ ),
    .B1(net153),
    .A1(\cs_registers_i/_1248_ ),
    .Y(\cs_registers_i/_1545_ ),
    .A2(net1294));
 sg13g2_nor2_2 \cs_registers_i/_4055_  (.A(crash_dump_o_3_),
    .B(net588),
    .Y(\cs_registers_i/_1546_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4056_  (.B1(\cs_registers_i/_1546_ ),
    .Y(\cs_registers_i/_0067_ ),
    .A2(\cs_registers_i/_1545_ ),
    .A1(net588));
 sg13g2_and2_1 \cs_registers_i/_4057_  (.A(\cs_registers_i/mstack_epc_q_4_ ),
    .B(net292),
    .X(\cs_registers_i/_1547_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4058_  (.B2(net1032),
    .C1(\cs_registers_i/_1547_ ),
    .B1(net153),
    .A1(\cs_registers_i/_1276_ ),
    .Y(\cs_registers_i/_1548_ ),
    .A2(net1293));
 sg13g2_nor2_2 \cs_registers_i/_4059_  (.A(crash_dump_o_4_),
    .B(net588),
    .Y(\cs_registers_i/_1549_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4060_  (.B1(\cs_registers_i/_1549_ ),
    .Y(\cs_registers_i/_0068_ ),
    .A2(\cs_registers_i/_1548_ ),
    .A1(net588));
 sg13g2_and2_1 \cs_registers_i/_4061_  (.A(\cs_registers_i/mstack_epc_q_5_ ),
    .B(net292),
    .X(\cs_registers_i/_1550_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4062_  (.B2(net1065),
    .C1(\cs_registers_i/_1550_ ),
    .B1(net153),
    .A1(\cs_registers_i/_1289_ ),
    .Y(\cs_registers_i/_1551_ ),
    .A2(net1293));
 sg13g2_nor2_2 \cs_registers_i/_4063_  (.A(crash_dump_o_5_),
    .B(net589),
    .Y(\cs_registers_i/_1552_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4064_  (.A1(net589),
    .A2(\cs_registers_i/_1551_ ),
    .Y(\cs_registers_i/_0069_ ),
    .B1(\cs_registers_i/_1552_ ));
 sg13g2_mux2_1 \cs_registers_i/_4065_  (.A0(\cs_registers_i/_1308_ ),
    .A1(net1064),
    .S(\cs_registers_i/_1417_ ),
    .X(\cs_registers_i/_1553_ ));
 sg13g2_nor4_1 \cs_registers_i/_4066_  (.A(net1349),
    .B(net1090),
    .C(\cs_registers_i/_1320_ ),
    .D(\cs_registers_i/_1430_ ),
    .Y(\cs_registers_i/_1554_ ));
 sg13g2_a21o_1 \cs_registers_i/_4067_  (.A2(\cs_registers_i/_1431_ ),
    .A1(net1349),
    .B1(\cs_registers_i/_1554_ ),
    .X(\cs_registers_i/_1555_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4068_  (.B2(net256),
    .C1(\cs_registers_i/_1555_ ),
    .B1(\cs_registers_i/_1553_ ),
    .A1(\cs_registers_i/mstack_epc_q_6_ ),
    .Y(\cs_registers_i/_1556_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_4069_  (.A(crash_dump_o_6_),
    .B(net591),
    .Y(\cs_registers_i/_1557_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4070_  (.A1(net591),
    .A2(\cs_registers_i/_1556_ ),
    .Y(\cs_registers_i/_0070_ ),
    .B1(\cs_registers_i/_1557_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4071_  (.A(net1086),
    .B_N(\cs_registers_i/_1346_ ),
    .Y(csr_rdata_7_));
 sg13g2_and2_1 \cs_registers_i/_4072_  (.A(\cs_registers_i/_1326_ ),
    .B(net1302),
    .X(\cs_registers_i/_1558_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4073_  (.A1(csr_op_1_),
    .A2(net155),
    .Y(\cs_registers_i/_1559_ ),
    .B1(\cs_registers_i/_1558_ ));
 sg13g2_nor2_1 \cs_registers_i/_4074_  (.A(net148),
    .B(\cs_registers_i/_1559_ ),
    .Y(\cs_registers_i/_1560_ ));
 sg13g2_a21o_1 \cs_registers_i/_4075_  (.A2(net294),
    .A1(\cs_registers_i/mstack_epc_q_7_ ),
    .B1(\cs_registers_i/_1558_ ),
    .X(\cs_registers_i/_1561_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4076_  (.B2(\cs_registers_i/_1560_ ),
    .C1(\cs_registers_i/_1561_ ),
    .B1(csr_rdata_7_),
    .A1(\cs_registers_i/_1327_ ),
    .Y(\cs_registers_i/_1562_ ),
    .A2(net155));
 sg13g2_nor2_2 \cs_registers_i/_4077_  (.A(crash_dump_o_7_),
    .B(net591),
    .Y(\cs_registers_i/_1563_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4078_  (.A1(net591),
    .A2(\cs_registers_i/_1562_ ),
    .Y(\cs_registers_i/_0071_ ),
    .B1(\cs_registers_i/_1563_ ));
 sg13g2_nand2_1 \cs_registers_i/_4079_  (.Y(\cs_registers_i/_1564_ ),
    .A(net1280),
    .B(net1205));
 sg13g2_inv_1 \cs_registers_i/_4080_  (.Y(\cs_registers_i/_1565_ ),
    .A(net1280));
 sg13g2_mux2_1 \cs_registers_i/_4081_  (.A0(net259),
    .A1(\cs_registers_i/_1352_ ),
    .S(\cs_registers_i/_1399_ ),
    .X(\cs_registers_i/_1566_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4082_  (.Y(\cs_registers_i/_1567_ ),
    .B1(\cs_registers_i/_1566_ ),
    .B2(net256),
    .A2(net155),
    .A1(\cs_registers_i/_1565_ ));
 sg13g2_or3_1 \cs_registers_i/_4083_  (.A(net1091),
    .B(\cs_registers_i/_1367_ ),
    .C(\cs_registers_i/_1567_ ),
    .X(\cs_registers_i/_1568_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4084_  (.Y(\cs_registers_i/_1569_ ),
    .B1(net290),
    .B2(\cs_registers_i/mstack_epc_q_8_ ),
    .A2(net1304),
    .A1(\cs_registers_i/_1352_ ));
 sg13g2_nand3_1 \cs_registers_i/_4085_  (.B(\cs_registers_i/_1568_ ),
    .C(\cs_registers_i/_1569_ ),
    .A(\cs_registers_i/_1564_ ),
    .Y(\cs_registers_i/_1570_ ));
 sg13g2_mux2_1 \cs_registers_i/_4086_  (.A0(crash_dump_o_8_),
    .A1(\cs_registers_i/_1570_ ),
    .S(net594),
    .X(\cs_registers_i/_0072_ ));
 sg13g2_nor2_1 \cs_registers_i/_4087_  (.A(net192),
    .B(\cs_registers_i/_1399_ ),
    .Y(\cs_registers_i/_1571_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4088_  (.Y(\cs_registers_i/_1572_ ),
    .B(\cs_registers_i/_1399_ ),
    .A_N(\cs_registers_i/_1373_ ));
 sg13g2_nand4_1 \cs_registers_i/_4089_  (.B(csr_op_1_),
    .C(csr_op_0_),
    .A(net193),
    .Y(\cs_registers_i/_1573_ ),
    .D(\cs_registers_i/_1417_ ));
 sg13g2_nand3_1 \cs_registers_i/_4090_  (.B(\cs_registers_i/_1572_ ),
    .C(\cs_registers_i/_1573_ ),
    .A(net257),
    .Y(\cs_registers_i/_1574_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4091_  (.A1(\cs_registers_i/_1394_ ),
    .A2(\cs_registers_i/_1571_ ),
    .Y(\cs_registers_i/_1575_ ),
    .B1(\cs_registers_i/_1574_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4092_  (.B2(net1030),
    .C1(\cs_registers_i/_1575_ ),
    .B1(\cs_registers_i/_1420_ ),
    .A1(\cs_registers_i/mstack_epc_q_9_ ),
    .Y(\cs_registers_i/_1576_ ),
    .A2(net295));
 sg13g2_nor2_2 \cs_registers_i/_4093_  (.A(crash_dump_o_9_),
    .B(net597),
    .Y(\cs_registers_i/_1577_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4094_  (.A1(net597),
    .A2(\cs_registers_i/_1576_ ),
    .Y(\cs_registers_i/_0073_ ),
    .B1(\cs_registers_i/_1577_ ));
 sg13g2_nand2_1 \cs_registers_i/_4095_  (.Y(\cs_registers_i/_1578_ ),
    .A(net256),
    .B(\cs_registers_i/_1399_ ));
 sg13g2_buf_8 fanout512 (.A(net518),
    .X(net512));
 sg13g2_buf_4 fanout511 (.X(net511),
    .A(net518));
 sg13g2_nand3_1 \cs_registers_i/_4098_  (.B(net722),
    .C(\cs_registers_i/_0599_ ),
    .A(net1117),
    .Y(\cs_registers_i/_1581_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4099_  (.Y(\cs_registers_i/_1582_ ),
    .B(net344),
    .A_N(net255));
 sg13g2_nand4_1 \cs_registers_i/_4100_  (.B(net1286),
    .C(\cs_registers_i/_1581_ ),
    .A(csr_mstatus_mie),
    .Y(\cs_registers_i/_1583_ ),
    .D(\cs_registers_i/_1582_ ));
 sg13g2_buf_8 fanout510 (.A(net518),
    .X(net510));
 sg13g2_nand2_1 \cs_registers_i/_4102_  (.Y(\cs_registers_i/_1585_ ),
    .A(net1286),
    .B(\cs_registers_i/_1582_ ));
 sg13g2_nor2_2 \cs_registers_i/_4103_  (.A(\cs_registers_i/_1581_ ),
    .B(\cs_registers_i/_1585_ ),
    .Y(\cs_registers_i/_1586_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4104_  (.Y(\cs_registers_i/_1587_ ),
    .B1(net1033),
    .B2(\cs_registers_i/_1586_ ),
    .A2(net346),
    .A1(\cs_registers_i/mstatus_q_4_ ));
 sg13g2_nand2_1 \cs_registers_i/_4105_  (.Y(\cs_registers_i/_0074_ ),
    .A(\cs_registers_i/_1583_ ),
    .B(\cs_registers_i/_1587_ ));
 sg13g2_mux2_1 \cs_registers_i/_4106_  (.A0(net1047),
    .A1(csr_mstatus_tw),
    .S(\cs_registers_i/_1581_ ),
    .X(\cs_registers_i/_0075_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4107_  (.B1(net1391),
    .Y(\cs_registers_i/_1588_ ),
    .A2(\cs_registers_i/_0600_ ),
    .A1(net722));
 sg13g2_and2_1 \cs_registers_i/_4108_  (.A(net2499),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0076_ ));
 sg13g2_buf_8 fanout509 (.A(net518),
    .X(net509));
 sg13g2_buf_8 fanout508 (.A(net518),
    .X(net508));
 sg13g2_nand2_2 \cs_registers_i/_4111_  (.Y(\cs_registers_i/_1591_ ),
    .A(net722),
    .B(\cs_registers_i/_0600_ ));
 sg13g2_buf_4 fanout507 (.X(net507),
    .A(net518));
 sg13g2_buf_4 fanout506 (.X(net506),
    .A(net518));
 sg13g2_buf_4 fanout505 (.X(net505),
    .A(net518));
 sg13g2_nand2b_1 \cs_registers_i/_4115_  (.Y(\cs_registers_i/_1595_ ),
    .B(net653),
    .A_N(csr_mtvec_10_));
 sg13g2_o21ai_1 \cs_registers_i/_4116_  (.B1(\cs_registers_i/_1595_ ),
    .Y(\cs_registers_i/_1596_ ),
    .A1(\cs_registers_i/_0653_ ),
    .A2(net651));
 sg13g2_nand2_1 \cs_registers_i/_4117_  (.Y(\cs_registers_i/_1597_ ),
    .A(boot_addr_i_10_),
    .B(net1388));
 sg13g2_o21ai_1 \cs_registers_i/_4118_  (.B1(\cs_registers_i/_1597_ ),
    .Y(\cs_registers_i/_0077_ ),
    .A1(net1389),
    .A2(\cs_registers_i/_1596_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4119_  (.Y(\cs_registers_i/_1598_ ),
    .B(net646),
    .A_N(csr_mtvec_11_));
 sg13g2_o21ai_1 \cs_registers_i/_4120_  (.B1(\cs_registers_i/_1598_ ),
    .Y(\cs_registers_i/_1599_ ),
    .A1(net1070),
    .A2(net646));
 sg13g2_buf_8 fanout504 (.A(net519),
    .X(net504));
 sg13g2_nand2_1 \cs_registers_i/_4122_  (.Y(\cs_registers_i/_1601_ ),
    .A(net1382),
    .B(boot_addr_i_11_));
 sg13g2_o21ai_1 \cs_registers_i/_4123_  (.B1(\cs_registers_i/_1601_ ),
    .Y(\cs_registers_i/_0078_ ),
    .A1(net1382),
    .A2(\cs_registers_i/_1599_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4124_  (.Y(\cs_registers_i/_1602_ ),
    .B(net651),
    .A_N(csr_mtvec_12_));
 sg13g2_o21ai_1 \cs_registers_i/_4125_  (.B1(\cs_registers_i/_1602_ ),
    .Y(\cs_registers_i/_1603_ ),
    .A1(net1029),
    .A2(net651));
 sg13g2_nand2_1 \cs_registers_i/_4126_  (.Y(\cs_registers_i/_1604_ ),
    .A(net1388),
    .B(boot_addr_i_12_));
 sg13g2_o21ai_1 \cs_registers_i/_4127_  (.B1(\cs_registers_i/_1604_ ),
    .Y(\cs_registers_i/_0079_ ),
    .A1(net1388),
    .A2(\cs_registers_i/_1603_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4128_  (.Y(\cs_registers_i/_1605_ ),
    .B(net647),
    .A_N(csr_mtvec_13_));
 sg13g2_o21ai_1 \cs_registers_i/_4129_  (.B1(\cs_registers_i/_1605_ ),
    .Y(\cs_registers_i/_1606_ ),
    .A1(net1057),
    .A2(net647));
 sg13g2_nand2_1 \cs_registers_i/_4130_  (.Y(\cs_registers_i/_1607_ ),
    .A(net1383),
    .B(boot_addr_i_13_));
 sg13g2_o21ai_1 \cs_registers_i/_4131_  (.B1(\cs_registers_i/_1607_ ),
    .Y(\cs_registers_i/_0080_ ),
    .A1(net1382),
    .A2(\cs_registers_i/_1606_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4132_  (.Y(\cs_registers_i/_1608_ ),
    .B(net646),
    .A_N(csr_mtvec_14_));
 sg13g2_o21ai_1 \cs_registers_i/_4133_  (.B1(\cs_registers_i/_1608_ ),
    .Y(\cs_registers_i/_1609_ ),
    .A1(net1056),
    .A2(net646));
 sg13g2_nand2_1 \cs_registers_i/_4134_  (.Y(\cs_registers_i/_1610_ ),
    .A(net1382),
    .B(boot_addr_i_14_));
 sg13g2_o21ai_1 \cs_registers_i/_4135_  (.B1(\cs_registers_i/_1610_ ),
    .Y(\cs_registers_i/_0081_ ),
    .A1(net1382),
    .A2(\cs_registers_i/_1609_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4136_  (.Y(\cs_registers_i/_1611_ ),
    .B(net647),
    .A_N(csr_mtvec_15_));
 sg13g2_o21ai_1 \cs_registers_i/_4137_  (.B1(\cs_registers_i/_1611_ ),
    .Y(\cs_registers_i/_1612_ ),
    .A1(net1068),
    .A2(net646));
 sg13g2_nand2_1 \cs_registers_i/_4138_  (.Y(\cs_registers_i/_1613_ ),
    .A(net1383),
    .B(boot_addr_i_15_));
 sg13g2_o21ai_1 \cs_registers_i/_4139_  (.B1(\cs_registers_i/_1613_ ),
    .Y(\cs_registers_i/_0082_ ),
    .A1(net1382),
    .A2(\cs_registers_i/_1612_ ));
 sg13g2_buf_8 fanout503 (.A(net519),
    .X(net503));
 sg13g2_nand2b_1 \cs_registers_i/_4141_  (.Y(\cs_registers_i/_1615_ ),
    .B(net652),
    .A_N(csr_mtvec_16_));
 sg13g2_o21ai_1 \cs_registers_i/_4142_  (.B1(\cs_registers_i/_1615_ ),
    .Y(\cs_registers_i/_1616_ ),
    .A1(net1055),
    .A2(net652));
 sg13g2_nand2_1 \cs_registers_i/_4143_  (.Y(\cs_registers_i/_1617_ ),
    .A(net1390),
    .B(boot_addr_i_16_));
 sg13g2_o21ai_1 \cs_registers_i/_4144_  (.B1(\cs_registers_i/_1617_ ),
    .Y(\cs_registers_i/_0083_ ),
    .A1(net1390),
    .A2(\cs_registers_i/_1616_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4145_  (.Y(\cs_registers_i/_1618_ ),
    .B(net649),
    .A_N(csr_mtvec_17_));
 sg13g2_o21ai_1 \cs_registers_i/_4146_  (.B1(\cs_registers_i/_1618_ ),
    .Y(\cs_registers_i/_1619_ ),
    .A1(net1053),
    .A2(net649));
 sg13g2_buf_8 fanout502 (.A(net519),
    .X(net502));
 sg13g2_nand2_1 \cs_registers_i/_4148_  (.Y(\cs_registers_i/_1621_ ),
    .A(net1385),
    .B(boot_addr_i_17_));
 sg13g2_o21ai_1 \cs_registers_i/_4149_  (.B1(\cs_registers_i/_1621_ ),
    .Y(\cs_registers_i/_0084_ ),
    .A1(net1385),
    .A2(\cs_registers_i/_1619_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4150_  (.Y(\cs_registers_i/_1622_ ),
    .B(net652),
    .A_N(csr_mtvec_18_));
 sg13g2_o21ai_1 \cs_registers_i/_4151_  (.B1(\cs_registers_i/_1622_ ),
    .Y(\cs_registers_i/_1623_ ),
    .A1(net1051),
    .A2(net651));
 sg13g2_nand2_1 \cs_registers_i/_4152_  (.Y(\cs_registers_i/_1624_ ),
    .A(net1388),
    .B(boot_addr_i_18_));
 sg13g2_o21ai_1 \cs_registers_i/_4153_  (.B1(\cs_registers_i/_1624_ ),
    .Y(\cs_registers_i/_0085_ ),
    .A1(net1389),
    .A2(\cs_registers_i/_1623_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4154_  (.Y(\cs_registers_i/_1625_ ),
    .B(net651),
    .A_N(csr_mtvec_19_));
 sg13g2_o21ai_1 \cs_registers_i/_4155_  (.B1(\cs_registers_i/_1625_ ),
    .Y(\cs_registers_i/_1626_ ),
    .A1(net1050),
    .A2(net651));
 sg13g2_nand2_1 \cs_registers_i/_4156_  (.Y(\cs_registers_i/_1627_ ),
    .A(net1386),
    .B(boot_addr_i_19_));
 sg13g2_o21ai_1 \cs_registers_i/_4157_  (.B1(\cs_registers_i/_1627_ ),
    .Y(\cs_registers_i/_0086_ ),
    .A1(net1388),
    .A2(\cs_registers_i/_1626_ ));
 sg13g2_and2_1 \cs_registers_i/_4158_  (.A(csr_mtvec_1_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0087_ ));
 sg13g2_buf_4 fanout501 (.X(net501),
    .A(net519));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(net519));
 sg13g2_nand2b_1 \cs_registers_i/_4161_  (.Y(\cs_registers_i/_1630_ ),
    .B(net650),
    .A_N(csr_mtvec_20_));
 sg13g2_o21ai_1 \cs_registers_i/_4162_  (.B1(\cs_registers_i/_1630_ ),
    .Y(\cs_registers_i/_1631_ ),
    .A1(net1049),
    .A2(net650));
 sg13g2_nand2_1 \cs_registers_i/_4163_  (.Y(\cs_registers_i/_1632_ ),
    .A(net1384),
    .B(boot_addr_i_20_));
 sg13g2_o21ai_1 \cs_registers_i/_4164_  (.B1(\cs_registers_i/_1632_ ),
    .Y(\cs_registers_i/_0088_ ),
    .A1(net1384),
    .A2(\cs_registers_i/_1631_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4165_  (.Y(\cs_registers_i/_1633_ ),
    .B(net649),
    .A_N(csr_mtvec_21_));
 sg13g2_o21ai_1 \cs_registers_i/_4166_  (.B1(\cs_registers_i/_1633_ ),
    .Y(\cs_registers_i/_1634_ ),
    .A1(net1047),
    .A2(net653));
 sg13g2_nand2_1 \cs_registers_i/_4167_  (.Y(\cs_registers_i/_1635_ ),
    .A(net1385),
    .B(boot_addr_i_21_));
 sg13g2_o21ai_1 \cs_registers_i/_4168_  (.B1(\cs_registers_i/_1635_ ),
    .Y(\cs_registers_i/_0089_ ),
    .A1(net1386),
    .A2(\cs_registers_i/_1634_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4169_  (.Y(\cs_registers_i/_1636_ ),
    .B(net650),
    .A_N(csr_mtvec_22_));
 sg13g2_o21ai_1 \cs_registers_i/_4170_  (.B1(\cs_registers_i/_1636_ ),
    .Y(\cs_registers_i/_1637_ ),
    .A1(net1027),
    .A2(net650));
 sg13g2_nand2_1 \cs_registers_i/_4171_  (.Y(\cs_registers_i/_1638_ ),
    .A(net1384),
    .B(boot_addr_i_22_));
 sg13g2_o21ai_1 \cs_registers_i/_4172_  (.B1(\cs_registers_i/_1638_ ),
    .Y(\cs_registers_i/_0090_ ),
    .A1(net1387),
    .A2(\cs_registers_i/_1637_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4173_  (.Y(\cs_registers_i/_1639_ ),
    .B(net652),
    .A_N(csr_mtvec_23_));
 sg13g2_o21ai_1 \cs_registers_i/_4174_  (.B1(\cs_registers_i/_1639_ ),
    .Y(\cs_registers_i/_1640_ ),
    .A1(net1046),
    .A2(net652));
 sg13g2_nand2_1 \cs_registers_i/_4175_  (.Y(\cs_registers_i/_1641_ ),
    .A(net1385),
    .B(boot_addr_i_23_));
 sg13g2_o21ai_1 \cs_registers_i/_4176_  (.B1(\cs_registers_i/_1641_ ),
    .Y(\cs_registers_i/_0091_ ),
    .A1(net1388),
    .A2(\cs_registers_i/_1640_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4177_  (.Y(\cs_registers_i/_1642_ ),
    .B(net649),
    .A_N(csr_mtvec_24_));
 sg13g2_o21ai_1 \cs_registers_i/_4178_  (.B1(\cs_registers_i/_1642_ ),
    .Y(\cs_registers_i/_1643_ ),
    .A1(net1044),
    .A2(net653));
 sg13g2_nand2_1 \cs_registers_i/_4179_  (.Y(\cs_registers_i/_1644_ ),
    .A(net1385),
    .B(boot_addr_i_24_));
 sg13g2_o21ai_1 \cs_registers_i/_4180_  (.B1(\cs_registers_i/_1644_ ),
    .Y(\cs_registers_i/_0092_ ),
    .A1(net1386),
    .A2(\cs_registers_i/_1643_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4181_  (.Y(\cs_registers_i/_1645_ ),
    .B(net652),
    .A_N(csr_mtvec_25_));
 sg13g2_o21ai_1 \cs_registers_i/_4182_  (.B1(\cs_registers_i/_1645_ ),
    .Y(\cs_registers_i/_1646_ ),
    .A1(net1043),
    .A2(net652));
 sg13g2_nand2_1 \cs_registers_i/_4183_  (.Y(\cs_registers_i/_1647_ ),
    .A(net1389),
    .B(boot_addr_i_25_));
 sg13g2_o21ai_1 \cs_registers_i/_4184_  (.B1(\cs_registers_i/_1647_ ),
    .Y(\cs_registers_i/_0093_ ),
    .A1(net1389),
    .A2(\cs_registers_i/_1646_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4185_  (.Y(\cs_registers_i/_1648_ ),
    .B(net649),
    .A_N(csr_mtvec_26_));
 sg13g2_o21ai_1 \cs_registers_i/_4186_  (.B1(\cs_registers_i/_1648_ ),
    .Y(\cs_registers_i/_1649_ ),
    .A1(net1066),
    .A2(net649));
 sg13g2_nand2_1 \cs_registers_i/_4187_  (.Y(\cs_registers_i/_1650_ ),
    .A(net1385),
    .B(boot_addr_i_26_));
 sg13g2_o21ai_1 \cs_registers_i/_4188_  (.B1(\cs_registers_i/_1650_ ),
    .Y(\cs_registers_i/_0094_ ),
    .A1(net1385),
    .A2(\cs_registers_i/_1649_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4189_  (.Y(\cs_registers_i/_1651_ ),
    .B(net650),
    .A_N(csr_mtvec_27_));
 sg13g2_o21ai_1 \cs_registers_i/_4190_  (.B1(\cs_registers_i/_1651_ ),
    .Y(\cs_registers_i/_1652_ ),
    .A1(net1026),
    .A2(net650));
 sg13g2_nand2_1 \cs_registers_i/_4191_  (.Y(\cs_registers_i/_1653_ ),
    .A(net1384),
    .B(boot_addr_i_27_));
 sg13g2_o21ai_1 \cs_registers_i/_4192_  (.B1(\cs_registers_i/_1653_ ),
    .Y(\cs_registers_i/_0095_ ),
    .A1(net1384),
    .A2(\cs_registers_i/_1652_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4193_  (.Y(\cs_registers_i/_1654_ ),
    .B(net650),
    .A_N(csr_mtvec_28_));
 sg13g2_o21ai_1 \cs_registers_i/_4194_  (.B1(\cs_registers_i/_1654_ ),
    .Y(\cs_registers_i/_1655_ ),
    .A1(net1042),
    .A2(net650));
 sg13g2_nand2_1 \cs_registers_i/_4195_  (.Y(\cs_registers_i/_1656_ ),
    .A(net1384),
    .B(boot_addr_i_28_));
 sg13g2_o21ai_1 \cs_registers_i/_4196_  (.B1(\cs_registers_i/_1656_ ),
    .Y(\cs_registers_i/_0096_ ),
    .A1(net1387),
    .A2(\cs_registers_i/_1655_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4197_  (.Y(\cs_registers_i/_1657_ ),
    .B(net649),
    .A_N(csr_mtvec_29_));
 sg13g2_o21ai_1 \cs_registers_i/_4198_  (.B1(\cs_registers_i/_1657_ ),
    .Y(\cs_registers_i/_1658_ ),
    .A1(net1040),
    .A2(net649));
 sg13g2_nand2_1 \cs_registers_i/_4199_  (.Y(\cs_registers_i/_1659_ ),
    .A(net1385),
    .B(boot_addr_i_29_));
 sg13g2_o21ai_1 \cs_registers_i/_4200_  (.B1(\cs_registers_i/_1659_ ),
    .Y(\cs_registers_i/_0097_ ),
    .A1(net1386),
    .A2(\cs_registers_i/_1658_ ));
 sg13g2_and2_1 \cs_registers_i/_4201_  (.A(csr_mtvec_2_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0098_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4202_  (.Y(\cs_registers_i/_1660_ ),
    .B(net646),
    .A_N(csr_mtvec_30_));
 sg13g2_o21ai_1 \cs_registers_i/_4203_  (.B1(\cs_registers_i/_1660_ ),
    .Y(\cs_registers_i/_1661_ ),
    .A1(net1037),
    .A2(net647));
 sg13g2_nand2_1 \cs_registers_i/_4204_  (.Y(\cs_registers_i/_1662_ ),
    .A(net1382),
    .B(boot_addr_i_30_));
 sg13g2_o21ai_1 \cs_registers_i/_4205_  (.B1(\cs_registers_i/_1662_ ),
    .Y(\cs_registers_i/_0099_ ),
    .A1(net1383),
    .A2(\cs_registers_i/_1661_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4206_  (.Y(\cs_registers_i/_1663_ ),
    .B(net651),
    .A_N(csr_mtvec_31_));
 sg13g2_o21ai_1 \cs_registers_i/_4207_  (.B1(\cs_registers_i/_1663_ ),
    .Y(\cs_registers_i/_1664_ ),
    .A1(net1035),
    .A2(net651));
 sg13g2_nand2_1 \cs_registers_i/_4208_  (.Y(\cs_registers_i/_1665_ ),
    .A(net1388),
    .B(boot_addr_i_31_));
 sg13g2_o21ai_1 \cs_registers_i/_4209_  (.B1(\cs_registers_i/_1665_ ),
    .Y(\cs_registers_i/_0100_ ),
    .A1(net1388),
    .A2(\cs_registers_i/_1664_ ));
 sg13g2_and2_1 \cs_registers_i/_4210_  (.A(csr_mtvec_3_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0101_ ));
 sg13g2_and2_1 \cs_registers_i/_4211_  (.A(csr_mtvec_4_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0102_ ));
 sg13g2_and2_1 \cs_registers_i/_4212_  (.A(csr_mtvec_5_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0103_ ));
 sg13g2_and2_1 \cs_registers_i/_4213_  (.A(csr_mtvec_6_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0104_ ));
 sg13g2_and2_1 \cs_registers_i/_4214_  (.A(csr_mtvec_7_),
    .B(\cs_registers_i/_1588_ ),
    .X(\cs_registers_i/_0105_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4215_  (.Y(\cs_registers_i/_1666_ ),
    .B(net646),
    .A_N(csr_mtvec_8_));
 sg13g2_o21ai_1 \cs_registers_i/_4216_  (.B1(\cs_registers_i/_1666_ ),
    .Y(\cs_registers_i/_1667_ ),
    .A1(net1025),
    .A2(net646));
 sg13g2_nand2_1 \cs_registers_i/_4217_  (.Y(\cs_registers_i/_1668_ ),
    .A(net1382),
    .B(boot_addr_i_8_));
 sg13g2_o21ai_1 \cs_registers_i/_4218_  (.B1(\cs_registers_i/_1668_ ),
    .Y(\cs_registers_i/_0106_ ),
    .A1(net1383),
    .A2(\cs_registers_i/_1667_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4219_  (.Y(\cs_registers_i/_1669_ ),
    .B(net648),
    .A_N(csr_mtvec_9_));
 sg13g2_o21ai_1 \cs_registers_i/_4220_  (.B1(\cs_registers_i/_1669_ ),
    .Y(\cs_registers_i/_1670_ ),
    .A1(net1030),
    .A2(net648));
 sg13g2_nand2_1 \cs_registers_i/_4221_  (.Y(\cs_registers_i/_1671_ ),
    .A(net1384),
    .B(boot_addr_i_9_));
 sg13g2_o21ai_1 \cs_registers_i/_4222_  (.B1(\cs_registers_i/_1671_ ),
    .Y(\cs_registers_i/_0107_ ),
    .A1(net1384),
    .A2(\cs_registers_i/_1670_ ));
 sg13g2_buf_4 fanout499 (.X(net499),
    .A(net519));
 sg13g2_nor2_1 \cs_registers_i/_4224_  (.A(net1084),
    .B(\cs_registers_i/_1242_ ),
    .Y(csr_rdata_31_));
 sg13g2_nor2b_1 \cs_registers_i/_4225_  (.A(net1084),
    .B_N(\cs_registers_i/_1221_ ),
    .Y(csr_rdata_30_));
 sg13g2_nor2_1 \cs_registers_i/_4226_  (.A(net1087),
    .B(\cs_registers_i/_0981_ ),
    .Y(csr_rdata_21_));
 sg13g2_nor2_1 \cs_registers_i/_4227_  (.A(net1085),
    .B(\cs_registers_i/_0959_ ),
    .Y(csr_rdata_20_));
 sg13g2_nor2_1 \cs_registers_i/_4228_  (.A(net1084),
    .B(\cs_registers_i/_0901_ ),
    .Y(csr_rdata_19_));
 sg13g2_nor2_1 \cs_registers_i/_4229_  (.A(net1084),
    .B(\cs_registers_i/_0881_ ),
    .Y(csr_rdata_18_));
 sg13g2_nor2_1 \cs_registers_i/_4230_  (.A(net1087),
    .B(\cs_registers_i/_0858_ ),
    .Y(csr_rdata_17_));
 sg13g2_nor2_1 \cs_registers_i/_4231_  (.A(net1087),
    .B(\cs_registers_i/_0832_ ),
    .Y(csr_rdata_16_));
 sg13g2_nor2_1 \cs_registers_i/_4232_  (.A(net1084),
    .B(\cs_registers_i/_0806_ ),
    .Y(csr_rdata_15_));
 sg13g2_buf_8 fanout498 (.A(net519),
    .X(net498));
 sg13g2_nor2_1 \cs_registers_i/_4234_  (.A(net1083),
    .B(\cs_registers_i/_0788_ ),
    .Y(csr_rdata_14_));
 sg13g2_nor2_1 \cs_registers_i/_4235_  (.A(net1084),
    .B(\cs_registers_i/_0762_ ),
    .Y(csr_rdata_13_));
 sg13g2_nor2_1 \cs_registers_i/_4236_  (.A(net1084),
    .B(\cs_registers_i/_0736_ ),
    .Y(csr_rdata_12_));
 sg13g2_nor2_1 \cs_registers_i/_4237_  (.A(net1083),
    .B(\cs_registers_i/_0696_ ),
    .Y(csr_rdata_11_));
 sg13g2_nor2_1 \cs_registers_i/_4238_  (.A(net1084),
    .B(\cs_registers_i/_0651_ ),
    .Y(csr_rdata_10_));
 sg13g2_nor2b_1 \cs_registers_i/_4239_  (.A(net1082),
    .B_N(\cs_registers_i/_1393_ ),
    .Y(csr_rdata_9_));
 sg13g2_nor2_1 \cs_registers_i/_4240_  (.A(net1082),
    .B(\cs_registers_i/_1367_ ),
    .Y(csr_rdata_8_));
 sg13g2_nor2_1 \cs_registers_i/_4241_  (.A(net1082),
    .B(\cs_registers_i/_1320_ ),
    .Y(csr_rdata_6_));
 sg13g2_nor2_1 \cs_registers_i/_4242_  (.A(net1082),
    .B(\cs_registers_i/_1302_ ),
    .Y(csr_rdata_5_));
 sg13g2_nor2_1 \cs_registers_i/_4243_  (.A(net1082),
    .B(\cs_registers_i/_1284_ ),
    .Y(csr_rdata_4_));
 sg13g2_nor2_1 \cs_registers_i/_4244_  (.A(net1082),
    .B(\cs_registers_i/_1270_ ),
    .Y(csr_rdata_3_));
 sg13g2_buf_4 fanout497 (.X(net497),
    .A(net519));
 sg13g2_nor2_1 \cs_registers_i/_4246_  (.A(net1082),
    .B(\cs_registers_i/_1201_ ),
    .Y(csr_rdata_2_));
 sg13g2_nor2_1 \cs_registers_i/_4247_  (.A(net1087),
    .B(\cs_registers_i/_1150_ ),
    .Y(csr_rdata_28_));
 sg13g2_nor2_1 \cs_registers_i/_4248_  (.A(net1082),
    .B(\cs_registers_i/_0930_ ),
    .Y(csr_rdata_1_));
 sg13g2_a21o_1 \cs_registers_i/_4249_  (.A2(\cs_registers_i/_0818_ ),
    .A1(hart_id_i_0_),
    .B1(\cs_registers_i/_1290_ ),
    .X(\cs_registers_i/_1675_ ));
 sg13g2_nand3_1 \cs_registers_i/_4250_  (.B(\cs_registers_i/_0923_ ),
    .C(\cs_registers_i/_1675_ ),
    .A(net54),
    .Y(\cs_registers_i/_1676_ ));
 sg13g2_nand2_1 \cs_registers_i/_4251_  (.Y(\cs_registers_i/_1677_ ),
    .A(csr_mtvec_0_),
    .B(\cs_registers_i/_0749_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4252_  (.Y(\cs_registers_i/_1678_ ),
    .B1(\cs_registers_i/_0678_ ),
    .B2(\cs_registers_i/mtval_q_0_ ),
    .A2(net1119),
    .A1(\cs_registers_i/mcountinhibit_0_ ));
 sg13g2_a21o_1 \cs_registers_i/_4253_  (.A2(\cs_registers_i/_1678_ ),
    .A1(\cs_registers_i/_1677_ ),
    .B1(net1172),
    .X(\cs_registers_i/_1679_ ));
 sg13g2_mux4_1 \cs_registers_i/_4254_  (.S0(net62),
    .A0(\cs_registers_i/dcsr_q_0_ ),
    .A1(\cs_registers_i/dscratch0_q_0_ ),
    .A2(csr_depc_0_),
    .A3(\cs_registers_i/dscratch1_q_0_ ),
    .S1(net1232),
    .X(\cs_registers_i/_1680_ ));
 sg13g2_nand2_1 \cs_registers_i/_4255_  (.Y(\cs_registers_i/_1681_ ),
    .A(net1150),
    .B(\cs_registers_i/_1680_ ));
 sg13g2_and2_1 \cs_registers_i/_4256_  (.A(crash_dump_o_0_),
    .B(net1231),
    .X(\cs_registers_i/_1682_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4257_  (.A1(net53),
    .A2(\cs_registers_i/mscratch_q_0_ ),
    .Y(\cs_registers_i/_1683_ ),
    .B1(\cs_registers_i/_1682_ ));
 sg13g2_nand3_1 \cs_registers_i/_4258_  (.B(net53),
    .C(\cs_registers_i/mcause_q_0_ ),
    .A(net76),
    .Y(\cs_registers_i/_1684_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4259_  (.B1(\cs_registers_i/_1684_ ),
    .Y(\cs_registers_i/_1685_ ),
    .A1(net64),
    .A2(\cs_registers_i/_1683_ ));
 sg13g2_mux4_1 \cs_registers_i/_4260_  (.S0(net62),
    .A0(\cs_registers_i/mcycle_counter_i.counter_val_o_0_ ),
    .A1(\cs_registers_i/mhpmcounter_1856_ ),
    .A2(\cs_registers_i/mcycle_counter_i.counter_val_o_32_ ),
    .A3(\cs_registers_i/mhpmcounter_1888_ ),
    .S1(net147),
    .X(\cs_registers_i/_1686_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4261_  (.Y(\cs_registers_i/_1687_ ),
    .B1(\cs_registers_i/_1686_ ),
    .B2(\cs_registers_i/_0877_ ),
    .A2(\cs_registers_i/_1685_ ),
    .A1(\cs_registers_i/_0605_ ));
 sg13g2_and4_2 \cs_registers_i/_4262_  (.A(\cs_registers_i/_1676_ ),
    .B(\cs_registers_i/_1679_ ),
    .C(\cs_registers_i/_1681_ ),
    .D(\cs_registers_i/_1687_ ),
    .X(\cs_registers_i/_1688_ ));
 sg13g2_nor2_1 \cs_registers_i/_4263_  (.A(net1083),
    .B(\cs_registers_i/_1688_ ),
    .Y(csr_rdata_0_));
 sg13g2_nor2_1 \cs_registers_i/_4264_  (.A(net1086),
    .B(\cs_registers_i/_1126_ ),
    .Y(csr_rdata_27_));
 sg13g2_nor2_1 \cs_registers_i/_4265_  (.A(net1085),
    .B(\cs_registers_i/_1098_ ),
    .Y(csr_rdata_26_));
 sg13g2_nor2_1 \cs_registers_i/_4266_  (.A(net1086),
    .B(\cs_registers_i/_1077_ ),
    .Y(csr_rdata_25_));
 sg13g2_nor2_1 \cs_registers_i/_4267_  (.A(net1085),
    .B(\cs_registers_i/_1050_ ),
    .Y(csr_rdata_24_));
 sg13g2_nor2_1 \cs_registers_i/_4268_  (.A(net1083),
    .B(\cs_registers_i/_1029_ ),
    .Y(csr_rdata_23_));
 sg13g2_nor2_1 \cs_registers_i/_4269_  (.A(net1087),
    .B(\cs_registers_i/_1007_ ),
    .Y(csr_rdata_22_));
 sg13g2_nand2_1 \cs_registers_i/_4270_  (.Y(\cs_registers_i/_1689_ ),
    .A(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .B(net1313));
 sg13g2_nand3_1 \cs_registers_i/_4271_  (.B(net1117),
    .C(\cs_registers_i/_0580_ ),
    .A(net60),
    .Y(\cs_registers_i/_1690_ ));
 sg13g2_buf_4 fanout496 (.X(net496),
    .A(net520));
 sg13g2_nand2_1 \cs_registers_i/_4273_  (.Y(\cs_registers_i/_1692_ ),
    .A(\cs_registers_i/_0002_ ),
    .B(net642));
 sg13g2_nor3_1 \cs_registers_i/_4274_  (.A(net197),
    .B(net1088),
    .C(\cs_registers_i/_1688_ ),
    .Y(\cs_registers_i/_1693_ ));
 sg13g2_a21o_2 \cs_registers_i/_4275_  (.A2(net259),
    .A1(net198),
    .B1(\cs_registers_i/_1693_ ),
    .X(\cs_registers_i/_1694_ ));
 sg13g2_or3_1 \cs_registers_i/_4276_  (.A(net1067),
    .B(net642),
    .C(net1063),
    .X(\cs_registers_i/_1695_ ));
 sg13g2_nand3_1 \cs_registers_i/_4277_  (.B(\cs_registers_i/_1692_ ),
    .C(\cs_registers_i/_1695_ ),
    .A(\cs_registers_i/_0655_ ),
    .Y(\cs_registers_i/_1696_ ));
 sg13g2_and2_1 \cs_registers_i/_4278_  (.A(\cs_registers_i/_1689_ ),
    .B(\cs_registers_i/_1696_ ),
    .X(\cs_registers_i/_0108_ ));
 sg13g2_buf_8 fanout495 (.A(net520),
    .X(net495));
 sg13g2_and2_1 \cs_registers_i/_4280_  (.A(\cs_registers_i/dcsr_q_10_ ),
    .B(net642),
    .X(\cs_registers_i/_0109_ ));
 sg13g2_and2_1 \cs_registers_i/_4281_  (.A(\cs_registers_i/dcsr_q_11_ ),
    .B(net644),
    .X(\cs_registers_i/_0110_ ));
 sg13g2_mux2_1 \cs_registers_i/_4282_  (.A0(net1057),
    .A1(\cs_registers_i/dcsr_q_13_ ),
    .S(net642),
    .X(\cs_registers_i/_0111_ ));
 sg13g2_and2_1 \cs_registers_i/_4283_  (.A(\cs_registers_i/dcsr_q_14_ ),
    .B(net643),
    .X(\cs_registers_i/_0112_ ));
 sg13g2_and2_1 \cs_registers_i/_4284_  (.A(\cs_registers_i/dcsr_q_16_ ),
    .B(net643),
    .X(\cs_registers_i/_0113_ ));
 sg13g2_and2_1 \cs_registers_i/_4285_  (.A(\cs_registers_i/dcsr_q_17_ ),
    .B(net644),
    .X(\cs_registers_i/_0114_ ));
 sg13g2_and2_1 \cs_registers_i/_4286_  (.A(\cs_registers_i/dcsr_q_18_ ),
    .B(net642),
    .X(\cs_registers_i/_0115_ ));
 sg13g2_and2_1 \cs_registers_i/_4287_  (.A(\cs_registers_i/dcsr_q_19_ ),
    .B(net644),
    .X(\cs_registers_i/_0116_ ));
 sg13g2_nand2_1 \cs_registers_i/_4288_  (.Y(\cs_registers_i/_1698_ ),
    .A(net2116),
    .B(net1312));
 sg13g2_nand2_1 \cs_registers_i/_4289_  (.Y(\cs_registers_i/_1699_ ),
    .A(\cs_registers_i/_0003_ ),
    .B(net643));
 sg13g2_nand3_1 \cs_registers_i/_4290_  (.B(\cs_registers_i/_1695_ ),
    .C(\cs_registers_i/_1699_ ),
    .A(\cs_registers_i/_0655_ ),
    .Y(\cs_registers_i/_1700_ ));
 sg13g2_and2_1 \cs_registers_i/_4291_  (.A(\cs_registers_i/_1698_ ),
    .B(\cs_registers_i/_1700_ ),
    .X(\cs_registers_i/_0117_ ));
 sg13g2_and2_1 \cs_registers_i/_4292_  (.A(\cs_registers_i/dcsr_q_20_ ),
    .B(net644),
    .X(\cs_registers_i/_0118_ ));
 sg13g2_and2_1 \cs_registers_i/_4293_  (.A(\cs_registers_i/dcsr_q_21_ ),
    .B(net644),
    .X(\cs_registers_i/_0119_ ));
 sg13g2_and2_1 \cs_registers_i/_4294_  (.A(\cs_registers_i/dcsr_q_22_ ),
    .B(net644),
    .X(\cs_registers_i/_0120_ ));
 sg13g2_buf_8 fanout494 (.A(net520),
    .X(net494));
 sg13g2_and2_1 \cs_registers_i/_4296_  (.A(\cs_registers_i/dcsr_q_23_ ),
    .B(net643),
    .X(\cs_registers_i/_0121_ ));
 sg13g2_and2_1 \cs_registers_i/_4297_  (.A(\cs_registers_i/dcsr_q_24_ ),
    .B(net645),
    .X(\cs_registers_i/_0122_ ));
 sg13g2_and2_1 \cs_registers_i/_4298_  (.A(\cs_registers_i/dcsr_q_25_ ),
    .B(net645),
    .X(\cs_registers_i/_0123_ ));
 sg13g2_and2_1 \cs_registers_i/_4299_  (.A(net2498),
    .B(net645),
    .X(\cs_registers_i/_0124_ ));
 sg13g2_and2_1 \cs_registers_i/_4300_  (.A(\cs_registers_i/dcsr_q_27_ ),
    .B(net644),
    .X(\cs_registers_i/_0125_ ));
 sg13g2_and2_1 \cs_registers_i/_4301_  (.A(\cs_registers_i/dcsr_q_28_ ),
    .B(net645),
    .X(\cs_registers_i/_0126_ ));
 sg13g2_and2_1 \cs_registers_i/_4302_  (.A(\cs_registers_i/dcsr_q_29_ ),
    .B(net645),
    .X(\cs_registers_i/_0127_ ));
 sg13g2_nor2_1 \cs_registers_i/_4303_  (.A(\cs_registers_i/_0004_ ),
    .B(net1313),
    .Y(\cs_registers_i/_1702_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4304_  (.B2(\cs_registers_i/_0581_ ),
    .C1(\cs_registers_i/_1702_ ),
    .B1(net1117),
    .A1(\cs_registers_i/dcsr_q_30_ ),
    .Y(\cs_registers_i/_0128_ ),
    .A2(net1313));
 sg13g2_and2_1 \cs_registers_i/_4305_  (.A(\cs_registers_i/dcsr_q_31_ ),
    .B(net645),
    .X(\cs_registers_i/_0129_ ));
 sg13g2_and2_1 \cs_registers_i/_4306_  (.A(\cs_registers_i/dcsr_q_3_ ),
    .B(net643),
    .X(\cs_registers_i/_0130_ ));
 sg13g2_and2_1 \cs_registers_i/_4307_  (.A(\cs_registers_i/dcsr_q_4_ ),
    .B(net643),
    .X(\cs_registers_i/_0131_ ));
 sg13g2_and2_1 \cs_registers_i/_4308_  (.A(\cs_registers_i/dcsr_q_5_ ),
    .B(net642),
    .X(\cs_registers_i/_0132_ ));
 sg13g2_mux2_1 \cs_registers_i/_4309_  (.A0(\cs_registers_i/dcsr_q_6_ ),
    .A1(debug_cause_0_),
    .S(net1313),
    .X(\cs_registers_i/_0133_ ));
 sg13g2_mux2_1 \cs_registers_i/_4310_  (.A0(\cs_registers_i/dcsr_q_7_ ),
    .A1(debug_cause_1_),
    .S(net1313),
    .X(\cs_registers_i/_0134_ ));
 sg13g2_mux2_1 \cs_registers_i/_4311_  (.A0(\cs_registers_i/dcsr_q_8_ ),
    .A1(debug_cause_2_),
    .S(net1313),
    .X(\cs_registers_i/_0135_ ));
 sg13g2_and2_1 \cs_registers_i/_4312_  (.A(\cs_registers_i/dcsr_q_9_ ),
    .B(net642),
    .X(\cs_registers_i/_0136_ ));
 sg13g2_mux2_1 \cs_registers_i/_4313_  (.A0(net1068),
    .A1(debug_ebreakm),
    .S(net642),
    .X(\cs_registers_i/_0137_ ));
 sg13g2_mux2_1 \cs_registers_i/_4314_  (.A0(net1029),
    .A1(debug_ebreaku),
    .S(net645),
    .X(\cs_registers_i/_0138_ ));
 sg13g2_mux2_1 \cs_registers_i/_4315_  (.A0(net1039),
    .A1(debug_single_step),
    .S(net644),
    .X(\cs_registers_i/_0139_ ));
 sg13g2_nand2_2 \cs_registers_i/_4316_  (.Y(\cs_registers_i/_1703_ ),
    .A(\cs_registers_i/_0581_ ),
    .B(\cs_registers_i/_1061_ ));
 sg13g2_buf_4 fanout493 (.X(net493),
    .A(net520));
 sg13g2_mux2_1 \cs_registers_i/_4318_  (.A0(net1063),
    .A1(\cs_registers_i/dscratch0_q_0_ ),
    .S(net637),
    .X(\cs_registers_i/_0140_ ));
 sg13g2_mux2_1 \cs_registers_i/_4319_  (.A0(net1059),
    .A1(\cs_registers_i/dscratch0_q_10_ ),
    .S(net637),
    .X(\cs_registers_i/_0141_ ));
 sg13g2_mux2_1 \cs_registers_i/_4320_  (.A0(net1071),
    .A1(\cs_registers_i/dscratch0_q_11_ ),
    .S(net639),
    .X(\cs_registers_i/_0142_ ));
 sg13g2_mux2_1 \cs_registers_i/_4321_  (.A0(net1029),
    .A1(\cs_registers_i/dscratch0_q_12_ ),
    .S(\cs_registers_i/_1703_ ),
    .X(\cs_registers_i/_0143_ ));
 sg13g2_mux2_1 \cs_registers_i/_4322_  (.A0(net1057),
    .A1(\cs_registers_i/dscratch0_q_13_ ),
    .S(net637),
    .X(\cs_registers_i/_0144_ ));
 sg13g2_mux2_1 \cs_registers_i/_4323_  (.A0(\cs_registers_i/_0790_ ),
    .A1(\cs_registers_i/dscratch0_q_14_ ),
    .S(net638),
    .X(\cs_registers_i/_0145_ ));
 sg13g2_mux2_1 \cs_registers_i/_4324_  (.A0(net1068),
    .A1(\cs_registers_i/dscratch0_q_15_ ),
    .S(net637),
    .X(\cs_registers_i/_0146_ ));
 sg13g2_mux2_1 \cs_registers_i/_4325_  (.A0(net1055),
    .A1(\cs_registers_i/dscratch0_q_16_ ),
    .S(net637),
    .X(\cs_registers_i/_0147_ ));
 sg13g2_mux2_1 \cs_registers_i/_4326_  (.A0(net1054),
    .A1(\cs_registers_i/dscratch0_q_17_ ),
    .S(net639),
    .X(\cs_registers_i/_0148_ ));
 sg13g2_mux2_1 \cs_registers_i/_4327_  (.A0(net1051),
    .A1(\cs_registers_i/dscratch0_q_18_ ),
    .S(net637),
    .X(\cs_registers_i/_0149_ ));
 sg13g2_buf_8 fanout492 (.A(net520),
    .X(net492));
 sg13g2_mux2_1 \cs_registers_i/_4329_  (.A0(\cs_registers_i/_0903_ ),
    .A1(\cs_registers_i/dscratch0_q_19_ ),
    .S(net639),
    .X(\cs_registers_i/_0150_ ));
 sg13g2_mux2_1 \cs_registers_i/_4330_  (.A0(\cs_registers_i/_0932_ ),
    .A1(\cs_registers_i/dscratch0_q_1_ ),
    .S(net638),
    .X(\cs_registers_i/_0151_ ));
 sg13g2_mux2_1 \cs_registers_i/_4331_  (.A0(\cs_registers_i/_0961_ ),
    .A1(\cs_registers_i/dscratch0_q_20_ ),
    .S(net639),
    .X(\cs_registers_i/_0152_ ));
 sg13g2_mux2_1 \cs_registers_i/_4332_  (.A0(net1048),
    .A1(\cs_registers_i/dscratch0_q_21_ ),
    .S(net640),
    .X(\cs_registers_i/_0153_ ));
 sg13g2_mux2_1 \cs_registers_i/_4333_  (.A0(\cs_registers_i/_1009_ ),
    .A1(\cs_registers_i/dscratch0_q_22_ ),
    .S(net640),
    .X(\cs_registers_i/_0154_ ));
 sg13g2_mux2_1 \cs_registers_i/_4334_  (.A0(net1046),
    .A1(\cs_registers_i/dscratch0_q_23_ ),
    .S(net638),
    .X(\cs_registers_i/_0155_ ));
 sg13g2_mux2_1 \cs_registers_i/_4335_  (.A0(net1045),
    .A1(\cs_registers_i/dscratch0_q_24_ ),
    .S(net639),
    .X(\cs_registers_i/_0156_ ));
 sg13g2_mux2_1 \cs_registers_i/_4336_  (.A0(\cs_registers_i/_1079_ ),
    .A1(\cs_registers_i/dscratch0_q_25_ ),
    .S(net641),
    .X(\cs_registers_i/_0157_ ));
 sg13g2_mux2_1 \cs_registers_i/_4337_  (.A0(\cs_registers_i/_1100_ ),
    .A1(\cs_registers_i/dscratch0_q_26_ ),
    .S(net641),
    .X(\cs_registers_i/_0158_ ));
 sg13g2_mux2_1 \cs_registers_i/_4338_  (.A0(\cs_registers_i/_1128_ ),
    .A1(\cs_registers_i/dscratch0_q_27_ ),
    .S(net639),
    .X(\cs_registers_i/_0159_ ));
 sg13g2_buf_8 fanout491 (.A(net520),
    .X(net491));
 sg13g2_mux2_1 \cs_registers_i/_4340_  (.A0(\cs_registers_i/_1152_ ),
    .A1(\cs_registers_i/dscratch0_q_28_ ),
    .S(net641),
    .X(\cs_registers_i/_0160_ ));
 sg13g2_mux2_1 \cs_registers_i/_4341_  (.A0(net1041),
    .A1(\cs_registers_i/dscratch0_q_29_ ),
    .S(net638),
    .X(\cs_registers_i/_0161_ ));
 sg13g2_mux2_1 \cs_registers_i/_4342_  (.A0(net1038),
    .A1(\cs_registers_i/dscratch0_q_2_ ),
    .S(net639),
    .X(\cs_registers_i/_0162_ ));
 sg13g2_mux2_1 \cs_registers_i/_4343_  (.A0(\cs_registers_i/_1224_ ),
    .A1(\cs_registers_i/dscratch0_q_30_ ),
    .S(net640),
    .X(\cs_registers_i/_0163_ ));
 sg13g2_mux2_1 \cs_registers_i/_4344_  (.A0(net1036),
    .A1(\cs_registers_i/dscratch0_q_31_ ),
    .S(net639),
    .X(\cs_registers_i/_0164_ ));
 sg13g2_mux2_1 \cs_registers_i/_4345_  (.A0(net1034),
    .A1(\cs_registers_i/dscratch0_q_3_ ),
    .S(net641),
    .X(\cs_registers_i/_0165_ ));
 sg13g2_mux2_1 \cs_registers_i/_4346_  (.A0(net1032),
    .A1(\cs_registers_i/dscratch0_q_4_ ),
    .S(net638),
    .X(\cs_registers_i/_0166_ ));
 sg13g2_mux2_1 \cs_registers_i/_4347_  (.A0(\cs_registers_i/_1304_ ),
    .A1(\cs_registers_i/dscratch0_q_5_ ),
    .S(net637),
    .X(\cs_registers_i/_0167_ ));
 sg13g2_mux2_1 \cs_registers_i/_4348_  (.A0(\cs_registers_i/_1322_ ),
    .A1(\cs_registers_i/dscratch0_q_6_ ),
    .S(net641),
    .X(\cs_registers_i/_0168_ ));
 sg13g2_mux2_1 \cs_registers_i/_4349_  (.A0(\cs_registers_i/_1348_ ),
    .A1(\cs_registers_i/dscratch0_q_7_ ),
    .S(net640),
    .X(\cs_registers_i/_0169_ ));
 sg13g2_mux2_1 \cs_registers_i/_4350_  (.A0(\cs_registers_i/_1369_ ),
    .A1(\cs_registers_i/dscratch0_q_8_ ),
    .S(net641),
    .X(\cs_registers_i/_0170_ ));
 sg13g2_mux2_1 \cs_registers_i/_4351_  (.A0(net1030),
    .A1(\cs_registers_i/dscratch0_q_9_ ),
    .S(net637),
    .X(\cs_registers_i/_0171_ ));
 sg13g2_nand2_2 \cs_registers_i/_4352_  (.Y(\cs_registers_i/_1707_ ),
    .A(\cs_registers_i/_0581_ ),
    .B(\cs_registers_i/_0948_ ));
 sg13g2_buf_8 fanout490 (.A(net520),
    .X(net490));
 sg13g2_mux2_1 \cs_registers_i/_4354_  (.A0(net1063),
    .A1(\cs_registers_i/dscratch1_q_0_ ),
    .S(net631),
    .X(\cs_registers_i/_0172_ ));
 sg13g2_mux2_1 \cs_registers_i/_4355_  (.A0(net1059),
    .A1(\cs_registers_i/dscratch1_q_10_ ),
    .S(net631),
    .X(\cs_registers_i/_0173_ ));
 sg13g2_mux2_1 \cs_registers_i/_4356_  (.A0(net1071),
    .A1(\cs_registers_i/dscratch1_q_11_ ),
    .S(net633),
    .X(\cs_registers_i/_0174_ ));
 sg13g2_mux2_1 \cs_registers_i/_4357_  (.A0(net1029),
    .A1(\cs_registers_i/dscratch1_q_12_ ),
    .S(net636),
    .X(\cs_registers_i/_0175_ ));
 sg13g2_mux2_1 \cs_registers_i/_4358_  (.A0(net1057),
    .A1(\cs_registers_i/dscratch1_q_13_ ),
    .S(net631),
    .X(\cs_registers_i/_0176_ ));
 sg13g2_mux2_1 \cs_registers_i/_4359_  (.A0(\cs_registers_i/_0790_ ),
    .A1(\cs_registers_i/dscratch1_q_14_ ),
    .S(net632),
    .X(\cs_registers_i/_0177_ ));
 sg13g2_mux2_1 \cs_registers_i/_4360_  (.A0(net1068),
    .A1(\cs_registers_i/dscratch1_q_15_ ),
    .S(net631),
    .X(\cs_registers_i/_0178_ ));
 sg13g2_mux2_1 \cs_registers_i/_4361_  (.A0(net1055),
    .A1(\cs_registers_i/dscratch1_q_16_ ),
    .S(net632),
    .X(\cs_registers_i/_0179_ ));
 sg13g2_mux2_1 \cs_registers_i/_4362_  (.A0(net1054),
    .A1(\cs_registers_i/dscratch1_q_17_ ),
    .S(net633),
    .X(\cs_registers_i/_0180_ ));
 sg13g2_mux2_1 \cs_registers_i/_4363_  (.A0(net1051),
    .A1(\cs_registers_i/dscratch1_q_18_ ),
    .S(net631),
    .X(\cs_registers_i/_0181_ ));
 sg13g2_buf_8 fanout489 (.A(net520),
    .X(net489));
 sg13g2_mux2_1 \cs_registers_i/_4365_  (.A0(\cs_registers_i/_0903_ ),
    .A1(\cs_registers_i/dscratch1_q_19_ ),
    .S(net633),
    .X(\cs_registers_i/_0182_ ));
 sg13g2_mux2_1 \cs_registers_i/_4366_  (.A0(\cs_registers_i/_0932_ ),
    .A1(\cs_registers_i/dscratch1_q_1_ ),
    .S(net632),
    .X(\cs_registers_i/_0183_ ));
 sg13g2_mux2_1 \cs_registers_i/_4367_  (.A0(\cs_registers_i/_0961_ ),
    .A1(\cs_registers_i/dscratch1_q_20_ ),
    .S(net635),
    .X(\cs_registers_i/_0184_ ));
 sg13g2_mux2_1 \cs_registers_i/_4368_  (.A0(net1048),
    .A1(\cs_registers_i/dscratch1_q_21_ ),
    .S(net633),
    .X(\cs_registers_i/_0185_ ));
 sg13g2_mux2_1 \cs_registers_i/_4369_  (.A0(\cs_registers_i/_1009_ ),
    .A1(\cs_registers_i/dscratch1_q_22_ ),
    .S(net633),
    .X(\cs_registers_i/_0186_ ));
 sg13g2_mux2_1 \cs_registers_i/_4370_  (.A0(net1046),
    .A1(\cs_registers_i/dscratch1_q_23_ ),
    .S(net632),
    .X(\cs_registers_i/_0187_ ));
 sg13g2_mux2_1 \cs_registers_i/_4371_  (.A0(net1045),
    .A1(\cs_registers_i/dscratch1_q_24_ ),
    .S(net633),
    .X(\cs_registers_i/_0188_ ));
 sg13g2_mux2_1 \cs_registers_i/_4372_  (.A0(\cs_registers_i/_1079_ ),
    .A1(\cs_registers_i/dscratch1_q_25_ ),
    .S(net635),
    .X(\cs_registers_i/_0189_ ));
 sg13g2_mux2_1 \cs_registers_i/_4373_  (.A0(\cs_registers_i/_1100_ ),
    .A1(\cs_registers_i/dscratch1_q_26_ ),
    .S(net635),
    .X(\cs_registers_i/_0190_ ));
 sg13g2_mux2_1 \cs_registers_i/_4374_  (.A0(\cs_registers_i/_1128_ ),
    .A1(\cs_registers_i/dscratch1_q_27_ ),
    .S(net633),
    .X(\cs_registers_i/_0191_ ));
 sg13g2_buf_8 fanout488 (.A(net521),
    .X(net488));
 sg13g2_mux2_1 \cs_registers_i/_4376_  (.A0(\cs_registers_i/_1152_ ),
    .A1(\cs_registers_i/dscratch1_q_28_ ),
    .S(net635),
    .X(\cs_registers_i/_0192_ ));
 sg13g2_mux2_1 \cs_registers_i/_4377_  (.A0(net1040),
    .A1(\cs_registers_i/dscratch1_q_29_ ),
    .S(net632),
    .X(\cs_registers_i/_0193_ ));
 sg13g2_mux2_1 \cs_registers_i/_4378_  (.A0(net1038),
    .A1(\cs_registers_i/dscratch1_q_2_ ),
    .S(net634),
    .X(\cs_registers_i/_0194_ ));
 sg13g2_mux2_1 \cs_registers_i/_4379_  (.A0(\cs_registers_i/_1224_ ),
    .A1(\cs_registers_i/dscratch1_q_30_ ),
    .S(net634),
    .X(\cs_registers_i/_0195_ ));
 sg13g2_mux2_1 \cs_registers_i/_4380_  (.A0(net1036),
    .A1(\cs_registers_i/dscratch1_q_31_ ),
    .S(net634),
    .X(\cs_registers_i/_0196_ ));
 sg13g2_mux2_1 \cs_registers_i/_4381_  (.A0(net1034),
    .A1(\cs_registers_i/dscratch1_q_3_ ),
    .S(net635),
    .X(\cs_registers_i/_0197_ ));
 sg13g2_mux2_1 \cs_registers_i/_4382_  (.A0(net1032),
    .A1(\cs_registers_i/dscratch1_q_4_ ),
    .S(net631),
    .X(\cs_registers_i/_0198_ ));
 sg13g2_mux2_1 \cs_registers_i/_4383_  (.A0(\cs_registers_i/_1304_ ),
    .A1(\cs_registers_i/dscratch1_q_5_ ),
    .S(net631),
    .X(\cs_registers_i/_0199_ ));
 sg13g2_mux2_1 \cs_registers_i/_4384_  (.A0(\cs_registers_i/_1322_ ),
    .A1(\cs_registers_i/dscratch1_q_6_ ),
    .S(net635),
    .X(\cs_registers_i/_0200_ ));
 sg13g2_mux2_1 \cs_registers_i/_4385_  (.A0(\cs_registers_i/_1348_ ),
    .A1(\cs_registers_i/dscratch1_q_7_ ),
    .S(net633),
    .X(\cs_registers_i/_0201_ ));
 sg13g2_mux2_1 \cs_registers_i/_4386_  (.A0(\cs_registers_i/_1369_ ),
    .A1(\cs_registers_i/dscratch1_q_8_ ),
    .S(net635),
    .X(\cs_registers_i/_0202_ ));
 sg13g2_mux2_1 \cs_registers_i/_4387_  (.A0(net1030),
    .A1(\cs_registers_i/dscratch1_q_9_ ),
    .S(net631),
    .X(\cs_registers_i/_0203_ ));
 sg13g2_or2_2 \cs_registers_i/_4388_  (.X(\id_stage_i.illegal_csr_insn_i ),
    .B(\cs_registers_i/_0568_ ),
    .A(\cs_registers_i/_0578_ ));
 sg13g2_and2_1 \cs_registers_i/_4389_  (.A(irq_fast_i_7_),
    .B(\cs_registers_i/mie_q_7_ ),
    .X(\id_stage_i.controller_i.irqs_i_7_ ));
 sg13g2_and2_1 \cs_registers_i/_4390_  (.A(irq_software_i),
    .B(\cs_registers_i/mie_q_18_ ),
    .X(\id_stage_i.controller_i.irqs_i_18_ ));
 sg13g2_and2_1 \cs_registers_i/_4391_  (.A(irq_fast_i_9_),
    .B(\cs_registers_i/mie_q_9_ ),
    .X(\id_stage_i.controller_i.irqs_i_9_ ));
 sg13g2_nor3_1 \cs_registers_i/_4392_  (.A(\id_stage_i.controller_i.irqs_i_7_ ),
    .B(\id_stage_i.controller_i.irqs_i_18_ ),
    .C(\id_stage_i.controller_i.irqs_i_9_ ),
    .Y(\cs_registers_i/_1711_ ));
 sg13g2_and2_1 \cs_registers_i/_4393_  (.A(irq_fast_i_3_),
    .B(\cs_registers_i/mie_q_3_ ),
    .X(\id_stage_i.controller_i.irqs_i_3_ ));
 sg13g2_and2_1 \cs_registers_i/_4394_  (.A(irq_timer_i),
    .B(\cs_registers_i/mie_q_17_ ),
    .X(\id_stage_i.controller_i.irqs_i_17_ ));
 sg13g2_nor2_1 \cs_registers_i/_4395_  (.A(\id_stage_i.controller_i.irqs_i_3_ ),
    .B(\id_stage_i.controller_i.irqs_i_17_ ),
    .Y(\cs_registers_i/_1712_ ));
 sg13g2_and2_2 \cs_registers_i/_4396_  (.A(irq_fast_i_4_),
    .B(\cs_registers_i/mie_q_4_ ),
    .X(\id_stage_i.controller_i.irqs_i_4_ ));
 sg13g2_and2_2 \cs_registers_i/_4397_  (.A(irq_fast_i_5_),
    .B(\cs_registers_i/mie_q_5_ ),
    .X(\id_stage_i.controller_i.irqs_i_5_ ));
 sg13g2_nor2_2 \cs_registers_i/_4398_  (.A(\id_stage_i.controller_i.irqs_i_4_ ),
    .B(\id_stage_i.controller_i.irqs_i_5_ ),
    .Y(\cs_registers_i/_1713_ ));
 sg13g2_and2_2 \cs_registers_i/_4399_  (.A(irq_fast_i_6_),
    .B(\cs_registers_i/mie_q_6_ ),
    .X(\id_stage_i.controller_i.irqs_i_6_ ));
 sg13g2_and2_1 \cs_registers_i/_4400_  (.A(irq_fast_i_0_),
    .B(\cs_registers_i/mie_q_0_ ),
    .X(\id_stage_i.controller_i.irqs_i_0_ ));
 sg13g2_nor2_2 \cs_registers_i/_4401_  (.A(\id_stage_i.controller_i.irqs_i_6_ ),
    .B(\id_stage_i.controller_i.irqs_i_0_ ),
    .Y(\cs_registers_i/_1714_ ));
 sg13g2_and2_2 \cs_registers_i/_4402_  (.A(irq_fast_i_8_),
    .B(\cs_registers_i/mie_q_8_ ),
    .X(\id_stage_i.controller_i.irqs_i_8_ ));
 sg13g2_and2_1 \cs_registers_i/_4403_  (.A(irq_fast_i_1_),
    .B(\cs_registers_i/mie_q_1_ ),
    .X(\id_stage_i.controller_i.irqs_i_1_ ));
 sg13g2_nor2_2 \cs_registers_i/_4404_  (.A(\id_stage_i.controller_i.irqs_i_8_ ),
    .B(\id_stage_i.controller_i.irqs_i_1_ ),
    .Y(\cs_registers_i/_1715_ ));
 sg13g2_and4_1 \cs_registers_i/_4405_  (.A(\cs_registers_i/_1712_ ),
    .B(\cs_registers_i/_1713_ ),
    .C(\cs_registers_i/_1714_ ),
    .D(\cs_registers_i/_1715_ ),
    .X(\cs_registers_i/_1716_ ));
 sg13g2_and2_1 \cs_registers_i/_4406_  (.A(irq_fast_i_2_),
    .B(\cs_registers_i/mie_q_2_ ),
    .X(\id_stage_i.controller_i.irqs_i_2_ ));
 sg13g2_and2_1 \cs_registers_i/_4407_  (.A(irq_fast_i_10_),
    .B(\cs_registers_i/mie_q_10_ ),
    .X(\id_stage_i.controller_i.irqs_i_10_ ));
 sg13g2_nor2_1 \cs_registers_i/_4408_  (.A(\id_stage_i.controller_i.irqs_i_2_ ),
    .B(\id_stage_i.controller_i.irqs_i_10_ ),
    .Y(\cs_registers_i/_1717_ ));
 sg13g2_and2_1 \cs_registers_i/_4409_  (.A(irq_fast_i_15_),
    .B(\cs_registers_i/mie_q_15_ ),
    .X(\id_stage_i.controller_i.irqs_i_15_ ));
 sg13g2_and2_1 \cs_registers_i/_4410_  (.A(irq_external_i),
    .B(\cs_registers_i/mie_q_16_ ),
    .X(\id_stage_i.controller_i.irqs_i_16_ ));
 sg13g2_nor2_1 \cs_registers_i/_4411_  (.A(\id_stage_i.controller_i.irqs_i_15_ ),
    .B(\id_stage_i.controller_i.irqs_i_16_ ),
    .Y(\cs_registers_i/_1718_ ));
 sg13g2_and2_1 \cs_registers_i/_4412_  (.A(irq_fast_i_11_),
    .B(\cs_registers_i/mie_q_11_ ),
    .X(\id_stage_i.controller_i.irqs_i_11_ ));
 sg13g2_and2_1 \cs_registers_i/_4413_  (.A(irq_fast_i_12_),
    .B(\cs_registers_i/mie_q_12_ ),
    .X(\id_stage_i.controller_i.irqs_i_12_ ));
 sg13g2_nor2_1 \cs_registers_i/_4414_  (.A(\id_stage_i.controller_i.irqs_i_11_ ),
    .B(\id_stage_i.controller_i.irqs_i_12_ ),
    .Y(\cs_registers_i/_1719_ ));
 sg13g2_and2_1 \cs_registers_i/_4415_  (.A(irq_fast_i_13_),
    .B(\cs_registers_i/mie_q_13_ ),
    .X(\id_stage_i.controller_i.irqs_i_13_ ));
 sg13g2_and2_1 \cs_registers_i/_4416_  (.A(irq_fast_i_14_),
    .B(\cs_registers_i/mie_q_14_ ),
    .X(\id_stage_i.controller_i.irqs_i_14_ ));
 sg13g2_nor2_1 \cs_registers_i/_4417_  (.A(\id_stage_i.controller_i.irqs_i_13_ ),
    .B(\id_stage_i.controller_i.irqs_i_14_ ),
    .Y(\cs_registers_i/_1720_ ));
 sg13g2_and4_1 \cs_registers_i/_4418_  (.A(\cs_registers_i/_1717_ ),
    .B(\cs_registers_i/_1718_ ),
    .C(\cs_registers_i/_1719_ ),
    .D(\cs_registers_i/_1720_ ),
    .X(\cs_registers_i/_1721_ ));
 sg13g2_nand3_1 \cs_registers_i/_4419_  (.B(\cs_registers_i/_1716_ ),
    .C(\cs_registers_i/_1721_ ),
    .A(\cs_registers_i/_1711_ ),
    .Y(irq_pending_o));
 sg13g2_nor2_1 \cs_registers_i/_4420_  (.A(net197),
    .B(\cs_registers_i/_1688_ ),
    .Y(\cs_registers_i/_1722_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4421_  (.Y(\cs_registers_i/_1723_ ),
    .B1(net290),
    .B2(\cs_registers_i/mstack_cause_q_0_ ),
    .A2(net1294),
    .A1(exc_cause_0_));
 sg13g2_inv_1 \cs_registers_i/_4422_  (.Y(\cs_registers_i/_1724_ ),
    .A(\cs_registers_i/_1723_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4423_  (.B2(\cs_registers_i/_1722_ ),
    .C1(\cs_registers_i/_1724_ ),
    .B1(net1079),
    .A1(net198),
    .Y(\cs_registers_i/_1725_ ),
    .A2(net1206));
 sg13g2_inv_1 \cs_registers_i/_4424_  (.Y(\cs_registers_i/_1726_ ),
    .A(\cs_registers_i/_1061_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4425_  (.B1(\cs_registers_i/_1411_ ),
    .Y(\cs_registers_i/_1727_ ),
    .A1(\cs_registers_i/_1726_ ),
    .A2(\cs_registers_i/_1410_ ));
 sg13g2_buf_8 fanout487 (.A(net521),
    .X(net487));
 sg13g2_nor2_2 \cs_registers_i/_4427_  (.A(\cs_registers_i/mcause_q_0_ ),
    .B(net586),
    .Y(\cs_registers_i/_1729_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4428_  (.A1(\cs_registers_i/_1725_ ),
    .A2(net586),
    .Y(\cs_registers_i/_0204_ ),
    .B1(\cs_registers_i/_1729_ ));
 sg13g2_nor2_1 \cs_registers_i/_4429_  (.A(alu_operand_a_ex_1_),
    .B(\cs_registers_i/_0930_ ),
    .Y(\cs_registers_i/_1730_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4430_  (.Y(\cs_registers_i/_1731_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_cause_q_1_ ),
    .A2(net1295),
    .A1(exc_cause_1_));
 sg13g2_inv_1 \cs_registers_i/_4431_  (.Y(\cs_registers_i/_1732_ ),
    .A(\cs_registers_i/_1731_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4432_  (.B2(\cs_registers_i/_1730_ ),
    .C1(\cs_registers_i/_1732_ ),
    .B1(net1079),
    .A1(alu_operand_a_ex_1_),
    .Y(\cs_registers_i/_1733_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4433_  (.A(\cs_registers_i/mcause_q_1_ ),
    .B(net587),
    .Y(\cs_registers_i/_1734_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4434_  (.A1(net587),
    .A2(\cs_registers_i/_1733_ ),
    .Y(\cs_registers_i/_0205_ ),
    .B1(\cs_registers_i/_1734_ ));
 sg13g2_nor2_1 \cs_registers_i/_4435_  (.A(net1410),
    .B(\cs_registers_i/_1201_ ),
    .Y(\cs_registers_i/_1735_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4436_  (.Y(\cs_registers_i/_1736_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_cause_q_2_ ),
    .A2(net1294),
    .A1(exc_cause_2_));
 sg13g2_inv_1 \cs_registers_i/_4437_  (.Y(\cs_registers_i/_1737_ ),
    .A(\cs_registers_i/_1736_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4438_  (.B2(\cs_registers_i/_1735_ ),
    .C1(\cs_registers_i/_1737_ ),
    .B1(net1079),
    .A1(net1410),
    .Y(\cs_registers_i/_1738_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4439_  (.A(\cs_registers_i/mcause_q_2_ ),
    .B(net587),
    .Y(\cs_registers_i/_1739_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4440_  (.A1(net587),
    .A2(\cs_registers_i/_1738_ ),
    .Y(\cs_registers_i/_0206_ ),
    .B1(\cs_registers_i/_1739_ ));
 sg13g2_nor2_1 \cs_registers_i/_4441_  (.A(alu_operand_a_ex_3_),
    .B(\cs_registers_i/_1270_ ),
    .Y(\cs_registers_i/_1740_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4442_  (.Y(\cs_registers_i/_1741_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_cause_q_3_ ),
    .A2(net1294),
    .A1(exc_cause_3_));
 sg13g2_inv_1 \cs_registers_i/_4443_  (.Y(\cs_registers_i/_1742_ ),
    .A(\cs_registers_i/_1741_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4444_  (.B2(\cs_registers_i/_1740_ ),
    .C1(\cs_registers_i/_1742_ ),
    .B1(net1079),
    .A1(alu_operand_a_ex_3_),
    .Y(\cs_registers_i/_1743_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4445_  (.A(\cs_registers_i/mcause_q_3_ ),
    .B(net586),
    .Y(\cs_registers_i/_1744_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4446_  (.A1(net586),
    .A2(\cs_registers_i/_1743_ ),
    .Y(\cs_registers_i/_0207_ ),
    .B1(\cs_registers_i/_1744_ ));
 sg13g2_nor2_1 \cs_registers_i/_4447_  (.A(net1406),
    .B(\cs_registers_i/_1284_ ),
    .Y(\cs_registers_i/_1745_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4448_  (.Y(\cs_registers_i/_1746_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_cause_q_4_ ),
    .A2(net1295),
    .A1(exc_cause_4_));
 sg13g2_inv_1 \cs_registers_i/_4449_  (.Y(\cs_registers_i/_1747_ ),
    .A(\cs_registers_i/_1746_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4450_  (.B2(\cs_registers_i/_1745_ ),
    .C1(\cs_registers_i/_1747_ ),
    .B1(net1079),
    .A1(net1406),
    .Y(\cs_registers_i/_1748_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4451_  (.A(\cs_registers_i/mcause_q_4_ ),
    .B(net586),
    .Y(\cs_registers_i/_1749_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4452_  (.A1(net586),
    .A2(\cs_registers_i/_1748_ ),
    .Y(\cs_registers_i/_0208_ ),
    .B1(\cs_registers_i/_1749_ ));
 sg13g2_nor2_1 \cs_registers_i/_4453_  (.A(net1405),
    .B(\cs_registers_i/_1302_ ),
    .Y(\cs_registers_i/_1750_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4454_  (.Y(\cs_registers_i/_1751_ ),
    .B1(net293),
    .B2(\cs_registers_i/mstack_cause_q_5_ ),
    .A2(net1295),
    .A1(exc_cause_5_));
 sg13g2_inv_1 \cs_registers_i/_4455_  (.Y(\cs_registers_i/_1752_ ),
    .A(\cs_registers_i/_1751_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4456_  (.B2(\cs_registers_i/_1750_ ),
    .C1(\cs_registers_i/_1752_ ),
    .B1(net1079),
    .A1(net1405),
    .Y(\cs_registers_i/_1753_ ),
    .A2(net1206));
 sg13g2_nor2_2 \cs_registers_i/_4457_  (.A(\cs_registers_i/mcause_q_5_ ),
    .B(net586),
    .Y(\cs_registers_i/_1754_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4458_  (.B1(\cs_registers_i/_1754_ ),
    .Y(\cs_registers_i/_0209_ ),
    .A2(\cs_registers_i/_1753_ ),
    .A1(net586));
 sg13g2_and2_1 \cs_registers_i/_4459_  (.A(\cs_registers_i/mstack_cause_q_6_ ),
    .B(net291),
    .X(\cs_registers_i/_1755_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4460_  (.B2(net1035),
    .C1(\cs_registers_i/_1755_ ),
    .B1(net153),
    .A1(exc_cause_6_),
    .Y(\cs_registers_i/_1756_ ),
    .A2(net1296));
 sg13g2_nor2_2 \cs_registers_i/_4461_  (.A(\cs_registers_i/mcause_q_6_ ),
    .B(net587),
    .Y(\cs_registers_i/_1757_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4462_  (.B1(\cs_registers_i/_1757_ ),
    .Y(\cs_registers_i/_0210_ ),
    .A2(\cs_registers_i/_1756_ ),
    .A1(net587));
 sg13g2_nand2_2 \cs_registers_i/_4463_  (.Y(\cs_registers_i/_1758_ ),
    .A(\cs_registers_i/_0580_ ),
    .B(\cs_registers_i/_0649_ ));
 sg13g2_mux2_1 \cs_registers_i/_4464_  (.A0(net1063),
    .A1(\cs_registers_i/mcountinhibit_0_ ),
    .S(\cs_registers_i/_1758_ ),
    .X(\cs_registers_i/_0211_ ));
 sg13g2_mux2_1 \cs_registers_i/_4465_  (.A0(net1038),
    .A1(\cs_registers_i/mcountinhibit_2_ ),
    .S(\cs_registers_i/_1758_ ),
    .X(\cs_registers_i/_0212_ ));
 sg13g2_nor2_1 \cs_registers_i/_4466_  (.A(\cs_registers_i/_0500_ ),
    .B(\cs_registers_i/_0527_ ),
    .Y(\cs_registers_i/_1759_ ));
 sg13g2_nand4_1 \cs_registers_i/_4467_  (.B(net1117),
    .C(\cs_registers_i/_1759_ ),
    .A(\cs_registers_i/_0552_ ),
    .Y(\cs_registers_i/_1760_ ),
    .D(net1156));
 sg13g2_nor3_2 \cs_registers_i/_4468_  (.A(\cs_registers_i/_0571_ ),
    .B(\cs_registers_i/_0578_ ),
    .C(\cs_registers_i/_1760_ ),
    .Y(\cs_registers_i/_1761_ ));
 sg13g2_buf_8 fanout486 (.A(net521),
    .X(net486));
 sg13g2_nand2b_2 \cs_registers_i/_4470_  (.Y(\cs_registers_i/_1763_ ),
    .B(net31),
    .A_N(\cs_registers_i/_0568_ ));
 sg13g2_buf_8 fanout485 (.A(net521),
    .X(net485));
 sg13g2_buf_8 fanout484 (.A(net521),
    .X(net484));
 sg13g2_nor2_1 \cs_registers_i/_4473_  (.A(net1245),
    .B(\cs_registers_i/_0601_ ),
    .Y(\cs_registers_i/_1766_ ));
 sg13g2_nand2_1 \cs_registers_i/_4474_  (.Y(\cs_registers_i/_1767_ ),
    .A(\cs_registers_i/_0525_ ),
    .B(\cs_registers_i/_1766_ ));
 sg13g2_nor2_1 \cs_registers_i/_4475_  (.A(\cs_registers_i/_1767_ ),
    .B(\cs_registers_i/_0876_ ),
    .Y(\cs_registers_i/_1768_ ));
 sg13g2_and2_2 \cs_registers_i/_4476_  (.A(\cs_registers_i/_0579_ ),
    .B(\cs_registers_i/_1768_ ),
    .X(\cs_registers_i/_1769_ ));
 sg13g2_buf_8 fanout483 (.A(net521),
    .X(net483));
 sg13g2_or4_2 \cs_registers_i/_4478_  (.A(\cs_registers_i/_0571_ ),
    .B(\cs_registers_i/_0578_ ),
    .C(\cs_registers_i/_1767_ ),
    .D(\cs_registers_i/_0876_ ),
    .X(\cs_registers_i/_1771_ ));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(net521));
 sg13g2_and3_1 \cs_registers_i/_4480_  (.X(\cs_registers_i/_1773_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_upd_0_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .C(net28));
 sg13g2_a21o_1 \cs_registers_i/_4481_  (.A2(net18),
    .A1(net1063),
    .B1(\cs_registers_i/_1773_ ),
    .X(\cs_registers_i/_1774_ ));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net521));
 sg13g2_o21ai_1 \cs_registers_i/_4483_  (.B1(net682),
    .Y(\cs_registers_i/_1776_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .A2(net17));
 sg13g2_a22oi_1 \cs_registers_i/_4484_  (.Y(\cs_registers_i/_1777_ ),
    .B1(\cs_registers_i/_1776_ ),
    .B2(\cs_registers_i/mcycle_counter_i.counter_val_o_0_ ),
    .A2(\cs_registers_i/_1774_ ),
    .A1(net682));
 sg13g2_inv_1 \cs_registers_i/_4485_  (.Y(\cs_registers_i/_0213_ ),
    .A(\cs_registers_i/_1777_ ));
 sg13g2_nor2b_2 \cs_registers_i/_4486_  (.A(\cs_registers_i/_0568_ ),
    .B_N(net30),
    .Y(\cs_registers_i/_1778_ ));
 sg13g2_buf_8 fanout480 (.A(net522),
    .X(net480));
 sg13g2_and4_1 \cs_registers_i/_4488_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_0_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_2_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .D(\cs_registers_i/mcycle_counter_i.counter_val_o_1_ ),
    .X(\cs_registers_i/_1780_ ));
 sg13g2_and4_1 \cs_registers_i/_4489_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_6_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_3_ ),
    .D(\cs_registers_i/mcycle_counter_i.counter_val_o_5_ ),
    .X(\cs_registers_i/_1781_ ));
 sg13g2_and2_2 \cs_registers_i/_4490_  (.A(\cs_registers_i/_1780_ ),
    .B(\cs_registers_i/_1781_ ),
    .X(\cs_registers_i/_1782_ ));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net522));
 sg13g2_and2_1 \cs_registers_i/_4492_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_7_ ),
    .B(\cs_registers_i/_1782_ ),
    .X(\cs_registers_i/_1784_ ));
 sg13g2_and2_1 \cs_registers_i/_4493_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_8_ ),
    .B(\cs_registers_i/_1784_ ),
    .X(\cs_registers_i/_1785_ ));
 sg13g2_and2_1 \cs_registers_i/_4494_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ),
    .B(\cs_registers_i/_1785_ ),
    .X(\cs_registers_i/_1786_ ));
 sg13g2_inv_1 \cs_registers_i/_4495_  (.Y(\cs_registers_i/_1787_ ),
    .A(\cs_registers_i/_1786_ ));
 sg13g2_nor3_1 \cs_registers_i/_4496_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .B(net18),
    .C(\cs_registers_i/_1787_ ),
    .Y(\cs_registers_i/_1788_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4497_  (.A1(net1059),
    .A2(net18),
    .Y(\cs_registers_i/_1789_ ),
    .B1(\cs_registers_i/_1788_ ));
 sg13g2_nor2_1 \cs_registers_i/_4498_  (.A(net17),
    .B(\cs_registers_i/_1786_ ),
    .Y(\cs_registers_i/_1790_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4499_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .Y(\cs_registers_i/_1791_ ),
    .A1(\cs_registers_i/_1778_ ),
    .A2(\cs_registers_i/_1790_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4500_  (.B1(\cs_registers_i/_1791_ ),
    .Y(\cs_registers_i/_0214_ ),
    .A1(\cs_registers_i/_1778_ ),
    .A2(\cs_registers_i/_1789_ ));
 sg13g2_buf_8 fanout478 (.A(net522),
    .X(net478));
 sg13g2_buf_8 fanout477 (.A(net522),
    .X(net477));
 sg13g2_nand3_1 \cs_registers_i/_4503_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_11_ ),
    .C(\cs_registers_i/_1786_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .Y(\cs_registers_i/_1794_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4504_  (.Y(\cs_registers_i/_1795_ ),
    .B(net25),
    .A_N(\cs_registers_i/_1794_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4505_  (.B1(\cs_registers_i/_1795_ ),
    .Y(\cs_registers_i/_1796_ ),
    .A1(net1070),
    .A2(net26));
 sg13g2_a21o_1 \cs_registers_i/_4506_  (.A2(\cs_registers_i/_1786_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .B1(\cs_registers_i/_1769_ ),
    .X(\cs_registers_i/_1797_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4507_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_11_ ),
    .Y(\cs_registers_i/_1798_ ),
    .A2(\cs_registers_i/_1797_ ),
    .A1(net681));
 sg13g2_a21oi_1 \cs_registers_i/_4508_  (.A1(net681),
    .A2(\cs_registers_i/_1796_ ),
    .Y(\cs_registers_i/_0215_ ),
    .B1(\cs_registers_i/_1798_ ));
 sg13g2_or2_1 \cs_registers_i/_4509_  (.X(\cs_registers_i/_1799_ ),
    .B(\cs_registers_i/_1795_ ),
    .A(\cs_registers_i/_0723_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4510_  (.B1(\cs_registers_i/_1799_ ),
    .Y(\cs_registers_i/_1800_ ),
    .A1(net1028),
    .A2(net26));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net522));
 sg13g2_a21o_1 \cs_registers_i/_4512_  (.A2(\cs_registers_i/_1794_ ),
    .A1(net29),
    .B1(\cs_registers_i/_1778_ ),
    .X(\cs_registers_i/_1802_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4513_  (.Y(\cs_registers_i/_0216_ ),
    .B1(\cs_registers_i/_1802_ ),
    .B2(\cs_registers_i/_0723_ ),
    .A2(\cs_registers_i/_1800_ ),
    .A1(net681));
 sg13g2_nand2_1 \cs_registers_i/_4514_  (.Y(\cs_registers_i/_1803_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_7_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ));
 sg13g2_nand4_1 \cs_registers_i/_4515_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_8_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_12_ ),
    .Y(\cs_registers_i/_1804_ ),
    .D(\cs_registers_i/mcycle_counter_i.counter_val_o_11_ ));
 sg13g2_nor2_1 \cs_registers_i/_4516_  (.A(\cs_registers_i/_1803_ ),
    .B(\cs_registers_i/_1804_ ),
    .Y(\cs_registers_i/_1805_ ));
 sg13g2_and3_1 \cs_registers_i/_4517_  (.X(\cs_registers_i/_1806_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_13_ ),
    .B(\cs_registers_i/_1782_ ),
    .C(\cs_registers_i/_1805_ ));
 sg13g2_nand2_1 \cs_registers_i/_4518_  (.Y(\cs_registers_i/_1807_ ),
    .A(net29),
    .B(\cs_registers_i/_1806_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4519_  (.B1(\cs_registers_i/_1807_ ),
    .Y(\cs_registers_i/_1808_ ),
    .A1(net1057),
    .A2(net26));
 sg13g2_a21o_1 \cs_registers_i/_4520_  (.A2(\cs_registers_i/_1805_ ),
    .A1(\cs_registers_i/_1782_ ),
    .B1(\cs_registers_i/_1769_ ),
    .X(\cs_registers_i/_1809_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4521_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_13_ ),
    .Y(\cs_registers_i/_1810_ ),
    .A2(\cs_registers_i/_1809_ ),
    .A1(net681));
 sg13g2_a21oi_1 \cs_registers_i/_4522_  (.A1(net681),
    .A2(\cs_registers_i/_1808_ ),
    .Y(\cs_registers_i/_0217_ ),
    .B1(\cs_registers_i/_1810_ ));
 sg13g2_buf_8 fanout475 (.A(net522),
    .X(net475));
 sg13g2_nand3_1 \cs_registers_i/_4524_  (.B(net28),
    .C(\cs_registers_i/_1806_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ),
    .Y(\cs_registers_i/_1812_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4525_  (.B1(\cs_registers_i/_1812_ ),
    .Y(\cs_registers_i/_1813_ ),
    .A1(\cs_registers_i/_0790_ ),
    .A2(net26));
 sg13g2_o21ai_1 \cs_registers_i/_4526_  (.B1(net681),
    .Y(\cs_registers_i/_1814_ ),
    .A1(net17),
    .A2(\cs_registers_i/_1806_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4527_  (.Y(\cs_registers_i/_0218_ ),
    .B1(\cs_registers_i/_1814_ ),
    .B2(\cs_registers_i/_0783_ ),
    .A2(\cs_registers_i/_1813_ ),
    .A1(net682));
 sg13g2_nand4_1 \cs_registers_i/_4528_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_15_ ),
    .C(net28),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ),
    .Y(\cs_registers_i/_1815_ ),
    .D(\cs_registers_i/_1806_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4529_  (.B1(\cs_registers_i/_1815_ ),
    .Y(\cs_registers_i/_1816_ ),
    .A1(net1069),
    .A2(net26));
 sg13g2_a21o_1 \cs_registers_i/_4530_  (.A2(\cs_registers_i/_1806_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ),
    .B1(\cs_registers_i/_1769_ ),
    .X(\cs_registers_i/_1817_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4531_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_15_ ),
    .Y(\cs_registers_i/_1818_ ),
    .A2(\cs_registers_i/_1817_ ),
    .A1(net681));
 sg13g2_a21oi_1 \cs_registers_i/_4532_  (.A1(net682),
    .A2(\cs_registers_i/_1816_ ),
    .Y(\cs_registers_i/_0219_ ),
    .B1(\cs_registers_i/_1818_ ));
 sg13g2_nand3_1 \cs_registers_i/_4533_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_13_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_15_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ),
    .Y(\cs_registers_i/_1819_ ));
 sg13g2_nor3_2 \cs_registers_i/_4534_  (.A(\cs_registers_i/_1803_ ),
    .B(\cs_registers_i/_1804_ ),
    .C(\cs_registers_i/_1819_ ),
    .Y(\cs_registers_i/_1820_ ));
 sg13g2_nand2_1 \cs_registers_i/_4535_  (.Y(\cs_registers_i/_1821_ ),
    .A(\cs_registers_i/_1782_ ),
    .B(\cs_registers_i/_1820_ ));
 sg13g2_nor2_1 \cs_registers_i/_4536_  (.A(net30),
    .B(\cs_registers_i/_1821_ ),
    .Y(\cs_registers_i/_1822_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4537_  (.Y(\cs_registers_i/_1823_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .B(\cs_registers_i/_1822_ ));
 sg13g2_nand3_1 \cs_registers_i/_4538_  (.B(\cs_registers_i/_1759_ ),
    .C(net1156),
    .A(\cs_registers_i/_0526_ ),
    .Y(\cs_registers_i/_1824_ ));
 sg13g2_nand2_2 \cs_registers_i/_4539_  (.Y(\cs_registers_i/_1825_ ),
    .A(net17),
    .B(net38));
 sg13g2_buf_8 fanout474 (.A(net522),
    .X(net474));
 sg13g2_nor2_2 \cs_registers_i/_4541_  (.A(\cs_registers_i/_0834_ ),
    .B(net628),
    .Y(\cs_registers_i/_1827_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4542_  (.A1(\cs_registers_i/_1823_ ),
    .A2(net628),
    .Y(\cs_registers_i/_0220_ ),
    .B1(\cs_registers_i/_1827_ ));
 sg13g2_nand2_1 \cs_registers_i/_4543_  (.Y(\cs_registers_i/_1828_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .B(\cs_registers_i/_1822_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4544_  (.Y(\cs_registers_i/_1829_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_17_ ),
    .B(\cs_registers_i/_1828_ ));
 sg13g2_mux2_1 \cs_registers_i/_4545_  (.A0(net1054),
    .A1(\cs_registers_i/_1829_ ),
    .S(net628),
    .X(\cs_registers_i/_0221_ ));
 sg13g2_nand3_1 \cs_registers_i/_4546_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_17_ ),
    .C(\cs_registers_i/_1822_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .Y(\cs_registers_i/_1830_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4547_  (.Y(\cs_registers_i/_1831_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_18_ ),
    .B(\cs_registers_i/_1830_ ));
 sg13g2_mux2_1 \cs_registers_i/_4548_  (.A0(net1052),
    .A1(\cs_registers_i/_1831_ ),
    .S(net627),
    .X(\cs_registers_i/_0222_ ));
 sg13g2_buf_8 fanout473 (.A(net522),
    .X(net473));
 sg13g2_or2_1 \cs_registers_i/_4550_  (.X(\cs_registers_i/_1833_ ),
    .B(\cs_registers_i/_1821_ ),
    .A(net30));
 sg13g2_nand3_1 \cs_registers_i/_4551_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_17_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_18_ ),
    .Y(\cs_registers_i/_1834_ ));
 sg13g2_nor2_2 \cs_registers_i/_4552_  (.A(\cs_registers_i/_1833_ ),
    .B(\cs_registers_i/_1834_ ),
    .Y(\cs_registers_i/_1835_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4553_  (.Y(\cs_registers_i/_1836_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .B(\cs_registers_i/_1835_ ));
 sg13g2_nor2_2 \cs_registers_i/_4554_  (.A(\cs_registers_i/_0903_ ),
    .B(net628),
    .Y(\cs_registers_i/_1837_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4555_  (.A1(net628),
    .A2(\cs_registers_i/_1836_ ),
    .Y(\cs_registers_i/_0223_ ),
    .B1(\cs_registers_i/_1837_ ));
 sg13g2_and2_1 \cs_registers_i/_4556_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_0_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .X(\cs_registers_i/_1838_ ));
 sg13g2_and2_1 \cs_registers_i/_4557_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_1_ ),
    .B(\cs_registers_i/_1838_ ),
    .X(\cs_registers_i/_1839_ ));
 sg13g2_nand2_1 \cs_registers_i/_4558_  (.Y(\cs_registers_i/_1840_ ),
    .A(\cs_registers_i/_1771_ ),
    .B(\cs_registers_i/_1839_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4559_  (.B1(\cs_registers_i/_1840_ ),
    .Y(\cs_registers_i/_1841_ ),
    .A1(\cs_registers_i/_0932_ ),
    .A2(net27));
 sg13g2_o21ai_1 \cs_registers_i/_4560_  (.B1(net679),
    .Y(\cs_registers_i/_1842_ ),
    .A1(net17),
    .A2(\cs_registers_i/_1838_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4561_  (.Y(\cs_registers_i/_0224_ ),
    .B1(\cs_registers_i/_1842_ ),
    .B2(\cs_registers_i/_0915_ ),
    .A2(\cs_registers_i/_1841_ ),
    .A1(net680));
 sg13g2_nand2_2 \cs_registers_i/_4562_  (.Y(\cs_registers_i/_1843_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .B(\cs_registers_i/_1835_ ));
 sg13g2_xor2_1 \cs_registers_i/_4563_  (.B(\cs_registers_i/_1843_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_20_ ),
    .X(\cs_registers_i/_1844_ ));
 sg13g2_nor2_2 \cs_registers_i/_4564_  (.A(\cs_registers_i/_0961_ ),
    .B(net626),
    .Y(\cs_registers_i/_1845_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4565_  (.A1(net630),
    .A2(\cs_registers_i/_1844_ ),
    .Y(\cs_registers_i/_0225_ ),
    .B1(\cs_registers_i/_1845_ ));
 sg13g2_nand3_1 \cs_registers_i/_4566_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .C(\cs_registers_i/_1835_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_20_ ),
    .Y(\cs_registers_i/_1846_ ));
 sg13g2_xor2_1 \cs_registers_i/_4567_  (.B(\cs_registers_i/_1846_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_21_ ),
    .X(\cs_registers_i/_1847_ ));
 sg13g2_nor2_1 \cs_registers_i/_4568_  (.A(net1048),
    .B(net626),
    .Y(\cs_registers_i/_1848_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4569_  (.A1(net630),
    .A2(\cs_registers_i/_1847_ ),
    .Y(\cs_registers_i/_0226_ ),
    .B1(\cs_registers_i/_1848_ ));
 sg13g2_nand3_1 \cs_registers_i/_4570_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_21_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_20_ ),
    .Y(\cs_registers_i/_1849_ ));
 sg13g2_nor3_2 \cs_registers_i/_4571_  (.A(\cs_registers_i/_1833_ ),
    .B(\cs_registers_i/_1834_ ),
    .C(\cs_registers_i/_1849_ ),
    .Y(\cs_registers_i/_1850_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4572_  (.Y(\cs_registers_i/_1851_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_22_ ),
    .B(\cs_registers_i/_1850_ ));
 sg13g2_nor2_2 \cs_registers_i/_4573_  (.A(\cs_registers_i/_1009_ ),
    .B(net626),
    .Y(\cs_registers_i/_1852_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4574_  (.A1(net626),
    .A2(\cs_registers_i/_1851_ ),
    .Y(\cs_registers_i/_0227_ ),
    .B1(\cs_registers_i/_1852_ ));
 sg13g2_nor3_1 \cs_registers_i/_4575_  (.A(\cs_registers_i/_0991_ ),
    .B(\cs_registers_i/_1834_ ),
    .C(\cs_registers_i/_1849_ ),
    .Y(\cs_registers_i/_1853_ ));
 sg13g2_nand4_1 \cs_registers_i/_4576_  (.B(\cs_registers_i/_1782_ ),
    .C(\cs_registers_i/_1820_ ),
    .A(net681),
    .Y(\cs_registers_i/_1854_ ),
    .D(\cs_registers_i/_1853_ ));
 sg13g2_xor2_1 \cs_registers_i/_4577_  (.B(\cs_registers_i/_1854_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_23_ ),
    .X(\cs_registers_i/_1855_ ));
 sg13g2_nor2_1 \cs_registers_i/_4578_  (.A(net1046),
    .B(net626),
    .Y(\cs_registers_i/_1856_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4579_  (.A1(net626),
    .A2(\cs_registers_i/_1855_ ),
    .Y(\cs_registers_i/_0228_ ),
    .B1(\cs_registers_i/_1856_ ));
 sg13g2_nand4_1 \cs_registers_i/_4580_  (.B(\cs_registers_i/_1782_ ),
    .C(\cs_registers_i/_1820_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_23_ ),
    .Y(\cs_registers_i/_1857_ ),
    .D(\cs_registers_i/_1853_ ));
 sg13g2_or2_2 \cs_registers_i/_4581_  (.X(\cs_registers_i/_1858_ ),
    .B(\cs_registers_i/_1857_ ),
    .A(net30));
 sg13g2_xor2_1 \cs_registers_i/_4582_  (.B(\cs_registers_i/_1858_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .X(\cs_registers_i/_1859_ ));
 sg13g2_nor2_2 \cs_registers_i/_4583_  (.A(net1045),
    .B(net627),
    .Y(\cs_registers_i/_1860_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4584_  (.A1(net629),
    .A2(\cs_registers_i/_1859_ ),
    .Y(\cs_registers_i/_0229_ ),
    .B1(\cs_registers_i/_1860_ ));
 sg13g2_inv_2 \cs_registers_i/_4585_  (.Y(\cs_registers_i/_1861_ ),
    .A(\cs_registers_i/_1858_ ));
 sg13g2_nand2_1 \cs_registers_i/_4586_  (.Y(\cs_registers_i/_1862_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .B(\cs_registers_i/_1861_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4587_  (.Y(\cs_registers_i/_1863_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_25_ ),
    .B(\cs_registers_i/_1862_ ));
 sg13g2_mux2_1 \cs_registers_i/_4588_  (.A0(\cs_registers_i/_1079_ ),
    .A1(\cs_registers_i/_1863_ ),
    .S(net627),
    .X(\cs_registers_i/_0230_ ));
 sg13g2_nand3_1 \cs_registers_i/_4589_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_25_ ),
    .C(\cs_registers_i/_1861_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .Y(\cs_registers_i/_1864_ ));
 sg13g2_xor2_1 \cs_registers_i/_4590_  (.B(\cs_registers_i/_1864_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_26_ ),
    .X(\cs_registers_i/_1865_ ));
 sg13g2_nor2_2 \cs_registers_i/_4591_  (.A(\cs_registers_i/_1100_ ),
    .B(net627),
    .Y(\cs_registers_i/_1866_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4592_  (.B1(\cs_registers_i/_1866_ ),
    .Y(\cs_registers_i/_0231_ ),
    .A2(\cs_registers_i/_1865_ ),
    .A1(net627));
 sg13g2_nand3_1 \cs_registers_i/_4593_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_25_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_26_ ),
    .Y(\cs_registers_i/_1867_ ));
 sg13g2_nor2_1 \cs_registers_i/_4594_  (.A(\cs_registers_i/_1858_ ),
    .B(\cs_registers_i/_1867_ ),
    .Y(\cs_registers_i/_1868_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4595_  (.Y(\cs_registers_i/_1869_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_27_ ),
    .B(\cs_registers_i/_1868_ ));
 sg13g2_nor2_2 \cs_registers_i/_4596_  (.A(\cs_registers_i/_1128_ ),
    .B(net628),
    .Y(\cs_registers_i/_1870_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4597_  (.A1(net629),
    .A2(\cs_registers_i/_1869_ ),
    .Y(\cs_registers_i/_0232_ ),
    .B1(\cs_registers_i/_1870_ ));
 sg13g2_nor2_1 \cs_registers_i/_4598_  (.A(\cs_registers_i/_1108_ ),
    .B(\cs_registers_i/_1867_ ),
    .Y(\cs_registers_i/_1871_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4599_  (.Y(\cs_registers_i/_1872_ ),
    .B(\cs_registers_i/_1871_ ),
    .A_N(\cs_registers_i/_1857_ ));
 sg13g2_and2_1 \cs_registers_i/_4600_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .B(\cs_registers_i/_1872_ ),
    .X(\cs_registers_i/_1873_ ));
 sg13g2_nor3_1 \cs_registers_i/_4601_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .B(net31),
    .C(\cs_registers_i/_1872_ ),
    .Y(\cs_registers_i/_1874_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4602_  (.B1(net26),
    .Y(\cs_registers_i/_1875_ ),
    .A1(\cs_registers_i/_1873_ ),
    .A2(\cs_registers_i/_1874_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4603_  (.A(net28),
    .B_N(net38),
    .Y(\cs_registers_i/_1876_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4604_  (.Y(\cs_registers_i/_1877_ ),
    .B1(\cs_registers_i/_1876_ ),
    .B2(\cs_registers_i/_1152_ ),
    .A2(\cs_registers_i/_1778_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ));
 sg13g2_nand2_1 \cs_registers_i/_4605_  (.Y(\cs_registers_i/_0233_ ),
    .A(\cs_registers_i/_1875_ ),
    .B(\cs_registers_i/_1877_ ));
 sg13g2_nand2_1 \cs_registers_i/_4606_  (.Y(\cs_registers_i/_1878_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .B(\cs_registers_i/_1871_ ));
 sg13g2_nor2_2 \cs_registers_i/_4607_  (.A(\cs_registers_i/_1858_ ),
    .B(\cs_registers_i/_1878_ ),
    .Y(\cs_registers_i/_1879_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4608_  (.Y(\cs_registers_i/_1880_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_29_ ),
    .B(\cs_registers_i/_1879_ ));
 sg13g2_nor2_2 \cs_registers_i/_4609_  (.A(net1041),
    .B(net627),
    .Y(\cs_registers_i/_1881_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4610_  (.A1(net627),
    .A2(\cs_registers_i/_1880_ ),
    .Y(\cs_registers_i/_0234_ ),
    .B1(\cs_registers_i/_1881_ ));
 sg13g2_nand2_1 \cs_registers_i/_4611_  (.Y(\cs_registers_i/_1882_ ),
    .A(net29),
    .B(\cs_registers_i/_1780_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4612_  (.B1(\cs_registers_i/_1882_ ),
    .Y(\cs_registers_i/_1883_ ),
    .A1(net1038),
    .A2(net27));
 sg13g2_o21ai_1 \cs_registers_i/_4613_  (.B1(net679),
    .Y(\cs_registers_i/_1884_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1839_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4614_  (.Y(\cs_registers_i/_0235_ ),
    .B1(\cs_registers_i/_1884_ ),
    .B2(\cs_registers_i/_1195_ ),
    .A2(\cs_registers_i/_1883_ ),
    .A1(net680));
 sg13g2_nand2_1 \cs_registers_i/_4615_  (.Y(\cs_registers_i/_1885_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_29_ ),
    .B(\cs_registers_i/_1879_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4616_  (.Y(\cs_registers_i/_1886_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_30_ ),
    .B(\cs_registers_i/_1885_ ));
 sg13g2_mux2_1 \cs_registers_i/_4617_  (.A0(\cs_registers_i/_1224_ ),
    .A1(\cs_registers_i/_1886_ ),
    .S(net627),
    .X(\cs_registers_i/_0236_ ));
 sg13g2_nand4_1 \cs_registers_i/_4618_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_29_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_30_ ),
    .Y(\cs_registers_i/_1887_ ),
    .D(\cs_registers_i/_1871_ ));
 sg13g2_nor2_1 \cs_registers_i/_4619_  (.A(\cs_registers_i/_1858_ ),
    .B(\cs_registers_i/_1887_ ),
    .Y(\cs_registers_i/_1888_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4620_  (.Y(\cs_registers_i/_1889_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_31_ ),
    .B(\cs_registers_i/_1888_ ));
 sg13g2_nor2_2 \cs_registers_i/_4621_  (.A(net1036),
    .B(net628),
    .Y(\cs_registers_i/_1890_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4622_  (.B1(\cs_registers_i/_1890_ ),
    .Y(\cs_registers_i/_0237_ ),
    .A2(\cs_registers_i/_1889_ ),
    .A1(net628));
 sg13g2_inv_2 \cs_registers_i/_4623_  (.Y(\cs_registers_i/_1891_ ),
    .A(\cs_registers_i/_0580_ ));
 sg13g2_nor2_1 \cs_registers_i/_4624_  (.A(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .B(\cs_registers_i/_1768_ ),
    .Y(\cs_registers_i/_1892_ ));
 sg13g2_nor3_2 \cs_registers_i/_4625_  (.A(\cs_registers_i/_1891_ ),
    .B(\cs_registers_i/_1760_ ),
    .C(\cs_registers_i/_1892_ ),
    .Y(\cs_registers_i/_1893_ ));
 sg13g2_inv_1 \cs_registers_i/_4626_  (.Y(\cs_registers_i/_1894_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_31_ ));
 sg13g2_nor3_2 \cs_registers_i/_4627_  (.A(\cs_registers_i/_1894_ ),
    .B(\cs_registers_i/_1857_ ),
    .C(\cs_registers_i/_1887_ ),
    .Y(\cs_registers_i/_1895_ ));
 sg13g2_and2_2 \cs_registers_i/_4628_  (.A(net25),
    .B(\cs_registers_i/_1895_ ),
    .X(\cs_registers_i/_1896_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4629_  (.B1(net626),
    .Y(\cs_registers_i/_1897_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1895_ ));
 sg13g2_mux2_1 \cs_registers_i/_4630_  (.A0(\cs_registers_i/_1896_ ),
    .A1(\cs_registers_i/_1897_ ),
    .S(\cs_registers_i/mcycle_counter_i.counter_val_o_32_ ),
    .X(\cs_registers_i/_1898_ ));
 sg13g2_a21o_1 \cs_registers_i/_4631_  (.A2(\cs_registers_i/_1893_ ),
    .A1(net1063),
    .B1(\cs_registers_i/_1898_ ),
    .X(\cs_registers_i/_0238_ ));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(net523));
 sg13g2_nand2_2 \cs_registers_i/_4633_  (.Y(\cs_registers_i/_1900_ ),
    .A(\cs_registers_i/_1778_ ),
    .B(net16));
 sg13g2_and3_2 \cs_registers_i/_4634_  (.X(\cs_registers_i/_1901_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_32_ ),
    .B(net25),
    .C(\cs_registers_i/_1895_ ));
 sg13g2_xor2_1 \cs_registers_i/_4635_  (.B(\cs_registers_i/_1901_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .X(\cs_registers_i/_1902_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4636_  (.Y(\cs_registers_i/_1903_ ),
    .B1(\cs_registers_i/_1900_ ),
    .B2(\cs_registers_i/_1902_ ),
    .A2(net33),
    .A1(net1067));
 sg13g2_inv_1 \cs_registers_i/_4637_  (.Y(\cs_registers_i/_0239_ ),
    .A(\cs_registers_i/_1903_ ));
 sg13g2_nor2_2 \cs_registers_i/_4638_  (.A(net25),
    .B(net38),
    .Y(\cs_registers_i/_1904_ ));
 sg13g2_nand2_2 \cs_registers_i/_4639_  (.Y(\cs_registers_i/_1905_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .B(\cs_registers_i/_1901_ ));
 sg13g2_xor2_1 \cs_registers_i/_4640_  (.B(\cs_registers_i/_1905_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .X(\cs_registers_i/_1906_ ));
 sg13g2_nand2_1 \cs_registers_i/_4641_  (.Y(\cs_registers_i/_1907_ ),
    .A(net1038),
    .B(\cs_registers_i/_1893_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4642_  (.B1(\cs_registers_i/_1907_ ),
    .Y(\cs_registers_i/_0240_ ),
    .A1(\cs_registers_i/_1904_ ),
    .A2(\cs_registers_i/_1906_ ));
 sg13g2_nand3_1 \cs_registers_i/_4643_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .C(\cs_registers_i/_1901_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .Y(\cs_registers_i/_1908_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4644_  (.Y(\cs_registers_i/_1909_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_35_ ),
    .B(\cs_registers_i/_1908_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4645_  (.Y(\cs_registers_i/_1910_ ),
    .B1(\cs_registers_i/_1900_ ),
    .B2(\cs_registers_i/_1909_ ),
    .A2(net32),
    .A1(net1034));
 sg13g2_inv_1 \cs_registers_i/_4646_  (.Y(\cs_registers_i/_0241_ ),
    .A(\cs_registers_i/_1910_ ));
 sg13g2_nand4_1 \cs_registers_i/_4647_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_35_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .Y(\cs_registers_i/_1911_ ),
    .D(\cs_registers_i/_1901_ ));
 sg13g2_xor2_1 \cs_registers_i/_4648_  (.B(\cs_registers_i/_1911_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_36_ ),
    .X(\cs_registers_i/_1912_ ));
 sg13g2_nand2_1 \cs_registers_i/_4649_  (.Y(\cs_registers_i/_1913_ ),
    .A(net1032),
    .B(\cs_registers_i/_1893_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4650_  (.B1(\cs_registers_i/_1913_ ),
    .Y(\cs_registers_i/_0242_ ),
    .A1(\cs_registers_i/_1904_ ),
    .A2(\cs_registers_i/_1912_ ));
 sg13g2_buf_8 fanout471 (.A(net523),
    .X(net471));
 sg13g2_nand4_1 \cs_registers_i/_4652_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_36_ ),
    .Y(\cs_registers_i/_1915_ ),
    .D(\cs_registers_i/mcycle_counter_i.counter_val_o_35_ ));
 sg13g2_inv_1 \cs_registers_i/_4653_  (.Y(\cs_registers_i/_1916_ ),
    .A(\cs_registers_i/_1915_ ));
 sg13g2_nand2_1 \cs_registers_i/_4654_  (.Y(\cs_registers_i/_1917_ ),
    .A(\cs_registers_i/_1901_ ),
    .B(\cs_registers_i/_1916_ ));
 sg13g2_nand3_1 \cs_registers_i/_4655_  (.B(\cs_registers_i/_1900_ ),
    .C(\cs_registers_i/_1917_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_37_ ),
    .Y(\cs_registers_i/_1918_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4656_  (.B1(\cs_registers_i/_1918_ ),
    .Y(\cs_registers_i/_1919_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_37_ ),
    .A2(\cs_registers_i/_1917_ ));
 sg13g2_a21o_1 \cs_registers_i/_4657_  (.A2(net34),
    .A1(net1065),
    .B1(\cs_registers_i/_1919_ ),
    .X(\cs_registers_i/_0243_ ));
 sg13g2_and3_1 \cs_registers_i/_4658_  (.X(\cs_registers_i/_1920_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_32_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_37_ ),
    .C(\cs_registers_i/_1916_ ));
 sg13g2_nand2_2 \cs_registers_i/_4659_  (.Y(\cs_registers_i/_1921_ ),
    .A(\cs_registers_i/_1896_ ),
    .B(\cs_registers_i/_1920_ ));
 sg13g2_xor2_1 \cs_registers_i/_4660_  (.B(\cs_registers_i/_1921_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_38_ ),
    .X(\cs_registers_i/_1922_ ));
 sg13g2_nand2_1 \cs_registers_i/_4661_  (.Y(\cs_registers_i/_1923_ ),
    .A(net1064),
    .B(net31));
 sg13g2_o21ai_1 \cs_registers_i/_4662_  (.B1(\cs_registers_i/_1923_ ),
    .Y(\cs_registers_i/_0244_ ),
    .A1(\cs_registers_i/_1904_ ),
    .A2(\cs_registers_i/_1922_ ));
 sg13g2_and2_1 \cs_registers_i/_4663_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_38_ ),
    .B(\cs_registers_i/_1920_ ),
    .X(\cs_registers_i/_1924_ ));
 sg13g2_and2_1 \cs_registers_i/_4664_  (.A(\cs_registers_i/_1895_ ),
    .B(\cs_registers_i/_1924_ ),
    .X(\cs_registers_i/_1925_ ));
 sg13g2_and2_2 \cs_registers_i/_4665_  (.A(net25),
    .B(\cs_registers_i/_1925_ ),
    .X(\cs_registers_i/_1926_ ));
 sg13g2_buf_8 fanout470 (.A(net523),
    .X(net470));
 sg13g2_o21ai_1 \cs_registers_i/_4667_  (.B1(net626),
    .Y(\cs_registers_i/_1928_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1925_ ));
 sg13g2_mux2_1 \cs_registers_i/_4668_  (.A0(net721),
    .A1(\cs_registers_i/_1928_ ),
    .S(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .X(\cs_registers_i/_1929_ ));
 sg13g2_a21o_1 \cs_registers_i/_4669_  (.A2(net33),
    .A1(\cs_registers_i/_1348_ ),
    .B1(\cs_registers_i/_1929_ ),
    .X(\cs_registers_i/_0245_ ));
 sg13g2_and2_1 \cs_registers_i/_4670_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_3_ ),
    .B(\cs_registers_i/_1780_ ),
    .X(\cs_registers_i/_1930_ ));
 sg13g2_nand2_1 \cs_registers_i/_4671_  (.Y(\cs_registers_i/_1931_ ),
    .A(net29),
    .B(\cs_registers_i/_1930_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4672_  (.B1(\cs_registers_i/_1931_ ),
    .Y(\cs_registers_i/_1932_ ),
    .A1(net1033),
    .A2(net27));
 sg13g2_o21ai_1 \cs_registers_i/_4673_  (.B1(net679),
    .Y(\cs_registers_i/_1933_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1780_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4674_  (.Y(\cs_registers_i/_0246_ ),
    .B1(\cs_registers_i/_1933_ ),
    .B2(\cs_registers_i/_1265_ ),
    .A2(\cs_registers_i/_1932_ ),
    .A1(net679));
 sg13g2_or2_2 \cs_registers_i/_4675_  (.X(\cs_registers_i/_1934_ ),
    .B(net25),
    .A(\cs_registers_i/_1760_ ));
 sg13g2_buf_8 fanout469 (.A(net523),
    .X(net469));
 sg13g2_inv_1 \cs_registers_i/_4677_  (.Y(\cs_registers_i/_1936_ ),
    .A(net720));
 sg13g2_nand2_2 \cs_registers_i/_4678_  (.Y(\cs_registers_i/_1937_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .B(net721));
 sg13g2_xor2_1 \cs_registers_i/_4679_  (.B(\cs_registers_i/_1937_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .X(\cs_registers_i/_1938_ ));
 sg13g2_nand2_1 \cs_registers_i/_4680_  (.Y(\cs_registers_i/_1939_ ),
    .A(net1025),
    .B(net30));
 sg13g2_o21ai_1 \cs_registers_i/_4681_  (.B1(\cs_registers_i/_1939_ ),
    .Y(\cs_registers_i/_0247_ ),
    .A1(\cs_registers_i/_1936_ ),
    .A2(\cs_registers_i/_1938_ ));
 sg13g2_nand3_1 \cs_registers_i/_4682_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .C(net721),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .Y(\cs_registers_i/_1940_ ));
 sg13g2_nand3_1 \cs_registers_i/_4683_  (.B(net720),
    .C(\cs_registers_i/_1940_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ),
    .Y(\cs_registers_i/_1941_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4684_  (.B1(\cs_registers_i/_1941_ ),
    .Y(\cs_registers_i/_1942_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ),
    .A2(\cs_registers_i/_1940_ ));
 sg13g2_a21o_1 \cs_registers_i/_4685_  (.A2(net33),
    .A1(\cs_registers_i/_1396_ ),
    .B1(\cs_registers_i/_1942_ ),
    .X(\cs_registers_i/_0248_ ));
 sg13g2_nand4_1 \cs_registers_i/_4686_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .Y(\cs_registers_i/_1943_ ),
    .D(net721));
 sg13g2_nand3_1 \cs_registers_i/_4687_  (.B(net720),
    .C(\cs_registers_i/_1943_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_42_ ),
    .Y(\cs_registers_i/_1944_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4688_  (.B1(\cs_registers_i/_1944_ ),
    .Y(\cs_registers_i/_1945_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_42_ ),
    .A2(\cs_registers_i/_1943_ ));
 sg13g2_a21o_1 \cs_registers_i/_4689_  (.A2(net33),
    .A1(net1059),
    .B1(\cs_registers_i/_1945_ ),
    .X(\cs_registers_i/_0249_ ));
 sg13g2_nand2_1 \cs_registers_i/_4690_  (.Y(\cs_registers_i/_1946_ ),
    .A(net1071),
    .B(net31));
 sg13g2_nand2_1 \cs_registers_i/_4691_  (.Y(\cs_registers_i/_1947_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ),
    .B(\cs_registers_i/_1900_ ));
 sg13g2_and4_1 \cs_registers_i/_4692_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_42_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .D(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ),
    .X(\cs_registers_i/_1948_ ));
 sg13g2_nand2_1 \cs_registers_i/_4693_  (.Y(\cs_registers_i/_1949_ ),
    .A(\cs_registers_i/_1926_ ),
    .B(\cs_registers_i/_1948_ ));
 sg13g2_mux2_1 \cs_registers_i/_4694_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ),
    .A1(\cs_registers_i/_1947_ ),
    .S(\cs_registers_i/_1949_ ),
    .X(\cs_registers_i/_1950_ ));
 sg13g2_nand2_1 \cs_registers_i/_4695_  (.Y(\cs_registers_i/_0250_ ),
    .A(\cs_registers_i/_1946_ ),
    .B(\cs_registers_i/_1950_ ));
 sg13g2_nand2_1 \cs_registers_i/_4696_  (.Y(\cs_registers_i/_1951_ ),
    .A(net1028),
    .B(net31));
 sg13g2_nand2_1 \cs_registers_i/_4697_  (.Y(\cs_registers_i/_1952_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_44_ ),
    .B(\cs_registers_i/_1934_ ));
 sg13g2_nand3_1 \cs_registers_i/_4698_  (.B(net721),
    .C(\cs_registers_i/_1948_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ),
    .Y(\cs_registers_i/_1953_ ));
 sg13g2_mux2_1 \cs_registers_i/_4699_  (.A0(\cs_registers_i/mcycle_counter_i.counter_val_o_44_ ),
    .A1(\cs_registers_i/_1952_ ),
    .S(\cs_registers_i/_1953_ ),
    .X(\cs_registers_i/_1954_ ));
 sg13g2_nand2_1 \cs_registers_i/_4700_  (.Y(\cs_registers_i/_0251_ ),
    .A(\cs_registers_i/_1951_ ),
    .B(\cs_registers_i/_1954_ ));
 sg13g2_and3_1 \cs_registers_i/_4701_  (.X(\cs_registers_i/_1955_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_44_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ),
    .C(\cs_registers_i/_1948_ ));
 sg13g2_nand2_2 \cs_registers_i/_4702_  (.Y(\cs_registers_i/_1956_ ),
    .A(net721),
    .B(\cs_registers_i/_1955_ ));
 sg13g2_xor2_1 \cs_registers_i/_4703_  (.B(\cs_registers_i/_1956_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_45_ ),
    .X(\cs_registers_i/_1957_ ));
 sg13g2_nand2_1 \cs_registers_i/_4704_  (.Y(\cs_registers_i/_1958_ ),
    .A(net1058),
    .B(\cs_registers_i/_1893_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4705_  (.B1(\cs_registers_i/_1958_ ),
    .Y(\cs_registers_i/_0252_ ),
    .A1(\cs_registers_i/_1904_ ),
    .A2(\cs_registers_i/_1957_ ));
 sg13g2_and2_1 \cs_registers_i/_4706_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_45_ ),
    .B(\cs_registers_i/_1955_ ),
    .X(\cs_registers_i/_1959_ ));
 sg13g2_nand2_1 \cs_registers_i/_4707_  (.Y(\cs_registers_i/_1960_ ),
    .A(\cs_registers_i/_1925_ ),
    .B(\cs_registers_i/_1959_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4708_  (.Y(\cs_registers_i/_1961_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .B(\cs_registers_i/_1960_ ));
 sg13g2_buf_8 fanout468 (.A(net523),
    .X(net468));
 sg13g2_and3_1 \cs_registers_i/_4710_  (.X(\cs_registers_i/_1963_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .B(net18),
    .C(net39));
 sg13g2_a221oi_1 \cs_registers_i/_4711_  (.B2(\cs_registers_i/_1961_ ),
    .C1(\cs_registers_i/_1963_ ),
    .B1(net28),
    .A1(net1056),
    .Y(\cs_registers_i/_1964_ ),
    .A2(net32));
 sg13g2_inv_1 \cs_registers_i/_4712_  (.Y(\cs_registers_i/_0253_ ),
    .A(\cs_registers_i/_1964_ ));
 sg13g2_and4_2 \cs_registers_i/_4713_  (.A(net25),
    .B(\cs_registers_i/_1895_ ),
    .C(\cs_registers_i/_1924_ ),
    .D(\cs_registers_i/_1959_ ),
    .X(\cs_registers_i/_1965_ ));
 sg13g2_nand2_1 \cs_registers_i/_4714_  (.Y(\cs_registers_i/_1966_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .B(\cs_registers_i/_1965_ ));
 sg13g2_nand3_1 \cs_registers_i/_4715_  (.B(\cs_registers_i/_1900_ ),
    .C(\cs_registers_i/_1966_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_47_ ),
    .Y(\cs_registers_i/_1967_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4716_  (.B1(\cs_registers_i/_1967_ ),
    .Y(\cs_registers_i/_1968_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_47_ ),
    .A2(\cs_registers_i/_1966_ ));
 sg13g2_a21o_1 \cs_registers_i/_4717_  (.A2(net33),
    .A1(net1069),
    .B1(\cs_registers_i/_1968_ ),
    .X(\cs_registers_i/_0254_ ));
 sg13g2_and2_1 \cs_registers_i/_4718_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_47_ ),
    .X(\cs_registers_i/_1969_ ));
 sg13g2_nand2_1 \cs_registers_i/_4719_  (.Y(\cs_registers_i/_1970_ ),
    .A(\cs_registers_i/_1965_ ),
    .B(\cs_registers_i/_1969_ ));
 sg13g2_and2_1 \cs_registers_i/_4720_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .B(\cs_registers_i/_1934_ ),
    .X(\cs_registers_i/_1971_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4721_  (.Y(\cs_registers_i/_1972_ ),
    .B1(\cs_registers_i/_1970_ ),
    .B2(\cs_registers_i/_1971_ ),
    .A2(net32),
    .A1(\cs_registers_i/_0834_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4722_  (.B1(\cs_registers_i/_1972_ ),
    .Y(\cs_registers_i/_0255_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .A2(\cs_registers_i/_1970_ ));
 sg13g2_nand3_1 \cs_registers_i/_4723_  (.B(\cs_registers_i/_1965_ ),
    .C(\cs_registers_i/_1969_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .Y(\cs_registers_i/_1973_ ));
 sg13g2_nand3_1 \cs_registers_i/_4724_  (.B(net720),
    .C(\cs_registers_i/_1973_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .Y(\cs_registers_i/_1974_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4725_  (.B1(\cs_registers_i/_1974_ ),
    .Y(\cs_registers_i/_1975_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .A2(\cs_registers_i/_1973_ ));
 sg13g2_a21o_1 \cs_registers_i/_4726_  (.A2(net33),
    .A1(net1054),
    .B1(\cs_registers_i/_1975_ ),
    .X(\cs_registers_i/_0256_ ));
 sg13g2_nand3_1 \cs_registers_i/_4727_  (.B(net27),
    .C(\cs_registers_i/_1930_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .Y(\cs_registers_i/_1976_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4728_  (.B1(\cs_registers_i/_1976_ ),
    .Y(\cs_registers_i/_1977_ ),
    .A1(net1032),
    .A2(net27));
 sg13g2_o21ai_1 \cs_registers_i/_4729_  (.B1(net679),
    .Y(\cs_registers_i/_1978_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1930_ ));
 sg13g2_inv_1 \cs_registers_i/_4730_  (.Y(\cs_registers_i/_1979_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4731_  (.Y(\cs_registers_i/_0257_ ),
    .B1(\cs_registers_i/_1978_ ),
    .B2(\cs_registers_i/_1979_ ),
    .A2(\cs_registers_i/_1977_ ),
    .A1(net679));
 sg13g2_nand4_1 \cs_registers_i/_4732_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .C(\cs_registers_i/_1965_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .Y(\cs_registers_i/_1980_ ),
    .D(\cs_registers_i/_1969_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4733_  (.Y(\cs_registers_i/_1981_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_50_ ),
    .B(\cs_registers_i/_1980_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4734_  (.Y(\cs_registers_i/_1982_ ),
    .B1(net720),
    .B2(\cs_registers_i/_1981_ ),
    .A2(net32),
    .A1(net1052));
 sg13g2_inv_1 \cs_registers_i/_4735_  (.Y(\cs_registers_i/_0258_ ),
    .A(\cs_registers_i/_1982_ ));
 sg13g2_and2_1 \cs_registers_i/_4736_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_50_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .X(\cs_registers_i/_1983_ ));
 sg13g2_nand4_1 \cs_registers_i/_4737_  (.B(\cs_registers_i/_1965_ ),
    .C(\cs_registers_i/_1969_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .Y(\cs_registers_i/_1984_ ),
    .D(\cs_registers_i/_1983_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4738_  (.Y(\cs_registers_i/_1985_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_51_ ),
    .B(\cs_registers_i/_1984_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4739_  (.Y(\cs_registers_i/_1986_ ),
    .B1(net720),
    .B2(\cs_registers_i/_1985_ ),
    .A2(net32),
    .A1(net1050));
 sg13g2_inv_1 \cs_registers_i/_4740_  (.Y(\cs_registers_i/_0259_ ),
    .A(\cs_registers_i/_1986_ ));
 sg13g2_and4_1 \cs_registers_i/_4741_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_51_ ),
    .C(\cs_registers_i/_1969_ ),
    .D(\cs_registers_i/_1983_ ),
    .X(\cs_registers_i/_1987_ ));
 sg13g2_nand2_2 \cs_registers_i/_4742_  (.Y(\cs_registers_i/_1988_ ),
    .A(\cs_registers_i/_1965_ ),
    .B(\cs_registers_i/_1987_ ));
 sg13g2_xor2_1 \cs_registers_i/_4743_  (.B(\cs_registers_i/_1988_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_52_ ),
    .X(\cs_registers_i/_1989_ ));
 sg13g2_nand2_1 \cs_registers_i/_4744_  (.Y(\cs_registers_i/_1990_ ),
    .A(net1049),
    .B(\cs_registers_i/_1893_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4745_  (.B1(\cs_registers_i/_1990_ ),
    .Y(\cs_registers_i/_0260_ ),
    .A1(\cs_registers_i/_1904_ ),
    .A2(\cs_registers_i/_1989_ ));
 sg13g2_nor2_2 \cs_registers_i/_4746_  (.A(net682),
    .B(net27),
    .Y(\cs_registers_i/_1991_ ));
 sg13g2_and2_1 \cs_registers_i/_4747_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_52_ ),
    .B(\cs_registers_i/_1987_ ),
    .X(\cs_registers_i/_1992_ ));
 sg13g2_nand3_1 \cs_registers_i/_4748_  (.B(\cs_registers_i/_1959_ ),
    .C(\cs_registers_i/_1992_ ),
    .A(net721),
    .Y(\cs_registers_i/_1993_ ));
 sg13g2_xor2_1 \cs_registers_i/_4749_  (.B(\cs_registers_i/_1993_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_53_ ),
    .X(\cs_registers_i/_1994_ ));
 sg13g2_nand2_1 \cs_registers_i/_4750_  (.Y(\cs_registers_i/_1995_ ),
    .A(net1048),
    .B(net30));
 sg13g2_o21ai_1 \cs_registers_i/_4751_  (.B1(\cs_registers_i/_1995_ ),
    .Y(\cs_registers_i/_0261_ ),
    .A1(\cs_registers_i/_1991_ ),
    .A2(\cs_registers_i/_1994_ ));
 sg13g2_nand4_1 \cs_registers_i/_4752_  (.B(net721),
    .C(\cs_registers_i/_1959_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_53_ ),
    .Y(\cs_registers_i/_1996_ ),
    .D(\cs_registers_i/_1992_ ));
 sg13g2_xor2_1 \cs_registers_i/_4753_  (.B(\cs_registers_i/_1996_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_54_ ),
    .X(\cs_registers_i/_1997_ ));
 sg13g2_nand2_1 \cs_registers_i/_4754_  (.Y(\cs_registers_i/_1998_ ),
    .A(net1027),
    .B(net30));
 sg13g2_o21ai_1 \cs_registers_i/_4755_  (.B1(\cs_registers_i/_1998_ ),
    .Y(\cs_registers_i/_0262_ ),
    .A1(\cs_registers_i/_1991_ ),
    .A2(\cs_registers_i/_1997_ ));
 sg13g2_nor3_1 \cs_registers_i/_4756_  (.A(net149),
    .B(\cs_registers_i/_1030_ ),
    .C(\cs_registers_i/_1760_ ),
    .Y(\cs_registers_i/_1999_ ));
 sg13g2_nand3_1 \cs_registers_i/_4757_  (.B(csr_op_1_),
    .C(csr_op_0_),
    .A(net150),
    .Y(\cs_registers_i/_2000_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4758_  (.A(\cs_registers_i/_1760_ ),
    .B_N(\cs_registers_i/_2000_ ),
    .Y(\cs_registers_i/_2001_ ));
 sg13g2_and3_1 \cs_registers_i/_4759_  (.X(\cs_registers_i/_2002_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_55_ ),
    .B(\cs_registers_i/_1760_ ),
    .C(\cs_registers_i/_1768_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4760_  (.B1(\cs_registers_i/_0579_ ),
    .Y(\cs_registers_i/_2003_ ),
    .A1(\cs_registers_i/_2001_ ),
    .A2(\cs_registers_i/_2002_ ));
 sg13g2_and4_1 \cs_registers_i/_4761_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_54_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_53_ ),
    .C(\cs_registers_i/_1959_ ),
    .D(\cs_registers_i/_1992_ ),
    .X(\cs_registers_i/_2004_ ));
 sg13g2_nand2_1 \cs_registers_i/_4762_  (.Y(\cs_registers_i/_2005_ ),
    .A(\cs_registers_i/_1925_ ),
    .B(\cs_registers_i/_2004_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4763_  (.Y(\cs_registers_i/_2006_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_55_ ),
    .B(\cs_registers_i/_2005_ ));
 sg13g2_nand2_2 \cs_registers_i/_4764_  (.Y(\cs_registers_i/_2007_ ),
    .A(net28),
    .B(\cs_registers_i/_2006_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4765_  (.B1(\cs_registers_i/_2007_ ),
    .Y(\cs_registers_i/_0263_ ),
    .A1(\cs_registers_i/_1999_ ),
    .A2(\cs_registers_i/_2003_ ));
 sg13g2_and2_1 \cs_registers_i/_4766_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_55_ ),
    .B(\cs_registers_i/_2004_ ),
    .X(\cs_registers_i/_2008_ ));
 sg13g2_nand4_1 \cs_registers_i/_4767_  (.B(\cs_registers_i/_1895_ ),
    .C(\cs_registers_i/_1924_ ),
    .A(net28),
    .Y(\cs_registers_i/_2009_ ),
    .D(\cs_registers_i/_2008_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4768_  (.Y(\cs_registers_i/_2010_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_56_ ),
    .B(\cs_registers_i/_2009_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4769_  (.Y(\cs_registers_i/_2011_ ),
    .B1(net720),
    .B2(\cs_registers_i/_2010_ ),
    .A2(net32),
    .A1(net1045));
 sg13g2_inv_1 \cs_registers_i/_4770_  (.Y(\cs_registers_i/_0264_ ),
    .A(\cs_registers_i/_2011_ ));
 sg13g2_nand4_1 \cs_registers_i/_4771_  (.B(\cs_registers_i/_1896_ ),
    .C(\cs_registers_i/_1924_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_56_ ),
    .Y(\cs_registers_i/_2012_ ),
    .D(\cs_registers_i/_2008_ ));
 sg13g2_nand3b_1 \cs_registers_i/_4772_  (.B(\cs_registers_i/_2012_ ),
    .C(\cs_registers_i/mcycle_counter_i.counter_val_o_57_ ),
    .Y(\cs_registers_i/_2013_ ),
    .A_N(\cs_registers_i/_1904_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4773_  (.B1(\cs_registers_i/_2013_ ),
    .Y(\cs_registers_i/_2014_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_57_ ),
    .A2(\cs_registers_i/_2012_ ));
 sg13g2_a21o_1 \cs_registers_i/_4774_  (.A2(net33),
    .A1(net1043),
    .B1(\cs_registers_i/_2014_ ),
    .X(\cs_registers_i/_0265_ ));
 sg13g2_nand2_1 \cs_registers_i/_4775_  (.Y(\cs_registers_i/_2015_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_56_ ),
    .B(\cs_registers_i/mcycle_counter_i.counter_val_o_57_ ));
 sg13g2_nor2_2 \cs_registers_i/_4776_  (.A(\cs_registers_i/_2009_ ),
    .B(\cs_registers_i/_2015_ ),
    .Y(\cs_registers_i/_2016_ ));
 sg13g2_nand2_2 \cs_registers_i/_4777_  (.Y(\cs_registers_i/_2017_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_58_ ),
    .B(\cs_registers_i/_1900_ ));
 sg13g2_inv_1 \cs_registers_i/_4778_  (.Y(\cs_registers_i/_2018_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_58_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4779_  (.Y(\cs_registers_i/_2019_ ),
    .B1(\cs_registers_i/_2016_ ),
    .B2(\cs_registers_i/_2018_ ),
    .A2(\cs_registers_i/_1778_ ),
    .A1(net1066));
 sg13g2_o21ai_1 \cs_registers_i/_4780_  (.B1(\cs_registers_i/_2019_ ),
    .Y(\cs_registers_i/_0266_ ),
    .A1(\cs_registers_i/_2016_ ),
    .A2(\cs_registers_i/_2017_ ));
 sg13g2_nand2_2 \cs_registers_i/_4781_  (.Y(\cs_registers_i/_2020_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_58_ ),
    .B(\cs_registers_i/_2016_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4782_  (.Y(\cs_registers_i/_2021_ ),
    .A(\cs_registers_i/_1113_ ),
    .B(\cs_registers_i/_2020_ ));
 sg13g2_nand2_1 \cs_registers_i/_4783_  (.Y(\cs_registers_i/_2022_ ),
    .A(net1026),
    .B(net30));
 sg13g2_o21ai_1 \cs_registers_i/_4784_  (.B1(\cs_registers_i/_2022_ ),
    .Y(\cs_registers_i/_0267_ ),
    .A1(\cs_registers_i/_1991_ ),
    .A2(\cs_registers_i/_2021_ ));
 sg13g2_nand3_1 \cs_registers_i/_4785_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_5_ ),
    .C(\cs_registers_i/_1930_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .Y(\cs_registers_i/_2023_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4786_  (.Y(\cs_registers_i/_2024_ ),
    .B(net27),
    .A_N(\cs_registers_i/_2023_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4787_  (.B1(\cs_registers_i/_2024_ ),
    .Y(\cs_registers_i/_2025_ ),
    .A1(net1065),
    .A2(net26));
 sg13g2_a21o_1 \cs_registers_i/_4788_  (.A2(\cs_registers_i/_1930_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .B1(net18),
    .X(\cs_registers_i/_2026_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4789_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_5_ ),
    .Y(\cs_registers_i/_2027_ ),
    .A2(\cs_registers_i/_2026_ ),
    .A1(net679));
 sg13g2_a21oi_1 \cs_registers_i/_4790_  (.A1(net679),
    .A2(\cs_registers_i/_2025_ ),
    .Y(\cs_registers_i/_0268_ ),
    .B1(\cs_registers_i/_2027_ ));
 sg13g2_nor3_2 \cs_registers_i/_4791_  (.A(\cs_registers_i/_2018_ ),
    .B(\cs_registers_i/_1113_ ),
    .C(\cs_registers_i/_2015_ ),
    .Y(\cs_registers_i/_2028_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4792_  (.Y(\cs_registers_i/_2029_ ),
    .B(\cs_registers_i/_2028_ ),
    .A_N(\cs_registers_i/_2009_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4793_  (.Y(\cs_registers_i/_2030_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_60_ ),
    .B(\cs_registers_i/_2029_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4794_  (.Y(\cs_registers_i/_2031_ ),
    .B1(\cs_registers_i/_1900_ ),
    .B2(\cs_registers_i/_2030_ ),
    .A2(net32),
    .A1(net1042));
 sg13g2_inv_1 \cs_registers_i/_4795_  (.Y(\cs_registers_i/_0269_ ),
    .A(\cs_registers_i/_2031_ ));
 sg13g2_nand2_1 \cs_registers_i/_4796_  (.Y(\cs_registers_i/_2032_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_60_ ),
    .B(\cs_registers_i/_2028_ ));
 sg13g2_or2_1 \cs_registers_i/_4797_  (.X(\cs_registers_i/_2033_ ),
    .B(\cs_registers_i/_2032_ ),
    .A(\cs_registers_i/_2009_ ));
 sg13g2_nand3_1 \cs_registers_i/_4798_  (.B(net720),
    .C(\cs_registers_i/_2033_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_61_ ),
    .Y(\cs_registers_i/_2034_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4799_  (.B1(\cs_registers_i/_2034_ ),
    .Y(\cs_registers_i/_2035_ ),
    .A1(\cs_registers_i/mcycle_counter_i.counter_val_o_61_ ),
    .A2(\cs_registers_i/_2033_ ));
 sg13g2_a21o_1 \cs_registers_i/_4800_  (.A2(net33),
    .A1(net1041),
    .B1(\cs_registers_i/_2035_ ),
    .X(\cs_registers_i/_0270_ ));
 sg13g2_nand3_1 \cs_registers_i/_4801_  (.B(\cs_registers_i/mcycle_counter_i.counter_val_o_61_ ),
    .C(\cs_registers_i/_2028_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_60_ ),
    .Y(\cs_registers_i/_2036_ ));
 sg13g2_inv_1 \cs_registers_i/_4802_  (.Y(\cs_registers_i/_2037_ ),
    .A(\cs_registers_i/_2036_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4803_  (.Y(\cs_registers_i/_2038_ ),
    .B(\cs_registers_i/_2037_ ),
    .A_N(\cs_registers_i/_2009_ ));
 sg13g2_and2_1 \cs_registers_i/_4804_  (.A(\cs_registers_i/_1900_ ),
    .B(\cs_registers_i/_2038_ ),
    .X(\cs_registers_i/_2039_ ));
 sg13g2_nor2_1 \cs_registers_i/_4805_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_62_ ),
    .B(\cs_registers_i/_2038_ ),
    .Y(\cs_registers_i/_2040_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4806_  (.B2(\cs_registers_i/mcycle_counter_i.counter_val_o_62_ ),
    .C1(\cs_registers_i/_2040_ ),
    .B1(\cs_registers_i/_2039_ ),
    .A1(net1037),
    .Y(\cs_registers_i/_2041_ ),
    .A2(net32));
 sg13g2_inv_1 \cs_registers_i/_4807_  (.Y(\cs_registers_i/_0271_ ),
    .A(\cs_registers_i/_2041_ ));
 sg13g2_nand4_1 \cs_registers_i/_4808_  (.B(\cs_registers_i/_1925_ ),
    .C(\cs_registers_i/_2008_ ),
    .A(\cs_registers_i/mcycle_counter_i.counter_val_o_62_ ),
    .Y(\cs_registers_i/_2042_ ),
    .D(\cs_registers_i/_2037_ ));
 sg13g2_a21o_1 \cs_registers_i/_4809_  (.A2(\cs_registers_i/_2042_ ),
    .A1(net28),
    .B1(\cs_registers_i/_1876_ ),
    .X(\cs_registers_i/_2043_ ));
 sg13g2_nor3_1 \cs_registers_i/_4810_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_63_ ),
    .B(net17),
    .C(\cs_registers_i/_2042_ ),
    .Y(\cs_registers_i/_2044_ ));
 sg13g2_a221oi_1 \cs_registers_i/_4811_  (.B2(\cs_registers_i/mcycle_counter_i.counter_val_o_63_ ),
    .C1(\cs_registers_i/_2044_ ),
    .B1(\cs_registers_i/_2043_ ),
    .A1(net1036),
    .Y(\cs_registers_i/_2045_ ),
    .A2(\cs_registers_i/_1893_ ));
 sg13g2_inv_1 \cs_registers_i/_4812_  (.Y(\cs_registers_i/_0272_ ),
    .A(\cs_registers_i/_2045_ ));
 sg13g2_nand2_2 \cs_registers_i/_4813_  (.Y(\cs_registers_i/_2046_ ),
    .A(net29),
    .B(\cs_registers_i/_1782_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4814_  (.B1(\cs_registers_i/_2046_ ),
    .Y(\cs_registers_i/_2047_ ),
    .A1(net1064),
    .A2(net25));
 sg13g2_nand2_1 \cs_registers_i/_4815_  (.Y(\cs_registers_i/_2048_ ),
    .A(net29),
    .B(\cs_registers_i/_2023_ ));
 sg13g2_a21oi_2 \cs_registers_i/_4816_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_6_ ),
    .Y(\cs_registers_i/_2049_ ),
    .A2(\cs_registers_i/_2048_ ),
    .A1(net680));
 sg13g2_a21oi_1 \cs_registers_i/_4817_  (.A1(\cs_registers_i/_1763_ ),
    .A2(\cs_registers_i/_2047_ ),
    .Y(\cs_registers_i/_0273_ ),
    .B1(\cs_registers_i/_2049_ ));
 sg13g2_nand2_1 \cs_registers_i/_4818_  (.Y(\cs_registers_i/_2050_ ),
    .A(net29),
    .B(\cs_registers_i/_1784_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4819_  (.B1(\cs_registers_i/_2050_ ),
    .Y(\cs_registers_i/_2051_ ),
    .A1(net1031),
    .A2(net27));
 sg13g2_o21ai_1 \cs_registers_i/_4820_  (.B1(net680),
    .Y(\cs_registers_i/_2052_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1782_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4821_  (.Y(\cs_registers_i/_0274_ ),
    .B1(\cs_registers_i/_2052_ ),
    .B2(\cs_registers_i/_1332_ ),
    .A2(\cs_registers_i/_2051_ ),
    .A1(net680));
 sg13g2_nand2_1 \cs_registers_i/_4822_  (.Y(\cs_registers_i/_2053_ ),
    .A(net29),
    .B(\cs_registers_i/_1785_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4823_  (.B1(\cs_registers_i/_2053_ ),
    .Y(\cs_registers_i/_2054_ ),
    .A1(net1025),
    .A2(net26));
 sg13g2_o21ai_1 \cs_registers_i/_4824_  (.B1(net680),
    .Y(\cs_registers_i/_2055_ ),
    .A1(net16),
    .A2(\cs_registers_i/_1784_ ));
 sg13g2_a22oi_1 \cs_registers_i/_4825_  (.Y(\cs_registers_i/_0275_ ),
    .B1(\cs_registers_i/_2055_ ),
    .B2(\cs_registers_i/_1360_ ),
    .A2(\cs_registers_i/_2054_ ),
    .A1(net680));
 sg13g2_inv_1 \cs_registers_i/_4826_  (.Y(\cs_registers_i/_2056_ ),
    .A(\cs_registers_i/_1785_ ));
 sg13g2_nor3_1 \cs_registers_i/_4827_  (.A(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ),
    .B(net17),
    .C(\cs_registers_i/_2056_ ),
    .Y(\cs_registers_i/_2057_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4828_  (.A1(\cs_registers_i/_1396_ ),
    .A2(net18),
    .Y(\cs_registers_i/_2058_ ),
    .B1(\cs_registers_i/_2057_ ));
 sg13g2_nor2_1 \cs_registers_i/_4829_  (.A(net17),
    .B(\cs_registers_i/_1785_ ),
    .Y(\cs_registers_i/_2059_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4830_  (.B1(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ),
    .Y(\cs_registers_i/_2060_ ),
    .A1(\cs_registers_i/_1778_ ),
    .A2(\cs_registers_i/_2059_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4831_  (.B1(\cs_registers_i/_2060_ ),
    .Y(\cs_registers_i/_0276_ ),
    .A1(\cs_registers_i/_1778_ ),
    .A2(\cs_registers_i/_2058_ ));
 sg13g2_nand4_1 \cs_registers_i/_4832_  (.B(\cs_registers_i/_1759_ ),
    .C(net1156),
    .A(\cs_registers_i/_1290_ ),
    .Y(\cs_registers_i/_2061_ ),
    .D(\cs_registers_i/_1766_ ));
 sg13g2_nor3_2 \cs_registers_i/_4833_  (.A(\cs_registers_i/_0571_ ),
    .B(\cs_registers_i/_0578_ ),
    .C(\cs_registers_i/_2061_ ),
    .Y(\cs_registers_i/_2062_ ));
 sg13g2_and2_2 \cs_registers_i/_4834_  (.A(perf_instr_ret_wb),
    .B(\cs_registers_i/minstret_counter_i.counter_inc_i_$_AND__Y_B ),
    .X(\cs_registers_i/_2063_ ));
 sg13g2_nand2b_1 \cs_registers_i/_4835_  (.Y(\cs_registers_i/_2064_ ),
    .B(\cs_registers_i/_2063_ ),
    .A_N(net733));
 sg13g2_mux2_1 \cs_registers_i/_4836_  (.A0(\cs_registers_i/minstret_counter_i.counter_val_upd_o_0_ ),
    .A1(\cs_registers_i/mhpmcounter_1856_ ),
    .S(\cs_registers_i/_2064_ ),
    .X(\cs_registers_i/_2065_ ));
 sg13g2_nand2_1 \cs_registers_i/_4837_  (.Y(\cs_registers_i/_2066_ ),
    .A(\cs_registers_i/_1290_ ),
    .B(\cs_registers_i/_1766_ ));
 sg13g2_nor4_2 \cs_registers_i/_4838_  (.A(\cs_registers_i/_0571_ ),
    .B(\cs_registers_i/_0578_ ),
    .C(\cs_registers_i/_0876_ ),
    .Y(\cs_registers_i/_2067_ ),
    .D(\cs_registers_i/_2066_ ));
 sg13g2_nand2_2 \cs_registers_i/_4839_  (.Y(\cs_registers_i/_2068_ ),
    .A(net39),
    .B(net19));
 sg13g2_mux2_1 \cs_registers_i/_4840_  (.A0(\cs_registers_i/_1694_ ),
    .A1(\cs_registers_i/_2065_ ),
    .S(net719),
    .X(\cs_registers_i/_0277_ ));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(net523));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(net523));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(net523));
 sg13g2_nand2_2 \cs_registers_i/_4844_  (.Y(\cs_registers_i/_2072_ ),
    .A(\cs_registers_i/mhpmcounter_1856_ ),
    .B(\cs_registers_i/_2063_ ));
 sg13g2_nor3_1 \cs_registers_i/_4845_  (.A(\cs_registers_i/mhpmcounter_1857_ ),
    .B(net21),
    .C(\cs_registers_i/_2072_ ),
    .Y(\cs_registers_i/_2073_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4846_  (.A1(net1067),
    .A2(net22),
    .Y(\cs_registers_i/_2074_ ),
    .B1(\cs_registers_i/_2073_ ));
 sg13g2_nor2b_2 \cs_registers_i/_4847_  (.A(net22),
    .B_N(\cs_registers_i/_2072_ ),
    .Y(\cs_registers_i/_2075_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4848_  (.B1(\cs_registers_i/mhpmcounter_1857_ ),
    .Y(\cs_registers_i/_2076_ ),
    .A1(net733),
    .A2(\cs_registers_i/_2075_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4849_  (.B1(\cs_registers_i/_2076_ ),
    .Y(\cs_registers_i/_0278_ ),
    .A1(net733),
    .A2(\cs_registers_i/_2074_ ));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(net524));
 sg13g2_and4_1 \cs_registers_i/_4851_  (.A(\cs_registers_i/mhpmcounter_1856_ ),
    .B(\cs_registers_i/mhpmcounter_1857_ ),
    .C(perf_instr_ret_wb),
    .D(\cs_registers_i/minstret_counter_i.counter_inc_i_$_AND__Y_B ),
    .X(\cs_registers_i/_2078_ ));
 sg13g2_nor2b_2 \cs_registers_i/_4852_  (.A(net733),
    .B_N(\cs_registers_i/_2078_ ),
    .Y(\cs_registers_i/_2079_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4853_  (.Y(\cs_registers_i/_2080_ ),
    .A(\cs_registers_i/mhpmcounter_1858_ ),
    .B(\cs_registers_i/_2079_ ));
 sg13g2_nor2_2 \cs_registers_i/_4854_  (.A(net1038),
    .B(net719),
    .Y(\cs_registers_i/_2081_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4855_  (.A1(net719),
    .A2(\cs_registers_i/_2080_ ),
    .Y(\cs_registers_i/_0279_ ),
    .B1(\cs_registers_i/_2081_ ));
 sg13g2_nand2_2 \cs_registers_i/_4856_  (.Y(\cs_registers_i/_2082_ ),
    .A(\cs_registers_i/mhpmcounter_1858_ ),
    .B(\cs_registers_i/_2078_ ));
 sg13g2_nor3_1 \cs_registers_i/_4857_  (.A(\cs_registers_i/mhpmcounter_1859_ ),
    .B(net21),
    .C(\cs_registers_i/_2082_ ),
    .Y(\cs_registers_i/_2083_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4858_  (.A1(net1034),
    .A2(net22),
    .Y(\cs_registers_i/_2084_ ),
    .B1(\cs_registers_i/_2083_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4859_  (.A(net23),
    .B_N(\cs_registers_i/_2082_ ),
    .Y(\cs_registers_i/_2085_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4860_  (.B1(\cs_registers_i/mhpmcounter_1859_ ),
    .Y(\cs_registers_i/_2086_ ),
    .A1(net734),
    .A2(\cs_registers_i/_2085_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4861_  (.B1(\cs_registers_i/_2086_ ),
    .Y(\cs_registers_i/_0280_ ),
    .A1(net734),
    .A2(\cs_registers_i/_2084_ ));
 sg13g2_inv_1 \cs_registers_i/_4862_  (.Y(\cs_registers_i/_2087_ ),
    .A(\cs_registers_i/_1286_ ));
 sg13g2_and2_1 \cs_registers_i/_4863_  (.A(net38),
    .B(net19),
    .X(\cs_registers_i/_2088_ ));
 sg13g2_inv_1 \cs_registers_i/_4864_  (.Y(\cs_registers_i/_2089_ ),
    .A(\cs_registers_i/mhpmcounter_1860_ ));
 sg13g2_nand3_1 \cs_registers_i/_4865_  (.B(\cs_registers_i/mhpmcounter_1859_ ),
    .C(\cs_registers_i/_2078_ ),
    .A(\cs_registers_i/mhpmcounter_1858_ ),
    .Y(\cs_registers_i/_2090_ ));
 sg13g2_nor2_1 \cs_registers_i/_4866_  (.A(net733),
    .B(\cs_registers_i/_2090_ ),
    .Y(\cs_registers_i/_2091_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4867_  (.Y(\cs_registers_i/_2092_ ),
    .A(\cs_registers_i/_2089_ ),
    .B(\cs_registers_i/_2091_ ));
 sg13g2_nor2_1 \cs_registers_i/_4868_  (.A(\cs_registers_i/_2088_ ),
    .B(\cs_registers_i/_2092_ ),
    .Y(\cs_registers_i/_2093_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4869_  (.A1(\cs_registers_i/_2087_ ),
    .A2(\cs_registers_i/_2088_ ),
    .Y(\cs_registers_i/_0281_ ),
    .B1(\cs_registers_i/_2093_ ));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(\id_stage_i.controller_i.instr_i_21_ ));
 sg13g2_nor4_1 \cs_registers_i/_4871_  (.A(\cs_registers_i/_2089_ ),
    .B(\cs_registers_i/mhpmcounter_1861_ ),
    .C(net21),
    .D(\cs_registers_i/_2090_ ),
    .Y(\cs_registers_i/_2095_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4872_  (.A1(net1065),
    .A2(net22),
    .Y(\cs_registers_i/_2096_ ),
    .B1(\cs_registers_i/_2095_ ));
 sg13g2_nor2_2 \cs_registers_i/_4873_  (.A(\cs_registers_i/_2089_ ),
    .B(\cs_registers_i/_2090_ ),
    .Y(\cs_registers_i/_2097_ ));
 sg13g2_nor2_1 \cs_registers_i/_4874_  (.A(net20),
    .B(\cs_registers_i/_2097_ ),
    .Y(\cs_registers_i/_2098_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4875_  (.B1(\cs_registers_i/mhpmcounter_1861_ ),
    .Y(\cs_registers_i/_2099_ ),
    .A1(net734),
    .A2(\cs_registers_i/_2098_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4876_  (.B1(\cs_registers_i/_2099_ ),
    .Y(\cs_registers_i/_0282_ ),
    .A1(net734),
    .A2(\cs_registers_i/_2096_ ));
 sg13g2_nand2_2 \cs_registers_i/_4877_  (.Y(\cs_registers_i/_2100_ ),
    .A(\cs_registers_i/mhpmcounter_1861_ ),
    .B(\cs_registers_i/_2097_ ));
 sg13g2_nor3_1 \cs_registers_i/_4878_  (.A(\cs_registers_i/mhpmcounter_1862_ ),
    .B(net20),
    .C(\cs_registers_i/_2100_ ),
    .Y(\cs_registers_i/_2101_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4879_  (.A1(net1064),
    .A2(net22),
    .Y(\cs_registers_i/_2102_ ),
    .B1(\cs_registers_i/_2101_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4880_  (.A(net22),
    .B_N(\cs_registers_i/_2100_ ),
    .Y(\cs_registers_i/_2103_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4881_  (.B1(\cs_registers_i/mhpmcounter_1862_ ),
    .Y(\cs_registers_i/_2104_ ),
    .A1(net734),
    .A2(\cs_registers_i/_2103_ ));
 sg13g2_o21ai_1 \cs_registers_i/_4882_  (.B1(\cs_registers_i/_2104_ ),
    .Y(\cs_registers_i/_0283_ ),
    .A1(net733),
    .A2(\cs_registers_i/_2102_ ));
 sg13g2_nand3_1 \cs_registers_i/_4883_  (.B(\cs_registers_i/mhpmcounter_1861_ ),
    .C(\cs_registers_i/_2097_ ),
    .A(\cs_registers_i/mhpmcounter_1862_ ),
    .Y(\cs_registers_i/_2105_ ));
 sg13g2_nor2_2 \cs_registers_i/_4884_  (.A(net735),
    .B(\cs_registers_i/_2105_ ),
    .Y(\cs_registers_i/_2106_ ));
 sg13g2_xor2_1 \cs_registers_i/_4885_  (.B(\cs_registers_i/_2106_ ),
    .A(\cs_registers_i/mhpmcounter_1863_ ),
    .X(\cs_registers_i/_2107_ ));
 sg13g2_nor2_1 \cs_registers_i/_4886_  (.A(\cs_registers_i/_0876_ ),
    .B(\cs_registers_i/_2066_ ),
    .Y(\cs_registers_i/_2108_ ));
 sg13g2_nand2_1 \cs_registers_i/_4887_  (.Y(\cs_registers_i/_2109_ ),
    .A(\cs_registers_i/_0579_ ),
    .B(\cs_registers_i/_2108_ ));
 sg13g2_nor2_2 \cs_registers_i/_4888_  (.A(net735),
    .B(net715),
    .Y(\cs_registers_i/_2110_ ));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(net463));
 sg13g2_mux2_1 \cs_registers_i/_4890_  (.A0(\cs_registers_i/_2107_ ),
    .A1(net1031),
    .S(net676),
    .X(\cs_registers_i/_0284_ ));
 sg13g2_nand2_1 \cs_registers_i/_4891_  (.Y(\cs_registers_i/_2112_ ),
    .A(\cs_registers_i/mhpmcounter_1863_ ),
    .B(\cs_registers_i/_2106_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4892_  (.Y(\cs_registers_i/_2113_ ),
    .A(\cs_registers_i/mhpmcounter_1864_ ),
    .B(\cs_registers_i/_2112_ ));
 sg13g2_mux2_1 \cs_registers_i/_4893_  (.A0(net1025),
    .A1(\cs_registers_i/_2113_ ),
    .S(net719),
    .X(\cs_registers_i/_0285_ ));
 sg13g2_and3_1 \cs_registers_i/_4894_  (.X(\cs_registers_i/_2114_ ),
    .A(\cs_registers_i/mhpmcounter_1864_ ),
    .B(\cs_registers_i/mhpmcounter_1863_ ),
    .C(\cs_registers_i/_2106_ ));
 sg13g2_xor2_1 \cs_registers_i/_4895_  (.B(\cs_registers_i/_2114_ ),
    .A(\cs_registers_i/mhpmcounter_1865_ ),
    .X(\cs_registers_i/_2115_ ));
 sg13g2_mux2_1 \cs_registers_i/_4896_  (.A0(\cs_registers_i/_2115_ ),
    .A1(\cs_registers_i/_1396_ ),
    .S(net676),
    .X(\cs_registers_i/_0286_ ));
 sg13g2_nand3_1 \cs_registers_i/_4897_  (.B(\cs_registers_i/mhpmcounter_1863_ ),
    .C(\cs_registers_i/mhpmcounter_1865_ ),
    .A(\cs_registers_i/mhpmcounter_1864_ ),
    .Y(\cs_registers_i/_2116_ ));
 sg13g2_nor3_2 \cs_registers_i/_4898_  (.A(net735),
    .B(\cs_registers_i/_2105_ ),
    .C(\cs_registers_i/_2116_ ),
    .Y(\cs_registers_i/_2117_ ));
 sg13g2_xor2_1 \cs_registers_i/_4899_  (.B(\cs_registers_i/_2117_ ),
    .A(\cs_registers_i/mhpmcounter_1866_ ),
    .X(\cs_registers_i/_2118_ ));
 sg13g2_mux2_1 \cs_registers_i/_4900_  (.A0(\cs_registers_i/_2118_ ),
    .A1(\cs_registers_i/_0653_ ),
    .S(net676),
    .X(\cs_registers_i/_0287_ ));
 sg13g2_nand2_1 \cs_registers_i/_4901_  (.Y(\cs_registers_i/_2119_ ),
    .A(\cs_registers_i/mhpmcounter_1866_ ),
    .B(\cs_registers_i/_2117_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4902_  (.Y(\cs_registers_i/_2120_ ),
    .A(\cs_registers_i/mhpmcounter_1867_ ),
    .B(\cs_registers_i/_2119_ ));
 sg13g2_mux2_1 \cs_registers_i/_4903_  (.A0(\cs_registers_i/_2120_ ),
    .A1(net1071),
    .S(net676),
    .X(\cs_registers_i/_0288_ ));
 sg13g2_and3_1 \cs_registers_i/_4904_  (.X(\cs_registers_i/_2121_ ),
    .A(\cs_registers_i/mhpmcounter_1866_ ),
    .B(\cs_registers_i/mhpmcounter_1867_ ),
    .C(\cs_registers_i/_2117_ ));
 sg13g2_xor2_1 \cs_registers_i/_4905_  (.B(\cs_registers_i/_2121_ ),
    .A(\cs_registers_i/mhpmcounter_1868_ ),
    .X(\cs_registers_i/_2122_ ));
 sg13g2_mux2_1 \cs_registers_i/_4906_  (.A0(\cs_registers_i/_2122_ ),
    .A1(net1028),
    .S(net676),
    .X(\cs_registers_i/_0289_ ));
 sg13g2_inv_1 \cs_registers_i/_4907_  (.Y(\cs_registers_i/_2123_ ),
    .A(\cs_registers_i/_2116_ ));
 sg13g2_nand4_1 \cs_registers_i/_4908_  (.B(\cs_registers_i/mhpmcounter_1866_ ),
    .C(\cs_registers_i/mhpmcounter_1867_ ),
    .A(\cs_registers_i/mhpmcounter_1868_ ),
    .Y(\cs_registers_i/_2124_ ),
    .D(\cs_registers_i/_2123_ ));
 sg13g2_nor3_2 \cs_registers_i/_4909_  (.A(net735),
    .B(\cs_registers_i/_2105_ ),
    .C(\cs_registers_i/_2124_ ),
    .Y(\cs_registers_i/_2125_ ));
 sg13g2_xor2_1 \cs_registers_i/_4910_  (.B(net714),
    .A(\cs_registers_i/mhpmcounter_1869_ ),
    .X(\cs_registers_i/_2126_ ));
 sg13g2_mux2_1 \cs_registers_i/_4911_  (.A0(\cs_registers_i/_2126_ ),
    .A1(net1058),
    .S(net677),
    .X(\cs_registers_i/_0290_ ));
 sg13g2_nand2_2 \cs_registers_i/_4912_  (.Y(\cs_registers_i/_2127_ ),
    .A(\cs_registers_i/mhpmcounter_1869_ ),
    .B(net714));
 sg13g2_xnor2_1 \cs_registers_i/_4913_  (.Y(\cs_registers_i/_2128_ ),
    .A(\cs_registers_i/mhpmcounter_1870_ ),
    .B(\cs_registers_i/_2127_ ));
 sg13g2_mux2_1 \cs_registers_i/_4914_  (.A0(\cs_registers_i/_2128_ ),
    .A1(net1056),
    .S(net676),
    .X(\cs_registers_i/_0291_ ));
 sg13g2_nand3_1 \cs_registers_i/_4915_  (.B(\cs_registers_i/mhpmcounter_1869_ ),
    .C(net714),
    .A(\cs_registers_i/mhpmcounter_1870_ ),
    .Y(\cs_registers_i/_2129_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4916_  (.Y(\cs_registers_i/_2130_ ),
    .A(\cs_registers_i/mhpmcounter_1871_ ),
    .B(\cs_registers_i/_2129_ ));
 sg13g2_mux2_1 \cs_registers_i/_4917_  (.A0(\cs_registers_i/_2130_ ),
    .A1(net1069),
    .S(net676),
    .X(\cs_registers_i/_0292_ ));
 sg13g2_nand4_1 \cs_registers_i/_4918_  (.B(\cs_registers_i/mhpmcounter_1869_ ),
    .C(\cs_registers_i/mhpmcounter_1871_ ),
    .A(\cs_registers_i/mhpmcounter_1870_ ),
    .Y(\cs_registers_i/_2131_ ),
    .D(net714));
 sg13g2_xnor2_1 \cs_registers_i/_4919_  (.Y(\cs_registers_i/_2132_ ),
    .A(\cs_registers_i/mhpmcounter_1872_ ),
    .B(\cs_registers_i/_2131_ ));
 sg13g2_mux2_1 \cs_registers_i/_4920_  (.A0(\cs_registers_i/_2132_ ),
    .A1(\cs_registers_i/_0834_ ),
    .S(net676),
    .X(\cs_registers_i/_0293_ ));
 sg13g2_nand4_1 \cs_registers_i/_4921_  (.B(\cs_registers_i/mhpmcounter_1870_ ),
    .C(\cs_registers_i/mhpmcounter_1869_ ),
    .A(\cs_registers_i/mhpmcounter_1872_ ),
    .Y(\cs_registers_i/_2133_ ),
    .D(\cs_registers_i/mhpmcounter_1871_ ));
 sg13g2_nor4_2 \cs_registers_i/_4922_  (.A(net735),
    .B(\cs_registers_i/_2105_ ),
    .C(\cs_registers_i/_2124_ ),
    .Y(\cs_registers_i/_2134_ ),
    .D(\cs_registers_i/_2133_ ));
 sg13g2_xor2_1 \cs_registers_i/_4923_  (.B(\cs_registers_i/_2134_ ),
    .A(\cs_registers_i/mhpmcounter_1873_ ),
    .X(\cs_registers_i/_2135_ ));
 sg13g2_mux2_1 \cs_registers_i/_4924_  (.A0(\cs_registers_i/_2135_ ),
    .A1(net1053),
    .S(net677),
    .X(\cs_registers_i/_0294_ ));
 sg13g2_nand2_1 \cs_registers_i/_4925_  (.Y(\cs_registers_i/_2136_ ),
    .A(\cs_registers_i/mhpmcounter_1873_ ),
    .B(\cs_registers_i/_2134_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4926_  (.Y(\cs_registers_i/_2137_ ),
    .A(\cs_registers_i/mhpmcounter_1874_ ),
    .B(\cs_registers_i/_2136_ ));
 sg13g2_mux2_1 \cs_registers_i/_4927_  (.A0(net1052),
    .A1(\cs_registers_i/_2137_ ),
    .S(net717),
    .X(\cs_registers_i/_0295_ ));
 sg13g2_nand3_1 \cs_registers_i/_4928_  (.B(\cs_registers_i/mhpmcounter_1873_ ),
    .C(\cs_registers_i/_2134_ ),
    .A(\cs_registers_i/mhpmcounter_1874_ ),
    .Y(\cs_registers_i/_2138_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4929_  (.Y(\cs_registers_i/_2139_ ),
    .A(\cs_registers_i/mhpmcounter_1875_ ),
    .B(\cs_registers_i/_2138_ ));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net463));
 sg13g2_mux2_1 \cs_registers_i/_4931_  (.A0(\cs_registers_i/_2139_ ),
    .A1(net1050),
    .S(net678),
    .X(\cs_registers_i/_0296_ ));
 sg13g2_nand4_1 \cs_registers_i/_4932_  (.B(\cs_registers_i/mhpmcounter_1873_ ),
    .C(\cs_registers_i/mhpmcounter_1875_ ),
    .A(\cs_registers_i/mhpmcounter_1874_ ),
    .Y(\cs_registers_i/_2141_ ),
    .D(\cs_registers_i/_2134_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4933_  (.Y(\cs_registers_i/_2142_ ),
    .A(\cs_registers_i/mhpmcounter_1876_ ),
    .B(\cs_registers_i/_2141_ ));
 sg13g2_mux2_1 \cs_registers_i/_4934_  (.A0(\cs_registers_i/_2142_ ),
    .A1(net1049),
    .S(\cs_registers_i/_2110_ ),
    .X(\cs_registers_i/_0297_ ));
 sg13g2_nand4_1 \cs_registers_i/_4935_  (.B(\cs_registers_i/mhpmcounter_1874_ ),
    .C(\cs_registers_i/mhpmcounter_1873_ ),
    .A(\cs_registers_i/mhpmcounter_1876_ ),
    .Y(\cs_registers_i/_2143_ ),
    .D(\cs_registers_i/mhpmcounter_1875_ ));
 sg13g2_nor2_1 \cs_registers_i/_4936_  (.A(\cs_registers_i/_2133_ ),
    .B(\cs_registers_i/_2143_ ),
    .Y(\cs_registers_i/_2144_ ));
 sg13g2_nand2_2 \cs_registers_i/_4937_  (.Y(\cs_registers_i/_2145_ ),
    .A(net714),
    .B(\cs_registers_i/_2144_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4938_  (.Y(\cs_registers_i/_2146_ ),
    .A(\cs_registers_i/mhpmcounter_1877_ ),
    .B(\cs_registers_i/_2145_ ));
 sg13g2_mux2_1 \cs_registers_i/_4939_  (.A0(\cs_registers_i/_2146_ ),
    .A1(net1047),
    .S(net677),
    .X(\cs_registers_i/_0298_ ));
 sg13g2_nand3_1 \cs_registers_i/_4940_  (.B(net714),
    .C(\cs_registers_i/_2144_ ),
    .A(\cs_registers_i/mhpmcounter_1877_ ),
    .Y(\cs_registers_i/_2147_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4941_  (.Y(\cs_registers_i/_2148_ ),
    .A(\cs_registers_i/mhpmcounter_1878_ ),
    .B(\cs_registers_i/_2147_ ));
 sg13g2_mux2_1 \cs_registers_i/_4942_  (.A0(\cs_registers_i/_2148_ ),
    .A1(net1027),
    .S(net677),
    .X(\cs_registers_i/_0299_ ));
 sg13g2_nand4_1 \cs_registers_i/_4943_  (.B(\cs_registers_i/mhpmcounter_1877_ ),
    .C(net714),
    .A(\cs_registers_i/mhpmcounter_1878_ ),
    .Y(\cs_registers_i/_2149_ ),
    .D(\cs_registers_i/_2144_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4944_  (.Y(\cs_registers_i/_2150_ ),
    .A(\cs_registers_i/mhpmcounter_1879_ ),
    .B(\cs_registers_i/_2149_ ));
 sg13g2_mux2_1 \cs_registers_i/_4945_  (.A0(\cs_registers_i/_2150_ ),
    .A1(\cs_registers_i/_1031_ ),
    .S(net677),
    .X(\cs_registers_i/_0300_ ));
 sg13g2_and4_1 \cs_registers_i/_4946_  (.A(\cs_registers_i/mhpmcounter_1878_ ),
    .B(\cs_registers_i/mhpmcounter_1877_ ),
    .C(\cs_registers_i/mhpmcounter_1879_ ),
    .D(\cs_registers_i/_2144_ ),
    .X(\cs_registers_i/_2151_ ));
 sg13g2_nand2_2 \cs_registers_i/_4947_  (.Y(\cs_registers_i/_2152_ ),
    .A(net714),
    .B(\cs_registers_i/_2151_ ));
 sg13g2_xor2_1 \cs_registers_i/_4948_  (.B(\cs_registers_i/_2152_ ),
    .A(\cs_registers_i/mhpmcounter_1880_ ),
    .X(\cs_registers_i/_2153_ ));
 sg13g2_nor2_1 \cs_registers_i/_4949_  (.A(net1044),
    .B(net718),
    .Y(\cs_registers_i/_2154_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4950_  (.A1(net718),
    .A2(\cs_registers_i/_2153_ ),
    .Y(\cs_registers_i/_0301_ ),
    .B1(\cs_registers_i/_2154_ ));
 sg13g2_and3_1 \cs_registers_i/_4951_  (.X(\cs_registers_i/_2155_ ),
    .A(\cs_registers_i/mhpmcounter_1880_ ),
    .B(\cs_registers_i/_2125_ ),
    .C(\cs_registers_i/_2151_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4952_  (.Y(\cs_registers_i/_2156_ ),
    .A(\cs_registers_i/mhpmcounter_1881_ ),
    .B(\cs_registers_i/_2155_ ));
 sg13g2_nor2_1 \cs_registers_i/_4953_  (.A(net1043),
    .B(net718),
    .Y(\cs_registers_i/_2157_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4954_  (.A1(net718),
    .A2(\cs_registers_i/_2156_ ),
    .Y(\cs_registers_i/_0302_ ),
    .B1(\cs_registers_i/_2157_ ));
 sg13g2_inv_1 \cs_registers_i/_4955_  (.Y(\cs_registers_i/_2158_ ),
    .A(\cs_registers_i/mhpmcounter_1882_ ));
 sg13g2_nand2_1 \cs_registers_i/_4956_  (.Y(\cs_registers_i/_2159_ ),
    .A(\cs_registers_i/mhpmcounter_1880_ ),
    .B(\cs_registers_i/mhpmcounter_1881_ ));
 sg13g2_nor2_2 \cs_registers_i/_4957_  (.A(\cs_registers_i/_2152_ ),
    .B(\cs_registers_i/_2159_ ),
    .Y(\cs_registers_i/_2160_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4958_  (.Y(\cs_registers_i/_2161_ ),
    .A(\cs_registers_i/_2158_ ),
    .B(\cs_registers_i/_2160_ ));
 sg13g2_mux2_1 \cs_registers_i/_4959_  (.A0(net1066),
    .A1(\cs_registers_i/_2161_ ),
    .S(net717),
    .X(\cs_registers_i/_0303_ ));
 sg13g2_nor3_2 \cs_registers_i/_4960_  (.A(\cs_registers_i/_2158_ ),
    .B(\cs_registers_i/_2152_ ),
    .C(\cs_registers_i/_2159_ ),
    .Y(\cs_registers_i/_2162_ ));
 sg13g2_xor2_1 \cs_registers_i/_4961_  (.B(\cs_registers_i/_2162_ ),
    .A(\cs_registers_i/mhpmcounter_1883_ ),
    .X(\cs_registers_i/_2163_ ));
 sg13g2_mux2_1 \cs_registers_i/_4962_  (.A0(\cs_registers_i/_2163_ ),
    .A1(net1026),
    .S(net677),
    .X(\cs_registers_i/_0304_ ));
 sg13g2_inv_1 \cs_registers_i/_4963_  (.Y(\cs_registers_i/_2164_ ),
    .A(\cs_registers_i/_2151_ ));
 sg13g2_nand4_1 \cs_registers_i/_4964_  (.B(\cs_registers_i/mhpmcounter_1880_ ),
    .C(\cs_registers_i/mhpmcounter_1881_ ),
    .A(\cs_registers_i/mhpmcounter_1882_ ),
    .Y(\cs_registers_i/_2165_ ),
    .D(\cs_registers_i/mhpmcounter_1883_ ));
 sg13g2_nor4_2 \cs_registers_i/_4965_  (.A(\cs_registers_i/_2105_ ),
    .B(\cs_registers_i/_2124_ ),
    .C(\cs_registers_i/_2164_ ),
    .Y(\cs_registers_i/_2166_ ),
    .D(\cs_registers_i/_2165_ ));
 sg13g2_buf_4 fanout460 (.X(net460),
    .A(net463));
 sg13g2_nor2b_2 \cs_registers_i/_4967_  (.A(net735),
    .B_N(net713),
    .Y(\cs_registers_i/_2168_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4968_  (.Y(\cs_registers_i/_2169_ ),
    .A(\cs_registers_i/mhpmcounter_1884_ ),
    .B(\cs_registers_i/_2168_ ));
 sg13g2_nor2_1 \cs_registers_i/_4969_  (.A(net1042),
    .B(net717),
    .Y(\cs_registers_i/_2170_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4970_  (.A1(net717),
    .A2(\cs_registers_i/_2169_ ),
    .Y(\cs_registers_i/_0305_ ),
    .B1(\cs_registers_i/_2170_ ));
 sg13g2_nand2_2 \cs_registers_i/_4971_  (.Y(\cs_registers_i/_2171_ ),
    .A(\cs_registers_i/mhpmcounter_1884_ ),
    .B(\cs_registers_i/_2168_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4972_  (.Y(\cs_registers_i/_2172_ ),
    .A(\cs_registers_i/mhpmcounter_1885_ ),
    .B(\cs_registers_i/_2171_ ));
 sg13g2_mux2_1 \cs_registers_i/_4973_  (.A0(\cs_registers_i/_2172_ ),
    .A1(net1041),
    .S(net677),
    .X(\cs_registers_i/_0306_ ));
 sg13g2_and3_1 \cs_registers_i/_4974_  (.X(\cs_registers_i/_2173_ ),
    .A(\cs_registers_i/mhpmcounter_1884_ ),
    .B(\cs_registers_i/mhpmcounter_1885_ ),
    .C(\cs_registers_i/_2168_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4975_  (.Y(\cs_registers_i/_2174_ ),
    .A(\cs_registers_i/mhpmcounter_1886_ ),
    .B(\cs_registers_i/_2173_ ));
 sg13g2_nor2_1 \cs_registers_i/_4976_  (.A(net1037),
    .B(net717),
    .Y(\cs_registers_i/_2175_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4977_  (.A1(net717),
    .A2(\cs_registers_i/_2174_ ),
    .Y(\cs_registers_i/_0307_ ),
    .B1(\cs_registers_i/_2175_ ));
 sg13g2_and4_1 \cs_registers_i/_4978_  (.A(\cs_registers_i/mhpmcounter_1886_ ),
    .B(\cs_registers_i/mhpmcounter_1884_ ),
    .C(\cs_registers_i/mhpmcounter_1885_ ),
    .D(\cs_registers_i/_2168_ ),
    .X(\cs_registers_i/_2176_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4979_  (.Y(\cs_registers_i/_2177_ ),
    .A(\cs_registers_i/mhpmcounter_1887_ ),
    .B(\cs_registers_i/_2176_ ));
 sg13g2_nor2_1 \cs_registers_i/_4980_  (.A(net1036),
    .B(net717),
    .Y(\cs_registers_i/_2178_ ));
 sg13g2_a21oi_1 \cs_registers_i/_4981_  (.A1(net717),
    .A2(\cs_registers_i/_2177_ ),
    .Y(\cs_registers_i/_0308_ ),
    .B1(\cs_registers_i/_2178_ ));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net463));
 sg13g2_and4_2 \cs_registers_i/_4983_  (.A(\cs_registers_i/mhpmcounter_1886_ ),
    .B(\cs_registers_i/mhpmcounter_1884_ ),
    .C(\cs_registers_i/mhpmcounter_1885_ ),
    .D(\cs_registers_i/mhpmcounter_1887_ ),
    .X(\cs_registers_i/_2180_ ));
 sg13g2_nand2_2 \cs_registers_i/_4984_  (.Y(\cs_registers_i/_2181_ ),
    .A(net712),
    .B(\cs_registers_i/_2180_ ));
 sg13g2_xnor2_1 \cs_registers_i/_4985_  (.Y(\cs_registers_i/_2182_ ),
    .A(\cs_registers_i/mhpmcounter_1888_ ),
    .B(\cs_registers_i/_2181_ ));
 sg13g2_nor2_1 \cs_registers_i/_4986_  (.A(\cs_registers_i/_2063_ ),
    .B(\cs_registers_i/_2108_ ),
    .Y(\cs_registers_i/_2183_ ));
 sg13g2_nor2b_1 \cs_registers_i/_4987_  (.A(\cs_registers_i/_2183_ ),
    .B_N(net733),
    .Y(\cs_registers_i/_2184_ ));
 sg13g2_buf_4 fanout458 (.X(net458),
    .A(net463));
 sg13g2_and3_1 \cs_registers_i/_4989_  (.X(\cs_registers_i/_2186_ ),
    .A(\cs_registers_i/mhpmcounter_1888_ ),
    .B(net39),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_4990_  (.B2(\cs_registers_i/_1694_ ),
    .C1(\cs_registers_i/_2186_ ),
    .B1(net13),
    .A1(net716),
    .Y(\cs_registers_i/_2187_ ),
    .A2(\cs_registers_i/_2182_ ));
 sg13g2_inv_1 \cs_registers_i/_4991_  (.Y(\cs_registers_i/_0309_ ),
    .A(\cs_registers_i/_2187_ ));
 sg13g2_nor2_2 \cs_registers_i/_4992_  (.A(net38),
    .B(net716),
    .Y(\cs_registers_i/_2188_ ));
 sg13g2_nor2b_2 \cs_registers_i/_4993_  (.A(net22),
    .B_N(net712),
    .Y(\cs_registers_i/_2189_ ));
 sg13g2_nand3_1 \cs_registers_i/_4994_  (.B(\cs_registers_i/_2180_ ),
    .C(\cs_registers_i/_2189_ ),
    .A(\cs_registers_i/mhpmcounter_1888_ ),
    .Y(\cs_registers_i/_2190_ ));
 sg13g2_xor2_1 \cs_registers_i/_4995_  (.B(\cs_registers_i/_2190_ ),
    .A(\cs_registers_i/mhpmcounter_1889_ ),
    .X(\cs_registers_i/_2191_ ));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net463));
 sg13g2_nand2_1 \cs_registers_i/_4997_  (.Y(\cs_registers_i/_2193_ ),
    .A(net1067),
    .B(net11));
 sg13g2_o21ai_1 \cs_registers_i/_4998_  (.B1(\cs_registers_i/_2193_ ),
    .Y(\cs_registers_i/_0310_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2191_ ));
 sg13g2_and4_1 \cs_registers_i/_4999_  (.A(\cs_registers_i/mhpmcounter_1888_ ),
    .B(\cs_registers_i/mhpmcounter_1889_ ),
    .C(\cs_registers_i/_2180_ ),
    .D(\cs_registers_i/_2189_ ),
    .X(\cs_registers_i/_2194_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5000_  (.Y(\cs_registers_i/_2195_ ),
    .A(\cs_registers_i/mhpmcounter_1890_ ),
    .B(\cs_registers_i/_2194_ ));
 sg13g2_buf_4 fanout456 (.X(net456),
    .A(net463));
 sg13g2_nand2_1 \cs_registers_i/_5002_  (.Y(\cs_registers_i/_2197_ ),
    .A(net1038),
    .B(net15));
 sg13g2_o21ai_1 \cs_registers_i/_5003_  (.B1(\cs_registers_i/_2197_ ),
    .Y(\cs_registers_i/_0311_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2195_ ));
 sg13g2_nand2_1 \cs_registers_i/_5004_  (.Y(\cs_registers_i/_2198_ ),
    .A(net1033),
    .B(net11));
 sg13g2_nand4_1 \cs_registers_i/_5005_  (.B(\cs_registers_i/mhpmcounter_1890_ ),
    .C(\cs_registers_i/mhpmcounter_1889_ ),
    .A(\cs_registers_i/mhpmcounter_1888_ ),
    .Y(\cs_registers_i/_2199_ ),
    .D(\cs_registers_i/_2180_ ));
 sg13g2_inv_1 \cs_registers_i/_5006_  (.Y(\cs_registers_i/_2200_ ),
    .A(\cs_registers_i/_2199_ ));
 sg13g2_nand2_2 \cs_registers_i/_5007_  (.Y(\cs_registers_i/_2201_ ),
    .A(\cs_registers_i/_2189_ ),
    .B(\cs_registers_i/_2200_ ));
 sg13g2_or2_1 \cs_registers_i/_5008_  (.X(\cs_registers_i/_2202_ ),
    .B(\cs_registers_i/_2201_ ),
    .A(\cs_registers_i/mhpmcounter_1891_ ));
 sg13g2_nand2b_2 \cs_registers_i/_5009_  (.Y(\cs_registers_i/_2203_ ),
    .B(net19),
    .A_N(net38));
 sg13g2_nand3_1 \cs_registers_i/_5010_  (.B(\cs_registers_i/_2203_ ),
    .C(\cs_registers_i/_2201_ ),
    .A(\cs_registers_i/mhpmcounter_1891_ ),
    .Y(\cs_registers_i/_2204_ ));
 sg13g2_nand3_1 \cs_registers_i/_5011_  (.B(\cs_registers_i/_2202_ ),
    .C(\cs_registers_i/_2204_ ),
    .A(\cs_registers_i/_2198_ ),
    .Y(\cs_registers_i/_0312_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5012_  (.B1(net733),
    .Y(\cs_registers_i/_2205_ ),
    .A1(\cs_registers_i/_2063_ ),
    .A2(net20));
 sg13g2_nand3_1 \cs_registers_i/_5013_  (.B(net712),
    .C(\cs_registers_i/_2200_ ),
    .A(\cs_registers_i/mhpmcounter_1891_ ),
    .Y(\cs_registers_i/_2206_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5014_  (.Y(\cs_registers_i/_2207_ ),
    .A(\cs_registers_i/mhpmcounter_1892_ ),
    .B(\cs_registers_i/_2206_ ));
 sg13g2_a22oi_1 \cs_registers_i/_5015_  (.Y(\cs_registers_i/_2208_ ),
    .B1(\cs_registers_i/_2207_ ),
    .B2(net716),
    .A2(net678),
    .A1(\cs_registers_i/mhpmcounter_1892_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5016_  (.B1(\cs_registers_i/_2208_ ),
    .Y(\cs_registers_i/_0313_ ),
    .A1(\cs_registers_i/_2087_ ),
    .A2(\cs_registers_i/_2205_ ));
 sg13g2_nand2_1 \cs_registers_i/_5017_  (.Y(\cs_registers_i/_2209_ ),
    .A(\cs_registers_i/mhpmcounter_1892_ ),
    .B(\cs_registers_i/mhpmcounter_1891_ ));
 sg13g2_nor2_2 \cs_registers_i/_5018_  (.A(\cs_registers_i/_2199_ ),
    .B(\cs_registers_i/_2209_ ),
    .Y(\cs_registers_i/_2210_ ));
 sg13g2_nand3_1 \cs_registers_i/_5019_  (.B(net712),
    .C(\cs_registers_i/_2210_ ),
    .A(net716),
    .Y(\cs_registers_i/_2211_ ));
 sg13g2_a21oi_2 \cs_registers_i/_5020_  (.B1(net21),
    .Y(\cs_registers_i/_2212_ ),
    .A2(\cs_registers_i/_2210_ ),
    .A1(net712));
 sg13g2_o21ai_1 \cs_registers_i/_5021_  (.B1(\cs_registers_i/mhpmcounter_1893_ ),
    .Y(\cs_registers_i/_2213_ ),
    .A1(\cs_registers_i/_2088_ ),
    .A2(\cs_registers_i/_2212_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5022_  (.B1(\cs_registers_i/_2213_ ),
    .Y(\cs_registers_i/_2214_ ),
    .A1(\cs_registers_i/mhpmcounter_1893_ ),
    .A2(\cs_registers_i/_2211_ ));
 sg13g2_a21o_1 \cs_registers_i/_5023_  (.A2(net14),
    .A1(net1065),
    .B1(\cs_registers_i/_2214_ ),
    .X(\cs_registers_i/_0314_ ));
 sg13g2_nand3_1 \cs_registers_i/_5024_  (.B(\cs_registers_i/_2189_ ),
    .C(\cs_registers_i/_2210_ ),
    .A(\cs_registers_i/mhpmcounter_1893_ ),
    .Y(\cs_registers_i/_2215_ ));
 sg13g2_nand3_1 \cs_registers_i/_5025_  (.B(\cs_registers_i/_2203_ ),
    .C(\cs_registers_i/_2215_ ),
    .A(\cs_registers_i/mhpmcounter_1894_ ),
    .Y(\cs_registers_i/_2216_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5026_  (.B1(\cs_registers_i/_2216_ ),
    .Y(\cs_registers_i/_2217_ ),
    .A1(\cs_registers_i/mhpmcounter_1894_ ),
    .A2(\cs_registers_i/_2215_ ));
 sg13g2_a21o_1 \cs_registers_i/_5027_  (.A2(net14),
    .A1(net1064),
    .B1(\cs_registers_i/_2217_ ),
    .X(\cs_registers_i/_0315_ ));
 sg13g2_and4_1 \cs_registers_i/_5028_  (.A(\cs_registers_i/mhpmcounter_1894_ ),
    .B(\cs_registers_i/mhpmcounter_1893_ ),
    .C(net712),
    .D(\cs_registers_i/_2210_ ),
    .X(\cs_registers_i/_2218_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5029_  (.B1(net719),
    .Y(\cs_registers_i/_2219_ ),
    .A1(net20),
    .A2(\cs_registers_i/_2218_ ));
 sg13g2_nand4_1 \cs_registers_i/_5030_  (.B(\cs_registers_i/mhpmcounter_1893_ ),
    .C(net712),
    .A(\cs_registers_i/mhpmcounter_1894_ ),
    .Y(\cs_registers_i/_2220_ ),
    .D(\cs_registers_i/_2210_ ));
 sg13g2_nor3_1 \cs_registers_i/_5031_  (.A(\cs_registers_i/mhpmcounter_1895_ ),
    .B(net20),
    .C(\cs_registers_i/_2220_ ),
    .Y(\cs_registers_i/_2221_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5032_  (.B2(\cs_registers_i/mhpmcounter_1895_ ),
    .C1(\cs_registers_i/_2221_ ),
    .B1(\cs_registers_i/_2219_ ),
    .A1(net1031),
    .Y(\cs_registers_i/_2222_ ),
    .A2(net14));
 sg13g2_inv_1 \cs_registers_i/_5033_  (.Y(\cs_registers_i/_0316_ ),
    .A(\cs_registers_i/_2222_ ));
 sg13g2_nand2_2 \cs_registers_i/_5034_  (.Y(\cs_registers_i/_2223_ ),
    .A(\cs_registers_i/mhpmcounter_1895_ ),
    .B(\cs_registers_i/_2218_ ));
 sg13g2_xor2_1 \cs_registers_i/_5035_  (.B(\cs_registers_i/_2223_ ),
    .A(\cs_registers_i/mhpmcounter_1896_ ),
    .X(\cs_registers_i/_2224_ ));
 sg13g2_a21o_1 \cs_registers_i/_5036_  (.A2(net22),
    .A1(\cs_registers_i/mhpmcounter_1896_ ),
    .B1(net13),
    .X(\cs_registers_i/_2225_ ));
 sg13g2_a22oi_1 \cs_registers_i/_5037_  (.Y(\cs_registers_i/_2226_ ),
    .B1(\cs_registers_i/_2225_ ),
    .B2(net1025),
    .A2(net678),
    .A1(\cs_registers_i/mhpmcounter_1896_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5038_  (.B1(\cs_registers_i/_2226_ ),
    .Y(\cs_registers_i/_0317_ ),
    .A1(net20),
    .A2(\cs_registers_i/_2224_ ));
 sg13g2_nand3_1 \cs_registers_i/_5039_  (.B(\cs_registers_i/mhpmcounter_1895_ ),
    .C(\cs_registers_i/_2218_ ),
    .A(\cs_registers_i/mhpmcounter_1896_ ),
    .Y(\cs_registers_i/_2227_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5040_  (.Y(\cs_registers_i/_2228_ ),
    .A(\cs_registers_i/mhpmcounter_1897_ ),
    .B(\cs_registers_i/_2227_ ));
 sg13g2_and3_1 \cs_registers_i/_5041_  (.X(\cs_registers_i/_2229_ ),
    .A(\cs_registers_i/mhpmcounter_1897_ ),
    .B(net39),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_5042_  (.B2(net716),
    .C1(\cs_registers_i/_2229_ ),
    .B1(\cs_registers_i/_2228_ ),
    .A1(net1030),
    .Y(\cs_registers_i/_2230_ ),
    .A2(net14));
 sg13g2_inv_1 \cs_registers_i/_5043_  (.Y(\cs_registers_i/_0318_ ),
    .A(\cs_registers_i/_2230_ ));
 sg13g2_nand3_1 \cs_registers_i/_5044_  (.B(\cs_registers_i/mhpmcounter_1895_ ),
    .C(\cs_registers_i/mhpmcounter_1897_ ),
    .A(\cs_registers_i/mhpmcounter_1896_ ),
    .Y(\cs_registers_i/_2231_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5045_  (.B1(net716),
    .Y(\cs_registers_i/_2232_ ),
    .A1(\cs_registers_i/_2220_ ),
    .A2(\cs_registers_i/_2231_ ));
 sg13g2_nand2_1 \cs_registers_i/_5046_  (.Y(\cs_registers_i/_2233_ ),
    .A(net719),
    .B(\cs_registers_i/_2232_ ));
 sg13g2_nor4_1 \cs_registers_i/_5047_  (.A(\cs_registers_i/mhpmcounter_1898_ ),
    .B(net20),
    .C(\cs_registers_i/_2220_ ),
    .D(\cs_registers_i/_2231_ ),
    .Y(\cs_registers_i/_2234_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5048_  (.B2(\cs_registers_i/mhpmcounter_1898_ ),
    .C1(\cs_registers_i/_2234_ ),
    .B1(\cs_registers_i/_2233_ ),
    .A1(net1059),
    .Y(\cs_registers_i/_2235_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5049_  (.Y(\cs_registers_i/_0319_ ),
    .A(\cs_registers_i/_2235_ ));
 sg13g2_nand3_1 \cs_registers_i/_5050_  (.B(\cs_registers_i/mhpmcounter_1894_ ),
    .C(\cs_registers_i/mhpmcounter_1893_ ),
    .A(\cs_registers_i/mhpmcounter_1898_ ),
    .Y(\cs_registers_i/_2236_ ));
 sg13g2_or4_1 \cs_registers_i/_5051_  (.A(\cs_registers_i/_2199_ ),
    .B(\cs_registers_i/_2209_ ),
    .C(\cs_registers_i/_2231_ ),
    .D(\cs_registers_i/_2236_ ),
    .X(\cs_registers_i/_2237_ ));
 sg13g2_inv_1 \cs_registers_i/_5052_  (.Y(\cs_registers_i/_2238_ ),
    .A(\cs_registers_i/_2237_ ));
 sg13g2_nand2_2 \cs_registers_i/_5053_  (.Y(\cs_registers_i/_2239_ ),
    .A(net713),
    .B(\cs_registers_i/_2238_ ));
 sg13g2_nand2b_2 \cs_registers_i/_5054_  (.Y(\cs_registers_i/_2240_ ),
    .B(net715),
    .A_N(\cs_registers_i/_2239_ ));
 sg13g2_a21oi_1 \cs_registers_i/_5055_  (.A1(net713),
    .A2(\cs_registers_i/_2238_ ),
    .Y(\cs_registers_i/_2241_ ),
    .B1(net19));
 sg13g2_o21ai_1 \cs_registers_i/_5056_  (.B1(\cs_registers_i/mhpmcounter_1899_ ),
    .Y(\cs_registers_i/_2242_ ),
    .A1(net678),
    .A2(\cs_registers_i/_2241_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5057_  (.B1(\cs_registers_i/_2242_ ),
    .Y(\cs_registers_i/_2243_ ),
    .A1(\cs_registers_i/mhpmcounter_1899_ ),
    .A2(\cs_registers_i/_2240_ ));
 sg13g2_a21o_1 \cs_registers_i/_5058_  (.A2(net14),
    .A1(net1071),
    .B1(\cs_registers_i/_2243_ ),
    .X(\cs_registers_i/_0320_ ));
 sg13g2_inv_1 \cs_registers_i/_5059_  (.Y(\cs_registers_i/_2244_ ),
    .A(\cs_registers_i/mhpmcounter_1899_ ));
 sg13g2_nor2_2 \cs_registers_i/_5060_  (.A(\cs_registers_i/_2244_ ),
    .B(\cs_registers_i/_2240_ ),
    .Y(\cs_registers_i/_2245_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5061_  (.Y(\cs_registers_i/_2246_ ),
    .A(\cs_registers_i/mhpmcounter_1900_ ),
    .B(\cs_registers_i/_2245_ ));
 sg13g2_nand2_1 \cs_registers_i/_5062_  (.Y(\cs_registers_i/_2247_ ),
    .A(net1028),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5063_  (.B1(\cs_registers_i/_2247_ ),
    .Y(\cs_registers_i/_0321_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2246_ ));
 sg13g2_nand2_1 \cs_registers_i/_5064_  (.Y(\cs_registers_i/_2248_ ),
    .A(\cs_registers_i/mhpmcounter_1900_ ),
    .B(\cs_registers_i/mhpmcounter_1899_ ));
 sg13g2_nor2_2 \cs_registers_i/_5065_  (.A(\cs_registers_i/_2239_ ),
    .B(\cs_registers_i/_2248_ ),
    .Y(\cs_registers_i/_2249_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5066_  (.Y(\cs_registers_i/_2250_ ),
    .A(\cs_registers_i/mhpmcounter_1901_ ),
    .B(\cs_registers_i/_2249_ ));
 sg13g2_a22oi_1 \cs_registers_i/_5067_  (.Y(\cs_registers_i/_2251_ ),
    .B1(net12),
    .B2(net1058),
    .A2(net678),
    .A1(\cs_registers_i/mhpmcounter_1901_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5068_  (.B1(\cs_registers_i/_2251_ ),
    .Y(\cs_registers_i/_0322_ ),
    .A1(net19),
    .A2(\cs_registers_i/_2250_ ));
 sg13g2_inv_1 \cs_registers_i/_5069_  (.Y(\cs_registers_i/_2252_ ),
    .A(\cs_registers_i/mhpmcounter_1901_ ));
 sg13g2_nor3_2 \cs_registers_i/_5070_  (.A(\cs_registers_i/_2252_ ),
    .B(\cs_registers_i/_2239_ ),
    .C(\cs_registers_i/_2248_ ),
    .Y(\cs_registers_i/_2253_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5071_  (.Y(\cs_registers_i/_2254_ ),
    .A(\cs_registers_i/mhpmcounter_1902_ ),
    .B(\cs_registers_i/_2253_ ));
 sg13g2_a22oi_1 \cs_registers_i/_5072_  (.Y(\cs_registers_i/_2255_ ),
    .B1(net11),
    .B2(net1056),
    .A2(net678),
    .A1(\cs_registers_i/mhpmcounter_1902_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5073_  (.B1(\cs_registers_i/_2255_ ),
    .Y(\cs_registers_i/_0323_ ),
    .A1(net19),
    .A2(\cs_registers_i/_2254_ ));
 sg13g2_nand4_1 \cs_registers_i/_5074_  (.B(\cs_registers_i/mhpmcounter_1900_ ),
    .C(\cs_registers_i/mhpmcounter_1899_ ),
    .A(\cs_registers_i/mhpmcounter_1902_ ),
    .Y(\cs_registers_i/_2256_ ),
    .D(\cs_registers_i/mhpmcounter_1901_ ));
 sg13g2_nor2_2 \cs_registers_i/_5075_  (.A(\cs_registers_i/_2240_ ),
    .B(\cs_registers_i/_2256_ ),
    .Y(\cs_registers_i/_2257_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5076_  (.Y(\cs_registers_i/_2258_ ),
    .A(\cs_registers_i/mhpmcounter_1903_ ),
    .B(\cs_registers_i/_2257_ ));
 sg13g2_nand2_1 \cs_registers_i/_5077_  (.Y(\cs_registers_i/_2259_ ),
    .A(net1069),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5078_  (.B1(\cs_registers_i/_2259_ ),
    .Y(\cs_registers_i/_0324_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2258_ ));
 sg13g2_inv_1 \cs_registers_i/_5079_  (.Y(\cs_registers_i/_2260_ ),
    .A(\cs_registers_i/mhpmcounter_1903_ ));
 sg13g2_nor3_2 \cs_registers_i/_5080_  (.A(\cs_registers_i/_2260_ ),
    .B(\cs_registers_i/_2237_ ),
    .C(\cs_registers_i/_2256_ ),
    .Y(\cs_registers_i/_2261_ ));
 sg13g2_and2_2 \cs_registers_i/_5081_  (.A(\cs_registers_i/_2189_ ),
    .B(\cs_registers_i/_2261_ ),
    .X(\cs_registers_i/_2262_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5082_  (.Y(\cs_registers_i/_2263_ ),
    .A(\cs_registers_i/mhpmcounter_1904_ ),
    .B(\cs_registers_i/_2262_ ));
 sg13g2_nand2_1 \cs_registers_i/_5083_  (.Y(\cs_registers_i/_2264_ ),
    .A(net1055),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5084_  (.B1(\cs_registers_i/_2264_ ),
    .Y(\cs_registers_i/_0325_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2263_ ));
 sg13g2_nand2_1 \cs_registers_i/_5085_  (.Y(\cs_registers_i/_2265_ ),
    .A(net1053),
    .B(net11));
 sg13g2_nand2_2 \cs_registers_i/_5086_  (.Y(\cs_registers_i/_2266_ ),
    .A(\cs_registers_i/mhpmcounter_1904_ ),
    .B(\cs_registers_i/_2262_ ));
 sg13g2_or2_1 \cs_registers_i/_5087_  (.X(\cs_registers_i/_2267_ ),
    .B(\cs_registers_i/_2266_ ),
    .A(\cs_registers_i/mhpmcounter_1905_ ));
 sg13g2_nand3_1 \cs_registers_i/_5088_  (.B(\cs_registers_i/_2203_ ),
    .C(\cs_registers_i/_2266_ ),
    .A(\cs_registers_i/mhpmcounter_1905_ ),
    .Y(\cs_registers_i/_2268_ ));
 sg13g2_nand3_1 \cs_registers_i/_5089_  (.B(\cs_registers_i/_2267_ ),
    .C(\cs_registers_i/_2268_ ),
    .A(\cs_registers_i/_2265_ ),
    .Y(\cs_registers_i/_0326_ ));
 sg13g2_nand4_1 \cs_registers_i/_5090_  (.B(\cs_registers_i/mhpmcounter_1905_ ),
    .C(net713),
    .A(\cs_registers_i/mhpmcounter_1904_ ),
    .Y(\cs_registers_i/_2269_ ),
    .D(\cs_registers_i/_2261_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5091_  (.Y(\cs_registers_i/_2270_ ),
    .A(\cs_registers_i/mhpmcounter_1906_ ),
    .B(\cs_registers_i/_2269_ ));
 sg13g2_and3_1 \cs_registers_i/_5092_  (.X(\cs_registers_i/_2271_ ),
    .A(\cs_registers_i/mhpmcounter_1906_ ),
    .B(net39),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_5093_  (.B2(net715),
    .C1(\cs_registers_i/_2271_ ),
    .B1(\cs_registers_i/_2270_ ),
    .A1(net1052),
    .Y(\cs_registers_i/_2272_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5094_  (.Y(\cs_registers_i/_0327_ ),
    .A(\cs_registers_i/_2272_ ));
 sg13g2_and4_1 \cs_registers_i/_5095_  (.A(\cs_registers_i/mhpmcounter_1906_ ),
    .B(\cs_registers_i/mhpmcounter_1904_ ),
    .C(\cs_registers_i/mhpmcounter_1905_ ),
    .D(\cs_registers_i/_2262_ ),
    .X(\cs_registers_i/_2273_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5096_  (.Y(\cs_registers_i/_2274_ ),
    .A(\cs_registers_i/mhpmcounter_1907_ ),
    .B(\cs_registers_i/_2273_ ));
 sg13g2_nand2_1 \cs_registers_i/_5097_  (.Y(\cs_registers_i/_2275_ ),
    .A(net1050),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5098_  (.B1(\cs_registers_i/_2275_ ),
    .Y(\cs_registers_i/_0328_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2274_ ));
 sg13g2_and4_1 \cs_registers_i/_5099_  (.A(\cs_registers_i/mhpmcounter_1906_ ),
    .B(\cs_registers_i/mhpmcounter_1904_ ),
    .C(\cs_registers_i/mhpmcounter_1905_ ),
    .D(\cs_registers_i/mhpmcounter_1907_ ),
    .X(\cs_registers_i/_2276_ ));
 sg13g2_nand2_2 \cs_registers_i/_5100_  (.Y(\cs_registers_i/_2277_ ),
    .A(\cs_registers_i/_2262_ ),
    .B(\cs_registers_i/_2276_ ));
 sg13g2_xor2_1 \cs_registers_i/_5101_  (.B(\cs_registers_i/_2277_ ),
    .A(\cs_registers_i/mhpmcounter_1908_ ),
    .X(\cs_registers_i/_2278_ ));
 sg13g2_nand2_1 \cs_registers_i/_5102_  (.Y(\cs_registers_i/_2279_ ),
    .A(net1049),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5103_  (.B1(\cs_registers_i/_2279_ ),
    .Y(\cs_registers_i/_0329_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2278_ ));
 sg13g2_nand3_1 \cs_registers_i/_5104_  (.B(\cs_registers_i/_2262_ ),
    .C(\cs_registers_i/_2276_ ),
    .A(\cs_registers_i/mhpmcounter_1908_ ),
    .Y(\cs_registers_i/_2280_ ));
 sg13g2_xor2_1 \cs_registers_i/_5105_  (.B(\cs_registers_i/_2280_ ),
    .A(\cs_registers_i/mhpmcounter_1909_ ),
    .X(\cs_registers_i/_2281_ ));
 sg13g2_nand2_1 \cs_registers_i/_5106_  (.Y(\cs_registers_i/_2282_ ),
    .A(net1047),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5107_  (.B1(\cs_registers_i/_2282_ ),
    .Y(\cs_registers_i/_0330_ ),
    .A1(net625),
    .A2(\cs_registers_i/_2281_ ));
 sg13g2_and3_1 \cs_registers_i/_5108_  (.X(\cs_registers_i/_2283_ ),
    .A(\cs_registers_i/mhpmcounter_1908_ ),
    .B(\cs_registers_i/mhpmcounter_1909_ ),
    .C(\cs_registers_i/_2276_ ));
 sg13g2_nand2_2 \cs_registers_i/_5109_  (.Y(\cs_registers_i/_2284_ ),
    .A(\cs_registers_i/_2262_ ),
    .B(\cs_registers_i/_2283_ ));
 sg13g2_xor2_1 \cs_registers_i/_5110_  (.B(\cs_registers_i/_2284_ ),
    .A(\cs_registers_i/mhpmcounter_1910_ ),
    .X(\cs_registers_i/_2285_ ));
 sg13g2_nand2_1 \cs_registers_i/_5111_  (.Y(\cs_registers_i/_2286_ ),
    .A(net1027),
    .B(net12));
 sg13g2_o21ai_1 \cs_registers_i/_5112_  (.B1(\cs_registers_i/_2286_ ),
    .Y(\cs_registers_i/_0331_ ),
    .A1(\cs_registers_i/_2188_ ),
    .A2(\cs_registers_i/_2285_ ));
 sg13g2_nand4_1 \cs_registers_i/_5113_  (.B(net712),
    .C(\cs_registers_i/_2261_ ),
    .A(\cs_registers_i/mhpmcounter_1910_ ),
    .Y(\cs_registers_i/_2287_ ),
    .D(\cs_registers_i/_2283_ ));
 sg13g2_a21o_1 \cs_registers_i/_5114_  (.A2(net2495),
    .A1(net715),
    .B1(net678),
    .X(\cs_registers_i/_2288_ ));
 sg13g2_nor3_1 \cs_registers_i/_5115_  (.A(\cs_registers_i/mhpmcounter_1911_ ),
    .B(net20),
    .C(net2495),
    .Y(\cs_registers_i/_2289_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5116_  (.B2(\cs_registers_i/mhpmcounter_1911_ ),
    .C1(\cs_registers_i/_2289_ ),
    .B1(\cs_registers_i/_2288_ ),
    .A1(\cs_registers_i/_1031_ ),
    .Y(\cs_registers_i/_2290_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5117_  (.Y(\cs_registers_i/_0332_ ),
    .A(\cs_registers_i/_2290_ ));
 sg13g2_nand2_1 \cs_registers_i/_5118_  (.Y(\cs_registers_i/_2291_ ),
    .A(net1044),
    .B(net11));
 sg13g2_nand2_1 \cs_registers_i/_5119_  (.Y(\cs_registers_i/_2292_ ),
    .A(\cs_registers_i/mhpmcounter_1912_ ),
    .B(\cs_registers_i/_2203_ ));
 sg13g2_nor2_2 \cs_registers_i/_5120_  (.A(net19),
    .B(\cs_registers_i/_2287_ ),
    .Y(\cs_registers_i/_2293_ ));
 sg13g2_nand2_2 \cs_registers_i/_5121_  (.Y(\cs_registers_i/_2294_ ),
    .A(\cs_registers_i/mhpmcounter_1911_ ),
    .B(\cs_registers_i/_2293_ ));
 sg13g2_mux2_1 \cs_registers_i/_5122_  (.A0(\cs_registers_i/mhpmcounter_1912_ ),
    .A1(\cs_registers_i/_2292_ ),
    .S(\cs_registers_i/_2294_ ),
    .X(\cs_registers_i/_2295_ ));
 sg13g2_nand2_1 \cs_registers_i/_5123_  (.Y(\cs_registers_i/_0333_ ),
    .A(\cs_registers_i/_2291_ ),
    .B(\cs_registers_i/_2295_ ));
 sg13g2_nand2_1 \cs_registers_i/_5124_  (.Y(\cs_registers_i/_2296_ ),
    .A(\cs_registers_i/mhpmcounter_1912_ ),
    .B(\cs_registers_i/mhpmcounter_1911_ ));
 sg13g2_nor2_2 \cs_registers_i/_5125_  (.A(net2495),
    .B(\cs_registers_i/_2296_ ),
    .Y(\cs_registers_i/_2297_ ));
 sg13g2_xor2_1 \cs_registers_i/_5126_  (.B(\cs_registers_i/_2297_ ),
    .A(\cs_registers_i/mhpmcounter_1913_ ),
    .X(\cs_registers_i/_2298_ ));
 sg13g2_and3_1 \cs_registers_i/_5127_  (.X(\cs_registers_i/_2299_ ),
    .A(\cs_registers_i/mhpmcounter_1913_ ),
    .B(net39),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_5128_  (.B2(net715),
    .C1(\cs_registers_i/_2299_ ),
    .B1(\cs_registers_i/_2298_ ),
    .A1(net1043),
    .Y(\cs_registers_i/_2300_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5129_  (.Y(\cs_registers_i/_0334_ ),
    .A(\cs_registers_i/_2300_ ));
 sg13g2_inv_1 \cs_registers_i/_5130_  (.Y(\cs_registers_i/_2301_ ),
    .A(\cs_registers_i/mhpmcounter_1914_ ));
 sg13g2_nand3_1 \cs_registers_i/_5131_  (.B(\cs_registers_i/mhpmcounter_1911_ ),
    .C(\cs_registers_i/mhpmcounter_1913_ ),
    .A(\cs_registers_i/mhpmcounter_1912_ ),
    .Y(\cs_registers_i/_2302_ ));
 sg13g2_nor2_2 \cs_registers_i/_5132_  (.A(net2495),
    .B(\cs_registers_i/_2302_ ),
    .Y(\cs_registers_i/_2303_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5133_  (.Y(\cs_registers_i/_2304_ ),
    .A(\cs_registers_i/_2301_ ),
    .B(\cs_registers_i/_2303_ ));
 sg13g2_and3_1 \cs_registers_i/_5134_  (.X(\cs_registers_i/_2305_ ),
    .A(\cs_registers_i/mhpmcounter_1914_ ),
    .B(net39),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_5135_  (.B2(net715),
    .C1(\cs_registers_i/_2305_ ),
    .B1(\cs_registers_i/_2304_ ),
    .A1(net1066),
    .Y(\cs_registers_i/_2306_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5136_  (.Y(\cs_registers_i/_0335_ ),
    .A(\cs_registers_i/_2306_ ));
 sg13g2_nor2_1 \cs_registers_i/_5137_  (.A(\cs_registers_i/_2301_ ),
    .B(\cs_registers_i/_2302_ ),
    .Y(\cs_registers_i/_2307_ ));
 sg13g2_nand2_2 \cs_registers_i/_5138_  (.Y(\cs_registers_i/_2308_ ),
    .A(\cs_registers_i/_2293_ ),
    .B(\cs_registers_i/_2307_ ));
 sg13g2_xor2_1 \cs_registers_i/_5139_  (.B(\cs_registers_i/_2308_ ),
    .A(\cs_registers_i/mhpmcounter_1915_ ),
    .X(\cs_registers_i/_2309_ ));
 sg13g2_nand2_1 \cs_registers_i/_5140_  (.Y(\cs_registers_i/_2310_ ),
    .A(net1026),
    .B(net11));
 sg13g2_o21ai_1 \cs_registers_i/_5141_  (.B1(\cs_registers_i/_2310_ ),
    .Y(\cs_registers_i/_0336_ ),
    .A1(\cs_registers_i/_2188_ ),
    .A2(\cs_registers_i/_2309_ ));
 sg13g2_nand2_1 \cs_registers_i/_5142_  (.Y(\cs_registers_i/_2311_ ),
    .A(\cs_registers_i/mhpmcounter_1915_ ),
    .B(\cs_registers_i/_2307_ ));
 sg13g2_nor2_2 \cs_registers_i/_5143_  (.A(net2495),
    .B(\cs_registers_i/_2311_ ),
    .Y(\cs_registers_i/_2312_ ));
 sg13g2_xor2_1 \cs_registers_i/_5144_  (.B(\cs_registers_i/_2312_ ),
    .A(\cs_registers_i/mhpmcounter_1916_ ),
    .X(\cs_registers_i/_2313_ ));
 sg13g2_and3_1 \cs_registers_i/_5145_  (.X(\cs_registers_i/_2314_ ),
    .A(\cs_registers_i/mhpmcounter_1916_ ),
    .B(net38),
    .C(net23));
 sg13g2_a221oi_1 \cs_registers_i/_5146_  (.B2(net715),
    .C1(\cs_registers_i/_2314_ ),
    .B1(\cs_registers_i/_2313_ ),
    .A1(net1042),
    .Y(\cs_registers_i/_2315_ ),
    .A2(net13));
 sg13g2_inv_1 \cs_registers_i/_5147_  (.Y(\cs_registers_i/_0337_ ),
    .A(\cs_registers_i/_2315_ ));
 sg13g2_nand3_1 \cs_registers_i/_5148_  (.B(\cs_registers_i/mhpmcounter_1915_ ),
    .C(\cs_registers_i/_2307_ ),
    .A(\cs_registers_i/mhpmcounter_1916_ ),
    .Y(\cs_registers_i/_2316_ ));
 sg13g2_nor2_2 \cs_registers_i/_5149_  (.A(net2495),
    .B(\cs_registers_i/_2316_ ),
    .Y(\cs_registers_i/_2317_ ));
 sg13g2_xnor2_1 \cs_registers_i/_5150_  (.Y(\cs_registers_i/_2318_ ),
    .A(\cs_registers_i/mhpmcounter_1917_ ),
    .B(\cs_registers_i/_2317_ ));
 sg13g2_nand3_1 \cs_registers_i/_5151_  (.B(net38),
    .C(net21),
    .A(\cs_registers_i/mhpmcounter_1917_ ),
    .Y(\cs_registers_i/_2319_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5152_  (.B1(\cs_registers_i/_2319_ ),
    .Y(\cs_registers_i/_2320_ ),
    .A1(net19),
    .A2(\cs_registers_i/_2318_ ));
 sg13g2_a21o_1 \cs_registers_i/_5153_  (.A2(net14),
    .A1(net1040),
    .B1(\cs_registers_i/_2320_ ),
    .X(\cs_registers_i/_0338_ ));
 sg13g2_nand2_1 \cs_registers_i/_5154_  (.Y(\cs_registers_i/_2321_ ),
    .A(net1037),
    .B(net11));
 sg13g2_o21ai_1 \cs_registers_i/_5155_  (.B1(\cs_registers_i/mhpmcounter_1918_ ),
    .Y(\cs_registers_i/_2322_ ),
    .A1(\cs_registers_i/_2061_ ),
    .A2(net715));
 sg13g2_inv_1 \cs_registers_i/_5156_  (.Y(\cs_registers_i/_2323_ ),
    .A(\cs_registers_i/_2316_ ));
 sg13g2_and3_1 \cs_registers_i/_5157_  (.X(\cs_registers_i/_2324_ ),
    .A(\cs_registers_i/mhpmcounter_1917_ ),
    .B(\cs_registers_i/_2293_ ),
    .C(\cs_registers_i/_2323_ ));
 sg13g2_mux2_1 \cs_registers_i/_5158_  (.A0(\cs_registers_i/_2322_ ),
    .A1(\cs_registers_i/mhpmcounter_1918_ ),
    .S(\cs_registers_i/_2324_ ),
    .X(\cs_registers_i/_2325_ ));
 sg13g2_nand2_1 \cs_registers_i/_5159_  (.Y(\cs_registers_i/_0339_ ),
    .A(\cs_registers_i/_2321_ ),
    .B(\cs_registers_i/_2325_ ));
 sg13g2_nand2_1 \cs_registers_i/_5160_  (.Y(\cs_registers_i/_2326_ ),
    .A(net1035),
    .B(net11));
 sg13g2_nand2_1 \cs_registers_i/_5161_  (.Y(\cs_registers_i/_2327_ ),
    .A(\cs_registers_i/mhpmcounter_1919_ ),
    .B(\cs_registers_i/_2203_ ));
 sg13g2_nand4_1 \cs_registers_i/_5162_  (.B(\cs_registers_i/mhpmcounter_1918_ ),
    .C(\cs_registers_i/_2293_ ),
    .A(\cs_registers_i/mhpmcounter_1917_ ),
    .Y(\cs_registers_i/_2328_ ),
    .D(\cs_registers_i/_2323_ ));
 sg13g2_mux2_1 \cs_registers_i/_5163_  (.A0(\cs_registers_i/mhpmcounter_1919_ ),
    .A1(\cs_registers_i/_2327_ ),
    .S(\cs_registers_i/_2328_ ),
    .X(\cs_registers_i/_2329_ ));
 sg13g2_nand2_1 \cs_registers_i/_5164_  (.Y(\cs_registers_i/_0340_ ),
    .A(\cs_registers_i/_2326_ ),
    .B(\cs_registers_i/_2329_ ));
 sg13g2_nand3_1 \cs_registers_i/_5165_  (.B(net722),
    .C(\cs_registers_i/_0599_ ),
    .A(net40),
    .Y(\cs_registers_i/_2330_ ));
 sg13g2_buf_4 fanout455 (.X(net455),
    .A(net463));
 sg13g2_buf_2 fanout454 (.A(\id_stage_i.controller_i.instr_i_21_ ),
    .X(net454));
 sg13g2_mux2_1 \cs_registers_i/_5168_  (.A0(net1055),
    .A1(\cs_registers_i/mie_q_0_ ),
    .S(net622),
    .X(\cs_registers_i/_0341_ ));
 sg13g2_mux2_1 \cs_registers_i/_5169_  (.A0(net1066),
    .A1(\cs_registers_i/mie_q_10_ ),
    .S(net621),
    .X(\cs_registers_i/_0342_ ));
 sg13g2_mux2_1 \cs_registers_i/_5170_  (.A0(net1026),
    .A1(\cs_registers_i/mie_q_11_ ),
    .S(net623),
    .X(\cs_registers_i/_0343_ ));
 sg13g2_mux2_1 \cs_registers_i/_5171_  (.A0(net1042),
    .A1(\cs_registers_i/mie_q_12_ ),
    .S(net622),
    .X(\cs_registers_i/_0344_ ));
 sg13g2_mux2_1 \cs_registers_i/_5172_  (.A0(net1040),
    .A1(\cs_registers_i/mie_q_13_ ),
    .S(net622),
    .X(\cs_registers_i/_0345_ ));
 sg13g2_mux2_1 \cs_registers_i/_5173_  (.A0(net1037),
    .A1(\cs_registers_i/mie_q_14_ ),
    .S(net624),
    .X(\cs_registers_i/_0346_ ));
 sg13g2_mux2_1 \cs_registers_i/_5174_  (.A0(net1035),
    .A1(\cs_registers_i/mie_q_15_ ),
    .S(net622),
    .X(\cs_registers_i/_0347_ ));
 sg13g2_mux2_1 \cs_registers_i/_5175_  (.A0(net1070),
    .A1(\cs_registers_i/mie_q_16_ ),
    .S(net624),
    .X(\cs_registers_i/_0348_ ));
 sg13g2_mux2_1 \cs_registers_i/_5176_  (.A0(net1031),
    .A1(\cs_registers_i/mie_q_17_ ),
    .S(net624),
    .X(\cs_registers_i/_0349_ ));
 sg13g2_mux2_1 \cs_registers_i/_5177_  (.A0(net1033),
    .A1(\cs_registers_i/mie_q_18_ ),
    .S(net624),
    .X(\cs_registers_i/_0350_ ));
 sg13g2_mux2_1 \cs_registers_i/_5178_  (.A0(net1053),
    .A1(\cs_registers_i/mie_q_1_ ),
    .S(net621),
    .X(\cs_registers_i/_0351_ ));
 sg13g2_mux2_1 \cs_registers_i/_5179_  (.A0(net1051),
    .A1(\cs_registers_i/mie_q_2_ ),
    .S(net621),
    .X(\cs_registers_i/_0352_ ));
 sg13g2_mux2_1 \cs_registers_i/_5180_  (.A0(net1050),
    .A1(\cs_registers_i/mie_q_3_ ),
    .S(net621),
    .X(\cs_registers_i/_0353_ ));
 sg13g2_mux2_1 \cs_registers_i/_5181_  (.A0(net1049),
    .A1(\cs_registers_i/mie_q_4_ ),
    .S(net623),
    .X(\cs_registers_i/_0354_ ));
 sg13g2_mux2_1 \cs_registers_i/_5182_  (.A0(net1047),
    .A1(\cs_registers_i/mie_q_5_ ),
    .S(net621),
    .X(\cs_registers_i/_0355_ ));
 sg13g2_mux2_1 \cs_registers_i/_5183_  (.A0(net1027),
    .A1(\cs_registers_i/mie_q_6_ ),
    .S(net623),
    .X(\cs_registers_i/_0356_ ));
 sg13g2_mux2_1 \cs_registers_i/_5184_  (.A0(net1046),
    .A1(\cs_registers_i/mie_q_7_ ),
    .S(net621),
    .X(\cs_registers_i/_0357_ ));
 sg13g2_mux2_1 \cs_registers_i/_5185_  (.A0(net1044),
    .A1(\cs_registers_i/mie_q_8_ ),
    .S(net621),
    .X(\cs_registers_i/_0358_ ));
 sg13g2_mux2_1 \cs_registers_i/_5186_  (.A0(net1043),
    .A1(\cs_registers_i/mie_q_9_ ),
    .S(net621),
    .X(\cs_registers_i/_0359_ ));
 sg13g2_nand3_1 \cs_registers_i/_5187_  (.B(net722),
    .C(net1149),
    .A(net1117),
    .Y(\cs_registers_i/_2333_ ));
 sg13g2_buf_4 fanout453 (.X(net453),
    .A(\id_stage_i.controller_i.instr_i_21_ ));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net453));
 sg13g2_mux2_1 \cs_registers_i/_5190_  (.A0(net1063),
    .A1(\cs_registers_i/mscratch_q_0_ ),
    .S(net617),
    .X(\cs_registers_i/_0360_ ));
 sg13g2_mux2_1 \cs_registers_i/_5191_  (.A0(net1059),
    .A1(\cs_registers_i/mscratch_q_10_ ),
    .S(net619),
    .X(\cs_registers_i/_0361_ ));
 sg13g2_mux2_1 \cs_registers_i/_5192_  (.A0(net1070),
    .A1(\cs_registers_i/mscratch_q_11_ ),
    .S(net616),
    .X(\cs_registers_i/_0362_ ));
 sg13g2_mux2_1 \cs_registers_i/_5193_  (.A0(net1028),
    .A1(\cs_registers_i/mscratch_q_12_ ),
    .S(net618),
    .X(\cs_registers_i/_0363_ ));
 sg13g2_mux2_1 \cs_registers_i/_5194_  (.A0(net1058),
    .A1(\cs_registers_i/mscratch_q_13_ ),
    .S(net616),
    .X(\cs_registers_i/_0364_ ));
 sg13g2_mux2_1 \cs_registers_i/_5195_  (.A0(net1056),
    .A1(\cs_registers_i/mscratch_q_14_ ),
    .S(net617),
    .X(\cs_registers_i/_0365_ ));
 sg13g2_mux2_1 \cs_registers_i/_5196_  (.A0(net1068),
    .A1(\cs_registers_i/mscratch_q_15_ ),
    .S(net620),
    .X(\cs_registers_i/_0366_ ));
 sg13g2_mux2_1 \cs_registers_i/_5197_  (.A0(net1055),
    .A1(\cs_registers_i/mscratch_q_16_ ),
    .S(net619),
    .X(\cs_registers_i/_0367_ ));
 sg13g2_mux2_1 \cs_registers_i/_5198_  (.A0(net1053),
    .A1(\cs_registers_i/mscratch_q_17_ ),
    .S(net618),
    .X(\cs_registers_i/_0368_ ));
 sg13g2_mux2_1 \cs_registers_i/_5199_  (.A0(net1051),
    .A1(\cs_registers_i/mscratch_q_18_ ),
    .S(net618),
    .X(\cs_registers_i/_0369_ ));
 sg13g2_buf_4 fanout451 (.X(net451),
    .A(net453));
 sg13g2_mux2_1 \cs_registers_i/_5201_  (.A0(net1050),
    .A1(\cs_registers_i/mscratch_q_19_ ),
    .S(net617),
    .X(\cs_registers_i/_0370_ ));
 sg13g2_mux2_1 \cs_registers_i/_5202_  (.A0(net1067),
    .A1(\cs_registers_i/mscratch_q_1_ ),
    .S(net617),
    .X(\cs_registers_i/_0371_ ));
 sg13g2_mux2_1 \cs_registers_i/_5203_  (.A0(net1049),
    .A1(\cs_registers_i/mscratch_q_20_ ),
    .S(net616),
    .X(\cs_registers_i/_0372_ ));
 sg13g2_mux2_1 \cs_registers_i/_5204_  (.A0(net1047),
    .A1(\cs_registers_i/mscratch_q_21_ ),
    .S(net618),
    .X(\cs_registers_i/_0373_ ));
 sg13g2_mux2_1 \cs_registers_i/_5205_  (.A0(net1027),
    .A1(\cs_registers_i/mscratch_q_22_ ),
    .S(net616),
    .X(\cs_registers_i/_0374_ ));
 sg13g2_mux2_1 \cs_registers_i/_5206_  (.A0(net1046),
    .A1(\cs_registers_i/mscratch_q_23_ ),
    .S(net616),
    .X(\cs_registers_i/_0375_ ));
 sg13g2_mux2_1 \cs_registers_i/_5207_  (.A0(net1044),
    .A1(\cs_registers_i/mscratch_q_24_ ),
    .S(net616),
    .X(\cs_registers_i/_0376_ ));
 sg13g2_mux2_1 \cs_registers_i/_5208_  (.A0(net1043),
    .A1(\cs_registers_i/mscratch_q_25_ ),
    .S(net618),
    .X(\cs_registers_i/_0377_ ));
 sg13g2_mux2_1 \cs_registers_i/_5209_  (.A0(net1066),
    .A1(\cs_registers_i/mscratch_q_26_ ),
    .S(net618),
    .X(\cs_registers_i/_0378_ ));
 sg13g2_mux2_1 \cs_registers_i/_5210_  (.A0(net1026),
    .A1(\cs_registers_i/mscratch_q_27_ ),
    .S(net618),
    .X(\cs_registers_i/_0379_ ));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(net453));
 sg13g2_mux2_1 \cs_registers_i/_5212_  (.A0(net1042),
    .A1(\cs_registers_i/mscratch_q_28_ ),
    .S(net618),
    .X(\cs_registers_i/_0380_ ));
 sg13g2_mux2_1 \cs_registers_i/_5213_  (.A0(net1040),
    .A1(\cs_registers_i/mscratch_q_29_ ),
    .S(net620),
    .X(\cs_registers_i/_0381_ ));
 sg13g2_mux2_1 \cs_registers_i/_5214_  (.A0(net1038),
    .A1(\cs_registers_i/mscratch_q_2_ ),
    .S(net616),
    .X(\cs_registers_i/_0382_ ));
 sg13g2_mux2_1 \cs_registers_i/_5215_  (.A0(net1037),
    .A1(\cs_registers_i/mscratch_q_30_ ),
    .S(net619),
    .X(\cs_registers_i/_0383_ ));
 sg13g2_mux2_1 \cs_registers_i/_5216_  (.A0(net1035),
    .A1(\cs_registers_i/mscratch_q_31_ ),
    .S(net619),
    .X(\cs_registers_i/_0384_ ));
 sg13g2_mux2_1 \cs_registers_i/_5217_  (.A0(net1033),
    .A1(\cs_registers_i/mscratch_q_3_ ),
    .S(net617),
    .X(\cs_registers_i/_0385_ ));
 sg13g2_mux2_1 \cs_registers_i/_5218_  (.A0(net1032),
    .A1(\cs_registers_i/mscratch_q_4_ ),
    .S(net617),
    .X(\cs_registers_i/_0386_ ));
 sg13g2_mux2_1 \cs_registers_i/_5219_  (.A0(net1065),
    .A1(\cs_registers_i/mscratch_q_5_ ),
    .S(net617),
    .X(\cs_registers_i/_0387_ ));
 sg13g2_mux2_1 \cs_registers_i/_5220_  (.A0(net1064),
    .A1(\cs_registers_i/mscratch_q_6_ ),
    .S(net617),
    .X(\cs_registers_i/_0388_ ));
 sg13g2_mux2_1 \cs_registers_i/_5221_  (.A0(net1031),
    .A1(\cs_registers_i/mscratch_q_7_ ),
    .S(net616),
    .X(\cs_registers_i/_0389_ ));
 sg13g2_mux2_1 \cs_registers_i/_5222_  (.A0(net1025),
    .A1(\cs_registers_i/mscratch_q_8_ ),
    .S(net620),
    .X(\cs_registers_i/_0390_ ));
 sg13g2_mux2_1 \cs_registers_i/_5223_  (.A0(net1030),
    .A1(\cs_registers_i/mscratch_q_9_ ),
    .S(net619),
    .X(\cs_registers_i/_0391_ ));
 sg13g2_mux2_1 \cs_registers_i/_5224_  (.A0(\cs_registers_i/mcause_q_0_ ),
    .A1(\cs_registers_i/mstack_cause_q_0_ ),
    .S(net1284),
    .X(\cs_registers_i/_0392_ ));
 sg13g2_mux2_1 \cs_registers_i/_5225_  (.A0(\cs_registers_i/mcause_q_1_ ),
    .A1(\cs_registers_i/mstack_cause_q_1_ ),
    .S(net1286),
    .X(\cs_registers_i/_0393_ ));
 sg13g2_mux2_1 \cs_registers_i/_5226_  (.A0(\cs_registers_i/mcause_q_2_ ),
    .A1(\cs_registers_i/mstack_cause_q_2_ ),
    .S(net1284),
    .X(\cs_registers_i/_0394_ ));
 sg13g2_mux2_1 \cs_registers_i/_5227_  (.A0(\cs_registers_i/mcause_q_3_ ),
    .A1(\cs_registers_i/mstack_cause_q_3_ ),
    .S(net1284),
    .X(\cs_registers_i/_0395_ ));
 sg13g2_mux2_1 \cs_registers_i/_5228_  (.A0(\cs_registers_i/mcause_q_4_ ),
    .A1(\cs_registers_i/mstack_cause_q_4_ ),
    .S(net1285),
    .X(\cs_registers_i/_0396_ ));
 sg13g2_mux2_1 \cs_registers_i/_5229_  (.A0(\cs_registers_i/mcause_q_5_ ),
    .A1(\cs_registers_i/mstack_cause_q_5_ ),
    .S(net1285),
    .X(\cs_registers_i/_0397_ ));
 sg13g2_mux2_1 \cs_registers_i/_5230_  (.A0(\cs_registers_i/mcause_q_6_ ),
    .A1(\cs_registers_i/mstack_cause_q_6_ ),
    .S(net1286),
    .X(\cs_registers_i/_0398_ ));
 sg13g2_mux2_1 \cs_registers_i/_5231_  (.A0(crash_dump_o_0_),
    .A1(\cs_registers_i/mstack_epc_q_0_ ),
    .S(net1285),
    .X(\cs_registers_i/_0399_ ));
 sg13g2_buf_4 fanout449 (.X(net449),
    .A(net453));
 sg13g2_mux2_1 \cs_registers_i/_5233_  (.A0(crash_dump_o_10_),
    .A1(\cs_registers_i/mstack_epc_q_10_ ),
    .S(net1289),
    .X(\cs_registers_i/_0400_ ));
 sg13g2_mux2_1 \cs_registers_i/_5234_  (.A0(crash_dump_o_11_),
    .A1(\cs_registers_i/mstack_epc_q_11_ ),
    .S(net1285),
    .X(\cs_registers_i/_0401_ ));
 sg13g2_mux2_1 \cs_registers_i/_5235_  (.A0(crash_dump_o_12_),
    .A1(\cs_registers_i/mstack_epc_q_12_ ),
    .S(net1289),
    .X(\cs_registers_i/_0402_ ));
 sg13g2_mux2_1 \cs_registers_i/_5236_  (.A0(crash_dump_o_13_),
    .A1(\cs_registers_i/mstack_epc_q_13_ ),
    .S(net1290),
    .X(\cs_registers_i/_0403_ ));
 sg13g2_mux2_1 \cs_registers_i/_5237_  (.A0(crash_dump_o_14_),
    .A1(\cs_registers_i/mstack_epc_q_14_ ),
    .S(net1284),
    .X(\cs_registers_i/_0404_ ));
 sg13g2_mux2_1 \cs_registers_i/_5238_  (.A0(crash_dump_o_15_),
    .A1(\cs_registers_i/mstack_epc_q_15_ ),
    .S(net1284),
    .X(\cs_registers_i/_0405_ ));
 sg13g2_mux2_1 \cs_registers_i/_5239_  (.A0(crash_dump_o_16_),
    .A1(\cs_registers_i/mstack_epc_q_16_ ),
    .S(net1287),
    .X(\cs_registers_i/_0406_ ));
 sg13g2_mux2_1 \cs_registers_i/_5240_  (.A0(crash_dump_o_17_),
    .A1(\cs_registers_i/mstack_epc_q_17_ ),
    .S(net1287),
    .X(\cs_registers_i/_0407_ ));
 sg13g2_mux2_1 \cs_registers_i/_5241_  (.A0(crash_dump_o_18_),
    .A1(\cs_registers_i/mstack_epc_q_18_ ),
    .S(net1289),
    .X(\cs_registers_i/_0408_ ));
 sg13g2_mux2_1 \cs_registers_i/_5242_  (.A0(crash_dump_o_19_),
    .A1(\cs_registers_i/mstack_epc_q_19_ ),
    .S(net1287),
    .X(\cs_registers_i/_0409_ ));
 sg13g2_buf_4 fanout448 (.X(net448),
    .A(net453));
 sg13g2_mux2_1 \cs_registers_i/_5244_  (.A0(crash_dump_o_1_),
    .A1(\cs_registers_i/mstack_epc_q_1_ ),
    .S(net1286),
    .X(\cs_registers_i/_0410_ ));
 sg13g2_mux2_1 \cs_registers_i/_5245_  (.A0(crash_dump_o_20_),
    .A1(\cs_registers_i/mstack_epc_q_20_ ),
    .S(net1287),
    .X(\cs_registers_i/_0411_ ));
 sg13g2_mux2_1 \cs_registers_i/_5246_  (.A0(crash_dump_o_21_),
    .A1(\cs_registers_i/mstack_epc_q_21_ ),
    .S(net1287),
    .X(\cs_registers_i/_0412_ ));
 sg13g2_mux2_1 \cs_registers_i/_5247_  (.A0(crash_dump_o_22_),
    .A1(\cs_registers_i/mstack_epc_q_22_ ),
    .S(net1287),
    .X(\cs_registers_i/_0413_ ));
 sg13g2_mux2_1 \cs_registers_i/_5248_  (.A0(crash_dump_o_23_),
    .A1(\cs_registers_i/mstack_epc_q_23_ ),
    .S(net1284),
    .X(\cs_registers_i/_0414_ ));
 sg13g2_mux2_1 \cs_registers_i/_5249_  (.A0(crash_dump_o_24_),
    .A1(\cs_registers_i/mstack_epc_q_24_ ),
    .S(net1289),
    .X(\cs_registers_i/_0415_ ));
 sg13g2_mux2_1 \cs_registers_i/_5250_  (.A0(crash_dump_o_25_),
    .A1(\cs_registers_i/mstack_epc_q_25_ ),
    .S(net1288),
    .X(\cs_registers_i/_0416_ ));
 sg13g2_mux2_1 \cs_registers_i/_5251_  (.A0(crash_dump_o_26_),
    .A1(\cs_registers_i/mstack_epc_q_26_ ),
    .S(net1287),
    .X(\cs_registers_i/_0417_ ));
 sg13g2_mux2_1 \cs_registers_i/_5252_  (.A0(crash_dump_o_27_),
    .A1(\cs_registers_i/mstack_epc_q_27_ ),
    .S(net1288),
    .X(\cs_registers_i/_0418_ ));
 sg13g2_mux2_1 \cs_registers_i/_5253_  (.A0(crash_dump_o_28_),
    .A1(\cs_registers_i/mstack_epc_q_28_ ),
    .S(net1287),
    .X(\cs_registers_i/_0419_ ));
 sg13g2_buf_4 fanout447 (.X(net447),
    .A(\id_stage_i.controller_i.instr_i_22_ ));
 sg13g2_mux2_1 \cs_registers_i/_5255_  (.A0(crash_dump_o_29_),
    .A1(\cs_registers_i/mstack_epc_q_29_ ),
    .S(net1290),
    .X(\cs_registers_i/_0420_ ));
 sg13g2_mux2_1 \cs_registers_i/_5256_  (.A0(crash_dump_o_2_),
    .A1(\cs_registers_i/mstack_epc_q_2_ ),
    .S(net1289),
    .X(\cs_registers_i/_0421_ ));
 sg13g2_mux2_1 \cs_registers_i/_5257_  (.A0(crash_dump_o_30_),
    .A1(\cs_registers_i/mstack_epc_q_30_ ),
    .S(net1288),
    .X(\cs_registers_i/_0422_ ));
 sg13g2_mux2_1 \cs_registers_i/_5258_  (.A0(crash_dump_o_31_),
    .A1(\cs_registers_i/mstack_epc_q_31_ ),
    .S(net1289),
    .X(\cs_registers_i/_0423_ ));
 sg13g2_mux2_1 \cs_registers_i/_5259_  (.A0(crash_dump_o_3_),
    .A1(\cs_registers_i/mstack_epc_q_3_ ),
    .S(net1284),
    .X(\cs_registers_i/_0424_ ));
 sg13g2_mux2_1 \cs_registers_i/_5260_  (.A0(crash_dump_o_4_),
    .A1(\cs_registers_i/mstack_epc_q_4_ ),
    .S(net1284),
    .X(\cs_registers_i/_0425_ ));
 sg13g2_mux2_1 \cs_registers_i/_5261_  (.A0(crash_dump_o_5_),
    .A1(\cs_registers_i/mstack_epc_q_5_ ),
    .S(net1285),
    .X(\cs_registers_i/_0426_ ));
 sg13g2_mux2_1 \cs_registers_i/_5262_  (.A0(crash_dump_o_6_),
    .A1(\cs_registers_i/mstack_epc_q_6_ ),
    .S(net1288),
    .X(\cs_registers_i/_0427_ ));
 sg13g2_mux2_1 \cs_registers_i/_5263_  (.A0(crash_dump_o_7_),
    .A1(\cs_registers_i/mstack_epc_q_7_ ),
    .S(net1288),
    .X(\cs_registers_i/_0428_ ));
 sg13g2_mux2_1 \cs_registers_i/_5264_  (.A0(crash_dump_o_8_),
    .A1(\cs_registers_i/mstack_epc_q_8_ ),
    .S(net1288),
    .X(\cs_registers_i/_0429_ ));
 sg13g2_mux2_1 \cs_registers_i/_5265_  (.A0(crash_dump_o_9_),
    .A1(\cs_registers_i/mstack_epc_q_9_ ),
    .S(net1289),
    .X(\cs_registers_i/_0430_ ));
 sg13g2_mux2_1 \cs_registers_i/_5266_  (.A0(\cs_registers_i/mstatus_q_2_ ),
    .A1(\cs_registers_i/mstack_q_0_ ),
    .S(net1286),
    .X(\cs_registers_i/_0431_ ));
 sg13g2_mux2_1 \cs_registers_i/_5267_  (.A0(\cs_registers_i/mstatus_q_3_ ),
    .A1(\cs_registers_i/mstack_q_1_ ),
    .S(net1286),
    .X(\cs_registers_i/_0432_ ));
 sg13g2_mux2_1 \cs_registers_i/_5268_  (.A0(\cs_registers_i/_0005_ ),
    .A1(net2496),
    .S(net1299),
    .X(\cs_registers_i/_0433_ ));
 sg13g2_nand2_1 \cs_registers_i/_5269_  (.Y(\cs_registers_i/_2341_ ),
    .A(\cs_registers_i/mstatus_q_3_ ),
    .B(\cs_registers_i/mstatus_q_2_ ));
 sg13g2_nor2_1 \cs_registers_i/_5270_  (.A(net1053),
    .B(\cs_registers_i/_1581_ ),
    .Y(\cs_registers_i/_2342_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5271_  (.B2(net345),
    .C1(\cs_registers_i/_2342_ ),
    .B1(\cs_registers_i/_2341_ ),
    .A1(\cs_registers_i/_0847_ ),
    .Y(\cs_registers_i/_0434_ ),
    .A2(\cs_registers_i/_1581_ ));
 sg13g2_or2_1 \cs_registers_i/_5272_  (.X(\cs_registers_i/_2343_ ),
    .B(net345),
    .A(\cs_registers_i/_0006_ ));
 sg13g2_nand3_1 \cs_registers_i/_5273_  (.B(net345),
    .C(net255),
    .A(\cs_registers_i/mstatus_q_2_ ),
    .Y(\cs_registers_i/_2344_ ));
 sg13g2_a21oi_1 \cs_registers_i/_5274_  (.A1(\cs_registers_i/_2343_ ),
    .A2(\cs_registers_i/_2344_ ),
    .Y(\cs_registers_i/_2345_ ),
    .B1(\cs_registers_i/_1399_ ));
 sg13g2_nor2_1 \cs_registers_i/_5275_  (.A(net255),
    .B(\cs_registers_i/_2343_ ),
    .Y(\cs_registers_i/_2346_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5276_  (.B1(\cs_registers_i/_1581_ ),
    .Y(\cs_registers_i/_2347_ ),
    .A1(\cs_registers_i/_2345_ ),
    .A2(\cs_registers_i/_2346_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5277_  (.B1(\cs_registers_i/_1586_ ),
    .Y(\cs_registers_i/_2348_ ),
    .A1(net1070),
    .A2(net1028));
 sg13g2_a22oi_1 \cs_registers_i/_5278_  (.Y(\cs_registers_i/_2349_ ),
    .B1(net290),
    .B2(\cs_registers_i/mstack_q_0_ ),
    .A2(net1299),
    .A1(\id_stage_i.controller_i.priv_mode_i_0_ ));
 sg13g2_and3_1 \cs_registers_i/_5279_  (.X(\cs_registers_i/_0435_ ),
    .A(\cs_registers_i/_2347_ ),
    .B(\cs_registers_i/_2348_ ),
    .C(\cs_registers_i/_2349_ ));
 sg13g2_or2_1 \cs_registers_i/_5280_  (.X(\cs_registers_i/_2350_ ),
    .B(net344),
    .A(\cs_registers_i/_0007_ ));
 sg13g2_nand3_1 \cs_registers_i/_5281_  (.B(net345),
    .C(net255),
    .A(\cs_registers_i/mstatus_q_3_ ),
    .Y(\cs_registers_i/_2351_ ));
 sg13g2_a21oi_1 \cs_registers_i/_5282_  (.A1(\cs_registers_i/_2350_ ),
    .A2(\cs_registers_i/_2351_ ),
    .Y(\cs_registers_i/_2352_ ),
    .B1(\cs_registers_i/_1399_ ));
 sg13g2_nor2_1 \cs_registers_i/_5283_  (.A(net255),
    .B(\cs_registers_i/_2350_ ),
    .Y(\cs_registers_i/_2353_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5284_  (.B1(\cs_registers_i/_1581_ ),
    .Y(\cs_registers_i/_2354_ ),
    .A1(\cs_registers_i/_2352_ ),
    .A2(\cs_registers_i/_2353_ ));
 sg13g2_a22oi_1 \cs_registers_i/_5285_  (.Y(\cs_registers_i/_2355_ ),
    .B1(net290),
    .B2(\cs_registers_i/mstack_q_1_ ),
    .A2(net1299),
    .A1(net2116));
 sg13g2_and3_1 \cs_registers_i/_5286_  (.X(\cs_registers_i/_0436_ ),
    .A(\cs_registers_i/_2348_ ),
    .B(\cs_registers_i/_2354_ ),
    .C(\cs_registers_i/_2355_ ));
 sg13g2_nand4_1 \cs_registers_i/_5287_  (.B(net1286),
    .C(\cs_registers_i/_1581_ ),
    .A(\cs_registers_i/mstatus_q_4_ ),
    .Y(\cs_registers_i/_2356_ ),
    .D(\cs_registers_i/_1582_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5288_  (.Y(\cs_registers_i/_2357_ ),
    .B(\id_stage_i.controller_i.nmi_mode_o ),
    .A_N(\cs_registers_i/mstack_q_2_ ));
 sg13g2_and2_1 \cs_registers_i/_5289_  (.A(net344),
    .B(\cs_registers_i/_2357_ ),
    .X(\cs_registers_i/_2358_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5290_  (.B2(net1031),
    .C1(\cs_registers_i/_2358_ ),
    .B1(\cs_registers_i/_1586_ ),
    .A1(csr_mstatus_mie),
    .Y(\cs_registers_i/_2359_ ),
    .A2(net1299));
 sg13g2_nand2_1 \cs_registers_i/_5291_  (.Y(\cs_registers_i/_0437_ ),
    .A(\cs_registers_i/_2356_ ),
    .B(\cs_registers_i/_2359_ ));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(net447));
 sg13g2_nand3_1 \cs_registers_i/_5293_  (.B(\cs_registers_i/_0948_ ),
    .C(net1148),
    .A(net722),
    .Y(\cs_registers_i/_2361_ ));
 sg13g2_buf_4 fanout445 (.X(net445),
    .A(net447));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(net447));
 sg13g2_buf_4 fanout443 (.X(net443),
    .A(net447));
 sg13g2_nand2b_1 \cs_registers_i/_5297_  (.Y(\cs_registers_i/_2365_ ),
    .B(net608),
    .A_N(\cs_registers_i/mtval_q_0_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5298_  (.B1(\cs_registers_i/_2365_ ),
    .Y(\cs_registers_i/_2366_ ),
    .A1(net1063),
    .A2(net608));
 sg13g2_buf_4 fanout442 (.X(net442),
    .A(net447));
 sg13g2_nand2_1 \cs_registers_i/_5300_  (.Y(\cs_registers_i/_2368_ ),
    .A(csr_mtval_0_),
    .B(net1295));
 sg13g2_o21ai_1 \cs_registers_i/_5301_  (.B1(\cs_registers_i/_2368_ ),
    .Y(\cs_registers_i/_0438_ ),
    .A1(net1299),
    .A2(\cs_registers_i/_2366_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5302_  (.Y(\cs_registers_i/_2369_ ),
    .B(net606),
    .A_N(\cs_registers_i/mtval_q_10_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5303_  (.B1(\cs_registers_i/_2369_ ),
    .Y(\cs_registers_i/_2370_ ),
    .A1(net1059),
    .A2(net606));
 sg13g2_nand2_1 \cs_registers_i/_5304_  (.Y(\cs_registers_i/_2371_ ),
    .A(csr_mtval_10_),
    .B(net1293));
 sg13g2_o21ai_1 \cs_registers_i/_5305_  (.B1(\cs_registers_i/_2371_ ),
    .Y(\cs_registers_i/_0439_ ),
    .A1(net1296),
    .A2(\cs_registers_i/_2370_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5306_  (.Y(\cs_registers_i/_2372_ ),
    .B(net609),
    .A_N(\cs_registers_i/mtval_q_11_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5307_  (.B1(\cs_registers_i/_2372_ ),
    .Y(\cs_registers_i/_2373_ ),
    .A1(net1070),
    .A2(net609));
 sg13g2_nand2_2 \cs_registers_i/_5308_  (.Y(\cs_registers_i/_2374_ ),
    .A(csr_mtval_11_),
    .B(net1292));
 sg13g2_o21ai_1 \cs_registers_i/_5309_  (.B1(\cs_registers_i/_2374_ ),
    .Y(\cs_registers_i/_0440_ ),
    .A1(net1298),
    .A2(\cs_registers_i/_2373_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5310_  (.Y(\cs_registers_i/_2375_ ),
    .B(net612),
    .A_N(\cs_registers_i/mtval_q_12_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5311_  (.B1(\cs_registers_i/_2375_ ),
    .Y(\cs_registers_i/_2376_ ),
    .A1(net1028),
    .A2(net612));
 sg13g2_nand2_2 \cs_registers_i/_5312_  (.Y(\cs_registers_i/_2377_ ),
    .A(csr_mtval_12_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5313_  (.B1(\cs_registers_i/_2377_ ),
    .Y(\cs_registers_i/_0441_ ),
    .A1(net1298),
    .A2(\cs_registers_i/_2376_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5314_  (.Y(\cs_registers_i/_2378_ ),
    .B(net610),
    .A_N(\cs_registers_i/mtval_q_13_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5315_  (.B1(\cs_registers_i/_2378_ ),
    .Y(\cs_registers_i/_2379_ ),
    .A1(net1057),
    .A2(net610));
 sg13g2_nand2_2 \cs_registers_i/_5316_  (.Y(\cs_registers_i/_2380_ ),
    .A(csr_mtval_13_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5317_  (.B1(\cs_registers_i/_2380_ ),
    .Y(\cs_registers_i/_0442_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2379_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5318_  (.Y(\cs_registers_i/_2381_ ),
    .B(net607),
    .A_N(\cs_registers_i/mtval_q_14_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5319_  (.B1(\cs_registers_i/_2381_ ),
    .Y(\cs_registers_i/_2382_ ),
    .A1(net1056),
    .A2(net607));
 sg13g2_nand2_1 \cs_registers_i/_5320_  (.Y(\cs_registers_i/_2383_ ),
    .A(csr_mtval_14_),
    .B(net1292));
 sg13g2_o21ai_1 \cs_registers_i/_5321_  (.B1(\cs_registers_i/_2383_ ),
    .Y(\cs_registers_i/_0443_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2382_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5322_  (.Y(\cs_registers_i/_2384_ ),
    .B(net610),
    .A_N(\cs_registers_i/mtval_q_15_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5323_  (.B1(\cs_registers_i/_2384_ ),
    .Y(\cs_registers_i/_2385_ ),
    .A1(net1068),
    .A2(net610));
 sg13g2_nand2_2 \cs_registers_i/_5324_  (.Y(\cs_registers_i/_2386_ ),
    .A(csr_mtval_15_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5325_  (.B1(\cs_registers_i/_2386_ ),
    .Y(\cs_registers_i/_0444_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2385_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5326_  (.Y(\cs_registers_i/_2387_ ),
    .B(net611),
    .A_N(\cs_registers_i/mtval_q_16_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5327_  (.B1(\cs_registers_i/_2387_ ),
    .Y(\cs_registers_i/_2388_ ),
    .A1(net1055),
    .A2(net611));
 sg13g2_nand2_1 \cs_registers_i/_5328_  (.Y(\cs_registers_i/_2389_ ),
    .A(csr_mtval_16_),
    .B(net1306));
 sg13g2_o21ai_1 \cs_registers_i/_5329_  (.B1(\cs_registers_i/_2389_ ),
    .Y(\cs_registers_i/_0445_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2388_ ));
 sg13g2_buf_4 fanout441 (.X(net441),
    .A(\id_stage_i.controller_i.instr_i_30_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5331_  (.Y(\cs_registers_i/_2391_ ),
    .B(net612),
    .A_N(\cs_registers_i/mtval_q_17_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5332_  (.B1(\cs_registers_i/_2391_ ),
    .Y(\cs_registers_i/_2392_ ),
    .A1(net1053),
    .A2(net612));
 sg13g2_buf_2 fanout440 (.A(\id_stage_i.controller_i.instr_is_compressed_i ),
    .X(net440));
 sg13g2_nand2_2 \cs_registers_i/_5334_  (.Y(\cs_registers_i/_2394_ ),
    .A(csr_mtval_17_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5335_  (.B1(\cs_registers_i/_2394_ ),
    .Y(\cs_registers_i/_0446_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2392_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5336_  (.Y(\cs_registers_i/_2395_ ),
    .B(net613),
    .A_N(\cs_registers_i/mtval_q_18_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5337_  (.B1(\cs_registers_i/_2395_ ),
    .Y(\cs_registers_i/_2396_ ),
    .A1(net1051),
    .A2(net613));
 sg13g2_nand2_2 \cs_registers_i/_5338_  (.Y(\cs_registers_i/_2397_ ),
    .A(csr_mtval_18_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5339_  (.B1(\cs_registers_i/_2397_ ),
    .Y(\cs_registers_i/_0447_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2396_ ));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(\id_stage_i.controller_i.instr_is_compressed_i ));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(\id_stage_i.controller_i.instr_is_compressed_i ));
 sg13g2_nand2b_1 \cs_registers_i/_5342_  (.Y(\cs_registers_i/_2400_ ),
    .B(net612),
    .A_N(\cs_registers_i/mtval_q_19_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5343_  (.B1(\cs_registers_i/_2400_ ),
    .Y(\cs_registers_i/_2401_ ),
    .A1(net1050),
    .A2(net612));
 sg13g2_nand2_2 \cs_registers_i/_5344_  (.Y(\cs_registers_i/_2402_ ),
    .A(csr_mtval_19_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5345_  (.B1(\cs_registers_i/_2402_ ),
    .Y(\cs_registers_i/_0448_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2401_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5346_  (.Y(\cs_registers_i/_2403_ ),
    .B(net608),
    .A_N(\cs_registers_i/mtval_q_1_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5347_  (.B1(\cs_registers_i/_2403_ ),
    .Y(\cs_registers_i/_2404_ ),
    .A1(net1067),
    .A2(net608));
 sg13g2_nand2_1 \cs_registers_i/_5348_  (.Y(\cs_registers_i/_2405_ ),
    .A(csr_mtval_1_),
    .B(net1299));
 sg13g2_o21ai_1 \cs_registers_i/_5349_  (.B1(\cs_registers_i/_2405_ ),
    .Y(\cs_registers_i/_0449_ ),
    .A1(net1299),
    .A2(\cs_registers_i/_2404_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5350_  (.Y(\cs_registers_i/_2406_ ),
    .B(net604),
    .A_N(\cs_registers_i/mtval_q_20_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5351_  (.B1(\cs_registers_i/_2406_ ),
    .Y(\cs_registers_i/_2407_ ),
    .A1(net1049),
    .A2(net605));
 sg13g2_nand2_1 \cs_registers_i/_5352_  (.Y(\cs_registers_i/_2408_ ),
    .A(csr_mtval_20_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5353_  (.B1(\cs_registers_i/_2408_ ),
    .Y(\cs_registers_i/_0450_ ),
    .A1(net1292),
    .A2(\cs_registers_i/_2407_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5354_  (.Y(\cs_registers_i/_2409_ ),
    .B(net612),
    .A_N(\cs_registers_i/mtval_q_21_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5355_  (.B1(\cs_registers_i/_2409_ ),
    .Y(\cs_registers_i/_2410_ ),
    .A1(net1047),
    .A2(net614));
 sg13g2_nand2_2 \cs_registers_i/_5356_  (.Y(\cs_registers_i/_2411_ ),
    .A(csr_mtval_21_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5357_  (.B1(\cs_registers_i/_2411_ ),
    .Y(\cs_registers_i/_0451_ ),
    .A1(net1298),
    .A2(\cs_registers_i/_2410_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5358_  (.Y(\cs_registers_i/_2412_ ),
    .B(net613),
    .A_N(\cs_registers_i/mtval_q_22_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5359_  (.B1(\cs_registers_i/_2412_ ),
    .Y(\cs_registers_i/_2413_ ),
    .A1(net1027),
    .A2(net613));
 sg13g2_nand2_2 \cs_registers_i/_5360_  (.Y(\cs_registers_i/_2414_ ),
    .A(csr_mtval_22_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5361_  (.B1(\cs_registers_i/_2414_ ),
    .Y(\cs_registers_i/_0452_ ),
    .A1(net1306),
    .A2(\cs_registers_i/_2413_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5362_  (.Y(\cs_registers_i/_2415_ ),
    .B(net612),
    .A_N(\cs_registers_i/mtval_q_23_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5363_  (.B1(\cs_registers_i/_2415_ ),
    .Y(\cs_registers_i/_2416_ ),
    .A1(net1046),
    .A2(net610));
 sg13g2_nand2_2 \cs_registers_i/_5364_  (.Y(\cs_registers_i/_2417_ ),
    .A(csr_mtval_23_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5365_  (.B1(\cs_registers_i/_2417_ ),
    .Y(\cs_registers_i/_0453_ ),
    .A1(net1298),
    .A2(\cs_registers_i/_2416_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5366_  (.Y(\cs_registers_i/_2418_ ),
    .B(net604),
    .A_N(\cs_registers_i/mtval_q_24_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5367_  (.B1(\cs_registers_i/_2418_ ),
    .Y(\cs_registers_i/_2419_ ),
    .A1(net1044),
    .A2(net605));
 sg13g2_nand2_1 \cs_registers_i/_5368_  (.Y(\cs_registers_i/_2420_ ),
    .A(csr_mtval_24_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5369_  (.B1(\cs_registers_i/_2420_ ),
    .Y(\cs_registers_i/_0454_ ),
    .A1(net1301),
    .A2(\cs_registers_i/_2419_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5370_  (.Y(\cs_registers_i/_2421_ ),
    .B(net613),
    .A_N(\cs_registers_i/mtval_q_25_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5371_  (.B1(\cs_registers_i/_2421_ ),
    .Y(\cs_registers_i/_2422_ ),
    .A1(net1043),
    .A2(net613));
 sg13g2_nand2_2 \cs_registers_i/_5372_  (.Y(\cs_registers_i/_2423_ ),
    .A(csr_mtval_25_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5373_  (.B1(\cs_registers_i/_2423_ ),
    .Y(\cs_registers_i/_0455_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2422_ ));
 sg13g2_buf_2 fanout437 (.A(\id_stage_i.controller_i.instr_valid_i ),
    .X(net437));
 sg13g2_nand2b_1 \cs_registers_i/_5375_  (.Y(\cs_registers_i/_2425_ ),
    .B(net614),
    .A_N(\cs_registers_i/mtval_q_26_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5376_  (.B1(\cs_registers_i/_2425_ ),
    .Y(\cs_registers_i/_2426_ ),
    .A1(net1066),
    .A2(net613));
 sg13g2_buf_2 fanout436 (.A(\id_stage_i.controller_i.instr_valid_i ),
    .X(net436));
 sg13g2_nand2_2 \cs_registers_i/_5378_  (.Y(\cs_registers_i/_2428_ ),
    .A(csr_mtval_26_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5379_  (.B1(\cs_registers_i/_2428_ ),
    .Y(\cs_registers_i/_0456_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2426_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5380_  (.Y(\cs_registers_i/_2429_ ),
    .B(net614),
    .A_N(\cs_registers_i/mtval_q_27_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5381_  (.B1(\cs_registers_i/_2429_ ),
    .Y(\cs_registers_i/_2430_ ),
    .A1(net1026),
    .A2(net613));
 sg13g2_nand2_1 \cs_registers_i/_5382_  (.Y(\cs_registers_i/_2431_ ),
    .A(csr_mtval_27_),
    .B(net1306));
 sg13g2_o21ai_1 \cs_registers_i/_5383_  (.B1(\cs_registers_i/_2431_ ),
    .Y(\cs_registers_i/_0457_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2430_ ));
 sg13g2_buf_2 fanout435 (.A(\if_stage_i.prefetch_buffer_i.fifo_busy_0_ ),
    .X(net435));
 sg13g2_buf_1 fanout434 (.A(net435),
    .X(net434));
 sg13g2_nand2b_1 \cs_registers_i/_5386_  (.Y(\cs_registers_i/_2434_ ),
    .B(net611),
    .A_N(\cs_registers_i/mtval_q_28_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5387_  (.B1(\cs_registers_i/_2434_ ),
    .Y(\cs_registers_i/_2435_ ),
    .A1(net1042),
    .A2(net611));
 sg13g2_nand2_2 \cs_registers_i/_5388_  (.Y(\cs_registers_i/_2436_ ),
    .A(csr_mtval_28_),
    .B(net1301));
 sg13g2_o21ai_1 \cs_registers_i/_5389_  (.B1(\cs_registers_i/_2436_ ),
    .Y(\cs_registers_i/_0458_ ),
    .A1(net1305),
    .A2(\cs_registers_i/_2435_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5390_  (.Y(\cs_registers_i/_2437_ ),
    .B(net610),
    .A_N(\cs_registers_i/mtval_q_29_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5391_  (.B1(\cs_registers_i/_2437_ ),
    .Y(\cs_registers_i/_2438_ ),
    .A1(net1040),
    .A2(net610));
 sg13g2_nand2_1 \cs_registers_i/_5392_  (.Y(\cs_registers_i/_2439_ ),
    .A(csr_mtval_29_),
    .B(net1292));
 sg13g2_o21ai_1 \cs_registers_i/_5393_  (.B1(\cs_registers_i/_2439_ ),
    .Y(\cs_registers_i/_0459_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2438_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5394_  (.Y(\cs_registers_i/_2440_ ),
    .B(net607),
    .A_N(\cs_registers_i/mtval_q_2_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5395_  (.B1(\cs_registers_i/_2440_ ),
    .Y(\cs_registers_i/_2441_ ),
    .A1(net1039),
    .A2(net606));
 sg13g2_nand2_1 \cs_registers_i/_5396_  (.Y(\cs_registers_i/_2442_ ),
    .A(csr_mtval_2_),
    .B(net1296));
 sg13g2_o21ai_1 \cs_registers_i/_5397_  (.B1(\cs_registers_i/_2442_ ),
    .Y(\cs_registers_i/_0460_ ),
    .A1(net1296),
    .A2(\cs_registers_i/_2441_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5398_  (.Y(\cs_registers_i/_2443_ ),
    .B(net610),
    .A_N(\cs_registers_i/mtval_q_30_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5399_  (.B1(\cs_registers_i/_2443_ ),
    .Y(\cs_registers_i/_2444_ ),
    .A1(net1037),
    .A2(net611));
 sg13g2_nand2_1 \cs_registers_i/_5400_  (.Y(\cs_registers_i/_2445_ ),
    .A(csr_mtval_30_),
    .B(net1291));
 sg13g2_o21ai_1 \cs_registers_i/_5401_  (.B1(\cs_registers_i/_2445_ ),
    .Y(\cs_registers_i/_0461_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2444_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5402_  (.Y(\cs_registers_i/_2446_ ),
    .B(net605),
    .A_N(\cs_registers_i/mtval_q_31_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5403_  (.B1(\cs_registers_i/_2446_ ),
    .Y(\cs_registers_i/_2447_ ),
    .A1(net1035),
    .A2(net605));
 sg13g2_nand2_1 \cs_registers_i/_5404_  (.Y(\cs_registers_i/_2448_ ),
    .A(csr_mtval_31_),
    .B(net1292));
 sg13g2_o21ai_1 \cs_registers_i/_5405_  (.B1(\cs_registers_i/_2448_ ),
    .Y(\cs_registers_i/_0462_ ),
    .A1(net1292),
    .A2(\cs_registers_i/_2447_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5406_  (.Y(\cs_registers_i/_2449_ ),
    .B(net604),
    .A_N(\cs_registers_i/mtval_q_3_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5407_  (.B1(\cs_registers_i/_2449_ ),
    .Y(\cs_registers_i/_2450_ ),
    .A1(net1033),
    .A2(net604));
 sg13g2_nand2_1 \cs_registers_i/_5408_  (.Y(\cs_registers_i/_2451_ ),
    .A(csr_mtval_3_),
    .B(net1293));
 sg13g2_o21ai_1 \cs_registers_i/_5409_  (.B1(\cs_registers_i/_2451_ ),
    .Y(\cs_registers_i/_0463_ ),
    .A1(net1293),
    .A2(\cs_registers_i/_2450_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5410_  (.Y(\cs_registers_i/_2452_ ),
    .B(net604),
    .A_N(\cs_registers_i/mtval_q_4_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5411_  (.B1(\cs_registers_i/_2452_ ),
    .Y(\cs_registers_i/_2453_ ),
    .A1(net1032),
    .A2(net604));
 sg13g2_nand2_1 \cs_registers_i/_5412_  (.Y(\cs_registers_i/_2454_ ),
    .A(csr_mtval_4_),
    .B(net1295));
 sg13g2_o21ai_1 \cs_registers_i/_5413_  (.B1(\cs_registers_i/_2454_ ),
    .Y(\cs_registers_i/_0464_ ),
    .A1(net1295),
    .A2(\cs_registers_i/_2453_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5414_  (.Y(\cs_registers_i/_2455_ ),
    .B(net604),
    .A_N(\cs_registers_i/mtval_q_5_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5415_  (.B1(\cs_registers_i/_2455_ ),
    .Y(\cs_registers_i/_2456_ ),
    .A1(net1065),
    .A2(net604));
 sg13g2_nand2_1 \cs_registers_i/_5416_  (.Y(\cs_registers_i/_2457_ ),
    .A(csr_mtval_5_),
    .B(net1295));
 sg13g2_o21ai_1 \cs_registers_i/_5417_  (.B1(\cs_registers_i/_2457_ ),
    .Y(\cs_registers_i/_0465_ ),
    .A1(net1295),
    .A2(\cs_registers_i/_2456_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5418_  (.Y(\cs_registers_i/_2458_ ),
    .B(net606),
    .A_N(\cs_registers_i/mtval_q_6_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5419_  (.B1(\cs_registers_i/_2458_ ),
    .Y(\cs_registers_i/_2459_ ),
    .A1(net1064),
    .A2(net607));
 sg13g2_nand2_2 \cs_registers_i/_5420_  (.Y(\cs_registers_i/_2460_ ),
    .A(csr_mtval_6_),
    .B(net1293));
 sg13g2_o21ai_1 \cs_registers_i/_5421_  (.B1(\cs_registers_i/_2460_ ),
    .Y(\cs_registers_i/_0466_ ),
    .A1(net1300),
    .A2(\cs_registers_i/_2459_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5422_  (.Y(\cs_registers_i/_2461_ ),
    .B(net609),
    .A_N(\cs_registers_i/mtval_q_7_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5423_  (.B1(\cs_registers_i/_2461_ ),
    .Y(\cs_registers_i/_2462_ ),
    .A1(net1031),
    .A2(net609));
 sg13g2_nand2_2 \cs_registers_i/_5424_  (.Y(\cs_registers_i/_2463_ ),
    .A(csr_mtval_7_),
    .B(net1293));
 sg13g2_o21ai_1 \cs_registers_i/_5425_  (.B1(\cs_registers_i/_2463_ ),
    .Y(\cs_registers_i/_0467_ ),
    .A1(net1298),
    .A2(\cs_registers_i/_2462_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5426_  (.Y(\cs_registers_i/_2464_ ),
    .B(net606),
    .A_N(\cs_registers_i/mtval_q_8_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5427_  (.B1(\cs_registers_i/_2464_ ),
    .Y(\cs_registers_i/_2465_ ),
    .A1(net1025),
    .A2(net606));
 sg13g2_nand2_1 \cs_registers_i/_5428_  (.Y(\cs_registers_i/_2466_ ),
    .A(csr_mtval_8_),
    .B(net1296));
 sg13g2_o21ai_1 \cs_registers_i/_5429_  (.B1(\cs_registers_i/_2466_ ),
    .Y(\cs_registers_i/_0468_ ),
    .A1(net1297),
    .A2(\cs_registers_i/_2465_ ));
 sg13g2_nand2b_1 \cs_registers_i/_5430_  (.Y(\cs_registers_i/_2467_ ),
    .B(net606),
    .A_N(\cs_registers_i/mtval_q_9_ ));
 sg13g2_o21ai_1 \cs_registers_i/_5431_  (.B1(\cs_registers_i/_2467_ ),
    .Y(\cs_registers_i/_2468_ ),
    .A1(net1030),
    .A2(net606));
 sg13g2_nand2_1 \cs_registers_i/_5432_  (.Y(\cs_registers_i/_2469_ ),
    .A(csr_mtval_9_),
    .B(net1296));
 sg13g2_o21ai_1 \cs_registers_i/_5433_  (.B1(\cs_registers_i/_2469_ ),
    .Y(\cs_registers_i/_0469_ ),
    .A1(net1296),
    .A2(\cs_registers_i/_2468_ ));
 sg13g2_nor2b_1 \cs_registers_i/_5434_  (.A(net257),
    .B_N(\cs_registers_i/_0008_ ),
    .Y(\cs_registers_i/_2470_ ));
 sg13g2_nor3_1 \cs_registers_i/_5435_  (.A(csr_restore_dret_id),
    .B(net345),
    .C(\cs_registers_i/_2470_ ),
    .Y(\cs_registers_i/_2471_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5436_  (.B2(\cs_registers_i/mstatus_q_2_ ),
    .C1(\cs_registers_i/_2471_ ),
    .B1(net346),
    .A1(csr_restore_dret_id),
    .Y(\cs_registers_i/_0470_ ),
    .A2(net2497));
 sg13g2_nor2b_1 \cs_registers_i/_5437_  (.A(net257),
    .B_N(\cs_registers_i/_0009_ ),
    .Y(\cs_registers_i/_2472_ ));
 sg13g2_nor3_1 \cs_registers_i/_5438_  (.A(csr_restore_dret_id),
    .B(net345),
    .C(\cs_registers_i/_2472_ ),
    .Y(\cs_registers_i/_2473_ ));
 sg13g2_a221oi_1 \cs_registers_i/_5439_  (.B2(\cs_registers_i/mstatus_q_3_ ),
    .C1(\cs_registers_i/_2473_ ),
    .B1(net346),
    .A1(\cs_registers_i/dcsr_q_1_ ),
    .Y(\cs_registers_i/_0471_ ),
    .A2(csr_restore_dret_id));
 sg13g2_mux2_1 \cs_registers_i/_5440_  (.A0(\id_stage_i.controller_i.priv_mode_i_1_ ),
    .A1(\cs_registers_i/mstatus_q_3_ ),
    .S(\cs_registers_i/mstatus_q_1_ ),
    .X(\g_no_pmp.unused_priv_lvl_ls_1_ ));
 sg13g2_mux2_1 \cs_registers_i/_5441_  (.A0(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .A1(\cs_registers_i/mstatus_q_2_ ),
    .S(\cs_registers_i/mstatus_q_1_ ),
    .X(\g_no_pmp.unused_priv_lvl_ls_0_ ));
 sg13g2_buf_2 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_dfrbp_1 \cs_registers_i/csr_depc_o[0]_reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0010_ ),
    .Q_N(\cs_registers_i/_2921_ ),
    .Q(csr_depc_0_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[10]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0011_ ),
    .Q(csr_depc_10_),
    .Q_N(\cs_registers_i/_2920_ ),
    .CLK(clknet_leaf_263_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[11]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0012_ ),
    .Q(csr_depc_11_),
    .Q_N(\cs_registers_i/_2919_ ),
    .CLK(clknet_leaf_259_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[12]_reg  (.RESET_B(net2421),
    .D(\cs_registers_i/_0013_ ),
    .Q(csr_depc_12_),
    .Q_N(\cs_registers_i/_2918_ ),
    .CLK(clknet_leaf_283_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[13]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0014_ ),
    .Q(csr_depc_13_),
    .Q_N(\cs_registers_i/_2917_ ),
    .CLK(clknet_leaf_261_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[14]_reg  (.RESET_B(net2401),
    .D(\cs_registers_i/_0015_ ),
    .Q(csr_depc_14_),
    .Q_N(\cs_registers_i/_2916_ ),
    .CLK(clknet_leaf_262_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[15]_reg  (.RESET_B(net2400),
    .D(\cs_registers_i/_0016_ ),
    .Q(csr_depc_15_),
    .Q_N(\cs_registers_i/_2915_ ),
    .CLK(clknet_leaf_264_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[16]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0017_ ),
    .Q(csr_depc_16_),
    .Q_N(\cs_registers_i/_2914_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[17]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0018_ ),
    .Q(csr_depc_17_),
    .Q_N(\cs_registers_i/_2913_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[18]_reg  (.RESET_B(net2421),
    .D(\cs_registers_i/_0019_ ),
    .Q(csr_depc_18_),
    .Q_N(\cs_registers_i/_2912_ ),
    .CLK(clknet_leaf_261_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[19]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0020_ ),
    .Q(csr_depc_19_),
    .Q_N(\cs_registers_i/_2911_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_depc_o[1]_reg  (.CLK(clknet_leaf_262_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0021_ ),
    .Q_N(\cs_registers_i/_2910_ ),
    .Q(csr_depc_1_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[20]_reg  (.RESET_B(net2408),
    .D(\cs_registers_i/_0022_ ),
    .Q(csr_depc_20_),
    .Q_N(\cs_registers_i/_2909_ ),
    .CLK(clknet_leaf_285_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[21]_reg  (.RESET_B(net2408),
    .D(\cs_registers_i/_0023_ ),
    .Q(csr_depc_21_),
    .Q_N(\cs_registers_i/_2908_ ),
    .CLK(clknet_leaf_284_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[22]_reg  (.RESET_B(net2417),
    .D(\cs_registers_i/_0024_ ),
    .Q(csr_depc_22_),
    .Q_N(\cs_registers_i/_2907_ ),
    .CLK(clknet_leaf_284_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[23]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0025_ ),
    .Q(csr_depc_23_),
    .Q_N(\cs_registers_i/_2906_ ),
    .CLK(clknet_leaf_261_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[24]_reg  (.RESET_B(net2417),
    .D(\cs_registers_i/_0026_ ),
    .Q(csr_depc_24_),
    .Q_N(\cs_registers_i/_2905_ ),
    .CLK(clknet_leaf_284_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_depc_o[25]_reg  (.CLK(clknet_leaf_285_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0027_ ),
    .Q_N(\cs_registers_i/_2904_ ),
    .Q(csr_depc_25_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[26]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0028_ ),
    .Q(csr_depc_26_),
    .Q_N(\cs_registers_i/_2903_ ),
    .CLK(clknet_leaf_283_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[27]_reg  (.RESET_B(net2403),
    .D(\cs_registers_i/_0029_ ),
    .Q(csr_depc_27_),
    .Q_N(\cs_registers_i/_2902_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[28]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0030_ ),
    .Q(csr_depc_28_),
    .Q_N(\cs_registers_i/_2901_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_depc_o[29]_reg  (.CLK(clknet_leaf_259_clk_i),
    .RESET_B(net2420),
    .D(\cs_registers_i/_0031_ ),
    .Q_N(\cs_registers_i/_2900_ ),
    .Q(csr_depc_29_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[2]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0032_ ),
    .Q(csr_depc_2_),
    .Q_N(\cs_registers_i/_2899_ ),
    .CLK(clknet_leaf_285_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[30]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0033_ ),
    .Q(csr_depc_30_),
    .Q_N(\cs_registers_i/_2898_ ),
    .CLK(clknet_leaf_285_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[31]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0034_ ),
    .Q(csr_depc_31_),
    .Q_N(\cs_registers_i/_2897_ ),
    .CLK(clknet_leaf_259_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[3]_reg  (.RESET_B(net2397),
    .D(\cs_registers_i/_0035_ ),
    .Q(csr_depc_3_),
    .Q_N(\cs_registers_i/_2896_ ),
    .CLK(clknet_leaf_256_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[4]_reg  (.RESET_B(net2395),
    .D(\cs_registers_i/_0036_ ),
    .Q(csr_depc_4_),
    .Q_N(\cs_registers_i/_2895_ ),
    .CLK(clknet_leaf_264_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[5]_reg  (.RESET_B(net2398),
    .D(\cs_registers_i/_0037_ ),
    .Q(csr_depc_5_),
    .Q_N(\cs_registers_i/_2894_ ),
    .CLK(clknet_leaf_264_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[6]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0038_ ),
    .Q(csr_depc_6_),
    .Q_N(\cs_registers_i/_2893_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[7]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0039_ ),
    .Q(csr_depc_7_),
    .Q_N(\cs_registers_i/_2892_ ),
    .CLK(clknet_leaf_258_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[8]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0040_ ),
    .Q(csr_depc_8_),
    .Q_N(\cs_registers_i/_2891_ ),
    .CLK(clknet_leaf_284_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_depc_o[9]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0041_ ),
    .Q(csr_depc_9_),
    .Q_N(\cs_registers_i/_2890_ ),
    .CLK(clknet_leaf_260_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[0]_reg  (.RESET_B(net2323),
    .D(\cs_registers_i/_0042_ ),
    .Q(crash_dump_o_0_),
    .Q_N(\cs_registers_i/_2889_ ),
    .CLK(clknet_leaf_254_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[10]_reg  (.RESET_B(net2435),
    .D(\cs_registers_i/_0043_ ),
    .Q(crash_dump_o_10_),
    .Q_N(\cs_registers_i/_2888_ ),
    .CLK(clknet_leaf_265_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[11]_reg  (.RESET_B(net2400),
    .D(\cs_registers_i/_0044_ ),
    .Q(crash_dump_o_11_),
    .Q_N(\cs_registers_i/_2887_ ),
    .CLK(clknet_leaf_253_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[12]_reg  (.RESET_B(net2420),
    .D(\cs_registers_i/_0045_ ),
    .Q(crash_dump_o_12_),
    .Q_N(\cs_registers_i/_2886_ ),
    .CLK(clknet_leaf_266_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[13]_reg  (.RESET_B(net2407),
    .D(\cs_registers_i/_0046_ ),
    .Q(crash_dump_o_13_),
    .Q_N(\cs_registers_i/_2885_ ),
    .CLK(clknet_leaf_267_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[14]_reg  (.RESET_B(net2397),
    .D(\cs_registers_i/_0047_ ),
    .Q(crash_dump_o_14_),
    .Q_N(\cs_registers_i/_2884_ ),
    .CLK(clknet_leaf_254_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[15]_reg  (.RESET_B(net2397),
    .D(\cs_registers_i/_0048_ ),
    .Q(crash_dump_o_15_),
    .Q_N(\cs_registers_i/_2883_ ),
    .CLK(clknet_leaf_253_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[16]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0049_ ),
    .Q(crash_dump_o_16_),
    .Q_N(\cs_registers_i/_2882_ ),
    .CLK(clknet_leaf_249_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[17]_reg  (.RESET_B(net2405),
    .D(\cs_registers_i/_0050_ ),
    .Q(crash_dump_o_17_),
    .Q_N(\cs_registers_i/_2881_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[18]_reg  (.RESET_B(net2420),
    .D(\cs_registers_i/_0051_ ),
    .Q(crash_dump_o_18_),
    .Q_N(\cs_registers_i/_2880_ ),
    .CLK(clknet_leaf_266_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[19]_reg  (.RESET_B(net2429),
    .D(\cs_registers_i/_0052_ ),
    .Q(crash_dump_o_19_),
    .Q_N(\cs_registers_i/_2879_ ),
    .CLK(clknet_leaf_249_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[1]_reg  (.RESET_B(net2399),
    .D(\cs_registers_i/_0053_ ),
    .Q(crash_dump_o_1_),
    .Q_N(\cs_registers_i/_2878_ ),
    .CLK(clknet_leaf_267_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[20]_reg  (.RESET_B(net2323),
    .D(\cs_registers_i/_0054_ ),
    .Q(crash_dump_o_20_),
    .Q_N(\cs_registers_i/_2877_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[21]_reg  (.RESET_B(net2348),
    .D(\cs_registers_i/_0055_ ),
    .Q(crash_dump_o_21_),
    .Q_N(\cs_registers_i/_2876_ ),
    .CLK(clknet_leaf_247_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[22]_reg  (.RESET_B(net2338),
    .D(\cs_registers_i/_0056_ ),
    .Q(crash_dump_o_22_),
    .Q_N(\cs_registers_i/_2875_ ),
    .CLK(clknet_leaf_247_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[23]_reg  (.RESET_B(net2397),
    .D(\cs_registers_i/_0057_ ),
    .Q(crash_dump_o_23_),
    .Q_N(\cs_registers_i/_2874_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[24]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0058_ ),
    .Q(crash_dump_o_24_),
    .Q_N(\cs_registers_i/_2873_ ),
    .CLK(clknet_leaf_265_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[25]_reg  (.RESET_B(net2429),
    .D(\cs_registers_i/_0059_ ),
    .Q(crash_dump_o_25_),
    .Q_N(\cs_registers_i/_2872_ ),
    .CLK(clknet_leaf_248_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[26]_reg  (.RESET_B(net2405),
    .D(\cs_registers_i/_0060_ ),
    .Q(crash_dump_o_26_),
    .Q_N(\cs_registers_i/_2871_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[27]_reg  (.RESET_B(net2403),
    .D(\cs_registers_i/_0061_ ),
    .Q(crash_dump_o_27_),
    .Q_N(\cs_registers_i/_2870_ ),
    .CLK(clknet_leaf_248_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[28]_reg  (.RESET_B(net2405),
    .D(\cs_registers_i/_0062_ ),
    .Q(crash_dump_o_28_),
    .Q_N(\cs_registers_i/_2869_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[29]_reg  (.RESET_B(net2421),
    .D(\cs_registers_i/_0063_ ),
    .Q(crash_dump_o_29_),
    .Q_N(\cs_registers_i/_2868_ ),
    .CLK(clknet_leaf_265_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[2]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0064_ ),
    .Q(crash_dump_o_2_),
    .Q_N(\cs_registers_i/_2867_ ),
    .CLK(clknet_leaf_263_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[30]_reg  (.RESET_B(net2404),
    .D(\cs_registers_i/_0065_ ),
    .Q(crash_dump_o_30_),
    .Q_N(\cs_registers_i/_2866_ ),
    .CLK(clknet_leaf_257_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[31]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0066_ ),
    .Q(crash_dump_o_31_),
    .Q_N(\cs_registers_i/_2865_ ),
    .CLK(clknet_leaf_264_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[3]_reg  (.RESET_B(net2323),
    .D(\cs_registers_i/_0067_ ),
    .Q(crash_dump_o_3_),
    .Q_N(\cs_registers_i/_2864_ ),
    .CLK(clknet_leaf_255_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[4]_reg  (.RESET_B(net2323),
    .D(\cs_registers_i/_0068_ ),
    .Q(crash_dump_o_4_),
    .Q_N(\cs_registers_i/_2863_ ),
    .CLK(clknet_leaf_254_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[5]_reg  (.RESET_B(net2397),
    .D(\cs_registers_i/_0069_ ),
    .Q(crash_dump_o_5_),
    .Q_N(\cs_registers_i/_2862_ ),
    .CLK(clknet_leaf_254_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[6]_reg  (.RESET_B(net2403),
    .D(\cs_registers_i/_0070_ ),
    .Q(crash_dump_o_6_),
    .Q_N(\cs_registers_i/_2861_ ),
    .CLK(clknet_leaf_257_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[7]_reg  (.RESET_B(net2403),
    .D(\cs_registers_i/_0071_ ),
    .Q(crash_dump_o_7_),
    .Q_N(\cs_registers_i/_2860_ ),
    .CLK(clknet_leaf_257_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[8]_reg  (.RESET_B(net2403),
    .D(\cs_registers_i/_0072_ ),
    .Q(crash_dump_o_8_),
    .Q_N(\cs_registers_i/_2859_ ),
    .CLK(clknet_leaf_257_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mepc_o[9]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0073_ ),
    .Q(crash_dump_o_9_),
    .Q_N(\cs_registers_i/_2858_ ),
    .CLK(clknet_leaf_263_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mstatus_mie_o_reg  (.RESET_B(net2375),
    .D(\cs_registers_i/_0074_ ),
    .Q(csr_mstatus_mie),
    .Q_N(\cs_registers_i/_2857_ ),
    .CLK(clknet_leaf_268_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mstatus_tw_o_reg  (.RESET_B(net2378),
    .D(\cs_registers_i/_0075_ ),
    .Q(csr_mstatus_tw),
    .Q_N(\cs_registers_i/_2856_ ),
    .CLK(clknet_leaf_275_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[0]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0076_ ),
    .Q_N(csr_mtvec_0_),
    .Q(\cs_registers_i/_0001_ ));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[10]_reg  (.RESET_B(net2420),
    .D(\cs_registers_i/_0077_ ),
    .Q(csr_mtvec_10_),
    .Q_N(\cs_registers_i/_2855_ ),
    .CLK(clknet_leaf_287_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[11]_reg  (.RESET_B(net2400),
    .D(\cs_registers_i/_0078_ ),
    .Q(csr_mtvec_11_),
    .Q_N(\cs_registers_i/_2854_ ),
    .CLK(clknet_leaf_228_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[12]_reg  (.RESET_B(net2417),
    .D(\cs_registers_i/_0079_ ),
    .Q(csr_mtvec_12_),
    .Q_N(\cs_registers_i/_2853_ ),
    .CLK(clknet_leaf_226_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[13]_reg  (.RESET_B(net2400),
    .D(\cs_registers_i/_0080_ ),
    .Q(csr_mtvec_13_),
    .Q_N(\cs_registers_i/_2852_ ),
    .CLK(clknet_leaf_228_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[14]_reg  (.RESET_B(net2400),
    .D(\cs_registers_i/_0081_ ),
    .Q(csr_mtvec_14_),
    .Q_N(\cs_registers_i/_2851_ ),
    .CLK(clknet_leaf_228_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[15]_reg  (.CLK(clknet_leaf_287_clk_i),
    .RESET_B(net2400),
    .D(\cs_registers_i/_0082_ ),
    .Q_N(\cs_registers_i/_2850_ ),
    .Q(csr_mtvec_15_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[16]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0083_ ),
    .Q(csr_mtvec_16_),
    .Q_N(\cs_registers_i/_2849_ ),
    .CLK(clknet_leaf_226_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[17]_reg  (.RESET_B(net2408),
    .D(\cs_registers_i/_0084_ ),
    .Q(csr_mtvec_17_),
    .Q_N(\cs_registers_i/_2848_ ),
    .CLK(clknet_leaf_220_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[18]_reg  (.RESET_B(net2418),
    .D(\cs_registers_i/_0085_ ),
    .Q(csr_mtvec_18_),
    .Q_N(\cs_registers_i/_2847_ ),
    .CLK(clknet_leaf_228_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[19]_reg  (.RESET_B(net2417),
    .D(\cs_registers_i/_0086_ ),
    .Q(csr_mtvec_19_),
    .Q_N(\cs_registers_i/_2846_ ),
    .CLK(clknet_leaf_225_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[1]_reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0087_ ),
    .Q_N(\cs_registers_i/_2845_ ),
    .Q(csr_mtvec_1_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[20]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0088_ ),
    .Q(csr_mtvec_20_),
    .Q_N(\cs_registers_i/_2844_ ),
    .CLK(clknet_leaf_224_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[21]_reg  (.RESET_B(net2408),
    .D(\cs_registers_i/_0089_ ),
    .Q(csr_mtvec_21_),
    .Q_N(\cs_registers_i/_2843_ ),
    .CLK(clknet_6_50_0_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[22]_reg  (.RESET_B(net2407),
    .D(\cs_registers_i/_0090_ ),
    .Q(csr_mtvec_22_),
    .Q_N(\cs_registers_i/_2842_ ),
    .CLK(clknet_leaf_224_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[23]_reg  (.RESET_B(net2416),
    .D(\cs_registers_i/_0091_ ),
    .Q(csr_mtvec_23_),
    .Q_N(\cs_registers_i/_2841_ ),
    .CLK(clknet_leaf_226_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[24]_reg  (.RESET_B(net2417),
    .D(\cs_registers_i/_0092_ ),
    .Q(csr_mtvec_24_),
    .Q_N(\cs_registers_i/_2840_ ),
    .CLK(clknet_leaf_224_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[25]_reg  (.CLK(clknet_leaf_292_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0093_ ),
    .Q_N(\cs_registers_i/_2839_ ),
    .Q(csr_mtvec_25_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[26]_reg  (.RESET_B(net2408),
    .D(\cs_registers_i/_0094_ ),
    .Q(csr_mtvec_26_),
    .Q_N(\cs_registers_i/_2838_ ),
    .CLK(clknet_leaf_220_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[27]_reg  (.RESET_B(net2406),
    .D(\cs_registers_i/_0095_ ),
    .Q(csr_mtvec_27_),
    .Q_N(\cs_registers_i/_2837_ ),
    .CLK(clknet_leaf_224_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[28]_reg  (.CLK(clknet_leaf_224_clk_i),
    .RESET_B(net2407),
    .D(\cs_registers_i/_0096_ ),
    .Q_N(\cs_registers_i/_2836_ ),
    .Q(csr_mtvec_28_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[29]_reg  (.CLK(clknet_leaf_224_clk_i),
    .RESET_B(net2407),
    .D(\cs_registers_i/_0097_ ),
    .Q_N(\cs_registers_i/_2835_ ),
    .Q(csr_mtvec_29_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[2]_reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0098_ ),
    .Q_N(\cs_registers_i/_2834_ ),
    .Q(csr_mtvec_2_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[30]_reg  (.RESET_B(net2401),
    .D(\cs_registers_i/_0099_ ),
    .Q(csr_mtvec_30_),
    .Q_N(\cs_registers_i/_2833_ ),
    .CLK(clknet_leaf_287_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[31]_reg  (.CLK(clknet_leaf_224_clk_i),
    .RESET_B(net2417),
    .D(\cs_registers_i/_0100_ ),
    .Q_N(\cs_registers_i/_2832_ ),
    .Q(csr_mtvec_31_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[3]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0101_ ),
    .Q_N(\cs_registers_i/_2831_ ),
    .Q(csr_mtvec_3_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[4]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0102_ ),
    .Q_N(\cs_registers_i/_2830_ ),
    .Q(csr_mtvec_4_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[5]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2411),
    .D(\cs_registers_i/_0103_ ),
    .Q_N(\cs_registers_i/_2829_ ),
    .Q(csr_mtvec_5_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[6]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0104_ ),
    .Q_N(\cs_registers_i/_2828_ ),
    .Q(csr_mtvec_6_));
 sg13g2_dfrbp_1 \cs_registers_i/csr_mtvec_o[7]_reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2411),
    .D(\cs_registers_i/_0105_ ),
    .Q_N(\cs_registers_i/_2827_ ),
    .Q(csr_mtvec_7_));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[8]_reg  (.RESET_B(net2401),
    .D(\cs_registers_i/_0106_ ),
    .Q(csr_mtvec_8_),
    .Q_N(\cs_registers_i/_2826_ ),
    .CLK(clknet_leaf_287_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/csr_mtvec_o[9]_reg  (.RESET_B(net2415),
    .D(\cs_registers_i/_0107_ ),
    .Q(csr_mtvec_9_),
    .Q_N(\cs_registers_i/_2825_ ),
    .CLK(clknet_leaf_226_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_0__reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0108_ ),
    .Q_N(\cs_registers_i/dcsr_q_0_ ),
    .Q(\cs_registers_i/_0002_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_10__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2373),
    .D(\cs_registers_i/_0109_ ),
    .Q_N(\cs_registers_i/_2824_ ),
    .Q(\cs_registers_i/dcsr_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_11__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0110_ ),
    .Q_N(\cs_registers_i/_2823_ ),
    .Q(\cs_registers_i/dcsr_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_13__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0111_ ),
    .Q_N(\cs_registers_i/_2822_ ),
    .Q(\cs_registers_i/dcsr_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_14__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0112_ ),
    .Q_N(\cs_registers_i/_2821_ ),
    .Q(\cs_registers_i/dcsr_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_16__reg  (.CLK(clknet_leaf_326_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0113_ ),
    .Q_N(\cs_registers_i/_2820_ ),
    .Q(\cs_registers_i/dcsr_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_17__reg  (.CLK(clknet_leaf_222_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0114_ ),
    .Q_N(\cs_registers_i/_2819_ ),
    .Q(\cs_registers_i/dcsr_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_18__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0115_ ),
    .Q_N(\cs_registers_i/_2818_ ),
    .Q(\cs_registers_i/dcsr_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_19__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0116_ ),
    .Q_N(\cs_registers_i/_2817_ ),
    .Q(\cs_registers_i/dcsr_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_1__reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2375),
    .D(\cs_registers_i/_0117_ ),
    .Q_N(\cs_registers_i/dcsr_q_1_ ),
    .Q(\cs_registers_i/_0003_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_20__reg  (.CLK(clknet_leaf_293_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0118_ ),
    .Q_N(\cs_registers_i/_2816_ ),
    .Q(\cs_registers_i/dcsr_q_20_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_21__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0119_ ),
    .Q_N(\cs_registers_i/_2815_ ),
    .Q(\cs_registers_i/dcsr_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_22__reg  (.CLK(clknet_leaf_290_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0120_ ),
    .Q_N(\cs_registers_i/_2814_ ),
    .Q(\cs_registers_i/dcsr_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_23__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0121_ ),
    .Q_N(\cs_registers_i/_2813_ ),
    .Q(\cs_registers_i/dcsr_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_24__reg  (.CLK(clknet_leaf_297_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0122_ ),
    .Q_N(\cs_registers_i/_2812_ ),
    .Q(\cs_registers_i/dcsr_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_25__reg  (.CLK(clknet_leaf_286_clk_i),
    .RESET_B(net2420),
    .D(\cs_registers_i/_0123_ ),
    .Q_N(\cs_registers_i/_2811_ ),
    .Q(\cs_registers_i/dcsr_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_26__reg  (.CLK(clknet_leaf_287_clk_i),
    .RESET_B(net2421),
    .D(\cs_registers_i/_0124_ ),
    .Q_N(\cs_registers_i/_2810_ ),
    .Q(\cs_registers_i/dcsr_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_27__reg  (.CLK(clknet_leaf_290_clk_i),
    .RESET_B(net2441),
    .D(\cs_registers_i/_0125_ ),
    .Q_N(\cs_registers_i/_2809_ ),
    .Q(\cs_registers_i/dcsr_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_28__reg  (.CLK(clknet_leaf_286_clk_i),
    .RESET_B(net2420),
    .D(\cs_registers_i/_0126_ ),
    .Q_N(\cs_registers_i/_2808_ ),
    .Q(\cs_registers_i/dcsr_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_29__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2421),
    .D(\cs_registers_i/_0127_ ),
    .Q_N(\cs_registers_i/_2807_ ),
    .Q(\cs_registers_i/dcsr_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_30__reg  (.CLK(clknet_leaf_278_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0128_ ),
    .Q_N(\cs_registers_i/dcsr_q_30_ ),
    .Q(\cs_registers_i/_0004_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_31__reg  (.CLK(clknet_leaf_223_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0129_ ),
    .Q_N(\cs_registers_i/_2806_ ),
    .Q(\cs_registers_i/dcsr_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_3__reg  (.CLK(clknet_leaf_321_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0130_ ),
    .Q_N(\cs_registers_i/_2805_ ),
    .Q(\cs_registers_i/dcsr_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_4__reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0131_ ),
    .Q_N(\cs_registers_i/_2804_ ),
    .Q(\cs_registers_i/dcsr_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_5__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0132_ ),
    .Q_N(\cs_registers_i/_2803_ ),
    .Q(\cs_registers_i/dcsr_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_6__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0133_ ),
    .Q_N(\cs_registers_i/_2802_ ),
    .Q(\cs_registers_i/dcsr_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_7__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0134_ ),
    .Q_N(\cs_registers_i/_2801_ ),
    .Q(\cs_registers_i/dcsr_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_8__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0135_ ),
    .Q_N(\cs_registers_i/_2800_ ),
    .Q(\cs_registers_i/dcsr_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dcsr_q_9__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2373),
    .D(\cs_registers_i/_0136_ ),
    .Q_N(\cs_registers_i/_2799_ ),
    .Q(\cs_registers_i/dcsr_q_9_ ));
 sg13g2_dfrbp_1 \cs_registers_i/debug_ebreakm_o_reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2373),
    .D(\cs_registers_i/_0137_ ),
    .Q_N(\cs_registers_i/_2798_ ),
    .Q(debug_ebreakm));
 sg13g2_dfrbp_1 \cs_registers_i/debug_ebreaku_o_reg  (.CLK(clknet_leaf_286_clk_i),
    .RESET_B(net2421),
    .D(\cs_registers_i/_0138_ ),
    .Q_N(\cs_registers_i/_2797_ ),
    .Q(debug_ebreaku));
 sg13g2_dfrbp_2 \cs_registers_i/debug_single_step_o_reg  (.RESET_B(net2443),
    .D(\cs_registers_i/_0139_ ),
    .Q(debug_single_step),
    .Q_N(\cs_registers_i/_2796_ ),
    .CLK(clknet_leaf_295_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_0__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0140_ ),
    .Q_N(\cs_registers_i/_2795_ ),
    .Q(\cs_registers_i/dscratch0_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_10__reg  (.CLK(clknet_leaf_326_clk_i),
    .RESET_B(net2374),
    .D(\cs_registers_i/_0141_ ),
    .Q_N(\cs_registers_i/_2794_ ),
    .Q(\cs_registers_i/dscratch0_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_11__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0142_ ),
    .Q_N(\cs_registers_i/_2793_ ),
    .Q(\cs_registers_i/dscratch0_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_12__reg  (.CLK(clknet_leaf_288_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0143_ ),
    .Q_N(\cs_registers_i/_2792_ ),
    .Q(\cs_registers_i/dscratch0_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_13__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0144_ ),
    .Q_N(\cs_registers_i/_2791_ ),
    .Q(\cs_registers_i/dscratch0_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_14__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0145_ ),
    .Q_N(\cs_registers_i/_2790_ ),
    .Q(\cs_registers_i/dscratch0_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_15__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2374),
    .D(\cs_registers_i/_0146_ ),
    .Q_N(\cs_registers_i/_2789_ ),
    .Q(\cs_registers_i/dscratch0_q_15_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_16__reg  (.CLK(clknet_leaf_326_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0147_ ),
    .Q_N(\cs_registers_i/_2788_ ),
    .Q(\cs_registers_i/dscratch0_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_17__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0148_ ),
    .Q_N(\cs_registers_i/_2787_ ),
    .Q(\cs_registers_i/dscratch0_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_18__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0149_ ),
    .Q_N(\cs_registers_i/_2786_ ),
    .Q(\cs_registers_i/dscratch0_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_19__reg  (.CLK(clknet_leaf_222_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0150_ ),
    .Q_N(\cs_registers_i/_2785_ ),
    .Q(\cs_registers_i/dscratch0_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_1__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0151_ ),
    .Q_N(\cs_registers_i/_2784_ ),
    .Q(\cs_registers_i/dscratch0_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_20__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0152_ ),
    .Q_N(\cs_registers_i/_2783_ ),
    .Q(\cs_registers_i/dscratch0_q_20_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_21__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0153_ ),
    .Q_N(\cs_registers_i/_2782_ ),
    .Q(\cs_registers_i/dscratch0_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_22__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0154_ ),
    .Q_N(\cs_registers_i/_2781_ ),
    .Q(\cs_registers_i/dscratch0_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_23__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0155_ ),
    .Q_N(\cs_registers_i/_2780_ ),
    .Q(\cs_registers_i/dscratch0_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_24__reg  (.CLK(clknet_leaf_297_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0156_ ),
    .Q_N(\cs_registers_i/_2779_ ),
    .Q(\cs_registers_i/dscratch0_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_25__reg  (.CLK(clknet_leaf_321_clk_i),
    .RESET_B(net2439),
    .D(\cs_registers_i/_0157_ ),
    .Q_N(\cs_registers_i/_2778_ ),
    .Q(\cs_registers_i/dscratch0_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_26__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0158_ ),
    .Q_N(\cs_registers_i/_2777_ ),
    .Q(\cs_registers_i/dscratch0_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_27__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2460),
    .D(\cs_registers_i/_0159_ ),
    .Q_N(\cs_registers_i/_2776_ ),
    .Q(\cs_registers_i/dscratch0_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_28__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0160_ ),
    .Q_N(\cs_registers_i/_2775_ ),
    .Q(\cs_registers_i/dscratch0_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_29__reg  (.CLK(clknet_leaf_303_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0161_ ),
    .Q_N(\cs_registers_i/_2774_ ),
    .Q(\cs_registers_i/dscratch0_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_2__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0162_ ),
    .Q_N(\cs_registers_i/_2773_ ),
    .Q(\cs_registers_i/dscratch0_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_30__reg  (.CLK(clknet_leaf_298_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0163_ ),
    .Q_N(\cs_registers_i/_2772_ ),
    .Q(\cs_registers_i/dscratch0_q_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_31__reg  (.CLK(clknet_leaf_223_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0164_ ),
    .Q_N(\cs_registers_i/_2771_ ),
    .Q(\cs_registers_i/dscratch0_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_3__reg  (.CLK(clknet_leaf_277_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0165_ ),
    .Q_N(\cs_registers_i/_2770_ ),
    .Q(\cs_registers_i/dscratch0_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_4__reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0166_ ),
    .Q_N(\cs_registers_i/_2769_ ),
    .Q(\cs_registers_i/dscratch0_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_5__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0167_ ),
    .Q_N(\cs_registers_i/_2768_ ),
    .Q(\cs_registers_i/dscratch0_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_6__reg  (.CLK(clknet_leaf_278_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0168_ ),
    .Q_N(\cs_registers_i/_2767_ ),
    .Q(\cs_registers_i/dscratch0_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_7__reg  (.CLK(clknet_leaf_298_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0169_ ),
    .Q_N(\cs_registers_i/_2766_ ),
    .Q(\cs_registers_i/dscratch0_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_8__reg  (.CLK(clknet_leaf_291_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0170_ ),
    .Q_N(\cs_registers_i/_2765_ ),
    .Q(\cs_registers_i/dscratch0_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch0_q_9__reg  (.CLK(clknet_leaf_326_clk_i),
    .RESET_B(net2374),
    .D(\cs_registers_i/_0171_ ),
    .Q_N(\cs_registers_i/_2764_ ),
    .Q(\cs_registers_i/dscratch0_q_9_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_0__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0172_ ),
    .Q_N(\cs_registers_i/_2763_ ),
    .Q(\cs_registers_i/dscratch1_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_10__reg  (.CLK(clknet_leaf_271_clk_i),
    .RESET_B(net2375),
    .D(\cs_registers_i/_0173_ ),
    .Q_N(\cs_registers_i/_2762_ ),
    .Q(\cs_registers_i/dscratch1_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_11__reg  (.CLK(clknet_leaf_298_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0174_ ),
    .Q_N(\cs_registers_i/_2761_ ),
    .Q(\cs_registers_i/dscratch1_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_12__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2422),
    .D(\cs_registers_i/_0175_ ),
    .Q_N(\cs_registers_i/_2760_ ),
    .Q(\cs_registers_i/dscratch1_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_13__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0176_ ),
    .Q_N(\cs_registers_i/_2759_ ),
    .Q(\cs_registers_i/dscratch1_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_14__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0177_ ),
    .Q_N(\cs_registers_i/_2758_ ),
    .Q(\cs_registers_i/dscratch1_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_15__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2375),
    .D(\cs_registers_i/_0178_ ),
    .Q_N(\cs_registers_i/_2757_ ),
    .Q(\cs_registers_i/dscratch1_q_15_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_16__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0179_ ),
    .Q_N(\cs_registers_i/_2756_ ),
    .Q(\cs_registers_i/dscratch1_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_17__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0180_ ),
    .Q_N(\cs_registers_i/_2755_ ),
    .Q(\cs_registers_i/dscratch1_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_18__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0181_ ),
    .Q_N(\cs_registers_i/_2754_ ),
    .Q(\cs_registers_i/dscratch1_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_19__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0182_ ),
    .Q_N(\cs_registers_i/_2753_ ),
    .Q(\cs_registers_i/dscratch1_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_1__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0183_ ),
    .Q_N(\cs_registers_i/_2752_ ),
    .Q(\cs_registers_i/dscratch1_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_20__reg  (.CLK(clknet_leaf_290_clk_i),
    .RESET_B(net2441),
    .D(\cs_registers_i/_0184_ ),
    .Q_N(\cs_registers_i/_2751_ ),
    .Q(\cs_registers_i/dscratch1_q_20_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_21__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2450),
    .D(\cs_registers_i/_0185_ ),
    .Q_N(\cs_registers_i/_2750_ ),
    .Q(\cs_registers_i/dscratch1_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_22__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net2449),
    .D(\cs_registers_i/_0186_ ),
    .Q_N(\cs_registers_i/_2749_ ),
    .Q(\cs_registers_i/dscratch1_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_23__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0187_ ),
    .Q_N(\cs_registers_i/_2748_ ),
    .Q(\cs_registers_i/dscratch1_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_24__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2450),
    .D(\cs_registers_i/_0188_ ),
    .Q_N(\cs_registers_i/_2747_ ),
    .Q(\cs_registers_i/dscratch1_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_25__reg  (.CLK(clknet_leaf_277_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0189_ ),
    .Q_N(\cs_registers_i/_2746_ ),
    .Q(\cs_registers_i/dscratch1_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_26__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0190_ ),
    .Q_N(\cs_registers_i/_2745_ ),
    .Q(\cs_registers_i/dscratch1_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_27__reg  (.CLK(clknet_leaf_296_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0191_ ),
    .Q_N(\cs_registers_i/_2744_ ),
    .Q(\cs_registers_i/dscratch1_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_28__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0192_ ),
    .Q_N(\cs_registers_i/_2743_ ),
    .Q(\cs_registers_i/dscratch1_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_29__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0193_ ),
    .Q_N(\cs_registers_i/_2742_ ),
    .Q(\cs_registers_i/dscratch1_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_2__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0194_ ),
    .Q_N(\cs_registers_i/_2741_ ),
    .Q(\cs_registers_i/dscratch1_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_30__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0195_ ),
    .Q_N(\cs_registers_i/_2740_ ),
    .Q(\cs_registers_i/dscratch1_q_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_31__reg  (.CLK(clknet_leaf_223_clk_i),
    .RESET_B(net2445),
    .D(\cs_registers_i/_0196_ ),
    .Q_N(\cs_registers_i/_2739_ ),
    .Q(\cs_registers_i/dscratch1_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_3__reg  (.CLK(clknet_leaf_276_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0197_ ),
    .Q_N(\cs_registers_i/_2738_ ),
    .Q(\cs_registers_i/dscratch1_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_4__reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0198_ ),
    .Q_N(\cs_registers_i/_2737_ ),
    .Q(\cs_registers_i/dscratch1_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_5__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0199_ ),
    .Q_N(\cs_registers_i/_2736_ ),
    .Q(\cs_registers_i/dscratch1_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_6__reg  (.CLK(clknet_leaf_278_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0200_ ),
    .Q_N(\cs_registers_i/_2735_ ),
    .Q(\cs_registers_i/dscratch1_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_7__reg  (.CLK(clknet_leaf_298_clk_i),
    .RESET_B(net2448),
    .D(\cs_registers_i/_0201_ ),
    .Q_N(\cs_registers_i/_2734_ ),
    .Q(\cs_registers_i/dscratch1_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_8__reg  (.CLK(clknet_leaf_289_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0202_ ),
    .Q_N(\cs_registers_i/_2733_ ),
    .Q(\cs_registers_i/dscratch1_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/dscratch1_q_9__reg  (.CLK(clknet_leaf_270_clk_i),
    .RESET_B(net2378),
    .D(\cs_registers_i/_0203_ ),
    .Q_N(\cs_registers_i/_2732_ ),
    .Q(\cs_registers_i/dscratch1_q_9_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcause_q_0__reg  (.RESET_B(net2395),
    .D(\cs_registers_i/_0204_ ),
    .Q(\cs_registers_i/mcause_q_0_ ),
    .Q_N(\cs_registers_i/_2731_ ),
    .CLK(clknet_leaf_259_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcause_q_1__reg  (.CLK(clknet_leaf_265_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0205_ ),
    .Q_N(\cs_registers_i/_2730_ ),
    .Q(\cs_registers_i/mcause_q_1_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcause_q_2__reg  (.RESET_B(net2399),
    .D(\cs_registers_i/_0206_ ),
    .Q(\cs_registers_i/mcause_q_2_ ),
    .Q_N(\cs_registers_i/_2729_ ),
    .CLK(clknet_leaf_263_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcause_q_3__reg  (.CLK(clknet_leaf_260_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0207_ ),
    .Q_N(\cs_registers_i/_2728_ ),
    .Q(\cs_registers_i/mcause_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcause_q_4__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2396),
    .D(\cs_registers_i/_0208_ ),
    .Q_N(\cs_registers_i/_2727_ ),
    .Q(\cs_registers_i/mcause_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcause_q_5__reg  (.CLK(clknet_leaf_259_clk_i),
    .RESET_B(net2396),
    .D(\cs_registers_i/_0209_ ),
    .Q_N(\cs_registers_i/_2726_ ),
    .Q(\cs_registers_i/mcause_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcause_q_6__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0210_ ),
    .Q_N(\cs_registers_i/_2725_ ),
    .Q(\cs_registers_i/mcause_q_6_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcountinhibit_0__reg  (.RESET_B(net2437),
    .D(\cs_registers_i/_0211_ ),
    .Q(\cs_registers_i/mcountinhibit_0_ ),
    .Q_N(\cs_registers_i/mcycle_counter_i.counter_inc_i ),
    .CLK(clknet_leaf_276_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcountinhibit_2__reg  (.CLK(clknet_leaf_277_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0212_ ),
    .Q_N(\cs_registers_i/minstret_counter_i.counter_inc_i_$_AND__Y_B ),
    .Q(\cs_registers_i/mcountinhibit_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_0__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0213_ ),
    .Q_N(\cs_registers_i/mcycle_counter_i.counter_upd_0_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_0_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_10__reg  (.RESET_B(net2439),
    .D(\cs_registers_i/_0214_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_10_ ),
    .Q_N(\cs_registers_i/_2724_ ),
    .CLK(clknet_leaf_321_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_11__reg  (.CLK(clknet_leaf_320_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0215_ ),
    .Q_N(\cs_registers_i/_2723_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_12__reg  (.CLK(clknet_leaf_320_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0216_ ),
    .Q_N(\cs_registers_i/_2722_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_13__reg  (.CLK(clknet_leaf_320_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0217_ ),
    .Q_N(\cs_registers_i/_2721_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_14__reg  (.CLK(clknet_leaf_319_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0218_ ),
    .Q_N(\cs_registers_i/_2720_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_15__reg  (.CLK(clknet_leaf_318_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0219_ ),
    .Q_N(\cs_registers_i/_2719_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_15_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_16__reg  (.RESET_B(net2458),
    .D(\cs_registers_i/_0220_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_16_ ),
    .Q_N(\cs_registers_i/_2718_ ),
    .CLK(clknet_leaf_298_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_17__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0221_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_17_ ),
    .Q_N(\cs_registers_i/_2717_ ),
    .CLK(clknet_leaf_299_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_18__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0222_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_18_ ),
    .Q_N(\cs_registers_i/_2716_ ),
    .CLK(clknet_leaf_299_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_19__reg  (.RESET_B(net2458),
    .D(\cs_registers_i/_0223_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_19_ ),
    .Q_N(\cs_registers_i/_2715_ ),
    .CLK(clknet_leaf_298_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_1__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0224_ ),
    .Q_N(\cs_registers_i/_2714_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_1_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_20__reg  (.RESET_B(net2460),
    .D(\cs_registers_i/_0225_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_20_ ),
    .Q_N(\cs_registers_i/_2713_ ),
    .CLK(clknet_leaf_301_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_21__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0226_ ),
    .Q_N(\cs_registers_i/_2712_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_22__reg  (.CLK(clknet_leaf_301_clk_i),
    .RESET_B(net2461),
    .D(\cs_registers_i/_0227_ ),
    .Q_N(\cs_registers_i/_2711_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_23__reg  (.CLK(clknet_leaf_302_clk_i),
    .RESET_B(net2454),
    .D(\cs_registers_i/_0228_ ),
    .Q_N(\cs_registers_i/_2710_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_23_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_24__reg  (.RESET_B(net2457),
    .D(\cs_registers_i/_0229_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_24_ ),
    .Q_N(\cs_registers_i/_2709_ ),
    .CLK(clknet_leaf_299_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_25__reg  (.RESET_B(net2457),
    .D(\cs_registers_i/_0230_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_25_ ),
    .Q_N(\cs_registers_i/_2708_ ),
    .CLK(clknet_leaf_299_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_26__reg  (.CLK(clknet_leaf_299_clk_i),
    .RESET_B(net2457),
    .D(\cs_registers_i/_0231_ ),
    .Q_N(\cs_registers_i/_2707_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_27__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2458),
    .D(\cs_registers_i/_0232_ ),
    .Q_N(\cs_registers_i/_2706_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_27_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_28__reg  (.RESET_B(net2454),
    .D(\cs_registers_i/_0233_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_28_ ),
    .Q_N(\cs_registers_i/_2705_ ),
    .CLK(clknet_leaf_318_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_29__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2457),
    .D(\cs_registers_i/_0234_ ),
    .Q_N(\cs_registers_i/_2704_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_2__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0235_ ),
    .Q_N(\cs_registers_i/_2703_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_30__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2458),
    .D(\cs_registers_i/_0236_ ),
    .Q_N(\cs_registers_i/_2702_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_31__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2458),
    .D(\cs_registers_i/_0237_ ),
    .Q_N(\cs_registers_i/_2701_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_32__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0238_ ),
    .Q_N(\cs_registers_i/_2700_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_32_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_33__reg  (.RESET_B(net2390),
    .D(\cs_registers_i/_0239_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_33_ ),
    .Q_N(\cs_registers_i/_2699_ ),
    .CLK(clknet_leaf_322_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_34__reg  (.RESET_B(net2390),
    .D(\cs_registers_i/_0240_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_34_ ),
    .Q_N(\cs_registers_i/_2698_ ),
    .CLK(clknet_leaf_322_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_35__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2387),
    .D(\cs_registers_i/_0241_ ),
    .Q_N(\cs_registers_i/_2697_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_35_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_36__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2388),
    .D(\cs_registers_i/_0242_ ),
    .Q_N(\cs_registers_i/_2696_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_36_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_37__reg  (.CLK(clknet_leaf_321_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0243_ ),
    .Q_N(\cs_registers_i/_2695_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_37_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_38__reg  (.CLK(clknet_leaf_322_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0244_ ),
    .Q_N(\cs_registers_i/_2694_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_38_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_39__reg  (.RESET_B(net2385),
    .D(\cs_registers_i/_0245_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_39_ ),
    .Q_N(\cs_registers_i/_2693_ ),
    .CLK(clknet_leaf_323_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_3__reg  (.CLK(clknet_leaf_325_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0246_ ),
    .Q_N(\cs_registers_i/_2692_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_3_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_40__reg  (.RESET_B(net2388),
    .D(\cs_registers_i/_0247_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_40_ ),
    .Q_N(\cs_registers_i/_2691_ ),
    .CLK(clknet_leaf_323_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_41__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0248_ ),
    .Q_N(\cs_registers_i/_2690_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_41_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_42__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2386),
    .D(\cs_registers_i/_0249_ ),
    .Q_N(\cs_registers_i/_2689_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_42_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_43__reg  (.CLK(clknet_leaf_316_clk_i),
    .RESET_B(net2390),
    .D(\cs_registers_i/_0250_ ),
    .Q_N(\cs_registers_i/_2688_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_43_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_44__reg  (.RESET_B(net2452),
    .D(\cs_registers_i/_0251_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_44_ ),
    .Q_N(\cs_registers_i/_2687_ ),
    .CLK(clknet_leaf_320_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_45__reg  (.CLK(clknet_leaf_316_clk_i),
    .RESET_B(net2390),
    .D(\cs_registers_i/_0252_ ),
    .Q_N(\cs_registers_i/_2686_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_45_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_46__reg  (.RESET_B(net2452),
    .D(\cs_registers_i/_0253_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_46_ ),
    .Q_N(\cs_registers_i/_2685_ ),
    .CLK(clknet_leaf_318_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_47__reg  (.CLK(clknet_leaf_316_clk_i),
    .RESET_B(net2390),
    .D(\cs_registers_i/_0254_ ),
    .Q_N(\cs_registers_i/_2684_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_47_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_48__reg  (.RESET_B(net2392),
    .D(\cs_registers_i/_0255_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_48_ ),
    .Q_N(\cs_registers_i/_2683_ ),
    .CLK(clknet_leaf_307_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_49__reg  (.RESET_B(net2392),
    .D(\cs_registers_i/_0256_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_49_ ),
    .Q_N(\cs_registers_i/_2682_ ),
    .CLK(clknet_leaf_300_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_4__reg  (.RESET_B(net2440),
    .D(\cs_registers_i/_0257_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_4_ ),
    .Q_N(\cs_registers_i/_2681_ ),
    .CLK(clknet_leaf_325_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_50__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2392),
    .D(\cs_registers_i/_0258_ ),
    .Q_N(\cs_registers_i/_2680_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_50_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_51__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2392),
    .D(\cs_registers_i/_0259_ ),
    .Q_N(\cs_registers_i/_2679_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_51_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_52__reg  (.CLK(clknet_leaf_317_clk_i),
    .RESET_B(net2390),
    .D(\cs_registers_i/_0260_ ),
    .Q_N(\cs_registers_i/_2678_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_52_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_53__reg  (.CLK(clknet_leaf_318_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0261_ ),
    .Q_N(\cs_registers_i/_2677_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_53_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_54__reg  (.CLK(clknet_leaf_318_clk_i),
    .RESET_B(net2452),
    .D(\cs_registers_i/_0262_ ),
    .Q_N(\cs_registers_i/_2676_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_54_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_55__reg  (.RESET_B(net2440),
    .D(\cs_registers_i/_0263_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_55_ ),
    .Q_N(\cs_registers_i/_2675_ ),
    .CLK(clknet_leaf_320_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_56__reg  (.CLK(clknet_leaf_306_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0264_ ),
    .Q_N(\cs_registers_i/_2674_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_56_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_57__reg  (.CLK(clknet_leaf_304_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0265_ ),
    .Q_N(\cs_registers_i/_2673_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_57_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_58__reg  (.CLK(clknet_leaf_304_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0266_ ),
    .Q_N(\cs_registers_i/_2672_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_58_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_59__reg  (.CLK(clknet_leaf_303_clk_i),
    .RESET_B(net2454),
    .D(\cs_registers_i/_0267_ ),
    .Q_N(\cs_registers_i/_2671_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_59_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_5__reg  (.RESET_B(net2439),
    .D(\cs_registers_i/_0268_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_5_ ),
    .Q_N(\cs_registers_i/_2670_ ),
    .CLK(clknet_leaf_325_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_60__reg  (.CLK(clknet_leaf_306_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0269_ ),
    .Q_N(\cs_registers_i/_2669_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_60_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_61__reg  (.CLK(clknet_leaf_304_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0270_ ),
    .Q_N(\cs_registers_i/_2668_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_61_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_62__reg  (.CLK(clknet_leaf_304_clk_i),
    .RESET_B(net2455),
    .D(\cs_registers_i/_0271_ ),
    .Q_N(\cs_registers_i/_2667_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_62_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_63__reg  (.CLK(clknet_leaf_303_clk_i),
    .RESET_B(net2454),
    .D(\cs_registers_i/_0272_ ),
    .Q_N(\cs_registers_i/_2666_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_63_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_6__reg  (.CLK(clknet_leaf_324_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0273_ ),
    .Q_N(\cs_registers_i/_2665_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_7__reg  (.CLK(clknet_leaf_324_clk_i),
    .RESET_B(net2439),
    .D(\cs_registers_i/_0274_ ),
    .Q_N(\cs_registers_i/_2664_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mcycle_counter_i.counter_val_o_8__reg  (.CLK(clknet_leaf_321_clk_i),
    .RESET_B(net2439),
    .D(\cs_registers_i/_0275_ ),
    .Q_N(\cs_registers_i/_2663_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_8_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mcycle_counter_i.counter_val_o_9__reg  (.RESET_B(net2453),
    .D(\cs_registers_i/_0276_ ),
    .Q(\cs_registers_i/mcycle_counter_i.counter_val_o_9_ ),
    .Q_N(\cs_registers_i/_2662_ ),
    .CLK(clknet_leaf_321_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1856__reg  (.CLK(clknet_leaf_327_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0277_ ),
    .Q_N(\cs_registers_i/minstret_counter_i.counter_val_upd_o_0_ ),
    .Q(\cs_registers_i/mhpmcounter_1856_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1857__reg  (.CLK(clknet_leaf_327_clk_i),
    .RESET_B(net2388),
    .D(\cs_registers_i/_0278_ ),
    .Q_N(\cs_registers_i/_2661_ ),
    .Q(\cs_registers_i/mhpmcounter_1857_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1858__reg  (.RESET_B(net2437),
    .D(\cs_registers_i/_0279_ ),
    .Q(\cs_registers_i/mhpmcounter_1858_ ),
    .Q_N(\cs_registers_i/_2660_ ),
    .CLK(clknet_leaf_327_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1859__reg  (.CLK(clknet_leaf_327_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0280_ ),
    .Q_N(\cs_registers_i/_2659_ ),
    .Q(\cs_registers_i/mhpmcounter_1859_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1860__reg  (.CLK(clknet_leaf_327_clk_i),
    .RESET_B(net2388),
    .D(\cs_registers_i/_0281_ ),
    .Q_N(\cs_registers_i/_2658_ ),
    .Q(\cs_registers_i/mhpmcounter_1860_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1861__reg  (.CLK(clknet_leaf_327_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0282_ ),
    .Q_N(\cs_registers_i/_2657_ ),
    .Q(\cs_registers_i/mhpmcounter_1861_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1862__reg  (.CLK(clknet_leaf_323_clk_i),
    .RESET_B(net2440),
    .D(\cs_registers_i/_0283_ ),
    .Q_N(\cs_registers_i/_2656_ ),
    .Q(\cs_registers_i/mhpmcounter_1862_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1863__reg  (.RESET_B(net2447),
    .D(\cs_registers_i/_0284_ ),
    .Q(\cs_registers_i/mhpmcounter_1863_ ),
    .Q_N(\cs_registers_i/_2655_ ),
    .CLK(clknet_leaf_324_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1864__reg  (.CLK(clknet_leaf_324_clk_i),
    .RESET_B(net2447),
    .D(\cs_registers_i/_0285_ ),
    .Q_N(\cs_registers_i/_2654_ ),
    .Q(\cs_registers_i/mhpmcounter_1864_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1865__reg  (.CLK(clknet_leaf_321_clk_i),
    .RESET_B(net2439),
    .D(\cs_registers_i/_0286_ ),
    .Q_N(\cs_registers_i/_2653_ ),
    .Q(\cs_registers_i/mhpmcounter_1865_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1866__reg  (.RESET_B(net2460),
    .D(\cs_registers_i/_0287_ ),
    .Q(\cs_registers_i/mhpmcounter_1866_ ),
    .Q_N(\cs_registers_i/_2652_ ),
    .CLK(clknet_leaf_319_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1867__reg  (.RESET_B(net2460),
    .D(\cs_registers_i/_0288_ ),
    .Q(\cs_registers_i/mhpmcounter_1867_ ),
    .Q_N(\cs_registers_i/_2651_ ),
    .CLK(clknet_leaf_319_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1868__reg  (.CLK(clknet_leaf_318_clk_i),
    .RESET_B(net2460),
    .D(\cs_registers_i/_0289_ ),
    .Q_N(\cs_registers_i/_2650_ ),
    .Q(\cs_registers_i/mhpmcounter_1868_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1869__reg  (.RESET_B(net2460),
    .D(\cs_registers_i/_0290_ ),
    .Q(\cs_registers_i/mhpmcounter_1869_ ),
    .Q_N(\cs_registers_i/_2649_ ),
    .CLK(clknet_leaf_303_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1870__reg  (.RESET_B(net2453),
    .D(\cs_registers_i/_0291_ ),
    .Q(\cs_registers_i/mhpmcounter_1870_ ),
    .Q_N(\cs_registers_i/_2648_ ),
    .CLK(clknet_leaf_303_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1871__reg  (.CLK(clknet_leaf_303_clk_i),
    .RESET_B(net2453),
    .D(\cs_registers_i/_0292_ ),
    .Q_N(\cs_registers_i/_2647_ ),
    .Q(\cs_registers_i/mhpmcounter_1871_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1872__reg  (.CLK(clknet_leaf_302_clk_i),
    .RESET_B(net2460),
    .D(\cs_registers_i/_0293_ ),
    .Q_N(\cs_registers_i/_2646_ ),
    .Q(\cs_registers_i/mhpmcounter_1872_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1873__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0294_ ),
    .Q(\cs_registers_i/mhpmcounter_1873_ ),
    .Q_N(\cs_registers_i/_2645_ ),
    .CLK(clknet_leaf_56_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1874__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0295_ ),
    .Q(\cs_registers_i/mhpmcounter_1874_ ),
    .Q_N(\cs_registers_i/_2644_ ),
    .CLK(clknet_leaf_297_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1875__reg  (.RESET_B(net2461),
    .D(\cs_registers_i/_0296_ ),
    .Q(\cs_registers_i/mhpmcounter_1875_ ),
    .Q_N(\cs_registers_i/_2643_ ),
    .CLK(clknet_leaf_297_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1876__reg  (.CLK(clknet_leaf_297_clk_i),
    .RESET_B(net2461),
    .D(\cs_registers_i/_0297_ ),
    .Q_N(\cs_registers_i/_2642_ ),
    .Q(\cs_registers_i/mhpmcounter_1876_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1877__reg  (.RESET_B(net2461),
    .D(\cs_registers_i/_0298_ ),
    .Q(\cs_registers_i/mhpmcounter_1877_ ),
    .Q_N(\cs_registers_i/_2641_ ),
    .CLK(clknet_leaf_56_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1878__reg  (.RESET_B(net2460),
    .D(\cs_registers_i/_0299_ ),
    .Q(\cs_registers_i/mhpmcounter_1878_ ),
    .Q_N(\cs_registers_i/_2640_ ),
    .CLK(clknet_leaf_297_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1879__reg  (.CLK(clknet_leaf_297_clk_i),
    .RESET_B(net2461),
    .D(\cs_registers_i/_0300_ ),
    .Q_N(\cs_registers_i/_2639_ ),
    .Q(\cs_registers_i/mhpmcounter_1879_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1880__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0301_ ),
    .Q(\cs_registers_i/mhpmcounter_1880_ ),
    .Q_N(\cs_registers_i/_2638_ ),
    .CLK(clknet_leaf_55_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1881__reg  (.RESET_B(net2462),
    .D(\cs_registers_i/_0302_ ),
    .Q(\cs_registers_i/mhpmcounter_1881_ ),
    .Q_N(\cs_registers_i/_2637_ ),
    .CLK(clknet_leaf_55_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1882__reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(net2463),
    .D(\cs_registers_i/_0303_ ),
    .Q_N(\cs_registers_i/_2636_ ),
    .Q(\cs_registers_i/mhpmcounter_1882_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1883__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net2463),
    .D(\cs_registers_i/_0304_ ),
    .Q_N(\cs_registers_i/_2635_ ),
    .Q(\cs_registers_i/mhpmcounter_1883_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1884__reg  (.RESET_B(net2457),
    .D(\cs_registers_i/_0305_ ),
    .Q(\cs_registers_i/mhpmcounter_1884_ ),
    .Q_N(\cs_registers_i/_2634_ ),
    .CLK(clknet_leaf_55_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1885__reg  (.RESET_B(net2457),
    .D(\cs_registers_i/_0306_ ),
    .Q(\cs_registers_i/mhpmcounter_1885_ ),
    .Q_N(\cs_registers_i/_2633_ ),
    .CLK(clknet_leaf_299_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1886__reg  (.RESET_B(net2457),
    .D(\cs_registers_i/_0307_ ),
    .Q(\cs_registers_i/mhpmcounter_1886_ ),
    .Q_N(\cs_registers_i/_2632_ ),
    .CLK(clknet_leaf_53_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1887__reg  (.CLK(clknet_leaf_299_clk_i),
    .RESET_B(net2457),
    .D(\cs_registers_i/_0308_ ),
    .Q_N(\cs_registers_i/_2631_ ),
    .Q(\cs_registers_i/mhpmcounter_1887_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1888__reg  (.RESET_B(net2391),
    .D(\cs_registers_i/_0309_ ),
    .Q(\cs_registers_i/mhpmcounter_1888_ ),
    .Q_N(\cs_registers_i/_2630_ ),
    .CLK(clknet_leaf_314_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1889__reg  (.CLK(clknet_leaf_314_clk_i),
    .RESET_B(net2387),
    .D(\cs_registers_i/_0310_ ),
    .Q_N(\cs_registers_i/_2629_ ),
    .Q(\cs_registers_i/mhpmcounter_1889_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1890__reg  (.CLK(clknet_leaf_315_clk_i),
    .RESET_B(net2388),
    .D(\cs_registers_i/_0311_ ),
    .Q_N(\cs_registers_i/_2628_ ),
    .Q(\cs_registers_i/mhpmcounter_1890_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1891__reg  (.CLK(clknet_leaf_328_clk_i),
    .RESET_B(net2388),
    .D(\cs_registers_i/_0312_ ),
    .Q_N(\cs_registers_i/_2627_ ),
    .Q(\cs_registers_i/mhpmcounter_1891_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1892__reg  (.RESET_B(net2388),
    .D(\cs_registers_i/_0313_ ),
    .Q(\cs_registers_i/mhpmcounter_1892_ ),
    .Q_N(\cs_registers_i/_2626_ ),
    .CLK(clknet_leaf_327_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1893__reg  (.RESET_B(net2387),
    .D(\cs_registers_i/_0314_ ),
    .Q(\cs_registers_i/mhpmcounter_1893_ ),
    .Q_N(\cs_registers_i/_2625_ ),
    .CLK(clknet_leaf_328_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1894__reg  (.RESET_B(net2387),
    .D(\cs_registers_i/_0315_ ),
    .Q(\cs_registers_i/mhpmcounter_1894_ ),
    .Q_N(\cs_registers_i/_2624_ ),
    .CLK(clknet_leaf_333_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1895__reg  (.RESET_B(net2387),
    .D(\cs_registers_i/_0316_ ),
    .Q(\cs_registers_i/mhpmcounter_1895_ ),
    .Q_N(\cs_registers_i/_2623_ ),
    .CLK(clknet_leaf_328_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1896__reg  (.RESET_B(net2387),
    .D(\cs_registers_i/_0317_ ),
    .Q(\cs_registers_i/mhpmcounter_1896_ ),
    .Q_N(\cs_registers_i/_2622_ ),
    .CLK(clknet_leaf_328_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1897__reg  (.CLK(clknet_leaf_328_clk_i),
    .RESET_B(net2387),
    .D(\cs_registers_i/_0318_ ),
    .Q_N(\cs_registers_i/_2621_ ),
    .Q(\cs_registers_i/mhpmcounter_1897_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1898__reg  (.CLK(clknet_leaf_328_clk_i),
    .RESET_B(net2387),
    .D(\cs_registers_i/_0319_ ),
    .Q_N(\cs_registers_i/_2620_ ),
    .Q(\cs_registers_i/mhpmcounter_1898_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1899__reg  (.RESET_B(net2390),
    .D(\cs_registers_i/_0320_ ),
    .Q(\cs_registers_i/mhpmcounter_1899_ ),
    .Q_N(\cs_registers_i/_2619_ ),
    .CLK(clknet_leaf_315_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1900__reg  (.RESET_B(net2391),
    .D(\cs_registers_i/_0321_ ),
    .Q(\cs_registers_i/mhpmcounter_1900_ ),
    .Q_N(\cs_registers_i/_2618_ ),
    .CLK(clknet_leaf_314_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1901__reg  (.RESET_B(net2391),
    .D(\cs_registers_i/_0322_ ),
    .Q(\cs_registers_i/mhpmcounter_1901_ ),
    .Q_N(\cs_registers_i/_2617_ ),
    .CLK(clknet_leaf_314_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1902__reg  (.RESET_B(net2391),
    .D(\cs_registers_i/_0323_ ),
    .Q(\cs_registers_i/mhpmcounter_1902_ ),
    .Q_N(\cs_registers_i/_2616_ ),
    .CLK(clknet_leaf_313_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1903__reg  (.CLK(clknet_leaf_313_clk_i),
    .RESET_B(net2391),
    .D(\cs_registers_i/_0324_ ),
    .Q_N(\cs_registers_i/_2615_ ),
    .Q(\cs_registers_i/mhpmcounter_1903_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1904__reg  (.RESET_B(net2392),
    .D(\cs_registers_i/_0325_ ),
    .Q(\cs_registers_i/mhpmcounter_1904_ ),
    .Q_N(\cs_registers_i/_2614_ ),
    .CLK(clknet_leaf_313_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1905__reg  (.RESET_B(net2392),
    .D(\cs_registers_i/_0326_ ),
    .Q(\cs_registers_i/mhpmcounter_1905_ ),
    .Q_N(\cs_registers_i/_2613_ ),
    .CLK(clknet_leaf_305_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1906__reg  (.RESET_B(net2392),
    .D(\cs_registers_i/_0327_ ),
    .Q(\cs_registers_i/mhpmcounter_1906_ ),
    .Q_N(\cs_registers_i/_2612_ ),
    .CLK(clknet_leaf_307_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1907__reg  (.CLK(clknet_leaf_317_clk_i),
    .RESET_B(net2392),
    .D(\cs_registers_i/_0328_ ),
    .Q_N(\cs_registers_i/_2611_ ),
    .Q(\cs_registers_i/mhpmcounter_1907_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1908__reg  (.CLK(clknet_leaf_313_clk_i),
    .RESET_B(net2391),
    .D(\cs_registers_i/_0329_ ),
    .Q_N(\cs_registers_i/_2610_ ),
    .Q(\cs_registers_i/mhpmcounter_1908_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1909__reg  (.CLK(clknet_leaf_316_clk_i),
    .RESET_B(net2390),
    .D(\cs_registers_i/_0330_ ),
    .Q_N(\cs_registers_i/_2609_ ),
    .Q(\cs_registers_i/mhpmcounter_1909_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1910__reg  (.CLK(clknet_leaf_313_clk_i),
    .RESET_B(net2391),
    .D(\cs_registers_i/_0331_ ),
    .Q_N(\cs_registers_i/_2608_ ),
    .Q(\cs_registers_i/mhpmcounter_1910_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1911__reg  (.RESET_B(net2455),
    .D(\cs_registers_i/_0332_ ),
    .Q(\cs_registers_i/mhpmcounter_1911_ ),
    .Q_N(\cs_registers_i/_2607_ ),
    .CLK(clknet_leaf_306_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1912__reg  (.RESET_B(net2455),
    .D(\cs_registers_i/_0333_ ),
    .Q(\cs_registers_i/mhpmcounter_1912_ ),
    .Q_N(\cs_registers_i/_2606_ ),
    .CLK(clknet_leaf_306_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1913__reg  (.RESET_B(net2456),
    .D(\cs_registers_i/_0334_ ),
    .Q(\cs_registers_i/mhpmcounter_1913_ ),
    .Q_N(\cs_registers_i/_2605_ ),
    .CLK(clknet_leaf_306_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1914__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2456),
    .D(\cs_registers_i/_0335_ ),
    .Q_N(\cs_registers_i/_2604_ ),
    .Q(\cs_registers_i/mhpmcounter_1914_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1915__reg  (.RESET_B(net2456),
    .D(\cs_registers_i/_0336_ ),
    .Q(\cs_registers_i/mhpmcounter_1915_ ),
    .Q_N(\cs_registers_i/_2603_ ),
    .CLK(clknet_leaf_308_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1916__reg  (.RESET_B(net2456),
    .D(\cs_registers_i/_0337_ ),
    .Q(\cs_registers_i/mhpmcounter_1916_ ),
    .Q_N(\cs_registers_i/_2602_ ),
    .CLK(clknet_leaf_305_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1917__reg  (.RESET_B(net2393),
    .D(\cs_registers_i/_0338_ ),
    .Q(\cs_registers_i/mhpmcounter_1917_ ),
    .Q_N(\cs_registers_i/_2601_ ),
    .CLK(clknet_leaf_305_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mhpmcounter_1918__reg  (.RESET_B(net2456),
    .D(\cs_registers_i/_0339_ ),
    .Q(\cs_registers_i/mhpmcounter_1918_ ),
    .Q_N(\cs_registers_i/_2600_ ),
    .CLK(clknet_leaf_306_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mhpmcounter_1919__reg  (.CLK(clknet_leaf_304_clk_i),
    .RESET_B(net2456),
    .D(\cs_registers_i/_0340_ ),
    .Q_N(\cs_registers_i/_2599_ ),
    .Q(\cs_registers_i/mhpmcounter_1919_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_0__reg  (.CLK(clknet_leaf_291_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0341_ ),
    .Q_N(\cs_registers_i/_2598_ ),
    .Q(\cs_registers_i/mie_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_10__reg  (.CLK(clknet_leaf_225_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0342_ ),
    .Q_N(\cs_registers_i/_2597_ ),
    .Q(\cs_registers_i/mie_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_11__reg  (.CLK(clknet_leaf_290_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0343_ ),
    .Q_N(\cs_registers_i/_2596_ ),
    .Q(\cs_registers_i/mie_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_12__reg  (.CLK(clknet_leaf_291_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0344_ ),
    .Q_N(\cs_registers_i/_2595_ ),
    .Q(\cs_registers_i/mie_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_13__reg  (.CLK(clknet_leaf_290_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0345_ ),
    .Q_N(\cs_registers_i/_2594_ ),
    .Q(\cs_registers_i/mie_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_14__reg  (.CLK(clknet_leaf_289_clk_i),
    .RESET_B(net2438),
    .D(\cs_registers_i/_0346_ ),
    .Q_N(\cs_registers_i/_2593_ ),
    .Q(\cs_registers_i/mie_q_14_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mie_q_15__reg  (.RESET_B(net2442),
    .D(\cs_registers_i/_0347_ ),
    .Q(\cs_registers_i/mie_q_15_ ),
    .Q_N(\cs_registers_i/_2592_ ),
    .CLK(clknet_leaf_291_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_16__reg  (.CLK(clknet_leaf_289_clk_i),
    .RESET_B(net2441),
    .D(\cs_registers_i/_0348_ ),
    .Q_N(\cs_registers_i/_2591_ ),
    .Q(\cs_registers_i/mie_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_17__reg  (.CLK(clknet_leaf_289_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0349_ ),
    .Q_N(\cs_registers_i/_2590_ ),
    .Q(\cs_registers_i/mie_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_18__reg  (.CLK(clknet_leaf_289_clk_i),
    .RESET_B(net2437),
    .D(\cs_registers_i/_0350_ ),
    .Q_N(\cs_registers_i/_2589_ ),
    .Q(\cs_registers_i/mie_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_1__reg  (.CLK(clknet_leaf_225_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0351_ ),
    .Q_N(\cs_registers_i/_2588_ ),
    .Q(\cs_registers_i/mie_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_2__reg  (.CLK(clknet_leaf_292_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0352_ ),
    .Q_N(\cs_registers_i/_2587_ ),
    .Q(\cs_registers_i/mie_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_3__reg  (.CLK(clknet_leaf_292_clk_i),
    .RESET_B(net2421),
    .D(\cs_registers_i/_0353_ ),
    .Q_N(\cs_registers_i/_2586_ ),
    .Q(\cs_registers_i/mie_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_4__reg  (.CLK(clknet_leaf_294_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0354_ ),
    .Q_N(\cs_registers_i/_2585_ ),
    .Q(\cs_registers_i/mie_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_5__reg  (.CLK(clknet_leaf_292_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0355_ ),
    .Q_N(\cs_registers_i/_2584_ ),
    .Q(\cs_registers_i/mie_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_6__reg  (.CLK(clknet_leaf_293_clk_i),
    .RESET_B(net2446),
    .D(\cs_registers_i/_0356_ ),
    .Q_N(\cs_registers_i/_2583_ ),
    .Q(\cs_registers_i/mie_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_7__reg  (.CLK(clknet_leaf_293_clk_i),
    .RESET_B(net2443),
    .D(\cs_registers_i/_0357_ ),
    .Q_N(\cs_registers_i/_2582_ ),
    .Q(\cs_registers_i/mie_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_8__reg  (.CLK(clknet_leaf_295_clk_i),
    .RESET_B(net2443),
    .D(\cs_registers_i/_0358_ ),
    .Q_N(\cs_registers_i/_2581_ ),
    .Q(\cs_registers_i/mie_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mie_q_9__reg  (.CLK(clknet_leaf_293_clk_i),
    .RESET_B(net2443),
    .D(\cs_registers_i/_0359_ ),
    .Q_N(\cs_registers_i/_2580_ ),
    .Q(\cs_registers_i/mie_q_9_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_0__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2411),
    .D(\cs_registers_i/_0360_ ),
    .Q_N(\cs_registers_i/_2579_ ),
    .Q(\cs_registers_i/mscratch_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_10__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0361_ ),
    .Q_N(\cs_registers_i/_2578_ ),
    .Q(\cs_registers_i/mscratch_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_11__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0362_ ),
    .Q_N(\cs_registers_i/_2577_ ),
    .Q(\cs_registers_i/mscratch_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_12__reg  (.CLK(clknet_leaf_288_clk_i),
    .RESET_B(net2421),
    .D(\cs_registers_i/_0363_ ),
    .Q_N(\cs_registers_i/_2576_ ),
    .Q(\cs_registers_i/mscratch_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_13__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0364_ ),
    .Q_N(\cs_registers_i/_2575_ ),
    .Q(\cs_registers_i/mscratch_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_14__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0365_ ),
    .Q_N(\cs_registers_i/_2574_ ),
    .Q(\cs_registers_i/mscratch_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_15__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0366_ ),
    .Q_N(\cs_registers_i/_2573_ ),
    .Q(\cs_registers_i/mscratch_q_15_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_16__reg  (.CLK(clknet_leaf_280_clk_i),
    .RESET_B(net2442),
    .D(\cs_registers_i/_0367_ ),
    .Q_N(\cs_registers_i/_2572_ ),
    .Q(\cs_registers_i/mscratch_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_17__reg  (.CLK(clknet_leaf_288_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0368_ ),
    .Q_N(\cs_registers_i/_2571_ ),
    .Q(\cs_registers_i/mscratch_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_18__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0369_ ),
    .Q_N(\cs_registers_i/_2570_ ),
    .Q(\cs_registers_i/mscratch_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_19__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0370_ ),
    .Q_N(\cs_registers_i/_2569_ ),
    .Q(\cs_registers_i/mscratch_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_1__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2373),
    .D(\cs_registers_i/_0371_ ),
    .Q_N(\cs_registers_i/_2568_ ),
    .Q(\cs_registers_i/mscratch_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_20__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0372_ ),
    .Q_N(\cs_registers_i/_2567_ ),
    .Q(\cs_registers_i/mscratch_q_20_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_21__reg  (.CLK(clknet_leaf_288_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0373_ ),
    .Q_N(\cs_registers_i/_2566_ ),
    .Q(\cs_registers_i/mscratch_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_22__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2379),
    .D(\cs_registers_i/_0374_ ),
    .Q_N(\cs_registers_i/_2565_ ),
    .Q(\cs_registers_i/mscratch_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_23__reg  (.CLK(clknet_leaf_272_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0375_ ),
    .Q_N(\cs_registers_i/_2564_ ),
    .Q(\cs_registers_i/mscratch_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_24__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0376_ ),
    .Q_N(\cs_registers_i/_2563_ ),
    .Q(\cs_registers_i/mscratch_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_25__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0377_ ),
    .Q_N(\cs_registers_i/_2562_ ),
    .Q(\cs_registers_i/mscratch_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_26__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0378_ ),
    .Q_N(\cs_registers_i/_2561_ ),
    .Q(\cs_registers_i/mscratch_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_27__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0379_ ),
    .Q_N(\cs_registers_i/_2560_ ),
    .Q(\cs_registers_i/mscratch_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_28__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0380_ ),
    .Q_N(\cs_registers_i/_2559_ ),
    .Q(\cs_registers_i/mscratch_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_29__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2380),
    .D(\cs_registers_i/_0381_ ),
    .Q_N(\cs_registers_i/_2558_ ),
    .Q(\cs_registers_i/mscratch_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_2__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2384),
    .D(\cs_registers_i/_0382_ ),
    .Q_N(\cs_registers_i/_2557_ ),
    .Q(\cs_registers_i/mscratch_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_30__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2444),
    .D(\cs_registers_i/_0383_ ),
    .Q_N(\cs_registers_i/_2556_ ),
    .Q(\cs_registers_i/mscratch_q_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_31__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0384_ ),
    .Q_N(\cs_registers_i/_2555_ ),
    .Q(\cs_registers_i/mscratch_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_3__reg  (.CLK(clknet_leaf_263_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0385_ ),
    .Q_N(\cs_registers_i/_2554_ ),
    .Q(\cs_registers_i/mscratch_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_4__reg  (.CLK(clknet_leaf_261_clk_i),
    .RESET_B(net2360),
    .D(\cs_registers_i/_0386_ ),
    .Q_N(\cs_registers_i/_2553_ ),
    .Q(\cs_registers_i/mscratch_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_5__reg  (.CLK(clknet_leaf_260_clk_i),
    .RESET_B(net2360),
    .D(\cs_registers_i/_0387_ ),
    .Q_N(\cs_registers_i/_2552_ ),
    .Q(\cs_registers_i/mscratch_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_6__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2373),
    .D(\cs_registers_i/_0388_ ),
    .Q_N(\cs_registers_i/_2551_ ),
    .Q(\cs_registers_i/mscratch_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_7__reg  (.CLK(clknet_leaf_273_clk_i),
    .RESET_B(net2385),
    .D(\cs_registers_i/_0389_ ),
    .Q_N(\cs_registers_i/_2550_ ),
    .Q(\cs_registers_i/mscratch_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_8__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0390_ ),
    .Q_N(\cs_registers_i/_2549_ ),
    .Q(\cs_registers_i/mscratch_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mscratch_q_9__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0391_ ),
    .Q_N(\cs_registers_i/_2548_ ),
    .Q(\cs_registers_i/mscratch_q_9_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_0__reg  (.CLK(clknet_leaf_259_clk_i),
    .RESET_B(net2396),
    .D(\cs_registers_i/_0392_ ),
    .Q_N(\cs_registers_i/_2547_ ),
    .Q(\cs_registers_i/mstack_cause_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_1__reg  (.CLK(clknet_leaf_263_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0393_ ),
    .Q_N(\cs_registers_i/_2546_ ),
    .Q(\cs_registers_i/mstack_cause_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_2__reg  (.CLK(clknet_leaf_263_clk_i),
    .RESET_B(net2399),
    .D(\cs_registers_i/_0394_ ),
    .Q_N(\cs_registers_i/_2545_ ),
    .Q(\cs_registers_i/mstack_cause_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_3__reg  (.CLK(clknet_leaf_260_clk_i),
    .RESET_B(net2400),
    .D(\cs_registers_i/_0395_ ),
    .Q_N(\cs_registers_i/_2544_ ),
    .Q(\cs_registers_i/mstack_cause_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_4__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2396),
    .D(\cs_registers_i/_0396_ ),
    .Q_N(\cs_registers_i/_2543_ ),
    .Q(\cs_registers_i/mstack_cause_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_5__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2396),
    .D(\cs_registers_i/_0397_ ),
    .Q_N(\cs_registers_i/_2542_ ),
    .Q(\cs_registers_i/mstack_cause_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_cause_q_6__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0398_ ),
    .Q_N(\cs_registers_i/_2541_ ),
    .Q(\cs_registers_i/mstack_cause_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_0__reg  (.CLK(clknet_leaf_254_clk_i),
    .RESET_B(net2323),
    .D(\cs_registers_i/_0399_ ),
    .Q_N(\cs_registers_i/_2540_ ),
    .Q(\cs_registers_i/mstack_epc_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_10__reg  (.CLK(clknet_leaf_266_clk_i),
    .RESET_B(net2435),
    .D(\cs_registers_i/_0400_ ),
    .Q_N(\cs_registers_i/_2539_ ),
    .Q(\cs_registers_i/mstack_epc_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_11__reg  (.CLK(clknet_leaf_264_clk_i),
    .RESET_B(net2400),
    .D(\cs_registers_i/_0401_ ),
    .Q_N(\cs_registers_i/_2538_ ),
    .Q(\cs_registers_i/mstack_epc_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_12__reg  (.CLK(clknet_leaf_266_clk_i),
    .RESET_B(net2420),
    .D(\cs_registers_i/_0402_ ),
    .Q_N(\cs_registers_i/_2537_ ),
    .Q(\cs_registers_i/mstack_epc_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_13__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2401),
    .D(\cs_registers_i/_0403_ ),
    .Q_N(\cs_registers_i/_2536_ ),
    .Q(\cs_registers_i/mstack_epc_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_14__reg  (.CLK(clknet_leaf_253_clk_i),
    .RESET_B(net2398),
    .D(\cs_registers_i/_0404_ ),
    .Q_N(\cs_registers_i/_2535_ ),
    .Q(\cs_registers_i/mstack_epc_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_15__reg  (.CLK(clknet_leaf_253_clk_i),
    .RESET_B(net2397),
    .D(\cs_registers_i/_0405_ ),
    .Q_N(\cs_registers_i/_2534_ ),
    .Q(\cs_registers_i/mstack_epc_q_15_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_16__reg  (.CLK(clknet_leaf_257_clk_i),
    .RESET_B(net2405),
    .D(\cs_registers_i/_0406_ ),
    .Q_N(\cs_registers_i/_2533_ ),
    .Q(\cs_registers_i/mstack_epc_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_17__reg  (.CLK(clknet_leaf_249_clk_i),
    .RESET_B(net2405),
    .D(\cs_registers_i/_0407_ ),
    .Q_N(\cs_registers_i/_2532_ ),
    .Q(\cs_registers_i/mstack_epc_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_18__reg  (.CLK(clknet_leaf_266_clk_i),
    .RESET_B(net2420),
    .D(\cs_registers_i/_0408_ ),
    .Q_N(\cs_registers_i/_2531_ ),
    .Q(\cs_registers_i/mstack_epc_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_19__reg  (.CLK(clknet_leaf_249_clk_i),
    .RESET_B(net2405),
    .D(\cs_registers_i/_0409_ ),
    .Q_N(\cs_registers_i/_2530_ ),
    .Q(\cs_registers_i/mstack_epc_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_1__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2402),
    .D(\cs_registers_i/_0410_ ),
    .Q_N(\cs_registers_i/_2529_ ),
    .Q(\cs_registers_i/mstack_epc_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_20__reg  (.CLK(clknet_leaf_249_clk_i),
    .RESET_B(net2338),
    .D(\cs_registers_i/_0411_ ),
    .Q_N(\cs_registers_i/_2528_ ),
    .Q(\cs_registers_i/mstack_epc_q_20_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_21__reg  (.CLK(clknet_leaf_249_clk_i),
    .RESET_B(net2429),
    .D(\cs_registers_i/_0412_ ),
    .Q_N(\cs_registers_i/_2527_ ),
    .Q(\cs_registers_i/mstack_epc_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_22__reg  (.CLK(clknet_leaf_247_clk_i),
    .RESET_B(net2338),
    .D(\cs_registers_i/_0413_ ),
    .Q_N(\cs_registers_i/_2526_ ),
    .Q(\cs_registers_i/mstack_epc_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_23__reg  (.CLK(clknet_leaf_255_clk_i),
    .RESET_B(net2323),
    .D(\cs_registers_i/_0414_ ),
    .Q_N(\cs_registers_i/_2525_ ),
    .Q(\cs_registers_i/mstack_epc_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_24__reg  (.CLK(clknet_leaf_265_clk_i),
    .RESET_B(net2435),
    .D(\cs_registers_i/_0415_ ),
    .Q_N(\cs_registers_i/_2524_ ),
    .Q(\cs_registers_i/mstack_epc_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_25__reg  (.CLK(clknet_leaf_247_clk_i),
    .RESET_B(net2429),
    .D(\cs_registers_i/_0416_ ),
    .Q_N(\cs_registers_i/_2523_ ),
    .Q(\cs_registers_i/mstack_epc_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_26__reg  (.CLK(clknet_leaf_248_clk_i),
    .RESET_B(net2404),
    .D(\cs_registers_i/_0417_ ),
    .Q_N(\cs_registers_i/_2522_ ),
    .Q(\cs_registers_i/mstack_epc_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_27__reg  (.CLK(clknet_leaf_248_clk_i),
    .RESET_B(net2403),
    .D(\cs_registers_i/_0418_ ),
    .Q_N(\cs_registers_i/_2521_ ),
    .Q(\cs_registers_i/mstack_epc_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_28__reg  (.CLK(clknet_leaf_248_clk_i),
    .RESET_B(net2429),
    .D(\cs_registers_i/_0419_ ),
    .Q_N(\cs_registers_i/_2520_ ),
    .Q(\cs_registers_i/mstack_epc_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_29__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2422),
    .D(\cs_registers_i/_0420_ ),
    .Q_N(\cs_registers_i/_2519_ ),
    .Q(\cs_registers_i/mstack_epc_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_2__reg  (.CLK(clknet_leaf_262_clk_i),
    .RESET_B(net2416),
    .D(\cs_registers_i/_0421_ ),
    .Q_N(\cs_registers_i/_2518_ ),
    .Q(\cs_registers_i/mstack_epc_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_30__reg  (.CLK(clknet_leaf_248_clk_i),
    .RESET_B(net2429),
    .D(\cs_registers_i/_0422_ ),
    .Q_N(\cs_registers_i/_2517_ ),
    .Q(\cs_registers_i/mstack_epc_q_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_31__reg  (.CLK(clknet_leaf_265_clk_i),
    .RESET_B(net2418),
    .D(\cs_registers_i/_0423_ ),
    .Q_N(\cs_registers_i/_2516_ ),
    .Q(\cs_registers_i/mstack_epc_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_3__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2397),
    .D(\cs_registers_i/_0424_ ),
    .Q_N(\cs_registers_i/_2515_ ),
    .Q(\cs_registers_i/mstack_epc_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_4__reg  (.CLK(clknet_leaf_253_clk_i),
    .RESET_B(net2395),
    .D(\cs_registers_i/_0425_ ),
    .Q_N(\cs_registers_i/_2514_ ),
    .Q(\cs_registers_i/mstack_epc_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_5__reg  (.CLK(clknet_leaf_253_clk_i),
    .RESET_B(net2395),
    .D(\cs_registers_i/_0426_ ),
    .Q_N(\cs_registers_i/_2513_ ),
    .Q(\cs_registers_i/mstack_epc_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_6__reg  (.CLK(clknet_leaf_257_clk_i),
    .RESET_B(net2403),
    .D(\cs_registers_i/_0427_ ),
    .Q_N(\cs_registers_i/_2512_ ),
    .Q(\cs_registers_i/mstack_epc_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_7__reg  (.CLK(clknet_6_56_0_clk_i),
    .RESET_B(net2403),
    .D(\cs_registers_i/_0428_ ),
    .Q_N(\cs_registers_i/_2511_ ),
    .Q(\cs_registers_i/mstack_epc_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_8__reg  (.CLK(clknet_leaf_258_clk_i),
    .RESET_B(net2409),
    .D(\cs_registers_i/_0429_ ),
    .Q_N(\cs_registers_i/_2510_ ),
    .Q(\cs_registers_i/mstack_epc_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_epc_q_9__reg  (.CLK(clknet_leaf_262_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0430_ ),
    .Q_N(\cs_registers_i/_2509_ ),
    .Q(\cs_registers_i/mstack_epc_q_9_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_q_0__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2376),
    .D(\cs_registers_i/_0431_ ),
    .Q_N(\cs_registers_i/_2508_ ),
    .Q(\cs_registers_i/mstack_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_q_1__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2376),
    .D(\cs_registers_i/_0432_ ),
    .Q_N(\cs_registers_i/_2507_ ),
    .Q(\cs_registers_i/mstack_q_1_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstack_q_2__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2375),
    .D(\cs_registers_i/_0433_ ),
    .Q_N(\cs_registers_i/mstack_q_2_ ),
    .Q(\cs_registers_i/_0005_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mstatus_q_1__reg  (.CLK(clknet_leaf_269_clk_i),
    .RESET_B(net2411),
    .D(\cs_registers_i/_0434_ ),
    .Q_N(\cs_registers_i/_2506_ ),
    .Q(\cs_registers_i/mstatus_q_1_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mstatus_q_2__reg  (.RESET_B(net2376),
    .D(\cs_registers_i/_0435_ ),
    .Q(\cs_registers_i/_0006_ ),
    .Q_N(\cs_registers_i/mstatus_q_2_ ),
    .CLK(clknet_leaf_269_clk_i));
 sg13g2_dfrbp_2 \cs_registers_i/mstatus_q_3__reg  (.RESET_B(net2376),
    .D(\cs_registers_i/_0436_ ),
    .Q(\cs_registers_i/_0007_ ),
    .Q_N(\cs_registers_i/mstatus_q_3_ ),
    .CLK(clknet_leaf_269_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mstatus_q_4__reg  (.CLK(clknet_leaf_268_clk_i),
    .RESET_B(net2375),
    .D(\cs_registers_i/_0437_ ),
    .Q_N(\cs_registers_i/_0000_ ),
    .Q(\cs_registers_i/mstatus_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_0__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0438_ ),
    .Q_N(\cs_registers_i/_2505_ ),
    .Q(\cs_registers_i/mtval_q_0_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_10__reg  (.CLK(clknet_leaf_261_clk_i),
    .RESET_B(net2401),
    .D(\cs_registers_i/_0439_ ),
    .Q_N(\cs_registers_i/_2504_ ),
    .Q(\cs_registers_i/mtval_q_10_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_11__reg  (.CLK(clknet_leaf_280_clk_i),
    .RESET_B(net2413),
    .D(\cs_registers_i/_0440_ ),
    .Q_N(\cs_registers_i/_2503_ ),
    .Q(\cs_registers_i/mtval_q_11_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_12__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0441_ ),
    .Q_N(\cs_registers_i/_2502_ ),
    .Q(\cs_registers_i/mtval_q_12_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_13__reg  (.CLK(clknet_leaf_282_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0442_ ),
    .Q_N(\cs_registers_i/_2501_ ),
    .Q(\cs_registers_i/mtval_q_13_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_14__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0443_ ),
    .Q_N(\cs_registers_i/_2500_ ),
    .Q(\cs_registers_i/mtval_q_14_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_15__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0444_ ),
    .Q_N(\cs_registers_i/_2499_ ),
    .Q(\cs_registers_i/mtval_q_15_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_16__reg  (.CLK(clknet_leaf_259_clk_i),
    .RESET_B(net2415),
    .D(\cs_registers_i/_0445_ ),
    .Q_N(\cs_registers_i/_2498_ ),
    .Q(\cs_registers_i/mtval_q_16_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_17__reg  (.CLK(clknet_leaf_282_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0446_ ),
    .Q_N(\cs_registers_i/_2497_ ),
    .Q(\cs_registers_i/mtval_q_17_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_18__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2419),
    .D(\cs_registers_i/_0447_ ),
    .Q_N(\cs_registers_i/_2496_ ),
    .Q(\cs_registers_i/mtval_q_18_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_19__reg  (.CLK(clknet_leaf_280_clk_i),
    .RESET_B(net2413),
    .D(\cs_registers_i/_0448_ ),
    .Q_N(\cs_registers_i/_2495_ ),
    .Q(\cs_registers_i/mtval_q_19_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_1__reg  (.CLK(clknet_leaf_267_clk_i),
    .RESET_B(net2402),
    .D(\cs_registers_i/_0449_ ),
    .Q_N(\cs_registers_i/_2494_ ),
    .Q(\cs_registers_i/mtval_q_1_ ));
 sg13g2_dfrbp_2 \cs_registers_i/mtval_q_20__reg  (.RESET_B(net2323),
    .D(\cs_registers_i/_0450_ ),
    .Q(\cs_registers_i/mtval_q_20_ ),
    .Q_N(\cs_registers_i/_2493_ ),
    .CLK(clknet_leaf_257_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_21__reg  (.CLK(clknet_leaf_279_clk_i),
    .RESET_B(net2414),
    .D(\cs_registers_i/_0451_ ),
    .Q_N(\cs_registers_i/_2492_ ),
    .Q(\cs_registers_i/mtval_q_21_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_22__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2424),
    .D(\cs_registers_i/_0452_ ),
    .Q_N(\cs_registers_i/_2491_ ),
    .Q(\cs_registers_i/mtval_q_22_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_23__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2413),
    .D(\cs_registers_i/_0453_ ),
    .Q_N(\cs_registers_i/_2490_ ),
    .Q(\cs_registers_i/mtval_q_23_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_24__reg  (.CLK(clknet_leaf_257_clk_i),
    .RESET_B(net2397),
    .D(\cs_registers_i/_0454_ ),
    .Q_N(\cs_registers_i/_2489_ ),
    .Q(\cs_registers_i/mtval_q_24_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_25__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2419),
    .D(\cs_registers_i/_0455_ ),
    .Q_N(\cs_registers_i/_2488_ ),
    .Q(\cs_registers_i/mtval_q_25_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_26__reg  (.CLK(clknet_leaf_283_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0456_ ),
    .Q_N(\cs_registers_i/_2487_ ),
    .Q(\cs_registers_i/mtval_q_26_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_27__reg  (.CLK(clknet_leaf_282_clk_i),
    .RESET_B(net2423),
    .D(\cs_registers_i/_0457_ ),
    .Q_N(\cs_registers_i/_2486_ ),
    .Q(\cs_registers_i/mtval_q_27_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_28__reg  (.CLK(clknet_leaf_284_clk_i),
    .RESET_B(net2415),
    .D(\cs_registers_i/_0458_ ),
    .Q_N(\cs_registers_i/_2485_ ),
    .Q(\cs_registers_i/mtval_q_28_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_29__reg  (.CLK(clknet_leaf_281_clk_i),
    .RESET_B(net2401),
    .D(\cs_registers_i/_0459_ ),
    .Q_N(\cs_registers_i/_2484_ ),
    .Q(\cs_registers_i/mtval_q_29_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_2__reg  (.CLK(clknet_leaf_262_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0460_ ),
    .Q_N(\cs_registers_i/_2483_ ),
    .Q(\cs_registers_i/mtval_q_2_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_30__reg  (.CLK(clknet_leaf_282_clk_i),
    .RESET_B(net2412),
    .D(\cs_registers_i/_0461_ ),
    .Q_N(\cs_registers_i/_2482_ ),
    .Q(\cs_registers_i/mtval_q_30_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_31__reg  (.CLK(clknet_leaf_255_clk_i),
    .RESET_B(net2323),
    .D(\cs_registers_i/_0462_ ),
    .Q_N(\cs_registers_i/_2481_ ),
    .Q(\cs_registers_i/mtval_q_31_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_3__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2395),
    .D(\cs_registers_i/_0463_ ),
    .Q_N(\cs_registers_i/_2480_ ),
    .Q(\cs_registers_i/mtval_q_3_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_4__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2395),
    .D(\cs_registers_i/_0464_ ),
    .Q_N(\cs_registers_i/_2479_ ),
    .Q(\cs_registers_i/mtval_q_4_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_5__reg  (.CLK(clknet_leaf_256_clk_i),
    .RESET_B(net2395),
    .D(\cs_registers_i/_0465_ ),
    .Q_N(\cs_registers_i/_2478_ ),
    .Q(\cs_registers_i/mtval_q_5_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_6__reg  (.CLK(clknet_leaf_261_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0466_ ),
    .Q_N(\cs_registers_i/_2477_ ),
    .Q(\cs_registers_i/mtval_q_6_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_7__reg  (.CLK(clknet_leaf_275_clk_i),
    .RESET_B(net2411),
    .D(\cs_registers_i/_0467_ ),
    .Q_N(\cs_registers_i/_2476_ ),
    .Q(\cs_registers_i/mtval_q_7_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_8__reg  (.CLK(clknet_leaf_261_clk_i),
    .RESET_B(net2401),
    .D(\cs_registers_i/_0468_ ),
    .Q_N(\cs_registers_i/_2475_ ),
    .Q(\cs_registers_i/mtval_q_8_ ));
 sg13g2_dfrbp_1 \cs_registers_i/mtval_q_9__reg  (.CLK(clknet_leaf_262_clk_i),
    .RESET_B(net2402),
    .D(\cs_registers_i/_0469_ ),
    .Q_N(\cs_registers_i/_2474_ ),
    .Q(\cs_registers_i/mtval_q_9_ ));
 sg13g2_dfrbp_2 \cs_registers_i/priv_mode_id_o[0]_reg  (.RESET_B(net2375),
    .D(\cs_registers_i/_0470_ ),
    .Q(\cs_registers_i/_0008_ ),
    .Q_N(\id_stage_i.controller_i.priv_mode_i_0_ ),
    .CLK(clknet_leaf_274_clk_i));
 sg13g2_dfrbp_1 \cs_registers_i/priv_mode_id_o[1]_reg  (.CLK(clknet_leaf_274_clk_i),
    .RESET_B(net2410),
    .D(\cs_registers_i/_0471_ ),
    .Q_N(\id_stage_i.controller_i.priv_mode_i_1_ ),
    .Q(\cs_registers_i/_0009_ ));
 sg13g2_dfrbp_2 debug_mode_reg (.RESET_B(net2364),
    .D(_00095_),
    .Q(debug_mode),
    .Q_N(\debug_single_step_$_AND__B_A ),
    .CLK(clknet_leaf_222_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_0__reg  (.CLK(clknet_leaf_219_clk_i),
    .RESET_B(net2324),
    .D(_00096_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_0__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_0_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_10__reg  (.CLK(clknet_leaf_214_clk_i),
    .RESET_B(net2305),
    .D(_00097_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_10__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_10_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_11__reg  (.CLK(clknet_leaf_185_clk_i),
    .RESET_B(net2342),
    .D(_00098_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_11__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_11_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_12__reg  (.CLK(clknet_leaf_214_clk_i),
    .RESET_B(net2304),
    .D(_00099_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_12__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_12_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_13__reg  (.CLK(clknet_leaf_219_clk_i),
    .RESET_B(net2326),
    .D(_00100_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_13__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_13_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_14__reg  (.CLK(clknet_leaf_219_clk_i),
    .RESET_B(net2326),
    .D(_00101_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_14__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_14_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_15__reg  (.CLK(clknet_leaf_213_clk_i),
    .RESET_B(net2304),
    .D(_00102_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_15__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_15_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_16__reg  (.CLK(clknet_leaf_185_clk_i),
    .RESET_B(net2342),
    .D(_00103_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_16__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_16_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_17__reg  (.CLK(clknet_leaf_189_clk_i),
    .RESET_B(net2338),
    .D(_00104_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_17__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_17_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_18__reg  (.CLK(clknet_leaf_185_clk_i),
    .RESET_B(net2336),
    .D(_00105_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_18__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_18_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_19__reg  (.CLK(clknet_leaf_189_clk_i),
    .RESET_B(net2338),
    .D(_00106_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_19__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_19_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_1__reg  (.CLK(clknet_leaf_189_clk_i),
    .RESET_B(net2339),
    .D(_00107_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_1__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_1_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_20__reg  (.CLK(clknet_leaf_219_clk_i),
    .RESET_B(net2324),
    .D(_00108_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_20__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_20_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_21__reg  (.CLK(clknet_leaf_183_clk_i),
    .RESET_B(net2336),
    .D(_00109_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_21__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_21_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_22__reg  (.CLK(clknet_leaf_184_clk_i),
    .RESET_B(net2336),
    .D(_00110_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_22__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_22_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_23__reg  (.CLK(clknet_leaf_215_clk_i),
    .RESET_B(net2304),
    .D(_00111_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_23__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_23_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_24__reg  (.CLK(clknet_leaf_213_clk_i),
    .RESET_B(net2304),
    .D(_00112_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_24__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_24_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_25__reg  (.CLK(clknet_leaf_219_clk_i),
    .RESET_B(net2308),
    .D(_00113_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_25__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_25_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_26__reg  (.CLK(clknet_leaf_216_clk_i),
    .RESET_B(net2304),
    .D(_00114_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_26__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_26_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_27__reg  (.CLK(clknet_leaf_213_clk_i),
    .RESET_B(net2307),
    .D(_00115_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_27__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_27_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_28__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2304),
    .D(_00116_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_28__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_28_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_29__reg  (.CLK(clknet_leaf_216_clk_i),
    .RESET_B(net2304),
    .D(_00117_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_29__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_29_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_2__reg  (.CLK(clknet_leaf_183_clk_i),
    .RESET_B(net2336),
    .D(_00118_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_2__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_2_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_30__reg  (.CLK(clknet_leaf_183_clk_i),
    .RESET_B(net2324),
    .D(_00119_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_30__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_30_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_31__reg  (.CLK(clknet_leaf_218_clk_i),
    .RESET_B(net2324),
    .D(_00120_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_31__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_31_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_32__reg  (.RESET_B(net2326),
    .D(_00121_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_32_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_1__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_218_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_33__reg  (.RESET_B(net2325),
    .D(_00122_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_33_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_218_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_34__reg  (.RESET_B(net2325),
    .D(_00123_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_34_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_3__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_218_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_35__reg  (.RESET_B(net2324),
    .D(_00124_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_35_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_4__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_217_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_36__reg  (.RESET_B(net2326),
    .D(_00125_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_36_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_5__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_196_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_37__reg  (.RESET_B(net2312),
    .D(_00126_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_37_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_6__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_38__reg  (.RESET_B(net2330),
    .D(_00127_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_38_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_7__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_214_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_39__reg  (.RESET_B(net2336),
    .D(_00128_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_39_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_8__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_3__reg  (.CLK(clknet_leaf_183_clk_i),
    .RESET_B(net2342),
    .D(_00129_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_3__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_3_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_40__reg  (.RESET_B(net2336),
    .D(_00130_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_40_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_9__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_41__reg  (.CLK(clknet_leaf_194_clk_i),
    .RESET_B(net2312),
    .D(_00131_),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_10__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_41_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_42__reg  (.RESET_B(net2308),
    .D(_00132_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_42_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_11__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_217_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_43__reg  (.RESET_B(net2336),
    .D(_00133_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_43_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_12__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_44__reg  (.RESET_B(net2326),
    .D(_00134_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_44_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_13__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_45__reg  (.RESET_B(net2326),
    .D(_00135_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_45_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_14__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_195_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_46__reg  (.RESET_B(net2339),
    .D(_00136_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_46_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_15__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_217_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_47__reg  (.RESET_B(net2306),
    .D(_00137_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_47_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_16__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_214_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_48__reg  (.RESET_B(net2325),
    .D(_00138_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_48_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_17__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_184_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_49__reg  (.RESET_B(net2325),
    .D(_00139_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_49_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_18__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_195_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_4__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2302),
    .D(_00140_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_4__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_4_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_50__reg  (.RESET_B(net2325),
    .D(_00141_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_50_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_19__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_184_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_51__reg  (.RESET_B(net2326),
    .D(_00142_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_51_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_20__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_217_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_52__reg  (.RESET_B(net2324),
    .D(_00143_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_52_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_21__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_219_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_53__reg  (.RESET_B(net2337),
    .D(_00144_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_53_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_22__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_184_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_54__reg  (.RESET_B(net2337),
    .D(_00145_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_54_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_23__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_184_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_55__reg  (.RESET_B(net2307),
    .D(_00146_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_55_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_24__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_215_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_56__reg  (.CLK(clknet_leaf_195_clk_i),
    .RESET_B(net2339),
    .D(_00147_),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_25__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_56_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_57__reg  (.RESET_B(net2308),
    .D(_00148_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_57_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_26__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_216_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_58__reg  (.RESET_B(net2308),
    .D(_00149_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_58_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_27__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_217_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_59__reg  (.RESET_B(net2306),
    .D(_00150_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_59_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_28__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_215_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_5__reg  (.CLK(clknet_leaf_215_clk_i),
    .RESET_B(net2304),
    .D(_00151_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_5__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_5_ ));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_60__reg  (.RESET_B(net2308),
    .D(_00152_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_60_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_29__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_196_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_61__reg  (.RESET_B(net2308),
    .D(_00153_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_61_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_30__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_196_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_62__reg  (.RESET_B(net2325),
    .D(_00154_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_62_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_31__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_184_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.alu_i.imd_val_q_i_63__reg  (.RESET_B(net2324),
    .D(_00155_),
    .Q(\ex_block_i.alu_i.imd_val_q_i_63_ ),
    .Q_N(\ex_block_i.alu_i.multdiv_operand_b_i_32__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .CLK(clknet_leaf_183_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_6__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2302),
    .D(_00156_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_6__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_6_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_7__reg  (.CLK(clknet_leaf_189_clk_i),
    .RESET_B(net2338),
    .D(_00157_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_7__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_7_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_8__reg  (.CLK(clknet_leaf_218_clk_i),
    .RESET_B(net2325),
    .D(_00158_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_8__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_8_ ));
 sg13g2_dfrbp_1 \ex_block_i.alu_i.imd_val_q_i_9__reg  (.CLK(clknet_leaf_214_clk_i),
    .RESET_B(net2305),
    .D(_00159_),
    .Q_N(\ex_block_i.alu_i.imd_val_q_i_9__$_NOT__A_Y ),
    .Q(\ex_block_i.alu_i.imd_val_q_i_9_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q_reg  (.CLK(clknet_leaf_197_clk_i),
    .RESET_B(net2312),
    .D(_00160_),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_change_sign_$_AND__Y_B ),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_by_zero_q ));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0__reg  (.RESET_B(net2309),
    .D(_00161_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_0_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_0__$_MUX__Y_A ),
    .CLK(clknet_leaf_209_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1__reg  (.RESET_B(net2309),
    .D(_00162_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_1_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .CLK(clknet_leaf_209_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2__reg  (.RESET_B(net2309),
    .D(_00163_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_2_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_A ),
    .CLK(clknet_leaf_209_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_3__reg  (.CLK(clknet_leaf_210_clk_i),
    .RESET_B(net2311),
    .D(_00164_),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_3__$_MUX__Y_A_$_XOR__Y_A ),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_3_ ));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4__reg  (.RESET_B(net2311),
    .D(_00165_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_4_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_A ),
    .CLK(clknet_leaf_211_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__reg  (.RESET_B(net2339),
    .D(_00166_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_0__$_NOT__A_Y ),
    .CLK(clknet_leaf_189_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__reg  (.RESET_B(net2342),
    .D(_00167_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q_1__$_NOT__A_Y ),
    .CLK(clknet_leaf_189_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66__reg  (.RESET_B(net2337),
    .D(_00168_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_66_ ),
    .Q_N(_09000_),
    .CLK(clknet_leaf_194_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67__reg  (.RESET_B(net2339),
    .D(_00169_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.imd_val_q_i_67_ ),
    .Q_N(_08999_),
    .CLK(clknet_leaf_189_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__reg  (.RESET_B(net2306),
    .D(_00170_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0__$_NOT__A_Y ),
    .CLK(clknet_leaf_205_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_1__reg  (.RESET_B(net2308),
    .D(_00171_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_1_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_212_clk_i));
 sg13g2_dfrbp_2 \ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2__reg  (.RESET_B(net2306),
    .D(_00172_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.div_valid_$_NOT__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_214_clk_i));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_0__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2303),
    .D(_00173_),
    .Q_N(_08998_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_0_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_10__reg  (.CLK(clknet_leaf_231_clk_i),
    .RESET_B(net2309),
    .D(_00174_),
    .Q_N(_08997_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_10_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_11__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2305),
    .D(_00175_),
    .Q_N(_08996_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_11_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_12__reg  (.CLK(clknet_leaf_246_clk_i),
    .RESET_B(net2302),
    .D(_00176_),
    .Q_N(_08995_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_12_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_13__reg  (.CLK(clknet_leaf_246_clk_i),
    .RESET_B(net2302),
    .D(_00177_),
    .Q_N(_08994_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_13_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_14__reg  (.CLK(clknet_leaf_237_clk_i),
    .RESET_B(net2302),
    .D(_00178_),
    .Q_N(_08993_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_14_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_15__reg  (.CLK(clknet_leaf_237_clk_i),
    .RESET_B(net2305),
    .D(_00179_),
    .Q_N(_08992_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_15_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_16__reg  (.CLK(clknet_leaf_231_clk_i),
    .RESET_B(net2309),
    .D(_00180_),
    .Q_N(_08991_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_16_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_17__reg  (.CLK(clknet_leaf_231_clk_i),
    .RESET_B(net2309),
    .D(_00181_),
    .Q_N(_08990_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_17_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_18__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2309),
    .D(_00182_),
    .Q_N(_08989_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_18_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_19__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2309),
    .D(_00183_),
    .Q_N(_08988_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_19_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_1__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2303),
    .D(_00184_),
    .Q_N(_08987_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_1_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_20__reg  (.CLK(clknet_leaf_210_clk_i),
    .RESET_B(net2312),
    .D(_00185_),
    .Q_N(_08986_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_20_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_21__reg  (.CLK(clknet_leaf_210_clk_i),
    .RESET_B(net2310),
    .D(_00186_),
    .Q_N(_08985_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_21_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_22__reg  (.CLK(clknet_leaf_210_clk_i),
    .RESET_B(net2312),
    .D(_00187_),
    .Q_N(_08984_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_22_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_23__reg  (.CLK(clknet_leaf_210_clk_i),
    .RESET_B(net2310),
    .D(_00188_),
    .Q_N(_08983_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_23_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_24__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2310),
    .D(_00189_),
    .Q_N(_08982_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_24_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_25__reg  (.CLK(clknet_leaf_231_clk_i),
    .RESET_B(net2310),
    .D(_00190_),
    .Q_N(_08981_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_25_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_26__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2306),
    .D(_00191_),
    .Q_N(_08980_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_26_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_27__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2310),
    .D(_00192_),
    .Q_N(_08979_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_27_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_28__reg  (.CLK(clknet_leaf_236_clk_i),
    .RESET_B(net2305),
    .D(_00193_),
    .Q_N(_08978_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_28_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_29__reg  (.CLK(clknet_leaf_236_clk_i),
    .RESET_B(net2305),
    .D(_00194_),
    .Q_N(_08977_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_29_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_2__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2303),
    .D(_00195_),
    .Q_N(_08976_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_2_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_30__reg  (.CLK(clknet_leaf_236_clk_i),
    .RESET_B(net2305),
    .D(_00196_),
    .Q_N(_08975_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_30_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31__reg  (.CLK(clknet_leaf_232_clk_i),
    .RESET_B(net2306),
    .D(_00197_),
    .Q_N(_08974_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_31_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_3__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2303),
    .D(_00198_),
    .Q_N(_08973_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_3_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_4__reg  (.CLK(clknet_leaf_246_clk_i),
    .RESET_B(net2302),
    .D(_00199_),
    .Q_N(_08972_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_4_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_5__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2302),
    .D(_00200_),
    .Q_N(_08971_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_5_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_6__reg  (.CLK(clknet_leaf_230_clk_i),
    .RESET_B(net2303),
    .D(_00201_),
    .Q_N(_08970_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_6_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_7__reg  (.CLK(clknet_leaf_246_clk_i),
    .RESET_B(net2302),
    .D(_00202_),
    .Q_N(_08969_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_7_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_8__reg  (.CLK(clknet_leaf_231_clk_i),
    .RESET_B(net2303),
    .D(_00203_),
    .Q_N(_08968_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_8_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_9__reg  (.CLK(clknet_leaf_236_clk_i),
    .RESET_B(net2305),
    .D(_00204_),
    .Q_N(_08967_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_numerator_q_9_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_0__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2330),
    .D(_00205_),
    .Q_N(_08966_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_0_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_10__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2330),
    .D(_00206_),
    .Q_N(_08965_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_10_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_11__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2328),
    .D(_00207_),
    .Q_N(_08964_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_11_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_12__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2327),
    .D(_00208_),
    .Q_N(_08963_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_12_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_13__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2312),
    .D(_00209_),
    .Q_N(_08962_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_13_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_14__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2327),
    .D(_00210_),
    .Q_N(_08961_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_14_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_15__reg  (.CLK(clknet_leaf_205_clk_i),
    .RESET_B(net2312),
    .D(_00211_),
    .Q_N(_08960_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_15_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_16__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2328),
    .D(_00212_),
    .Q_N(_08959_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_16_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_17__reg  (.CLK(clknet_leaf_204_clk_i),
    .RESET_B(net2330),
    .D(_00213_),
    .Q_N(_08958_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_17_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_18__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2328),
    .D(_00214_),
    .Q_N(_08957_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_18_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_19__reg  (.CLK(clknet_leaf_211_clk_i),
    .RESET_B(net2330),
    .D(_00215_),
    .Q_N(_08956_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_19_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_1__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2328),
    .D(_00216_),
    .Q_N(_08955_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_1_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_20__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2313),
    .D(_00217_),
    .Q_N(_08954_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_20_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_21__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2327),
    .D(_00218_),
    .Q_N(_08953_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_21_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_22__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2314),
    .D(_00219_),
    .Q_N(_08952_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_22_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_23__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2314),
    .D(_00220_),
    .Q_N(_08951_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_23_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_24__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2313),
    .D(_00221_),
    .Q_N(_08950_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_24_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_25__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2314),
    .D(_00222_),
    .Q_N(_08949_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_25_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_26__reg  (.CLK(clknet_leaf_197_clk_i),
    .RESET_B(net2313),
    .D(_00223_),
    .Q_N(_08948_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_26_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_27__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2314),
    .D(_00224_),
    .Q_N(_08947_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_27_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_28__reg  (.CLK(clknet_leaf_211_clk_i),
    .RESET_B(net2311),
    .D(_00225_),
    .Q_N(_08946_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_28_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_29__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2313),
    .D(_00226_),
    .Q_N(_08945_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_29_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_2__reg  (.CLK(clknet_leaf_198_clk_i),
    .RESET_B(net2336),
    .D(_00227_),
    .Q_N(_08944_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_2_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_30__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2313),
    .D(_00228_),
    .Q_N(_08943_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_30_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_31__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2327),
    .D(_00229_),
    .Q_N(_08942_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_31_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_3__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2331),
    .D(_00230_),
    .Q_N(_08941_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_3_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_4__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2327),
    .D(_00231_),
    .Q_N(_08940_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_4_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_5__reg  (.CLK(clknet_leaf_212_clk_i),
    .RESET_B(net2312),
    .D(_00232_),
    .Q_N(_08939_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_5_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_6__reg  (.CLK(clknet_leaf_199_clk_i),
    .RESET_B(net2330),
    .D(_00233_),
    .Q_N(_08938_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_6_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_7__reg  (.CLK(clknet_leaf_211_clk_i),
    .RESET_B(net2316),
    .D(_00234_),
    .Q_N(_08937_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_7_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_8__reg  (.CLK(clknet_leaf_204_clk_i),
    .RESET_B(net2331),
    .D(_00235_),
    .Q_N(_08936_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_8_ ));
 sg13g2_dfrbp_1 \ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_9__reg  (.CLK(clknet_leaf_197_clk_i),
    .RESET_B(net2331),
    .D(_00236_),
    .Q_N(_09095_),
    .Q(\ex_block_i.gen_multdiv_fast.multdiv_i.op_quotient_q_9_ ));
 sg13g2_dfrbp_1 \id_stage_i.branch_jump_set_done_q_reg  (.CLK(clknet_leaf_221_clk_i),
    .RESET_B(net2360),
    .D(\id_stage_i.branch_jump_set_done_d ),
    .Q_N(\id_stage_i.branch_set_$_AND__Y_B ),
    .Q(\id_stage_i.branch_jump_set_done_q ));
 sg13g2_dfrbp_1 \id_stage_i.branch_set_raw_reg  (.CLK(clknet_leaf_221_clk_i),
    .RESET_B(net2395),
    .D(\id_stage_i.branch_set_raw_d ),
    .Q_N(_08935_),
    .Q(\id_stage_i.branch_set_raw ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.ctrl_fsm_cs_0__reg  (.CLK(clknet_leaf_174_clk_i),
    .RESET_B(net2364),
    .D(_00237_),
    .Q_N(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs_0_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.ctrl_fsm_cs_1__reg  (.RESET_B(net2362),
    .D(_00238_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs_1_ ),
    .Q_N(\id_stage_i.controller_i.debug_mode_d_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_174_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.ctrl_fsm_cs_2__reg  (.RESET_B(net2363),
    .D(_00239_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs_2_ ),
    .Q_N(\id_stage_i.controller_i.ctrl_fsm_cs_2__$_NOT__A_Y ),
    .CLK(clknet_leaf_174_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.ctrl_fsm_cs_3__reg  (.RESET_B(net2364),
    .D(_00240_),
    .Q(\id_stage_i.controller_i.ctrl_fsm_cs_3_ ),
    .Q_N(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .CLK(clknet_leaf_174_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.do_single_step_q_reg  (.CLK(clknet_leaf_222_clk_i),
    .RESET_B(net2375),
    .D(\id_stage_i.controller_i.do_single_step_d ),
    .Q_N(_09096_),
    .Q(\id_stage_i.controller_i.do_single_step_q ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.enter_debug_mode_prio_q_reg  (.CLK(clknet_leaf_222_clk_i),
    .RESET_B(net2364),
    .D(\id_stage_i.controller_i.enter_debug_mode_prio_d ),
    .Q_N(_09097_),
    .Q(\id_stage_i.controller_i.enter_debug_mode_prio_q ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.exc_req_q_reg  (.CLK(clknet_leaf_221_clk_i),
    .RESET_B(net2360),
    .D(\id_stage_i.controller_i.exc_req_d ),
    .Q_N(_09098_),
    .Q(\id_stage_i.controller_i.exc_req_q ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.illegal_insn_q_reg  (.CLK(clknet_leaf_221_clk_i),
    .RESET_B(net2360),
    .D(\id_stage_i.controller_i.illegal_insn_d ),
    .Q_N(_08934_),
    .Q(\id_stage_i.controller_i.illegal_insn_q ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_0__reg  (.CLK(clknet_leaf_179_clk_i),
    .RESET_B(net2269),
    .D(_00241_),
    .Q_N(_08933_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_0_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_10__reg  (.CLK(clknet_leaf_167_clk_i),
    .RESET_B(net2263),
    .D(_00242_),
    .Q_N(_08932_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_10_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_11__reg  (.CLK(clknet_leaf_178_clk_i),
    .RESET_B(net2270),
    .D(_00243_),
    .Q_N(_08931_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_11_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_compressed_i_12__reg  (.RESET_B(net2263),
    .D(_00244_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_12_ ),
    .Q_N(_08930_),
    .CLK(clknet_leaf_180_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_13__reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2362),
    .D(_00245_),
    .Q_N(_08929_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_13_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_14__reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2266),
    .D(_00246_),
    .Q_N(_08928_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_14_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_15__reg  (.CLK(clknet_leaf_179_clk_i),
    .RESET_B(net2269),
    .D(_00247_),
    .Q_N(_08927_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_15_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_1__reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2362),
    .D(_00248_),
    .Q_N(_08926_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_1_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_2__reg  (.CLK(clknet_leaf_179_clk_i),
    .RESET_B(net2269),
    .D(_00249_),
    .Q_N(_08925_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_2_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_3__reg  (.CLK(clknet_leaf_178_clk_i),
    .RESET_B(net2361),
    .D(_00250_),
    .Q_N(_08924_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_3_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_4__reg  (.CLK(clknet_leaf_179_clk_i),
    .RESET_B(net2270),
    .D(_00251_),
    .Q_N(_08923_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_4_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_5__reg  (.CLK(clknet_leaf_167_clk_i),
    .RESET_B(net2263),
    .D(_00252_),
    .Q_N(_08922_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_5_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_6__reg  (.CLK(clknet_leaf_179_clk_i),
    .RESET_B(net2269),
    .D(_00253_),
    .Q_N(_08921_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_6_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_7__reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2269),
    .D(_00254_),
    .Q_N(_08920_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_7_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_compressed_i_8__reg  (.RESET_B(net2363),
    .D(_00255_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_8_ ),
    .Q_N(_08919_),
    .CLK(clknet_leaf_167_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_compressed_i_9__reg  (.CLK(clknet_leaf_178_clk_i),
    .RESET_B(net2270),
    .D(_00256_),
    .Q_N(_08918_),
    .Q(\id_stage_i.controller_i.instr_compressed_i_9_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_fetch_err_i_reg  (.CLK(clknet_leaf_176_clk_i),
    .RESET_B(net2360),
    .D(_00257_),
    .Q_N(\id_stage_i.instr_perf_count_id_o_$_AND__Y_B ),
    .Q(\id_stage_i.controller_i.instr_fetch_err_i ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_fetch_err_plus2_i_reg  (.RESET_B(net2363),
    .D(_00258_),
    .Q(\id_stage_i.controller_i.instr_fetch_err_plus2_i ),
    .Q_N(_08917_),
    .CLK(clknet_leaf_169_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_0__reg  (.RESET_B(net2269),
    .D(_00259_),
    .Q(\id_stage_i.controller_i.instr_i_0_ ),
    .Q_N(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y ),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_10__reg  (.RESET_B(net2265),
    .D(_00260_),
    .Q(\id_stage_i.controller_i.instr_i_10_ ),
    .Q_N(_08916_),
    .CLK(clknet_leaf_167_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_11__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2264),
    .D(_00261_),
    .Q_N(_08915_),
    .Q(\id_stage_i.controller_i.instr_i_11_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_12__reg  (.RESET_B(net2254),
    .D(_00262_),
    .Q(\id_stage_i.controller_i.instr_i_12_ ),
    .Q_N(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .CLK(clknet_6_53_0_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_13__reg  (.CLK(clknet_leaf_186_clk_i),
    .RESET_B(net2268),
    .D(_00263_),
    .Q_N(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .Q(\id_stage_i.controller_i.instr_i_13_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_14__reg  (.CLK(clknet_leaf_187_clk_i),
    .RESET_B(net2266),
    .D(_00264_),
    .Q_N(\id_stage_i.alu_op_b_mux_sel_dec_$_MUX__Y_B_$_OR__Y_A_$_AND__Y_A ),
    .Q(\id_stage_i.controller_i.instr_i_14_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_15__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2263),
    .D(_00265_),
    .Q_N(_08914_),
    .Q(\id_stage_i.controller_i.instr_i_15_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_16__reg  (.RESET_B(net2266),
    .D(_00266_),
    .Q(\id_stage_i.controller_i.instr_i_16_ ),
    .Q_N(_08913_),
    .CLK(clknet_leaf_169_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_17__reg  (.RESET_B(net2266),
    .D(_00267_),
    .Q(\id_stage_i.controller_i.instr_i_17_ ),
    .Q_N(_08912_),
    .CLK(clknet_leaf_169_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_18__reg  (.RESET_B(net2270),
    .D(_00268_),
    .Q(\id_stage_i.controller_i.instr_i_18_ ),
    .Q_N(_08911_),
    .CLK(clknet_leaf_177_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_19__reg  (.RESET_B(net2265),
    .D(_00269_),
    .Q(\id_stage_i.controller_i.instr_i_19_ ),
    .Q_N(_08910_),
    .CLK(clknet_leaf_167_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_1__reg  (.RESET_B(net2361),
    .D(_00270_),
    .Q(\id_stage_i.controller_i.instr_i_1_ ),
    .Q_N(\id_stage_i.controller_i.instr_i_1__$_NOT__A_1_Y ),
    .CLK(clknet_leaf_177_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_20__reg  (.RESET_B(net2361),
    .D(_00271_),
    .Q(\id_stage_i.controller_i.instr_i_20_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .CLK(clknet_leaf_180_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_21__reg  (.RESET_B(net2269),
    .D(_00272_),
    .Q(\id_stage_i.controller_i.instr_i_21_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_178_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_22__reg  (.RESET_B(net2268),
    .D(_00273_),
    .Q(\id_stage_i.controller_i.instr_i_22_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .CLK(clknet_leaf_187_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_23__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2263),
    .D(_00274_),
    .Q_N(_08909_),
    .Q(\id_stage_i.controller_i.instr_i_23_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_24__reg  (.RESET_B(net2266),
    .D(_00275_),
    .Q(\id_stage_i.controller_i.instr_i_24_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__B_A ),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_25__reg  (.RESET_B(net2266),
    .D(_00276_),
    .Q(\id_stage_i.controller_i.instr_i_25_ ),
    .Q_N(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .CLK(clknet_leaf_187_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_26__reg  (.RESET_B(net2268),
    .D(_00277_),
    .Q(\id_stage_i.controller_i.instr_i_26_ ),
    .Q_N(\ex_block_i.gen_multdiv_fast.multdiv_i.operator_i_0__$_MUX__Y_A_$_MUX__Y_S_$_OR__Y_B ),
    .CLK(clknet_leaf_186_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_27__reg  (.RESET_B(net2268),
    .D(_00278_),
    .Q(\id_stage_i.controller_i.instr_i_27_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .CLK(clknet_leaf_187_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_28__reg  (.RESET_B(net2269),
    .D(_00279_),
    .Q(\id_stage_i.controller_i.instr_i_28_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B ),
    .CLK(clknet_leaf_177_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_29__reg  (.RESET_B(net2361),
    .D(_00280_),
    .Q(\id_stage_i.controller_i.instr_i_29_ ),
    .Q_N(\id_stage_i.controller_i.csr_pipe_flush_i_$_MUX__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .CLK(clknet_leaf_177_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_2__reg  (.RESET_B(net2271),
    .D(_00281_),
    .Q(\id_stage_i.controller_i.instr_i_2_ ),
    .Q_N(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_B_$_OR__Y_A ),
    .CLK(clknet_leaf_179_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_30__reg  (.CLK(clknet_leaf_187_clk_i),
    .RESET_B(net2268),
    .D(_00282_),
    .Q_N(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__A_B_$_NOT__Y_A_$_OR__Y_B_$_OR__Y_A ),
    .Q(\id_stage_i.controller_i.instr_i_30_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_31__reg  (.CLK(clknet_leaf_151_clk_i),
    .RESET_B(net2263),
    .D(_00283_),
    .Q_N(_08908_),
    .Q(\id_stage_i.controller_i.instr_i_31_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_3__reg  (.RESET_B(net2270),
    .D(_00284_),
    .Q(\id_stage_i.controller_i.instr_i_3_ ),
    .Q_N(\id_stage_i.controller_i.instr_i_0__$_NOT__A_1_Y_$_OR__A_Y_$_OR__A_1_B_$_OR__Y_B ),
    .CLK(clknet_leaf_179_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_4__reg  (.RESET_B(net2271),
    .D(_00285_),
    .Q(\id_stage_i.controller_i.instr_i_4_ ),
    .Q_N(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A ),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_5__reg  (.RESET_B(net2271),
    .D(_00286_),
    .Q(\id_stage_i.controller_i.instr_i_5_ ),
    .Q_N(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_6__reg  (.RESET_B(net2271),
    .D(_00287_),
    .Q(\id_stage_i.controller_i.instr_i_6_ ),
    .Q_N(\id_stage_i.decoder_i.csr_op_0__$_MUX__Y_S_$_OR__Y_B_$_OR__Y_B ),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_7__reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2361),
    .D(_00288_),
    .Q_N(_08907_),
    .Q(\id_stage_i.controller_i.instr_i_7_ ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.instr_i_8__reg  (.RESET_B(net2266),
    .D(_00289_),
    .Q(\id_stage_i.controller_i.instr_i_8_ ),
    .Q_N(_08906_),
    .CLK(clknet_leaf_181_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_i_9__reg  (.CLK(clknet_leaf_178_clk_i),
    .RESET_B(net2270),
    .D(_00290_),
    .Q_N(_08905_),
    .Q(\id_stage_i.controller_i.instr_i_9_ ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_is_compressed_i_reg  (.CLK(clknet_leaf_177_clk_i),
    .RESET_B(net2270),
    .D(_00291_),
    .Q_N(\id_stage_i.imm_b_2__$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_AND__Y_A ),
    .Q(\id_stage_i.controller_i.instr_is_compressed_i ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.instr_valid_i_reg  (.CLK(clknet_leaf_175_clk_i),
    .RESET_B(net2365),
    .D(\if_stage_i.instr_valid_id_d ),
    .Q_N(\id_in_ready_$_AND__Y_A_$_AND__Y_A_$_AND__A_Y_$_AND__A_B ),
    .Q(\id_stage_i.controller_i.instr_valid_i ));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.load_err_q_reg  (.CLK(clknet_leaf_175_clk_i),
    .RESET_B(net2360),
    .D(\id_stage_i.controller_i.load_err_i ),
    .Q_N(_08904_),
    .Q(\id_stage_i.controller_i.load_err_q ));
 sg13g2_dfrbp_2 \id_stage_i.controller_i.nmi_mode_o_reg  (.RESET_B(net2364),
    .D(_00292_),
    .Q(\id_stage_i.controller_i.nmi_mode_o ),
    .Q_N(\id_stage_i.controller_i.handle_irq_$_AND__Y_A_$_AND__Y_B ),
    .CLK(clknet_leaf_222_clk_i));
 sg13g2_dfrbp_1 \id_stage_i.controller_i.store_err_q_reg  (.CLK(clknet_leaf_175_clk_i),
    .RESET_B(net2360),
    .D(\id_stage_i.controller_i.store_err_i ),
    .Q_N(_08903_),
    .Q(\id_stage_i.controller_i.store_err_q ));
 sg13g2_dfrbp_1 \id_stage_i.decoder_i.illegal_c_insn_i_reg  (.CLK(clknet_leaf_180_clk_i),
    .RESET_B(net2264),
    .D(_00293_),
    .Q_N(_08902_),
    .Q(\id_stage_i.decoder_i.illegal_c_insn_i ));
 sg13g2_dfrbp_2 \id_stage_i.id_fsm_q_reg  (.RESET_B(net2271),
    .D(_00294_),
    .Q(\id_stage_i.id_fsm_q ),
    .Q_N(\ex_block_i.alu_i.instr_first_cycle_i_$_AND__Y_B ),
    .CLK(clknet_leaf_176_clk_i));
 sg13g2_dfrbp_2 \if_stage_i.prefetch_buffer_i.branch_discard_q_0__reg  (.RESET_B(net2417),
    .D(\if_stage_i.prefetch_buffer_i.branch_discard_s_0_ ),
    .Q(\if_stage_i.prefetch_buffer_i.branch_discard_q_0_ ),
    .Q_N(\if_stage_i.prefetch_buffer_i.fifo_i.in_valid_i_$_AND__Y_B ),
    .CLK(clknet_leaf_186_clk_i));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.branch_discard_q_1__reg  (.CLK(clknet_leaf_186_clk_i),
    .RESET_B(net2435),
    .D(\if_stage_i.prefetch_buffer_i.branch_discard_s_1_ ),
    .Q_N(_09099_),
    .Q(\if_stage_i.prefetch_buffer_i.branch_discard_q_1_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.discard_req_q_reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2430),
    .D(\if_stage_i.prefetch_buffer_i.discard_req_d ),
    .Q_N(_08901_),
    .Q(\if_stage_i.prefetch_buffer_i.discard_req_q ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_10__reg  (.CLK(clknet_leaf_207_clk_i),
    .RESET_B(net2427),
    .D(_00295_),
    .Q_N(_08900_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_10_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_11__reg  (.CLK(clknet_leaf_207_clk_i),
    .RESET_B(net2426),
    .D(_00296_),
    .Q_N(_08899_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_11_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_12__reg  (.CLK(clknet_leaf_208_clk_i),
    .RESET_B(net2344),
    .D(_00297_),
    .Q_N(_08898_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_12_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_13__reg  (.CLK(clknet_leaf_208_clk_i),
    .RESET_B(net2426),
    .D(_00298_),
    .Q_N(_08897_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_13_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_14__reg  (.CLK(clknet_leaf_208_clk_i),
    .RESET_B(net2426),
    .D(_00299_),
    .Q_N(_08896_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_14_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_15__reg  (.CLK(clknet_leaf_208_clk_i),
    .RESET_B(net2344),
    .D(_00300_),
    .Q_N(_08895_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_15_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_16__reg  (.CLK(clknet_leaf_209_clk_i),
    .RESET_B(net2426),
    .D(_00301_),
    .Q_N(_08894_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_16_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_17__reg  (.CLK(clknet_leaf_209_clk_i),
    .RESET_B(net2428),
    .D(_00302_),
    .Q_N(_08893_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_17_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_18__reg  (.CLK(clknet_leaf_207_clk_i),
    .RESET_B(net2428),
    .D(_00303_),
    .Q_N(_08892_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_18_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_19__reg  (.CLK(clknet_leaf_207_clk_i),
    .RESET_B(net2427),
    .D(_00304_),
    .Q_N(_08891_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_19_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_20__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2428),
    .D(_00305_),
    .Q_N(_08890_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_20_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_21__reg  (.CLK(clknet_leaf_199_clk_i),
    .RESET_B(net2427),
    .D(_00306_),
    .Q_N(_08889_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_21_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_22__reg  (.CLK(clknet_leaf_199_clk_i),
    .RESET_B(net2427),
    .D(_00307_),
    .Q_N(_08888_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_22_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_23__reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2430),
    .D(_00308_),
    .Q_N(_08887_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_23_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_24__reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2427),
    .D(_00309_),
    .Q_N(_08886_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_24_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_25__reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2427),
    .D(_00310_),
    .Q_N(_08885_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_25_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_26__reg  (.CLK(clknet_leaf_233_clk_i),
    .RESET_B(net2346),
    .D(_00311_),
    .Q_N(_08884_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_26_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_27__reg  (.CLK(clknet_leaf_201_clk_i),
    .RESET_B(net2428),
    .D(_00312_),
    .Q_N(_08883_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_27_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_28__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2428),
    .D(_00313_),
    .Q_N(_08882_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_28_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_29__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2428),
    .D(_00314_),
    .Q_N(_08881_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_29_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_2__reg  (.CLK(clknet_leaf_209_clk_i),
    .RESET_B(net2426),
    .D(_00315_),
    .Q_N(_08880_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_2_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_30__reg  (.CLK(clknet_leaf_199_clk_i),
    .RESET_B(net2428),
    .D(_00316_),
    .Q_N(_08879_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_30_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_31__reg  (.CLK(clknet_leaf_200_clk_i),
    .RESET_B(net2430),
    .D(_00317_),
    .Q_N(_08878_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_31_ ));
 sg13g2_dfrbp_2 \if_stage_i.prefetch_buffer_i.fetch_addr_q_3__reg  (.RESET_B(net2426),
    .D(_00318_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_3_ ),
    .Q_N(_08877_),
    .CLK(clknet_leaf_208_clk_i));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_4__reg  (.CLK(clknet_leaf_233_clk_i),
    .RESET_B(net2344),
    .D(_00319_),
    .Q_N(_08876_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_4_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_5__reg  (.CLK(clknet_leaf_208_clk_i),
    .RESET_B(net2426),
    .D(_00320_),
    .Q_N(_08875_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_5_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_6__reg  (.CLK(clknet_leaf_209_clk_i),
    .RESET_B(net2426),
    .D(_00321_),
    .Q_N(_08874_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_6_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_7__reg  (.CLK(clknet_leaf_206_clk_i),
    .RESET_B(net2429),
    .D(_00322_),
    .Q_N(_08873_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_7_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_8__reg  (.CLK(clknet_leaf_207_clk_i),
    .RESET_B(net2427),
    .D(_00323_),
    .Q_N(_08872_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_8_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fetch_addr_q_9__reg  (.CLK(clknet_leaf_203_clk_i),
    .RESET_B(net2427),
    .D(_00324_),
    .Q_N(_09100_),
    .Q(\if_stage_i.prefetch_buffer_i.fetch_addr_q_9_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_busy_0__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2373),
    .D(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_1_ ),
    .Q_N(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_1__$_AND__Y_A ),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_busy_0_ ));
 sg13g2_dfrbp_2 \if_stage_i.prefetch_buffer_i.fifo_busy_1__reg  (.RESET_B(net2373),
    .D(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_2_ ),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_busy_1_ ),
    .Q_N(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_2__$_AND__Y_A ),
    .CLK(clknet_leaf_151_clk_i));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.err_q_0__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2373),
    .D(_00325_),
    .Q_N(\if_stage_i.prefetch_buffer_i.fifo_i.err_plus2_$_AND__Y_B ),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_0_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.err_q_1__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2374),
    .D(_00326_),
    .Q_N(_08871_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_1_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.err_q_2__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2374),
    .D(_00327_),
    .Q_N(_08870_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.err_q_2_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2368),
    .D(_00328_),
    .Q_N(_08869_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_0_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_10__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2350),
    .D(_00329_),
    .Q_N(_08868_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_10_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_11__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00330_),
    .Q_N(_08867_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_11_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_12__reg  (.CLK(clknet_leaf_149_clk_i),
    .RESET_B(net2366),
    .D(_00331_),
    .Q_N(_08866_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_12_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_13__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2366),
    .D(_00332_),
    .Q_N(_08865_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_13_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_14__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2358),
    .D(_00333_),
    .Q_N(_08864_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_14_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_15__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2366),
    .D(_00334_),
    .Q_N(_08863_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_15_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2368),
    .D(_00335_),
    .Q_N(_08862_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_16_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17__reg  (.CLK(clknet_6_27_0_clk_i),
    .RESET_B(net2368),
    .D(_00336_),
    .Q_N(_08861_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_17_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_18__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2355),
    .D(_00337_),
    .Q_N(_08860_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_18_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_19__reg  (.CLK(clknet_leaf_136_clk_i),
    .RESET_B(net2383),
    .D(_00338_),
    .Q_N(_08859_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_19_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1__reg  (.CLK(clknet_leaf_149_clk_i),
    .RESET_B(net2368),
    .D(_00339_),
    .Q_N(_08858_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_1_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_20__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2383),
    .D(_00340_),
    .Q_N(_08857_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_20_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_21__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2355),
    .D(_00341_),
    .Q_N(_08856_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_21_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_22__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2383),
    .D(_00342_),
    .Q_N(_08855_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_22_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2371),
    .D(_00343_),
    .Q_N(_08854_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_23_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_24__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2355),
    .D(_00344_),
    .Q_N(_08853_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_24_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_25__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2389),
    .D(_00345_),
    .Q_N(_08852_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_25_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_26__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2355),
    .D(_00346_),
    .Q_N(_08851_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_26_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_27__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2354),
    .D(_00347_),
    .Q_N(_08850_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_27_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_28__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2371),
    .D(_00348_),
    .Q_N(_08849_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_28_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_29__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2371),
    .D(_00349_),
    .Q_N(_08848_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_29_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_2__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2353),
    .D(_00350_),
    .Q_N(_08847_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_2_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_30__reg  (.CLK(clknet_leaf_137_clk_i),
    .RESET_B(net2354),
    .D(_00351_),
    .Q_N(_08846_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_30_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_31__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2389),
    .D(_00352_),
    .Q_N(_08845_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_31_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_32__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2368),
    .D(_00353_),
    .Q_N(_08844_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_32_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_33__reg  (.CLK(clknet_leaf_149_clk_i),
    .RESET_B(net2368),
    .D(_00354_),
    .Q_N(_08843_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_33_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_34__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2353),
    .D(_00355_),
    .Q_N(_08842_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_34_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_35__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2353),
    .D(_00356_),
    .Q_N(_08841_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_35_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_36__reg  (.CLK(clknet_leaf_144_clk_i),
    .RESET_B(net2367),
    .D(_00357_),
    .Q_N(_08840_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_36_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_37__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00358_),
    .Q_N(_08839_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_37_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_38__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00359_),
    .Q_N(_08838_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_38_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_39__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2370),
    .D(_00360_),
    .Q_N(_08837_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_39_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_3__reg  (.CLK(clknet_leaf_144_clk_i),
    .RESET_B(net2353),
    .D(_00361_),
    .Q_N(_08836_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_3_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_40__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2367),
    .D(_00362_),
    .Q_N(_08835_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_40_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_41__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2370),
    .D(_00363_),
    .Q_N(_08834_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_41_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_42__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2350),
    .D(_00364_),
    .Q_N(_08833_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_42_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_43__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00365_),
    .Q_N(_08832_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_43_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_44__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2366),
    .D(_00366_),
    .Q_N(_08831_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_44_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_45__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2366),
    .D(_00367_),
    .Q_N(_08830_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_45_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_46__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2358),
    .D(_00368_),
    .Q_N(_08829_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_46_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_47__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2366),
    .D(_00369_),
    .Q_N(_08828_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_47_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_48__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2368),
    .D(_00370_),
    .Q_N(_08827_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_48_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_49__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2372),
    .D(_00371_),
    .Q_N(_08826_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_49_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_4__reg  (.CLK(clknet_leaf_144_clk_i),
    .RESET_B(net2367),
    .D(_00372_),
    .Q_N(_08825_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_4_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_50__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2355),
    .D(_00373_),
    .Q_N(_08824_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_50_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_51__reg  (.CLK(clknet_leaf_136_clk_i),
    .RESET_B(net2383),
    .D(_00374_),
    .Q_N(_08823_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_51_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_52__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2383),
    .D(_00375_),
    .Q_N(_08822_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_52_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_53__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2355),
    .D(_00376_),
    .Q_N(_08821_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_53_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_54__reg  (.CLK(clknet_leaf_136_clk_i),
    .RESET_B(net2383),
    .D(_00377_),
    .Q_N(_08820_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_54_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_55__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2370),
    .D(_00378_),
    .Q_N(_08819_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_55_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_56__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2370),
    .D(_00379_),
    .Q_N(_08818_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_56_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_57__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2389),
    .D(_00380_),
    .Q_N(_08817_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_57_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_58__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2355),
    .D(_00381_),
    .Q_N(_08816_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_58_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_59__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2354),
    .D(_00382_),
    .Q_N(_08815_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_59_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_5__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00383_),
    .Q_N(_08814_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_5_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_60__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2371),
    .D(_00384_),
    .Q_N(_08813_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_60_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_61__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2389),
    .D(_00385_),
    .Q_N(_08812_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_61_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_62__reg  (.CLK(clknet_leaf_137_clk_i),
    .RESET_B(net2354),
    .D(_00386_),
    .Q_N(_08811_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_62_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_63__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2389),
    .D(_00387_),
    .Q_N(_08810_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_63_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_64__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2369),
    .D(_00388_),
    .Q_N(_08809_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_64_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_65__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2368),
    .D(_00389_),
    .Q_N(_08808_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_65_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_66__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2353),
    .D(_00390_),
    .Q_N(_08807_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_66_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_67__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2353),
    .D(_00391_),
    .Q_N(_08806_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_67_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_68__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2367),
    .D(_00392_),
    .Q_N(_08805_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_68_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_69__reg  (.CLK(clknet_leaf_144_clk_i),
    .RESET_B(net2357),
    .D(_00393_),
    .Q_N(_08804_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_69_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_6__reg  (.CLK(clknet_leaf_188_clk_i),
    .RESET_B(net2352),
    .D(_00394_),
    .Q_N(_08803_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_6_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_70__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2352),
    .D(_00395_),
    .Q_N(_08802_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_70_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_71__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2370),
    .D(_00396_),
    .Q_N(_08801_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_71_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_72__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2355),
    .D(_00397_),
    .Q_N(_08800_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_72_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_73__reg  (.CLK(clknet_leaf_140_clk_i),
    .RESET_B(net2370),
    .D(_00398_),
    .Q_N(_08799_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_73_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_74__reg  (.CLK(clknet_leaf_142_clk_i),
    .RESET_B(net2350),
    .D(_00399_),
    .Q_N(_08798_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_74_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_75__reg  (.CLK(clknet_leaf_143_clk_i),
    .RESET_B(net2352),
    .D(_00400_),
    .Q_N(_08797_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_75_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_76__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2366),
    .D(_00401_),
    .Q_N(_08796_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_76_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_77__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2353),
    .D(_00402_),
    .Q_N(_08795_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_77_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_78__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2358),
    .D(_00403_),
    .Q_N(_08794_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_78_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_79__reg  (.CLK(clknet_leaf_146_clk_i),
    .RESET_B(net2366),
    .D(_00404_),
    .Q_N(_08793_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_79_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_7__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2369),
    .D(_00405_),
    .Q_N(_08792_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_7_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_80__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2369),
    .D(_00406_),
    .Q_N(_08791_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_80_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_81__reg  (.CLK(clknet_leaf_148_clk_i),
    .RESET_B(net2372),
    .D(_00407_),
    .Q_N(_08790_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_81_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_82__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2354),
    .D(_00408_),
    .Q_N(_08789_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_82_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_83__reg  (.CLK(clknet_leaf_136_clk_i),
    .RESET_B(net2383),
    .D(_00409_),
    .Q_N(_08788_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_83_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_84__reg  (.CLK(clknet_leaf_135_clk_i),
    .RESET_B(net2383),
    .D(_00410_),
    .Q_N(_08787_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_84_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_85__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2356),
    .D(_00411_),
    .Q_N(_08786_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_85_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_86__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2394),
    .D(_00412_),
    .Q_N(_08785_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_86_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_87__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2370),
    .D(_00413_),
    .Q_N(_08784_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_87_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_88__reg  (.CLK(clknet_leaf_137_clk_i),
    .RESET_B(net2354),
    .D(_00414_),
    .Q_N(_08783_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_88_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_89__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2389),
    .D(_00415_),
    .Q_N(_08782_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_89_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_8__reg  (.CLK(clknet_leaf_144_clk_i),
    .RESET_B(net2367),
    .D(_00416_),
    .Q_N(_08781_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_8_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_90__reg  (.CLK(clknet_leaf_141_clk_i),
    .RESET_B(net2356),
    .D(_00417_),
    .Q_N(_08780_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_90_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_91__reg  (.CLK(clknet_leaf_137_clk_i),
    .RESET_B(net2354),
    .D(_00418_),
    .Q_N(_08779_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_91_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_92__reg  (.CLK(clknet_leaf_139_clk_i),
    .RESET_B(net2354),
    .D(_00419_),
    .Q_N(_08778_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_92_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_93__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2356),
    .D(_00420_),
    .Q_N(_08777_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_93_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_94__reg  (.CLK(clknet_leaf_137_clk_i),
    .RESET_B(net2356),
    .D(_00421_),
    .Q_N(_08776_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_94_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_95__reg  (.CLK(clknet_leaf_138_clk_i),
    .RESET_B(net2389),
    .D(_00422_),
    .Q_N(_08775_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_95_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_9__reg  (.CLK(clknet_leaf_145_clk_i),
    .RESET_B(net2370),
    .D(_00423_),
    .Q_N(_09101_),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.rdata_q_9_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.fifo_i.valid_q_0__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2363),
    .D(\if_stage_i.prefetch_buffer_i.fifo_i.valid_d_0_ ),
    .Q_N(\if_stage_i.prefetch_buffer_i.fifo_i.lowest_free_entry_0_ ),
    .Q(\if_stage_i.prefetch_buffer_i.fifo_i.valid_q_0_ ));
 sg13g2_dfrbp_2 \if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0__reg  (.RESET_B(net2417),
    .D(\if_stage_i.prefetch_buffer_i.rdata_outstanding_s_0_ ),
    .Q(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_0_ ),
    .Q_N(_09102_),
    .CLK(clknet_leaf_186_clk_i));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1__reg  (.CLK(clknet_leaf_186_clk_i),
    .RESET_B(net2435),
    .D(\if_stage_i.prefetch_buffer_i.rdata_outstanding_s_1_ ),
    .Q_N(\if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__Y_B ),
    .Q(\if_stage_i.prefetch_buffer_i.rdata_outstanding_q_1_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_10__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2433),
    .D(_00424_),
    .Q_N(_08774_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_10_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_11__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2430),
    .D(_00425_),
    .Q_N(_08773_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_11_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_12__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00426_),
    .Q_N(_08772_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_12_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_13__reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2464),
    .D(_00427_),
    .Q_N(_08771_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_13_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_14__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2433),
    .D(_00428_),
    .Q_N(_08770_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_14_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_15__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2430),
    .D(_00429_),
    .Q_N(_08769_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_15_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_16__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00430_),
    .Q_N(_08768_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_16_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_17__reg  (.CLK(clknet_leaf_200_clk_i),
    .RESET_B(net2432),
    .D(_00431_),
    .Q_N(_08767_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_17_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_18__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00432_),
    .Q_N(_08766_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_18_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_19__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00433_),
    .Q_N(_08765_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_19_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_20__reg  (.CLK(clknet_leaf_201_clk_i),
    .RESET_B(net2431),
    .D(_00434_),
    .Q_N(_08764_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_20_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_21__reg  (.CLK(clknet_leaf_193_clk_i),
    .RESET_B(net2464),
    .D(_00435_),
    .Q_N(_08763_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_21_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_22__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00436_),
    .Q_N(_08762_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_22_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_23__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2432),
    .D(_00437_),
    .Q_N(_08761_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_23_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_24__reg  (.CLK(clknet_leaf_192_clk_i),
    .RESET_B(net2431),
    .D(_00438_),
    .Q_N(_08760_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_24_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_25__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2433),
    .D(_00439_),
    .Q_N(_08759_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_25_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_26__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2433),
    .D(_00440_),
    .Q_N(_08758_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_26_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_27__reg  (.CLK(clknet_leaf_201_clk_i),
    .RESET_B(net2430),
    .D(_00441_),
    .Q_N(_08757_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_27_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_28__reg  (.CLK(clknet_leaf_192_clk_i),
    .RESET_B(net2431),
    .D(_00442_),
    .Q_N(_08756_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_28_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_29__reg  (.CLK(clknet_leaf_191_clk_i),
    .RESET_B(net2432),
    .D(_00443_),
    .Q_N(_08755_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_29_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_2__reg  (.CLK(clknet_leaf_200_clk_i),
    .RESET_B(net2431),
    .D(_00444_),
    .Q_N(_08754_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_2_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_30__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2433),
    .D(_00445_),
    .Q_N(_08753_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_30_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_31__reg  (.CLK(clknet_leaf_192_clk_i),
    .RESET_B(net2433),
    .D(_00446_),
    .Q_N(_08752_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_31_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_3__reg  (.CLK(clknet_leaf_201_clk_i),
    .RESET_B(net2430),
    .D(_00447_),
    .Q_N(_08751_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_3_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_4__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2433),
    .D(_00448_),
    .Q_N(_08750_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_4_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_5__reg  (.CLK(clknet_leaf_201_clk_i),
    .RESET_B(net2431),
    .D(_00449_),
    .Q_N(_08749_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_5_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_6__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2434),
    .D(_00450_),
    .Q_N(_08748_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_6_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_7__reg  (.CLK(clknet_leaf_200_clk_i),
    .RESET_B(net2431),
    .D(_00451_),
    .Q_N(_08747_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_7_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_8__reg  (.CLK(clknet_leaf_190_clk_i),
    .RESET_B(net2434),
    .D(_00452_),
    .Q_N(_08746_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_8_ ));
 sg13g2_dfrbp_1 \if_stage_i.prefetch_buffer_i.stored_addr_q_9__reg  (.CLK(clknet_leaf_202_clk_i),
    .RESET_B(net2431),
    .D(_00453_),
    .Q_N(_09103_),
    .Q(\if_stage_i.prefetch_buffer_i.stored_addr_q_9_ ));
 sg13g2_dfrbp_2 \if_stage_i.prefetch_buffer_i.valid_req_q_reg  (.RESET_B(net2430),
    .D(\if_stage_i.prefetch_buffer_i.valid_req_d ),
    .Q(\if_stage_i.prefetch_buffer_i.valid_req_q ),
    .Q_N(\if_stage_i.prefetch_buffer_i.valid_new_req_$_AND__A_B ),
    .CLK(clknet_leaf_193_clk_i));
 sg13g2_dfrbp_1 \load_store_unit_i.data_sign_ext_q_reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2262),
    .D(_00454_),
    .Q_N(_08745_),
    .Q(\load_store_unit_i.data_sign_ext_q ));
 sg13g2_dfrbp_1 \load_store_unit_i.data_type_q_0__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2359),
    .D(_00455_),
    .Q_N(\load_store_unit_i.data_type_q_0__$_NOT__A_Y ),
    .Q(\load_store_unit_i.data_type_q_0_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.data_type_q_1__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2359),
    .D(_00456_),
    .Q_N(\load_store_unit_i.data_type_q_1__$_NOT__A_Y ),
    .Q(\load_store_unit_i.data_type_q_1_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.data_we_q_reg  (.CLK(clknet_leaf_175_clk_i),
    .RESET_B(net2361),
    .D(_00457_),
    .Q_N(\load_store_unit_i.lsu_rdata_valid_o_$_AND__Y_B ),
    .Q(\load_store_unit_i.data_we_q ));
 sg13g2_dfrbp_2 \load_store_unit_i.handle_misaligned_q_reg  (.RESET_B(net2271),
    .D(_00458_),
    .Q(\load_store_unit_i.handle_misaligned_q ),
    .Q_N(\data_be_o_$_MUX__Y_A ),
    .CLK(clknet_leaf_176_clk_i));
 sg13g2_dfrbp_1 \load_store_unit_i.ls_fsm_cs_0__reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2362),
    .D(_00459_),
    .Q_N(\load_store_unit_i.ls_fsm_cs_0__$_NOT__A_Y ),
    .Q(\load_store_unit_i.ls_fsm_cs_0_ ));
 sg13g2_dfrbp_2 \load_store_unit_i.ls_fsm_cs_1__reg  (.RESET_B(net2362),
    .D(_00460_),
    .Q(\load_store_unit_i.ls_fsm_cs_1_ ),
    .Q_N(\load_store_unit_i.ls_fsm_cs_1__$_NOT__A_Y ),
    .CLK(clknet_leaf_176_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.ls_fsm_cs_2__reg  (.RESET_B(net2362),
    .D(_00461_),
    .Q(\load_store_unit_i.ls_fsm_cs_2_ ),
    .Q_N(\load_store_unit_i.busy_o_$_OR__Y_A_$_OR__A_B ),
    .CLK(clknet_leaf_173_clk_i));
 sg13g2_dfrbp_1 \load_store_unit_i.lsu_err_q_reg  (.CLK(clknet_leaf_174_clk_i),
    .RESET_B(net2361),
    .D(_00462_),
    .Q_N(\load_store_unit_i.lsu_err_q_$_NOT__A_Y ),
    .Q(\load_store_unit_i.lsu_err_q ));
 sg13g2_dfrbp_1 \load_store_unit_i.pmp_err_q_reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2361),
    .D(_00463_),
    .Q_N(_08744_),
    .Q(\load_store_unit_i.pmp_err_q ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_offset_q_0__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2359),
    .D(_00464_),
    .Q_N(\load_store_unit_i.rdata_offset_q_0__$_NOT__A_Y ),
    .Q(\load_store_unit_i.rdata_offset_q_0_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_offset_q_1__reg  (.CLK(clknet_6_16_0_clk_i),
    .RESET_B(net2358),
    .D(_00465_),
    .Q_N(\load_store_unit_i.rdata_offset_q_1__$_NOT__A_Y ),
    .Q(\load_store_unit_i.rdata_offset_q_1_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_0__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net2350),
    .D(_00466_),
    .Q_N(_08743_),
    .Q(\load_store_unit_i.rdata_q_0_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_10__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net2349),
    .D(_00467_),
    .Q_N(_08742_),
    .Q(\load_store_unit_i.rdata_q_10_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_11__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2262),
    .D(_00468_),
    .Q_N(_08741_),
    .Q(\load_store_unit_i.rdata_q_11_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_12__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2358),
    .D(_00469_),
    .Q_N(_08740_),
    .Q(\load_store_unit_i.rdata_q_12_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_13__reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net2358),
    .D(_00470_),
    .Q_N(_08739_),
    .Q(\load_store_unit_i.rdata_q_13_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_14__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net2349),
    .D(_00471_),
    .Q_N(_08738_),
    .Q(\load_store_unit_i.rdata_q_14_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_15__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net2349),
    .D(_00472_),
    .Q_N(_08737_),
    .Q(\load_store_unit_i.rdata_q_15_ ));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_16__reg  (.RESET_B(net2350),
    .D(_00473_),
    .Q(\load_store_unit_i.rdata_q_16_ ),
    .Q_N(_08736_),
    .CLK(clknet_leaf_91_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_17__reg  (.RESET_B(net2358),
    .D(_00474_),
    .Q(\load_store_unit_i.rdata_q_17_ ),
    .Q_N(_08735_),
    .CLK(clknet_leaf_107_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_18__reg  (.RESET_B(net2349),
    .D(_00475_),
    .Q(\load_store_unit_i.rdata_q_18_ ),
    .Q_N(_08734_),
    .CLK(clknet_leaf_86_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_19__reg  (.RESET_B(net2359),
    .D(_00476_),
    .Q(\load_store_unit_i.rdata_q_19_ ),
    .Q_N(_08733_),
    .CLK(clknet_leaf_92_clk_i));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_1__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2359),
    .D(_00477_),
    .Q_N(_08732_),
    .Q(\load_store_unit_i.rdata_q_1_ ));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_20__reg  (.RESET_B(net2359),
    .D(_00478_),
    .Q(\load_store_unit_i.rdata_q_20_ ),
    .Q_N(_08731_),
    .CLK(clknet_leaf_92_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_21__reg  (.RESET_B(net2350),
    .D(_00479_),
    .Q(\load_store_unit_i.rdata_q_21_ ),
    .Q_N(_08730_),
    .CLK(clknet_leaf_92_clk_i));
 sg13g2_dfrbp_2 \load_store_unit_i.rdata_q_22__reg  (.RESET_B(net2349),
    .D(_00480_),
    .Q(\load_store_unit_i.rdata_q_22_ ),
    .Q_N(_08729_),
    .CLK(clknet_leaf_86_clk_i));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_23__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net2349),
    .D(_00481_),
    .Q_N(_08728_),
    .Q(\load_store_unit_i.rdata_q_23_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_2__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net2351),
    .D(_00482_),
    .Q_N(_08727_),
    .Q(\load_store_unit_i.rdata_q_2_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_3__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2359),
    .D(_00483_),
    .Q_N(_08726_),
    .Q(\load_store_unit_i.rdata_q_3_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_4__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net2359),
    .D(_00484_),
    .Q_N(_08725_),
    .Q(\load_store_unit_i.rdata_q_4_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_5__reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net2351),
    .D(_00485_),
    .Q_N(_08724_),
    .Q(\load_store_unit_i.rdata_q_5_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_6__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net2350),
    .D(_00486_),
    .Q_N(_08723_),
    .Q(\load_store_unit_i.rdata_q_6_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_7__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net2351),
    .D(_00487_),
    .Q_N(_08722_),
    .Q(\load_store_unit_i.rdata_q_7_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_8__reg  (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net2350),
    .D(_00488_),
    .Q_N(_08721_),
    .Q(\load_store_unit_i.rdata_q_8_ ));
 sg13g2_dfrbp_1 \load_store_unit_i.rdata_q_9__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net2358),
    .D(_00489_),
    .Q_N(_08720_),
    .Q(\load_store_unit_i.rdata_q_9_ ));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(net435));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(net435));
 sg13g2_nor2b_1 \register_file_i/_4036_  (.A(net536),
    .B_N(net525),
    .Y(\register_file_i/_0994_ ));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(net435));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net435));
 sg13g2_buf_2 fanout429 (.A(_01167_),
    .X(net429));
 sg13g2_buf_2 fanout428 (.A(_01167_),
    .X(net428));
 sg13g2_buf_2 fanout427 (.A(_04045_),
    .X(net427));
 sg13g2_mux2_1 \register_file_i/_4042_  (.A0(\register_file_i/rf_reg_927_ ),
    .A1(\register_file_i/rf_reg_959_ ),
    .S(net2050),
    .X(\register_file_i/_1000_ ));
 sg13g2_buf_2 fanout426 (.A(net427),
    .X(net426));
 sg13g2_mux2_1 \register_file_i/_4044_  (.A0(\register_file_i/rf_reg_991_ ),
    .A1(\register_file_i/rf_reg_1023_ ),
    .S(net2051),
    .X(\register_file_i/_1002_ ));
 sg13g2_and2_2 \register_file_i/_4045_  (.A(net525),
    .B(net531),
    .X(\register_file_i/_1003_ ));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(net427));
 sg13g2_buf_4 fanout424 (.X(net424),
    .A(net427));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(net427));
 sg13g2_a22oi_1 \register_file_i/_4049_  (.Y(\register_file_i/_1007_ ),
    .B1(\register_file_i/_1002_ ),
    .B2(net1826),
    .A2(\register_file_i/_1000_ ),
    .A1(net1843));
 sg13g2_nor2b_1 \register_file_i/_4050_  (.A(net530),
    .B_N(net531),
    .Y(\register_file_i/_1008_ ));
 sg13g2_buf_2 fanout422 (.A(_04116_),
    .X(net422));
 sg13g2_buf_2 fanout421 (.A(_04116_),
    .X(net421));
 sg13g2_mux2_1 \register_file_i/_4053_  (.A0(\register_file_i/rf_reg_863_ ),
    .A1(\register_file_i/rf_reg_895_ ),
    .S(net2049),
    .X(\register_file_i/_1011_ ));
 sg13g2_buf_2 fanout420 (.A(_04116_),
    .X(net420));
 sg13g2_mux2_1 \register_file_i/_4055_  (.A0(\register_file_i/rf_reg_799_ ),
    .A1(\register_file_i/rf_reg_831_ ),
    .S(net2049),
    .X(\register_file_i/_1013_ ));
 sg13g2_nor2_1 \register_file_i/_4056_  (.A(net525),
    .B(net531),
    .Y(\register_file_i/_1014_ ));
 sg13g2_buf_2 fanout419 (.A(_04116_),
    .X(net419));
 sg13g2_buf_1 fanout418 (.A(_08409_),
    .X(net418));
 sg13g2_a22oi_1 \register_file_i/_4059_  (.Y(\register_file_i/_1017_ ),
    .B1(\register_file_i/_1013_ ),
    .B2(net1807),
    .A2(\register_file_i/_1011_ ),
    .A1(net1818));
 sg13g2_nand2_2 \register_file_i/_4060_  (.Y(\register_file_i/_1018_ ),
    .A(\id_stage_i.controller_i.instr_i_19_ ),
    .B(net2009));
 sg13g2_buf_1 fanout417 (.A(net418),
    .X(net417));
 sg13g2_a21o_1 \register_file_i/_4062_  (.A2(\register_file_i/_1017_ ),
    .A1(\register_file_i/_1007_ ),
    .B1(net1929),
    .X(\register_file_i/_1020_ ));
 sg13g2_nor2_1 \register_file_i/_4063_  (.A(\id_stage_i.controller_i.instr_i_19_ ),
    .B(net2009),
    .Y(\register_file_i/_1021_ ));
 sg13g2_buf_2 fanout416 (.A(net418),
    .X(net416));
 sg13g2_buf_2 fanout415 (.A(net418),
    .X(net415));
 sg13g2_buf_4 fanout414 (.X(net414),
    .A(net418));
 sg13g2_buf_4 fanout413 (.X(net413),
    .A(net418));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_01153_));
 sg13g2_mux2_1 \register_file_i/_4069_  (.A0(\register_file_i/rf_reg_63_ ),
    .A1(\register_file_i/rf_reg_127_ ),
    .S(net532),
    .X(\register_file_i/_1027_ ));
 sg13g2_buf_4 fanout411 (.X(net411),
    .A(_01394_));
 sg13g2_nor2b_1 \register_file_i/_4071_  (.A(net2084),
    .B_N(net531),
    .Y(\register_file_i/_1029_ ));
 sg13g2_buf_4 fanout410 (.X(net410),
    .A(_01394_));
 sg13g2_a22oi_1 \register_file_i/_4073_  (.Y(\register_file_i/_1031_ ),
    .B1(net1702),
    .B2(\register_file_i/rf_reg_95_ ),
    .A2(\register_file_i/_1027_ ),
    .A1(net2078));
 sg13g2_buf_1 fanout409 (.A(_01832_),
    .X(net409));
 sg13g2_buf_2 fanout408 (.A(_01832_),
    .X(net408));
 sg13g2_mux2_1 \register_file_i/_4076_  (.A0(\register_file_i/rf_reg_223_ ),
    .A1(\register_file_i/rf_reg_255_ ),
    .S(net2079),
    .X(\register_file_i/_1034_ ));
 sg13g2_buf_4 fanout407 (.X(net407),
    .A(net408));
 sg13g2_mux2_1 \register_file_i/_4078_  (.A0(\register_file_i/rf_reg_159_ ),
    .A1(\register_file_i/rf_reg_191_ ),
    .S(net2079),
    .X(\register_file_i/_1036_ ));
 sg13g2_buf_2 fanout406 (.A(net408),
    .X(net406));
 sg13g2_a22oi_1 \register_file_i/_4080_  (.Y(\register_file_i/_1038_ ),
    .B1(\register_file_i/_1036_ ),
    .B2(net1851),
    .A2(\register_file_i/_1034_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4081_  (.B1(\register_file_i/_1038_ ),
    .Y(\register_file_i/_1039_ ),
    .A1(net527),
    .A2(\register_file_i/_1031_ ));
 sg13g2_nand2_1 \register_file_i/_4082_  (.Y(\register_file_i/_1040_ ),
    .A(net1922),
    .B(\register_file_i/_1039_ ));
 sg13g2_inv_1 \register_file_i/_4083_  (.Y(\register_file_i/_1041_ ),
    .A(\id_stage_i.controller_i.instr_i_19_ ));
 sg13g2_nor3_2 \register_file_i/_4084_  (.A(\register_file_i/_1041_ ),
    .B(net2009),
    .C(net530),
    .Y(\register_file_i/_1042_ ));
 sg13g2_buf_2 fanout405 (.A(net408),
    .X(net405));
 sg13g2_buf_4 fanout404 (.X(net404),
    .A(net408));
 sg13g2_buf_2 fanout403 (.A(net408),
    .X(net403));
 sg13g2_buf_2 fanout402 (.A(net409),
    .X(net402));
 sg13g2_mux4_1 \register_file_i/_4089_  (.S0(net2038),
    .A0(\register_file_i/rf_reg_543_ ),
    .A1(\register_file_i/rf_reg_575_ ),
    .A2(\register_file_i/rf_reg_607_ ),
    .A3(\register_file_i/rf_reg_639_ ),
    .S1(net538),
    .X(\register_file_i/_1047_ ));
 sg13g2_inv_1 \register_file_i/_4090_  (.Y(\register_file_i/_1048_ ),
    .A(net525));
 sg13g2_nor3_2 \register_file_i/_4091_  (.A(\register_file_i/_1041_ ),
    .B(net2009),
    .C(\register_file_i/_1048_ ),
    .Y(\register_file_i/_1049_ ));
 sg13g2_buf_2 fanout401 (.A(net409),
    .X(net401));
 sg13g2_buf_2 fanout400 (.A(net409),
    .X(net400));
 sg13g2_mux4_1 \register_file_i/_4094_  (.S0(net2039),
    .A0(\register_file_i/rf_reg_671_ ),
    .A1(\register_file_i/rf_reg_703_ ),
    .A2(\register_file_i/rf_reg_735_ ),
    .A3(\register_file_i/rf_reg_767_ ),
    .S1(net538),
    .X(\register_file_i/_1052_ ));
 sg13g2_buf_4 fanout399 (.X(net399),
    .A(net408));
 sg13g2_buf_4 fanout398 (.X(net398),
    .A(net408));
 sg13g2_mux2_1 \register_file_i/_4097_  (.A0(\register_file_i/rf_reg_479_ ),
    .A1(\register_file_i/rf_reg_511_ ),
    .S(net2038),
    .X(\register_file_i/_1055_ ));
 sg13g2_buf_4 fanout397 (.X(net397),
    .A(_01199_));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_01199_));
 sg13g2_mux2_1 \register_file_i/_4100_  (.A0(\register_file_i/rf_reg_415_ ),
    .A1(\register_file_i/rf_reg_447_ ),
    .S(net2036),
    .X(\register_file_i/_1058_ ));
 sg13g2_a22oi_1 \register_file_i/_4101_  (.Y(\register_file_i/_1059_ ),
    .B1(net1840),
    .B2(\register_file_i/_1058_ ),
    .A2(\register_file_i/_1055_ ),
    .A1(net1823));
 sg13g2_buf_2 fanout395 (.A(_01582_),
    .X(net395));
 sg13g2_mux2_1 \register_file_i/_4103_  (.A0(\register_file_i/rf_reg_351_ ),
    .A1(\register_file_i/rf_reg_383_ ),
    .S(net2036),
    .X(\register_file_i/_1061_ ));
 sg13g2_buf_2 fanout394 (.A(_07476_),
    .X(net394));
 sg13g2_mux2_1 \register_file_i/_4105_  (.A0(\register_file_i/rf_reg_287_ ),
    .A1(\register_file_i/rf_reg_319_ ),
    .S(net2040),
    .X(\register_file_i/_1063_ ));
 sg13g2_buf_2 fanout393 (.A(net394),
    .X(net393));
 sg13g2_a22oi_1 \register_file_i/_4107_  (.Y(\register_file_i/_1065_ ),
    .B1(\register_file_i/_1063_ ),
    .B2(net1803),
    .A2(net1811),
    .A1(\register_file_i/_1061_ ));
 sg13g2_nand2_2 \register_file_i/_4108_  (.Y(\register_file_i/_1066_ ),
    .A(\register_file_i/_1041_ ),
    .B(net2009));
 sg13g2_buf_2 fanout392 (.A(net394),
    .X(net392));
 sg13g2_a21oi_1 \register_file_i/_4110_  (.A1(\register_file_i/_1059_ ),
    .A2(\register_file_i/_1065_ ),
    .Y(\register_file_i/_1068_ ),
    .B1(net1791));
 sg13g2_a221oi_1 \register_file_i/_4111_  (.B2(\register_file_i/_1052_ ),
    .C1(\register_file_i/_1068_ ),
    .B1(net1697),
    .A1(net1796),
    .Y(\register_file_i/_1069_ ),
    .A2(\register_file_i/_1047_ ));
 sg13g2_nand3_1 \register_file_i/_4112_  (.B(\register_file_i/_1040_ ),
    .C(\register_file_i/_1069_ ),
    .A(\register_file_i/_1020_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_31_ ));
 sg13g2_mux2_1 \register_file_i/_4113_  (.A0(\register_file_i/rf_reg_926_ ),
    .A1(\register_file_i/rf_reg_958_ ),
    .S(net2045),
    .X(\register_file_i/_1070_ ));
 sg13g2_mux2_1 \register_file_i/_4114_  (.A0(\register_file_i/rf_reg_990_ ),
    .A1(\register_file_i/rf_reg_1022_ ),
    .S(net2049),
    .X(\register_file_i/_1071_ ));
 sg13g2_a22oi_1 \register_file_i/_4115_  (.Y(\register_file_i/_1072_ ),
    .B1(\register_file_i/_1071_ ),
    .B2(net1826),
    .A2(\register_file_i/_1070_ ),
    .A1(net1843));
 sg13g2_buf_2 fanout391 (.A(_07480_),
    .X(net391));
 sg13g2_mux2_1 \register_file_i/_4117_  (.A0(\register_file_i/rf_reg_862_ ),
    .A1(\register_file_i/rf_reg_894_ ),
    .S(net2048),
    .X(\register_file_i/_1074_ ));
 sg13g2_mux2_1 \register_file_i/_4118_  (.A0(\register_file_i/rf_reg_798_ ),
    .A1(\register_file_i/rf_reg_830_ ),
    .S(net2045),
    .X(\register_file_i/_1075_ ));
 sg13g2_a22oi_1 \register_file_i/_4119_  (.Y(\register_file_i/_1076_ ),
    .B1(\register_file_i/_1075_ ),
    .B2(net1802),
    .A2(\register_file_i/_1074_ ),
    .A1(net1813));
 sg13g2_a21o_1 \register_file_i/_4120_  (.A2(\register_file_i/_1076_ ),
    .A1(\register_file_i/_1072_ ),
    .B1(net1929),
    .X(\register_file_i/_1077_ ));
 sg13g2_mux2_1 \register_file_i/_4121_  (.A0(\register_file_i/rf_reg_62_ ),
    .A1(\register_file_i/rf_reg_126_ ),
    .S(net533),
    .X(\register_file_i/_1078_ ));
 sg13g2_buf_2 fanout390 (.A(_07480_),
    .X(net390));
 sg13g2_a22oi_1 \register_file_i/_4123_  (.Y(\register_file_i/_1080_ ),
    .B1(\register_file_i/_1078_ ),
    .B2(net2079),
    .A2(net1702),
    .A1(\register_file_i/rf_reg_94_ ));
 sg13g2_mux2_1 \register_file_i/_4124_  (.A0(\register_file_i/rf_reg_222_ ),
    .A1(\register_file_i/rf_reg_254_ ),
    .S(net2078),
    .X(\register_file_i/_1081_ ));
 sg13g2_mux2_1 \register_file_i/_4125_  (.A0(\register_file_i/rf_reg_158_ ),
    .A1(\register_file_i/rf_reg_190_ ),
    .S(net2079),
    .X(\register_file_i/_1082_ ));
 sg13g2_a22oi_1 \register_file_i/_4126_  (.Y(\register_file_i/_1083_ ),
    .B1(\register_file_i/_1082_ ),
    .B2(net1851),
    .A2(\register_file_i/_1081_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4127_  (.B1(\register_file_i/_1083_ ),
    .Y(\register_file_i/_1084_ ),
    .A1(net527),
    .A2(\register_file_i/_1080_ ));
 sg13g2_nand2_1 \register_file_i/_4128_  (.Y(\register_file_i/_1085_ ),
    .A(net1923),
    .B(\register_file_i/_1084_ ));
 sg13g2_mux4_1 \register_file_i/_4129_  (.S0(net2043),
    .A0(\register_file_i/rf_reg_542_ ),
    .A1(\register_file_i/rf_reg_574_ ),
    .A2(\register_file_i/rf_reg_606_ ),
    .A3(\register_file_i/rf_reg_638_ ),
    .S1(net538),
    .X(\register_file_i/_1086_ ));
 sg13g2_buf_2 fanout389 (.A(_07586_),
    .X(net389));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(_07586_));
 sg13g2_mux4_1 \register_file_i/_4132_  (.S0(net2043),
    .A0(\register_file_i/rf_reg_670_ ),
    .A1(\register_file_i/rf_reg_702_ ),
    .A2(\register_file_i/rf_reg_734_ ),
    .A3(\register_file_i/rf_reg_766_ ),
    .S1(net540),
    .X(\register_file_i/_1089_ ));
 sg13g2_buf_2 fanout387 (.A(_01803_),
    .X(net387));
 sg13g2_mux2_1 \register_file_i/_4134_  (.A0(\register_file_i/rf_reg_414_ ),
    .A1(\register_file_i/rf_reg_446_ ),
    .S(net2047),
    .X(\register_file_i/_1091_ ));
 sg13g2_mux2_1 \register_file_i/_4135_  (.A0(\register_file_i/rf_reg_478_ ),
    .A1(\register_file_i/rf_reg_510_ ),
    .S(net2038),
    .X(\register_file_i/_1092_ ));
 sg13g2_buf_1 fanout386 (.A(_07542_),
    .X(net386));
 sg13g2_a22oi_1 \register_file_i/_4137_  (.Y(\register_file_i/_1094_ ),
    .B1(\register_file_i/_1092_ ),
    .B2(net1824),
    .A2(\register_file_i/_1091_ ),
    .A1(net1840));
 sg13g2_buf_2 fanout385 (.A(_07542_),
    .X(net385));
 sg13g2_mux2_1 \register_file_i/_4139_  (.A0(\register_file_i/rf_reg_350_ ),
    .A1(\register_file_i/rf_reg_382_ ),
    .S(net2047),
    .X(\register_file_i/_1096_ ));
 sg13g2_mux2_1 \register_file_i/_4140_  (.A0(\register_file_i/rf_reg_286_ ),
    .A1(\register_file_i/rf_reg_318_ ),
    .S(net2047),
    .X(\register_file_i/_1097_ ));
 sg13g2_a22oi_1 \register_file_i/_4141_  (.Y(\register_file_i/_1098_ ),
    .B1(\register_file_i/_1097_ ),
    .B2(net1802),
    .A2(\register_file_i/_1096_ ),
    .A1(net1813));
 sg13g2_a21oi_1 \register_file_i/_4142_  (.A1(\register_file_i/_1094_ ),
    .A2(\register_file_i/_1098_ ),
    .Y(\register_file_i/_1099_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4143_  (.B2(net1697),
    .C1(\register_file_i/_1099_ ),
    .B1(\register_file_i/_1089_ ),
    .A1(net1796),
    .Y(\register_file_i/_1100_ ),
    .A2(\register_file_i/_1086_ ));
 sg13g2_nand3_1 \register_file_i/_4144_  (.B(\register_file_i/_1085_ ),
    .C(\register_file_i/_1100_ ),
    .A(\register_file_i/_1077_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_30_ ));
 sg13g2_mux2_1 \register_file_i/_4145_  (.A0(\register_file_i/rf_reg_917_ ),
    .A1(\register_file_i/rf_reg_949_ ),
    .S(net2081),
    .X(\register_file_i/_1101_ ));
 sg13g2_mux2_1 \register_file_i/_4146_  (.A0(\register_file_i/rf_reg_981_ ),
    .A1(\register_file_i/rf_reg_1013_ ),
    .S(net2050),
    .X(\register_file_i/_1102_ ));
 sg13g2_a22oi_1 \register_file_i/_4147_  (.Y(\register_file_i/_1103_ ),
    .B1(\register_file_i/_1102_ ),
    .B2(net1826),
    .A2(\register_file_i/_1101_ ),
    .A1(net1843));
 sg13g2_mux2_1 \register_file_i/_4148_  (.A0(\register_file_i/rf_reg_853_ ),
    .A1(\register_file_i/rf_reg_885_ ),
    .S(net2049),
    .X(\register_file_i/_1104_ ));
 sg13g2_mux2_1 \register_file_i/_4149_  (.A0(\register_file_i/rf_reg_789_ ),
    .A1(\register_file_i/rf_reg_821_ ),
    .S(net2049),
    .X(\register_file_i/_1105_ ));
 sg13g2_a22oi_1 \register_file_i/_4150_  (.Y(\register_file_i/_1106_ ),
    .B1(\register_file_i/_1105_ ),
    .B2(net1807),
    .A2(\register_file_i/_1104_ ),
    .A1(net1818));
 sg13g2_a21o_1 \register_file_i/_4151_  (.A2(\register_file_i/_1106_ ),
    .A1(\register_file_i/_1103_ ),
    .B1(net1929),
    .X(\register_file_i/_1107_ ));
 sg13g2_mux2_1 \register_file_i/_4152_  (.A0(\register_file_i/rf_reg_53_ ),
    .A1(\register_file_i/rf_reg_117_ ),
    .S(net533),
    .X(\register_file_i/_1108_ ));
 sg13g2_a22oi_1 \register_file_i/_4153_  (.Y(\register_file_i/_1109_ ),
    .B1(\register_file_i/_1108_ ),
    .B2(net2077),
    .A2(net1702),
    .A1(\register_file_i/rf_reg_85_ ));
 sg13g2_mux2_1 \register_file_i/_4154_  (.A0(\register_file_i/rf_reg_213_ ),
    .A1(\register_file_i/rf_reg_245_ ),
    .S(net2077),
    .X(\register_file_i/_1110_ ));
 sg13g2_mux2_1 \register_file_i/_4155_  (.A0(\register_file_i/rf_reg_149_ ),
    .A1(\register_file_i/rf_reg_181_ ),
    .S(net2045),
    .X(\register_file_i/_1111_ ));
 sg13g2_a22oi_1 \register_file_i/_4156_  (.Y(\register_file_i/_1112_ ),
    .B1(\register_file_i/_1111_ ),
    .B2(net1852),
    .A2(\register_file_i/_1110_ ),
    .A1(net1825));
 sg13g2_o21ai_1 \register_file_i/_4157_  (.B1(\register_file_i/_1112_ ),
    .Y(\register_file_i/_1113_ ),
    .A1(net526),
    .A2(\register_file_i/_1109_ ));
 sg13g2_nand2_1 \register_file_i/_4158_  (.Y(\register_file_i/_1114_ ),
    .A(net1922),
    .B(\register_file_i/_1113_ ));
 sg13g2_mux4_1 \register_file_i/_4159_  (.S0(net2038),
    .A0(\register_file_i/rf_reg_533_ ),
    .A1(\register_file_i/rf_reg_565_ ),
    .A2(\register_file_i/rf_reg_597_ ),
    .A3(\register_file_i/rf_reg_629_ ),
    .S1(net538),
    .X(\register_file_i/_1115_ ));
 sg13g2_mux4_1 \register_file_i/_4160_  (.S0(net2039),
    .A0(\register_file_i/rf_reg_661_ ),
    .A1(\register_file_i/rf_reg_693_ ),
    .A2(\register_file_i/rf_reg_725_ ),
    .A3(\register_file_i/rf_reg_757_ ),
    .S1(net540),
    .X(\register_file_i/_1116_ ));
 sg13g2_buf_1 fanout384 (.A(_01542_),
    .X(net384));
 sg13g2_mux2_1 \register_file_i/_4162_  (.A0(\register_file_i/rf_reg_405_ ),
    .A1(\register_file_i/rf_reg_437_ ),
    .S(net2036),
    .X(\register_file_i/_1118_ ));
 sg13g2_mux2_1 \register_file_i/_4163_  (.A0(\register_file_i/rf_reg_469_ ),
    .A1(\register_file_i/rf_reg_501_ ),
    .S(net2036),
    .X(\register_file_i/_1119_ ));
 sg13g2_a22oi_1 \register_file_i/_4164_  (.Y(\register_file_i/_1120_ ),
    .B1(\register_file_i/_1119_ ),
    .B2(net1824),
    .A2(\register_file_i/_1118_ ),
    .A1(net1841));
 sg13g2_mux2_1 \register_file_i/_4165_  (.A0(\register_file_i/rf_reg_341_ ),
    .A1(\register_file_i/rf_reg_373_ ),
    .S(net2036),
    .X(\register_file_i/_1121_ ));
 sg13g2_mux2_1 \register_file_i/_4166_  (.A0(\register_file_i/rf_reg_277_ ),
    .A1(\register_file_i/rf_reg_309_ ),
    .S(net2036),
    .X(\register_file_i/_1122_ ));
 sg13g2_a22oi_1 \register_file_i/_4167_  (.Y(\register_file_i/_1123_ ),
    .B1(\register_file_i/_1122_ ),
    .B2(net1803),
    .A2(\register_file_i/_1121_ ),
    .A1(net1814));
 sg13g2_a21oi_1 \register_file_i/_4168_  (.A1(\register_file_i/_1120_ ),
    .A2(\register_file_i/_1123_ ),
    .Y(\register_file_i/_1124_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4169_  (.B2(net1697),
    .C1(\register_file_i/_1124_ ),
    .B1(\register_file_i/_1116_ ),
    .A1(net1795),
    .Y(\register_file_i/_1125_ ),
    .A2(\register_file_i/_1115_ ));
 sg13g2_nand3_1 \register_file_i/_4170_  (.B(\register_file_i/_1114_ ),
    .C(\register_file_i/_1125_ ),
    .A(\register_file_i/_1107_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_21_ ));
 sg13g2_buf_2 fanout383 (.A(_01542_),
    .X(net383));
 sg13g2_mux2_1 \register_file_i/_4172_  (.A0(\register_file_i/rf_reg_916_ ),
    .A1(\register_file_i/rf_reg_948_ ),
    .S(net2050),
    .X(\register_file_i/_1127_ ));
 sg13g2_mux2_1 \register_file_i/_4173_  (.A0(\register_file_i/rf_reg_980_ ),
    .A1(\register_file_i/rf_reg_1012_ ),
    .S(net2050),
    .X(\register_file_i/_1128_ ));
 sg13g2_a22oi_1 \register_file_i/_4174_  (.Y(\register_file_i/_1129_ ),
    .B1(\register_file_i/_1128_ ),
    .B2(net1826),
    .A2(\register_file_i/_1127_ ),
    .A1(net1843));
 sg13g2_mux2_1 \register_file_i/_4175_  (.A0(\register_file_i/rf_reg_852_ ),
    .A1(\register_file_i/rf_reg_884_ ),
    .S(net2049),
    .X(\register_file_i/_1130_ ));
 sg13g2_mux2_1 \register_file_i/_4176_  (.A0(\register_file_i/rf_reg_788_ ),
    .A1(\register_file_i/rf_reg_820_ ),
    .S(net2050),
    .X(\register_file_i/_1131_ ));
 sg13g2_a22oi_1 \register_file_i/_4177_  (.Y(\register_file_i/_1132_ ),
    .B1(\register_file_i/_1131_ ),
    .B2(net1802),
    .A2(\register_file_i/_1130_ ),
    .A1(net1813));
 sg13g2_a21o_1 \register_file_i/_4178_  (.A2(\register_file_i/_1132_ ),
    .A1(\register_file_i/_1129_ ),
    .B1(net1929),
    .X(\register_file_i/_1133_ ));
 sg13g2_mux2_1 \register_file_i/_4179_  (.A0(\register_file_i/rf_reg_52_ ),
    .A1(\register_file_i/rf_reg_116_ ),
    .S(net533),
    .X(\register_file_i/_1134_ ));
 sg13g2_a22oi_1 \register_file_i/_4180_  (.Y(\register_file_i/_1135_ ),
    .B1(\register_file_i/_1134_ ),
    .B2(net2079),
    .A2(net1702),
    .A1(\register_file_i/rf_reg_84_ ));
 sg13g2_mux2_1 \register_file_i/_4181_  (.A0(\register_file_i/rf_reg_212_ ),
    .A1(\register_file_i/rf_reg_244_ ),
    .S(net2081),
    .X(\register_file_i/_1136_ ));
 sg13g2_mux2_1 \register_file_i/_4182_  (.A0(\register_file_i/rf_reg_148_ ),
    .A1(\register_file_i/rf_reg_180_ ),
    .S(net2081),
    .X(\register_file_i/_1137_ ));
 sg13g2_a22oi_1 \register_file_i/_4183_  (.Y(\register_file_i/_1138_ ),
    .B1(\register_file_i/_1137_ ),
    .B2(net1852),
    .A2(\register_file_i/_1136_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4184_  (.B1(\register_file_i/_1138_ ),
    .Y(\register_file_i/_1139_ ),
    .A1(net526),
    .A2(\register_file_i/_1135_ ));
 sg13g2_nand2_1 \register_file_i/_4185_  (.Y(\register_file_i/_1140_ ),
    .A(net1922),
    .B(\register_file_i/_1139_ ));
 sg13g2_mux4_1 \register_file_i/_4186_  (.S0(net2038),
    .A0(\register_file_i/rf_reg_532_ ),
    .A1(\register_file_i/rf_reg_564_ ),
    .A2(\register_file_i/rf_reg_596_ ),
    .A3(\register_file_i/rf_reg_628_ ),
    .S1(net538),
    .X(\register_file_i/_1141_ ));
 sg13g2_mux4_1 \register_file_i/_4187_  (.S0(net2039),
    .A0(\register_file_i/rf_reg_660_ ),
    .A1(\register_file_i/rf_reg_692_ ),
    .A2(\register_file_i/rf_reg_724_ ),
    .A3(\register_file_i/rf_reg_756_ ),
    .S1(net540),
    .X(\register_file_i/_1142_ ));
 sg13g2_mux2_1 \register_file_i/_4188_  (.A0(\register_file_i/rf_reg_404_ ),
    .A1(\register_file_i/rf_reg_436_ ),
    .S(net2039),
    .X(\register_file_i/_1143_ ));
 sg13g2_mux2_1 \register_file_i/_4189_  (.A0(\register_file_i/rf_reg_468_ ),
    .A1(\register_file_i/rf_reg_500_ ),
    .S(net2038),
    .X(\register_file_i/_1144_ ));
 sg13g2_a22oi_1 \register_file_i/_4190_  (.Y(\register_file_i/_1145_ ),
    .B1(\register_file_i/_1144_ ),
    .B2(net1824),
    .A2(\register_file_i/_1143_ ),
    .A1(net1841));
 sg13g2_mux2_1 \register_file_i/_4191_  (.A0(\register_file_i/rf_reg_340_ ),
    .A1(\register_file_i/rf_reg_372_ ),
    .S(net2038),
    .X(\register_file_i/_1146_ ));
 sg13g2_buf_2 fanout382 (.A(_01542_),
    .X(net382));
 sg13g2_mux2_1 \register_file_i/_4193_  (.A0(\register_file_i/rf_reg_276_ ),
    .A1(\register_file_i/rf_reg_308_ ),
    .S(net2038),
    .X(\register_file_i/_1148_ ));
 sg13g2_a22oi_1 \register_file_i/_4194_  (.Y(\register_file_i/_1149_ ),
    .B1(\register_file_i/_1148_ ),
    .B2(net1800),
    .A2(\register_file_i/_1146_ ),
    .A1(net1814));
 sg13g2_a21oi_1 \register_file_i/_4195_  (.A1(\register_file_i/_1145_ ),
    .A2(\register_file_i/_1149_ ),
    .Y(\register_file_i/_1150_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4196_  (.B2(net1697),
    .C1(\register_file_i/_1150_ ),
    .B1(\register_file_i/_1142_ ),
    .A1(net1795),
    .Y(\register_file_i/_1151_ ),
    .A2(\register_file_i/_1141_ ));
 sg13g2_nand3_1 \register_file_i/_4197_  (.B(\register_file_i/_1140_ ),
    .C(\register_file_i/_1151_ ),
    .A(\register_file_i/_1133_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_mux2_1 \register_file_i/_4198_  (.A0(\register_file_i/rf_reg_915_ ),
    .A1(\register_file_i/rf_reg_947_ ),
    .S(net2048),
    .X(\register_file_i/_1152_ ));
 sg13g2_mux2_1 \register_file_i/_4199_  (.A0(\register_file_i/rf_reg_979_ ),
    .A1(\register_file_i/rf_reg_1011_ ),
    .S(net2047),
    .X(\register_file_i/_1153_ ));
 sg13g2_a22oi_1 \register_file_i/_4200_  (.Y(\register_file_i/_1154_ ),
    .B1(\register_file_i/_1153_ ),
    .B2(net1826),
    .A2(\register_file_i/_1152_ ),
    .A1(net1843));
 sg13g2_mux2_1 \register_file_i/_4201_  (.A0(\register_file_i/rf_reg_851_ ),
    .A1(\register_file_i/rf_reg_883_ ),
    .S(net2048),
    .X(\register_file_i/_1155_ ));
 sg13g2_mux2_1 \register_file_i/_4202_  (.A0(\register_file_i/rf_reg_787_ ),
    .A1(\register_file_i/rf_reg_819_ ),
    .S(net2048),
    .X(\register_file_i/_1156_ ));
 sg13g2_a22oi_1 \register_file_i/_4203_  (.Y(\register_file_i/_1157_ ),
    .B1(\register_file_i/_1156_ ),
    .B2(net1802),
    .A2(\register_file_i/_1155_ ),
    .A1(net1813));
 sg13g2_a21o_1 \register_file_i/_4204_  (.A2(\register_file_i/_1157_ ),
    .A1(\register_file_i/_1154_ ),
    .B1(net1928),
    .X(\register_file_i/_1158_ ));
 sg13g2_mux2_1 \register_file_i/_4205_  (.A0(\register_file_i/rf_reg_51_ ),
    .A1(\register_file_i/rf_reg_115_ ),
    .S(net533),
    .X(\register_file_i/_1159_ ));
 sg13g2_a22oi_1 \register_file_i/_4206_  (.Y(\register_file_i/_1160_ ),
    .B1(\register_file_i/_1159_ ),
    .B2(net2077),
    .A2(net1702),
    .A1(\register_file_i/rf_reg_83_ ));
 sg13g2_buf_2 fanout381 (.A(net384),
    .X(net381));
 sg13g2_mux2_1 \register_file_i/_4208_  (.A0(\register_file_i/rf_reg_211_ ),
    .A1(\register_file_i/rf_reg_243_ ),
    .S(net2081),
    .X(\register_file_i/_1162_ ));
 sg13g2_mux2_1 \register_file_i/_4209_  (.A0(\register_file_i/rf_reg_147_ ),
    .A1(\register_file_i/rf_reg_179_ ),
    .S(net2051),
    .X(\register_file_i/_1163_ ));
 sg13g2_a22oi_1 \register_file_i/_4210_  (.Y(\register_file_i/_1164_ ),
    .B1(\register_file_i/_1163_ ),
    .B2(net1852),
    .A2(\register_file_i/_1162_ ),
    .A1(net1835));
 sg13g2_o21ai_1 \register_file_i/_4211_  (.B1(\register_file_i/_1164_ ),
    .Y(\register_file_i/_1165_ ),
    .A1(net526),
    .A2(\register_file_i/_1160_ ));
 sg13g2_nand2_1 \register_file_i/_4212_  (.Y(\register_file_i/_1166_ ),
    .A(net1922),
    .B(\register_file_i/_1165_ ));
 sg13g2_buf_4 fanout380 (.X(net380),
    .A(net384));
 sg13g2_mux4_1 \register_file_i/_4214_  (.S0(net2035),
    .A0(\register_file_i/rf_reg_531_ ),
    .A1(\register_file_i/rf_reg_563_ ),
    .A2(\register_file_i/rf_reg_595_ ),
    .A3(\register_file_i/rf_reg_627_ ),
    .S1(net542),
    .X(\register_file_i/_1168_ ));
 sg13g2_mux4_1 \register_file_i/_4215_  (.S0(net2039),
    .A0(\register_file_i/rf_reg_659_ ),
    .A1(\register_file_i/rf_reg_691_ ),
    .A2(\register_file_i/rf_reg_723_ ),
    .A3(\register_file_i/rf_reg_755_ ),
    .S1(net540),
    .X(\register_file_i/_1169_ ));
 sg13g2_mux2_1 \register_file_i/_4216_  (.A0(\register_file_i/rf_reg_403_ ),
    .A1(\register_file_i/rf_reg_435_ ),
    .S(net2037),
    .X(\register_file_i/_1170_ ));
 sg13g2_mux2_1 \register_file_i/_4217_  (.A0(\register_file_i/rf_reg_467_ ),
    .A1(\register_file_i/rf_reg_499_ ),
    .S(net2036),
    .X(\register_file_i/_1171_ ));
 sg13g2_a22oi_1 \register_file_i/_4218_  (.Y(\register_file_i/_1172_ ),
    .B1(\register_file_i/_1171_ ),
    .B2(net1823),
    .A2(\register_file_i/_1170_ ),
    .A1(net1841));
 sg13g2_mux2_1 \register_file_i/_4219_  (.A0(\register_file_i/rf_reg_339_ ),
    .A1(\register_file_i/rf_reg_371_ ),
    .S(net2036),
    .X(\register_file_i/_1173_ ));
 sg13g2_mux2_1 \register_file_i/_4220_  (.A0(\register_file_i/rf_reg_275_ ),
    .A1(\register_file_i/rf_reg_307_ ),
    .S(net2040),
    .X(\register_file_i/_1174_ ));
 sg13g2_a22oi_1 \register_file_i/_4221_  (.Y(\register_file_i/_1175_ ),
    .B1(\register_file_i/_1174_ ),
    .B2(net1800),
    .A2(\register_file_i/_1173_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4222_  (.A1(\register_file_i/_1172_ ),
    .A2(\register_file_i/_1175_ ),
    .Y(\register_file_i/_1176_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4223_  (.B2(net1696),
    .C1(\register_file_i/_1176_ ),
    .B1(\register_file_i/_1169_ ),
    .A1(net1795),
    .Y(\register_file_i/_1177_ ),
    .A2(\register_file_i/_1168_ ));
 sg13g2_nand3_1 \register_file_i/_4224_  (.B(\register_file_i/_1166_ ),
    .C(\register_file_i/_1177_ ),
    .A(\register_file_i/_1158_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_19_ ));
 sg13g2_mux2_1 \register_file_i/_4225_  (.A0(\register_file_i/rf_reg_914_ ),
    .A1(\register_file_i/rf_reg_946_ ),
    .S(net2043),
    .X(\register_file_i/_1178_ ));
 sg13g2_mux2_1 \register_file_i/_4226_  (.A0(\register_file_i/rf_reg_978_ ),
    .A1(\register_file_i/rf_reg_1010_ ),
    .S(net2042),
    .X(\register_file_i/_1179_ ));
 sg13g2_a22oi_1 \register_file_i/_4227_  (.Y(\register_file_i/_1180_ ),
    .B1(\register_file_i/_1179_ ),
    .B2(net1825),
    .A2(\register_file_i/_1178_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4228_  (.A0(\register_file_i/rf_reg_850_ ),
    .A1(\register_file_i/rf_reg_882_ ),
    .S(net2043),
    .X(\register_file_i/_1181_ ));
 sg13g2_buf_4 fanout379 (.X(net379),
    .A(net384));
 sg13g2_mux2_1 \register_file_i/_4230_  (.A0(\register_file_i/rf_reg_786_ ),
    .A1(\register_file_i/rf_reg_818_ ),
    .S(net2043),
    .X(\register_file_i/_1183_ ));
 sg13g2_a22oi_1 \register_file_i/_4231_  (.Y(\register_file_i/_1184_ ),
    .B1(\register_file_i/_1183_ ),
    .B2(net1801),
    .A2(\register_file_i/_1181_ ),
    .A1(net1812));
 sg13g2_a21o_1 \register_file_i/_4232_  (.A2(\register_file_i/_1184_ ),
    .A1(\register_file_i/_1180_ ),
    .B1(net1928),
    .X(\register_file_i/_1185_ ));
 sg13g2_mux2_1 \register_file_i/_4233_  (.A0(\register_file_i/rf_reg_50_ ),
    .A1(\register_file_i/rf_reg_114_ ),
    .S(net532),
    .X(\register_file_i/_1186_ ));
 sg13g2_a22oi_1 \register_file_i/_4234_  (.Y(\register_file_i/_1187_ ),
    .B1(\register_file_i/_1186_ ),
    .B2(net2077),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_82_ ));
 sg13g2_mux2_1 \register_file_i/_4235_  (.A0(\register_file_i/rf_reg_210_ ),
    .A1(\register_file_i/rf_reg_242_ ),
    .S(net2077),
    .X(\register_file_i/_1188_ ));
 sg13g2_mux2_1 \register_file_i/_4236_  (.A0(\register_file_i/rf_reg_146_ ),
    .A1(\register_file_i/rf_reg_178_ ),
    .S(net2045),
    .X(\register_file_i/_1189_ ));
 sg13g2_a22oi_1 \register_file_i/_4237_  (.Y(\register_file_i/_1190_ ),
    .B1(\register_file_i/_1189_ ),
    .B2(net1851),
    .A2(\register_file_i/_1188_ ),
    .A1(net1825));
 sg13g2_o21ai_1 \register_file_i/_4238_  (.B1(\register_file_i/_1190_ ),
    .Y(\register_file_i/_1191_ ),
    .A1(net526),
    .A2(\register_file_i/_1187_ ));
 sg13g2_nand2_1 \register_file_i/_4239_  (.Y(\register_file_i/_1192_ ),
    .A(net1922),
    .B(\register_file_i/_1191_ ));
 sg13g2_mux4_1 \register_file_i/_4240_  (.S0(net2034),
    .A0(\register_file_i/rf_reg_530_ ),
    .A1(\register_file_i/rf_reg_562_ ),
    .A2(\register_file_i/rf_reg_594_ ),
    .A3(\register_file_i/rf_reg_626_ ),
    .S1(net542),
    .X(\register_file_i/_1193_ ));
 sg13g2_buf_4 fanout378 (.X(net378),
    .A(net384));
 sg13g2_mux4_1 \register_file_i/_4242_  (.S0(net2035),
    .A0(\register_file_i/rf_reg_658_ ),
    .A1(\register_file_i/rf_reg_690_ ),
    .A2(\register_file_i/rf_reg_722_ ),
    .A3(\register_file_i/rf_reg_754_ ),
    .S1(net540),
    .X(\register_file_i/_1195_ ));
 sg13g2_mux2_1 \register_file_i/_4243_  (.A0(\register_file_i/rf_reg_402_ ),
    .A1(\register_file_i/rf_reg_434_ ),
    .S(net2032),
    .X(\register_file_i/_1196_ ));
 sg13g2_buf_1 fanout377 (.A(net382),
    .X(net377));
 sg13g2_mux2_1 \register_file_i/_4245_  (.A0(\register_file_i/rf_reg_466_ ),
    .A1(\register_file_i/rf_reg_498_ ),
    .S(net2032),
    .X(\register_file_i/_1198_ ));
 sg13g2_a22oi_1 \register_file_i/_4246_  (.Y(\register_file_i/_1199_ ),
    .B1(\register_file_i/_1198_ ),
    .B2(net1823),
    .A2(\register_file_i/_1196_ ),
    .A1(net1840));
 sg13g2_mux2_1 \register_file_i/_4247_  (.A0(\register_file_i/rf_reg_338_ ),
    .A1(\register_file_i/rf_reg_370_ ),
    .S(net2037),
    .X(\register_file_i/_1200_ ));
 sg13g2_mux2_1 \register_file_i/_4248_  (.A0(\register_file_i/rf_reg_274_ ),
    .A1(\register_file_i/rf_reg_306_ ),
    .S(net2032),
    .X(\register_file_i/_1201_ ));
 sg13g2_a22oi_1 \register_file_i/_4249_  (.Y(\register_file_i/_1202_ ),
    .B1(\register_file_i/_1201_ ),
    .B2(net1800),
    .A2(\register_file_i/_1200_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4250_  (.A1(\register_file_i/_1199_ ),
    .A2(\register_file_i/_1202_ ),
    .Y(\register_file_i/_1203_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4251_  (.B2(net1696),
    .C1(\register_file_i/_1203_ ),
    .B1(\register_file_i/_1195_ ),
    .A1(net1795),
    .Y(\register_file_i/_1204_ ),
    .A2(\register_file_i/_1193_ ));
 sg13g2_nand3_1 \register_file_i/_4252_  (.B(\register_file_i/_1192_ ),
    .C(\register_file_i/_1204_ ),
    .A(\register_file_i/_1185_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_18_ ));
 sg13g2_mux2_1 \register_file_i/_4253_  (.A0(\register_file_i/rf_reg_913_ ),
    .A1(\register_file_i/rf_reg_945_ ),
    .S(net2050),
    .X(\register_file_i/_1205_ ));
 sg13g2_mux2_1 \register_file_i/_4254_  (.A0(\register_file_i/rf_reg_977_ ),
    .A1(\register_file_i/rf_reg_1009_ ),
    .S(net2050),
    .X(\register_file_i/_1206_ ));
 sg13g2_a22oi_1 \register_file_i/_4255_  (.Y(\register_file_i/_1207_ ),
    .B1(\register_file_i/_1206_ ),
    .B2(net1826),
    .A2(\register_file_i/_1205_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4256_  (.A0(\register_file_i/rf_reg_849_ ),
    .A1(\register_file_i/rf_reg_881_ ),
    .S(net2049),
    .X(\register_file_i/_1208_ ));
 sg13g2_mux2_1 \register_file_i/_4257_  (.A0(\register_file_i/rf_reg_785_ ),
    .A1(\register_file_i/rf_reg_817_ ),
    .S(net2049),
    .X(\register_file_i/_1209_ ));
 sg13g2_a22oi_1 \register_file_i/_4258_  (.Y(\register_file_i/_1210_ ),
    .B1(\register_file_i/_1209_ ),
    .B2(net1801),
    .A2(\register_file_i/_1208_ ),
    .A1(net1812));
 sg13g2_a21o_1 \register_file_i/_4259_  (.A2(\register_file_i/_1210_ ),
    .A1(\register_file_i/_1207_ ),
    .B1(net1928),
    .X(\register_file_i/_1211_ ));
 sg13g2_mux2_1 \register_file_i/_4260_  (.A0(\register_file_i/rf_reg_49_ ),
    .A1(\register_file_i/rf_reg_113_ ),
    .S(net532),
    .X(\register_file_i/_1212_ ));
 sg13g2_a22oi_1 \register_file_i/_4261_  (.Y(\register_file_i/_1213_ ),
    .B1(\register_file_i/_1212_ ),
    .B2(net2077),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_81_ ));
 sg13g2_mux2_1 \register_file_i/_4262_  (.A0(\register_file_i/rf_reg_209_ ),
    .A1(\register_file_i/rf_reg_241_ ),
    .S(net2081),
    .X(\register_file_i/_1214_ ));
 sg13g2_mux2_1 \register_file_i/_4263_  (.A0(\register_file_i/rf_reg_145_ ),
    .A1(\register_file_i/rf_reg_177_ ),
    .S(net2081),
    .X(\register_file_i/_1215_ ));
 sg13g2_a22oi_1 \register_file_i/_4264_  (.Y(\register_file_i/_1216_ ),
    .B1(\register_file_i/_1215_ ),
    .B2(net1852),
    .A2(\register_file_i/_1214_ ),
    .A1(net1835));
 sg13g2_o21ai_1 \register_file_i/_4265_  (.B1(\register_file_i/_1216_ ),
    .Y(\register_file_i/_1217_ ),
    .A1(net526),
    .A2(\register_file_i/_1213_ ));
 sg13g2_nand2_1 \register_file_i/_4266_  (.Y(\register_file_i/_1218_ ),
    .A(net1922),
    .B(\register_file_i/_1217_ ));
 sg13g2_buf_2 fanout376 (.A(net382),
    .X(net376));
 sg13g2_mux4_1 \register_file_i/_4268_  (.S0(net2034),
    .A0(\register_file_i/rf_reg_529_ ),
    .A1(\register_file_i/rf_reg_561_ ),
    .A2(\register_file_i/rf_reg_593_ ),
    .A3(\register_file_i/rf_reg_625_ ),
    .S1(net541),
    .X(\register_file_i/_1220_ ));
 sg13g2_mux4_1 \register_file_i/_4269_  (.S0(net2039),
    .A0(\register_file_i/rf_reg_657_ ),
    .A1(\register_file_i/rf_reg_689_ ),
    .A2(\register_file_i/rf_reg_721_ ),
    .A3(\register_file_i/rf_reg_753_ ),
    .S1(net540),
    .X(\register_file_i/_1221_ ));
 sg13g2_mux2_1 \register_file_i/_4270_  (.A0(\register_file_i/rf_reg_401_ ),
    .A1(\register_file_i/rf_reg_433_ ),
    .S(net2037),
    .X(\register_file_i/_1222_ ));
 sg13g2_mux2_1 \register_file_i/_4271_  (.A0(\register_file_i/rf_reg_465_ ),
    .A1(\register_file_i/rf_reg_497_ ),
    .S(net2037),
    .X(\register_file_i/_1223_ ));
 sg13g2_a22oi_1 \register_file_i/_4272_  (.Y(\register_file_i/_1224_ ),
    .B1(\register_file_i/_1223_ ),
    .B2(net1823),
    .A2(\register_file_i/_1222_ ),
    .A1(net1841));
 sg13g2_mux2_1 \register_file_i/_4273_  (.A0(\register_file_i/rf_reg_337_ ),
    .A1(\register_file_i/rf_reg_369_ ),
    .S(net2037),
    .X(\register_file_i/_1225_ ));
 sg13g2_mux2_1 \register_file_i/_4274_  (.A0(\register_file_i/rf_reg_273_ ),
    .A1(\register_file_i/rf_reg_305_ ),
    .S(net2037),
    .X(\register_file_i/_1226_ ));
 sg13g2_a22oi_1 \register_file_i/_4275_  (.Y(\register_file_i/_1227_ ),
    .B1(\register_file_i/_1226_ ),
    .B2(net1800),
    .A2(\register_file_i/_1225_ ),
    .A1(net1811));
 sg13g2_buf_2 fanout375 (.A(net382),
    .X(net375));
 sg13g2_a21oi_1 \register_file_i/_4277_  (.A1(\register_file_i/_1224_ ),
    .A2(\register_file_i/_1227_ ),
    .Y(\register_file_i/_1229_ ),
    .B1(net1791));
 sg13g2_a221oi_1 \register_file_i/_4278_  (.B2(net1696),
    .C1(\register_file_i/_1229_ ),
    .B1(\register_file_i/_1221_ ),
    .A1(net1796),
    .Y(\register_file_i/_1230_ ),
    .A2(\register_file_i/_1220_ ));
 sg13g2_nand3_1 \register_file_i/_4279_  (.B(\register_file_i/_1218_ ),
    .C(\register_file_i/_1230_ ),
    .A(\register_file_i/_1211_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_17_ ));
 sg13g2_mux2_1 \register_file_i/_4280_  (.A0(\register_file_i/rf_reg_912_ ),
    .A1(\register_file_i/rf_reg_944_ ),
    .S(net2045),
    .X(\register_file_i/_1231_ ));
 sg13g2_mux2_1 \register_file_i/_4281_  (.A0(\register_file_i/rf_reg_976_ ),
    .A1(\register_file_i/rf_reg_1008_ ),
    .S(net2045),
    .X(\register_file_i/_1232_ ));
 sg13g2_a22oi_1 \register_file_i/_4282_  (.Y(\register_file_i/_1233_ ),
    .B1(\register_file_i/_1232_ ),
    .B2(net1825),
    .A2(\register_file_i/_1231_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4283_  (.A0(\register_file_i/rf_reg_848_ ),
    .A1(\register_file_i/rf_reg_880_ ),
    .S(net2045),
    .X(\register_file_i/_1234_ ));
 sg13g2_mux2_1 \register_file_i/_4284_  (.A0(\register_file_i/rf_reg_784_ ),
    .A1(\register_file_i/rf_reg_816_ ),
    .S(net2045),
    .X(\register_file_i/_1235_ ));
 sg13g2_a22oi_1 \register_file_i/_4285_  (.Y(\register_file_i/_1236_ ),
    .B1(\register_file_i/_1235_ ),
    .B2(net1801),
    .A2(\register_file_i/_1234_ ),
    .A1(net1812));
 sg13g2_a21o_1 \register_file_i/_4286_  (.A2(\register_file_i/_1236_ ),
    .A1(\register_file_i/_1233_ ),
    .B1(net1928),
    .X(\register_file_i/_1237_ ));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(net382));
 sg13g2_mux2_1 \register_file_i/_4288_  (.A0(\register_file_i/rf_reg_48_ ),
    .A1(\register_file_i/rf_reg_112_ ),
    .S(net534),
    .X(\register_file_i/_1239_ ));
 sg13g2_a22oi_1 \register_file_i/_4289_  (.Y(\register_file_i/_1240_ ),
    .B1(\register_file_i/_1239_ ),
    .B2(net2076),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_80_ ));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(net382));
 sg13g2_mux2_1 \register_file_i/_4291_  (.A0(\register_file_i/rf_reg_208_ ),
    .A1(\register_file_i/rf_reg_240_ ),
    .S(net2076),
    .X(\register_file_i/_1242_ ));
 sg13g2_mux2_1 \register_file_i/_4292_  (.A0(\register_file_i/rf_reg_144_ ),
    .A1(\register_file_i/rf_reg_176_ ),
    .S(net2044),
    .X(\register_file_i/_1243_ ));
 sg13g2_a22oi_1 \register_file_i/_4293_  (.Y(\register_file_i/_1244_ ),
    .B1(\register_file_i/_1243_ ),
    .B2(net1851),
    .A2(\register_file_i/_1242_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4294_  (.B1(\register_file_i/_1244_ ),
    .Y(\register_file_i/_1245_ ),
    .A1(net526),
    .A2(\register_file_i/_1240_ ));
 sg13g2_nand2_1 \register_file_i/_4295_  (.Y(\register_file_i/_1246_ ),
    .A(net1922),
    .B(\register_file_i/_1245_ ));
 sg13g2_mux4_1 \register_file_i/_4296_  (.S0(net2033),
    .A0(\register_file_i/rf_reg_528_ ),
    .A1(\register_file_i/rf_reg_560_ ),
    .A2(\register_file_i/rf_reg_592_ ),
    .A3(\register_file_i/rf_reg_624_ ),
    .S1(net541),
    .X(\register_file_i/_1247_ ));
 sg13g2_mux4_1 \register_file_i/_4297_  (.S0(net2035),
    .A0(\register_file_i/rf_reg_656_ ),
    .A1(\register_file_i/rf_reg_688_ ),
    .A2(\register_file_i/rf_reg_720_ ),
    .A3(\register_file_i/rf_reg_752_ ),
    .S1(net540),
    .X(\register_file_i/_1248_ ));
 sg13g2_mux2_1 \register_file_i/_4298_  (.A0(\register_file_i/rf_reg_400_ ),
    .A1(\register_file_i/rf_reg_432_ ),
    .S(net2032),
    .X(\register_file_i/_1249_ ));
 sg13g2_mux2_1 \register_file_i/_4299_  (.A0(\register_file_i/rf_reg_464_ ),
    .A1(\register_file_i/rf_reg_496_ ),
    .S(net2032),
    .X(\register_file_i/_1250_ ));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net382));
 sg13g2_a22oi_1 \register_file_i/_4301_  (.Y(\register_file_i/_1252_ ),
    .B1(\register_file_i/_1250_ ),
    .B2(net1824),
    .A2(\register_file_i/_1249_ ),
    .A1(net1840));
 sg13g2_mux2_1 \register_file_i/_4302_  (.A0(\register_file_i/rf_reg_336_ ),
    .A1(\register_file_i/rf_reg_368_ ),
    .S(net2037),
    .X(\register_file_i/_1253_ ));
 sg13g2_mux2_1 \register_file_i/_4303_  (.A0(\register_file_i/rf_reg_272_ ),
    .A1(\register_file_i/rf_reg_304_ ),
    .S(net2037),
    .X(\register_file_i/_1254_ ));
 sg13g2_a22oi_1 \register_file_i/_4304_  (.Y(\register_file_i/_1255_ ),
    .B1(\register_file_i/_1254_ ),
    .B2(net1800),
    .A2(\register_file_i/_1253_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4305_  (.A1(\register_file_i/_1252_ ),
    .A2(\register_file_i/_1255_ ),
    .Y(\register_file_i/_1256_ ),
    .B1(net1791));
 sg13g2_a221oi_1 \register_file_i/_4306_  (.B2(net1696),
    .C1(\register_file_i/_1256_ ),
    .B1(\register_file_i/_1248_ ),
    .A1(net1796),
    .Y(\register_file_i/_1257_ ),
    .A2(\register_file_i/_1247_ ));
 sg13g2_nand3_1 \register_file_i/_4307_  (.B(\register_file_i/_1246_ ),
    .C(\register_file_i/_1257_ ),
    .A(\register_file_i/_1237_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_16_ ));
 sg13g2_mux2_1 \register_file_i/_4308_  (.A0(\register_file_i/rf_reg_911_ ),
    .A1(\register_file_i/rf_reg_943_ ),
    .S(net2044),
    .X(\register_file_i/_1258_ ));
 sg13g2_buf_2 fanout371 (.A(net382),
    .X(net371));
 sg13g2_mux2_1 \register_file_i/_4310_  (.A0(\register_file_i/rf_reg_975_ ),
    .A1(\register_file_i/rf_reg_1007_ ),
    .S(net2044),
    .X(\register_file_i/_1260_ ));
 sg13g2_a22oi_1 \register_file_i/_4311_  (.Y(\register_file_i/_1261_ ),
    .B1(\register_file_i/_1260_ ),
    .B2(net1825),
    .A2(\register_file_i/_1258_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4312_  (.A0(\register_file_i/rf_reg_847_ ),
    .A1(\register_file_i/rf_reg_879_ ),
    .S(net2044),
    .X(\register_file_i/_1262_ ));
 sg13g2_mux2_1 \register_file_i/_4313_  (.A0(\register_file_i/rf_reg_783_ ),
    .A1(\register_file_i/rf_reg_815_ ),
    .S(net2046),
    .X(\register_file_i/_1263_ ));
 sg13g2_a22oi_1 \register_file_i/_4314_  (.Y(\register_file_i/_1264_ ),
    .B1(\register_file_i/_1263_ ),
    .B2(net1807),
    .A2(\register_file_i/_1262_ ),
    .A1(net1818));
 sg13g2_a21o_1 \register_file_i/_4315_  (.A2(\register_file_i/_1264_ ),
    .A1(\register_file_i/_1261_ ),
    .B1(net1928),
    .X(\register_file_i/_1265_ ));
 sg13g2_mux2_1 \register_file_i/_4316_  (.A0(\register_file_i/rf_reg_47_ ),
    .A1(\register_file_i/rf_reg_111_ ),
    .S(net534),
    .X(\register_file_i/_1266_ ));
 sg13g2_a22oi_1 \register_file_i/_4317_  (.Y(\register_file_i/_1267_ ),
    .B1(\register_file_i/_1266_ ),
    .B2(net2076),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_79_ ));
 sg13g2_mux2_1 \register_file_i/_4318_  (.A0(\register_file_i/rf_reg_207_ ),
    .A1(\register_file_i/rf_reg_239_ ),
    .S(net2076),
    .X(\register_file_i/_1268_ ));
 sg13g2_mux2_1 \register_file_i/_4319_  (.A0(\register_file_i/rf_reg_143_ ),
    .A1(\register_file_i/rf_reg_175_ ),
    .S(net2077),
    .X(\register_file_i/_1269_ ));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(net382));
 sg13g2_a22oi_1 \register_file_i/_4321_  (.Y(\register_file_i/_1271_ ),
    .B1(\register_file_i/_1269_ ),
    .B2(net1851),
    .A2(\register_file_i/_1268_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4322_  (.B1(\register_file_i/_1271_ ),
    .Y(\register_file_i/_1272_ ),
    .A1(net526),
    .A2(\register_file_i/_1267_ ));
 sg13g2_nand2_1 \register_file_i/_4323_  (.Y(\register_file_i/_1273_ ),
    .A(net1922),
    .B(\register_file_i/_1272_ ));
 sg13g2_mux4_1 \register_file_i/_4324_  (.S0(net2032),
    .A0(\register_file_i/rf_reg_527_ ),
    .A1(\register_file_i/rf_reg_559_ ),
    .A2(\register_file_i/rf_reg_591_ ),
    .A3(\register_file_i/rf_reg_623_ ),
    .S1(net541),
    .X(\register_file_i/_1274_ ));
 sg13g2_mux4_1 \register_file_i/_4325_  (.S0(net2035),
    .A0(\register_file_i/rf_reg_655_ ),
    .A1(\register_file_i/rf_reg_687_ ),
    .A2(\register_file_i/rf_reg_719_ ),
    .A3(\register_file_i/rf_reg_751_ ),
    .S1(net540),
    .X(\register_file_i/_1275_ ));
 sg13g2_mux2_1 \register_file_i/_4326_  (.A0(\register_file_i/rf_reg_399_ ),
    .A1(\register_file_i/rf_reg_431_ ),
    .S(net2031),
    .X(\register_file_i/_1276_ ));
 sg13g2_mux2_1 \register_file_i/_4327_  (.A0(\register_file_i/rf_reg_463_ ),
    .A1(\register_file_i/rf_reg_495_ ),
    .S(net2031),
    .X(\register_file_i/_1277_ ));
 sg13g2_a22oi_1 \register_file_i/_4328_  (.Y(\register_file_i/_1278_ ),
    .B1(\register_file_i/_1277_ ),
    .B2(net1823),
    .A2(\register_file_i/_1276_ ),
    .A1(net1840));
 sg13g2_mux2_1 \register_file_i/_4329_  (.A0(\register_file_i/rf_reg_335_ ),
    .A1(\register_file_i/rf_reg_367_ ),
    .S(net2032),
    .X(\register_file_i/_1279_ ));
 sg13g2_mux2_1 \register_file_i/_4330_  (.A0(\register_file_i/rf_reg_271_ ),
    .A1(\register_file_i/rf_reg_303_ ),
    .S(net2032),
    .X(\register_file_i/_1280_ ));
 sg13g2_buf_2 fanout369 (.A(net383),
    .X(net369));
 sg13g2_a22oi_1 \register_file_i/_4332_  (.Y(\register_file_i/_1282_ ),
    .B1(\register_file_i/_1280_ ),
    .B2(net1800),
    .A2(\register_file_i/_1279_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4333_  (.A1(\register_file_i/_1278_ ),
    .A2(\register_file_i/_1282_ ),
    .Y(\register_file_i/_1283_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4334_  (.B2(net1696),
    .C1(\register_file_i/_1283_ ),
    .B1(\register_file_i/_1275_ ),
    .A1(net1795),
    .Y(\register_file_i/_1284_ ),
    .A2(\register_file_i/_1274_ ));
 sg13g2_nand3_1 \register_file_i/_4335_  (.B(\register_file_i/_1273_ ),
    .C(\register_file_i/_1284_ ),
    .A(\register_file_i/_1265_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_mux2_1 \register_file_i/_4336_  (.A0(\register_file_i/rf_reg_910_ ),
    .A1(\register_file_i/rf_reg_942_ ),
    .S(net2044),
    .X(\register_file_i/_1285_ ));
 sg13g2_mux2_1 \register_file_i/_4337_  (.A0(\register_file_i/rf_reg_974_ ),
    .A1(\register_file_i/rf_reg_1006_ ),
    .S(net2044),
    .X(\register_file_i/_1286_ ));
 sg13g2_a22oi_1 \register_file_i/_4338_  (.Y(\register_file_i/_1287_ ),
    .B1(\register_file_i/_1286_ ),
    .B2(net1825),
    .A2(\register_file_i/_1285_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4339_  (.A0(\register_file_i/rf_reg_846_ ),
    .A1(\register_file_i/rf_reg_878_ ),
    .S(net2044),
    .X(\register_file_i/_1288_ ));
 sg13g2_mux2_1 \register_file_i/_4340_  (.A0(\register_file_i/rf_reg_782_ ),
    .A1(\register_file_i/rf_reg_814_ ),
    .S(net2044),
    .X(\register_file_i/_1289_ ));
 sg13g2_a22oi_1 \register_file_i/_4341_  (.Y(\register_file_i/_1290_ ),
    .B1(\register_file_i/_1289_ ),
    .B2(net1801),
    .A2(\register_file_i/_1288_ ),
    .A1(net1812));
 sg13g2_a21o_1 \register_file_i/_4342_  (.A2(\register_file_i/_1290_ ),
    .A1(\register_file_i/_1287_ ),
    .B1(net1928),
    .X(\register_file_i/_1291_ ));
 sg13g2_mux2_1 \register_file_i/_4343_  (.A0(\register_file_i/rf_reg_46_ ),
    .A1(\register_file_i/rf_reg_110_ ),
    .S(net534),
    .X(\register_file_i/_1292_ ));
 sg13g2_a22oi_1 \register_file_i/_4344_  (.Y(\register_file_i/_1293_ ),
    .B1(\register_file_i/_1292_ ),
    .B2(net2076),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_78_ ));
 sg13g2_mux2_1 \register_file_i/_4345_  (.A0(\register_file_i/rf_reg_206_ ),
    .A1(\register_file_i/rf_reg_238_ ),
    .S(net2076),
    .X(\register_file_i/_1294_ ));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(net383));
 sg13g2_mux2_1 \register_file_i/_4347_  (.A0(\register_file_i/rf_reg_142_ ),
    .A1(\register_file_i/rf_reg_174_ ),
    .S(net2046),
    .X(\register_file_i/_1296_ ));
 sg13g2_a22oi_1 \register_file_i/_4348_  (.Y(\register_file_i/_1297_ ),
    .B1(\register_file_i/_1296_ ),
    .B2(net1851),
    .A2(\register_file_i/_1294_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4349_  (.B1(\register_file_i/_1297_ ),
    .Y(\register_file_i/_1298_ ),
    .A1(net526),
    .A2(\register_file_i/_1293_ ));
 sg13g2_nand2_1 \register_file_i/_4350_  (.Y(\register_file_i/_1299_ ),
    .A(net1923),
    .B(\register_file_i/_1298_ ));
 sg13g2_mux4_1 \register_file_i/_4351_  (.S0(net2033),
    .A0(\register_file_i/rf_reg_526_ ),
    .A1(\register_file_i/rf_reg_558_ ),
    .A2(\register_file_i/rf_reg_590_ ),
    .A3(\register_file_i/rf_reg_622_ ),
    .S1(net541),
    .X(\register_file_i/_1300_ ));
 sg13g2_mux4_1 \register_file_i/_4352_  (.S0(net2034),
    .A0(\register_file_i/rf_reg_654_ ),
    .A1(\register_file_i/rf_reg_686_ ),
    .A2(\register_file_i/rf_reg_718_ ),
    .A3(\register_file_i/rf_reg_750_ ),
    .S1(net539),
    .X(\register_file_i/_1301_ ));
 sg13g2_mux2_1 \register_file_i/_4353_  (.A0(\register_file_i/rf_reg_398_ ),
    .A1(\register_file_i/rf_reg_430_ ),
    .S(net2031),
    .X(\register_file_i/_1302_ ));
 sg13g2_mux2_1 \register_file_i/_4354_  (.A0(\register_file_i/rf_reg_462_ ),
    .A1(\register_file_i/rf_reg_494_ ),
    .S(net2031),
    .X(\register_file_i/_1303_ ));
 sg13g2_a22oi_1 \register_file_i/_4355_  (.Y(\register_file_i/_1304_ ),
    .B1(\register_file_i/_1303_ ),
    .B2(net1823),
    .A2(\register_file_i/_1302_ ),
    .A1(net1840));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(net383));
 sg13g2_buf_4 fanout366 (.X(net366),
    .A(net383));
 sg13g2_mux2_1 \register_file_i/_4358_  (.A0(\register_file_i/rf_reg_334_ ),
    .A1(\register_file_i/rf_reg_366_ ),
    .S(net2031),
    .X(\register_file_i/_1307_ ));
 sg13g2_mux2_1 \register_file_i/_4359_  (.A0(\register_file_i/rf_reg_270_ ),
    .A1(\register_file_i/rf_reg_302_ ),
    .S(net2031),
    .X(\register_file_i/_1308_ ));
 sg13g2_a22oi_1 \register_file_i/_4360_  (.Y(\register_file_i/_1309_ ),
    .B1(\register_file_i/_1308_ ),
    .B2(net1800),
    .A2(\register_file_i/_1307_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4361_  (.A1(\register_file_i/_1304_ ),
    .A2(\register_file_i/_1309_ ),
    .Y(\register_file_i/_1310_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4362_  (.B2(net1696),
    .C1(\register_file_i/_1310_ ),
    .B1(\register_file_i/_1301_ ),
    .A1(net1795),
    .Y(\register_file_i/_1311_ ),
    .A2(\register_file_i/_1300_ ));
 sg13g2_nand3_1 \register_file_i/_4363_  (.B(\register_file_i/_1299_ ),
    .C(\register_file_i/_1311_ ),
    .A(\register_file_i/_1291_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_14_ ));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net383));
 sg13g2_mux2_1 \register_file_i/_4365_  (.A0(\register_file_i/rf_reg_909_ ),
    .A1(\register_file_i/rf_reg_941_ ),
    .S(net2027),
    .X(\register_file_i/_1313_ ));
 sg13g2_mux2_1 \register_file_i/_4366_  (.A0(\register_file_i/rf_reg_973_ ),
    .A1(\register_file_i/rf_reg_1005_ ),
    .S(net2027),
    .X(\register_file_i/_1314_ ));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net383));
 sg13g2_a22oi_1 \register_file_i/_4368_  (.Y(\register_file_i/_1316_ ),
    .B1(\register_file_i/_1314_ ),
    .B2(net1822),
    .A2(\register_file_i/_1313_ ),
    .A1(net1838));
 sg13g2_buf_4 fanout363 (.X(net363),
    .A(net383));
 sg13g2_mux2_1 \register_file_i/_4370_  (.A0(\register_file_i/rf_reg_845_ ),
    .A1(\register_file_i/rf_reg_877_ ),
    .S(net2027),
    .X(\register_file_i/_1318_ ));
 sg13g2_mux2_1 \register_file_i/_4371_  (.A0(\register_file_i/rf_reg_781_ ),
    .A1(\register_file_i/rf_reg_813_ ),
    .S(net2027),
    .X(\register_file_i/_1319_ ));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net383));
 sg13g2_a22oi_1 \register_file_i/_4373_  (.Y(\register_file_i/_1321_ ),
    .B1(\register_file_i/_1319_ ),
    .B2(net1801),
    .A2(\register_file_i/_1318_ ),
    .A1(net1812));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net384));
 sg13g2_a21o_1 \register_file_i/_4375_  (.A2(\register_file_i/_1321_ ),
    .A1(\register_file_i/_1316_ ),
    .B1(net1928),
    .X(\register_file_i/_1323_ ));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net1616));
 sg13g2_buf_4 fanout359 (.X(net359),
    .A(net1615));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(net1616));
 sg13g2_mux2_1 \register_file_i/_4379_  (.A0(\register_file_i/rf_reg_45_ ),
    .A1(\register_file_i/rf_reg_109_ ),
    .S(net534),
    .X(\register_file_i/_1327_ ));
 sg13g2_a22oi_1 \register_file_i/_4380_  (.Y(\register_file_i/_1328_ ),
    .B1(\register_file_i/_1327_ ),
    .B2(net2076),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_77_ ));
 sg13g2_mux2_1 \register_file_i/_4381_  (.A0(\register_file_i/rf_reg_205_ ),
    .A1(\register_file_i/rf_reg_237_ ),
    .S(net2078),
    .X(\register_file_i/_1329_ ));
 sg13g2_mux2_1 \register_file_i/_4382_  (.A0(\register_file_i/rf_reg_141_ ),
    .A1(\register_file_i/rf_reg_173_ ),
    .S(net2076),
    .X(\register_file_i/_1330_ ));
 sg13g2_a22oi_1 \register_file_i/_4383_  (.Y(\register_file_i/_1331_ ),
    .B1(\register_file_i/_1330_ ),
    .B2(net1851),
    .A2(\register_file_i/_1329_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4384_  (.B1(\register_file_i/_1331_ ),
    .Y(\register_file_i/_1332_ ),
    .A1(net528),
    .A2(\register_file_i/_1328_ ));
 sg13g2_nand2_1 \register_file_i/_4385_  (.Y(\register_file_i/_1333_ ),
    .A(net1923),
    .B(\register_file_i/_1332_ ));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(net1615));
 sg13g2_mux4_1 \register_file_i/_4387_  (.S0(net2016),
    .A0(\register_file_i/rf_reg_525_ ),
    .A1(\register_file_i/rf_reg_557_ ),
    .A2(\register_file_i/rf_reg_589_ ),
    .A3(\register_file_i/rf_reg_621_ ),
    .S1(net541),
    .X(\register_file_i/_1335_ ));
 sg13g2_mux4_1 \register_file_i/_4388_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_653_ ),
    .A1(\register_file_i/rf_reg_685_ ),
    .A2(\register_file_i/rf_reg_717_ ),
    .A3(\register_file_i/rf_reg_749_ ),
    .S1(net539),
    .X(\register_file_i/_1336_ ));
 sg13g2_buf_2 fanout356 (.A(net1616),
    .X(net356));
 sg13g2_mux2_1 \register_file_i/_4390_  (.A0(\register_file_i/rf_reg_397_ ),
    .A1(\register_file_i/rf_reg_429_ ),
    .S(net2031),
    .X(\register_file_i/_1338_ ));
 sg13g2_mux2_1 \register_file_i/_4391_  (.A0(\register_file_i/rf_reg_461_ ),
    .A1(\register_file_i/rf_reg_493_ ),
    .S(net2031),
    .X(\register_file_i/_1339_ ));
 sg13g2_a22oi_1 \register_file_i/_4392_  (.Y(\register_file_i/_1340_ ),
    .B1(\register_file_i/_1339_ ),
    .B2(net1823),
    .A2(\register_file_i/_1338_ ),
    .A1(net1840));
 sg13g2_mux2_1 \register_file_i/_4393_  (.A0(\register_file_i/rf_reg_333_ ),
    .A1(\register_file_i/rf_reg_365_ ),
    .S(net2014),
    .X(\register_file_i/_1341_ ));
 sg13g2_mux2_1 \register_file_i/_4394_  (.A0(\register_file_i/rf_reg_269_ ),
    .A1(\register_file_i/rf_reg_301_ ),
    .S(net2014),
    .X(\register_file_i/_1342_ ));
 sg13g2_a22oi_1 \register_file_i/_4395_  (.Y(\register_file_i/_1343_ ),
    .B1(\register_file_i/_1342_ ),
    .B2(net1800),
    .A2(\register_file_i/_1341_ ),
    .A1(net1811));
 sg13g2_a21oi_1 \register_file_i/_4396_  (.A1(\register_file_i/_1340_ ),
    .A2(\register_file_i/_1343_ ),
    .Y(\register_file_i/_1344_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4397_  (.B2(net1693),
    .C1(\register_file_i/_1344_ ),
    .B1(\register_file_i/_1336_ ),
    .A1(net1792),
    .Y(\register_file_i/_1345_ ),
    .A2(\register_file_i/_1335_ ));
 sg13g2_nand3_1 \register_file_i/_4398_  (.B(\register_file_i/_1333_ ),
    .C(\register_file_i/_1345_ ),
    .A(\register_file_i/_1323_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_mux2_1 \register_file_i/_4399_  (.A0(\register_file_i/rf_reg_908_ ),
    .A1(\register_file_i/rf_reg_940_ ),
    .S(net2053),
    .X(\register_file_i/_1346_ ));
 sg13g2_mux2_1 \register_file_i/_4400_  (.A0(\register_file_i/rf_reg_972_ ),
    .A1(\register_file_i/rf_reg_1004_ ),
    .S(net2053),
    .X(\register_file_i/_1347_ ));
 sg13g2_a22oi_1 \register_file_i/_4401_  (.Y(\register_file_i/_1348_ ),
    .B1(\register_file_i/_1347_ ),
    .B2(net1828),
    .A2(\register_file_i/_1346_ ),
    .A1(net1845));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net1616));
 sg13g2_mux2_1 \register_file_i/_4403_  (.A0(\register_file_i/rf_reg_844_ ),
    .A1(\register_file_i/rf_reg_876_ ),
    .S(net2055),
    .X(\register_file_i/_1350_ ));
 sg13g2_mux2_1 \register_file_i/_4404_  (.A0(\register_file_i/rf_reg_780_ ),
    .A1(\register_file_i/rf_reg_812_ ),
    .S(net2053),
    .X(\register_file_i/_1351_ ));
 sg13g2_a22oi_1 \register_file_i/_4405_  (.Y(\register_file_i/_1352_ ),
    .B1(\register_file_i/_1351_ ),
    .B2(net1804),
    .A2(\register_file_i/_1350_ ),
    .A1(net1815));
 sg13g2_a21o_1 \register_file_i/_4406_  (.A2(\register_file_i/_1352_ ),
    .A1(\register_file_i/_1348_ ),
    .B1(net1927),
    .X(\register_file_i/_1353_ ));
 sg13g2_mux2_1 \register_file_i/_4407_  (.A0(\register_file_i/rf_reg_44_ ),
    .A1(\register_file_i/rf_reg_108_ ),
    .S(net534),
    .X(\register_file_i/_1354_ ));
 sg13g2_buf_4 fanout354 (.X(net354),
    .A(net1616));
 sg13g2_a22oi_1 \register_file_i/_4409_  (.Y(\register_file_i/_1356_ ),
    .B1(\register_file_i/_1354_ ),
    .B2(net2062),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_76_ ));
 sg13g2_mux2_1 \register_file_i/_4410_  (.A0(\register_file_i/rf_reg_204_ ),
    .A1(\register_file_i/rf_reg_236_ ),
    .S(net2062),
    .X(\register_file_i/_1357_ ));
 sg13g2_mux2_1 \register_file_i/_4411_  (.A0(\register_file_i/rf_reg_140_ ),
    .A1(\register_file_i/rf_reg_172_ ),
    .S(net2062),
    .X(\register_file_i/_1358_ ));
 sg13g2_a22oi_1 \register_file_i/_4412_  (.Y(\register_file_i/_1359_ ),
    .B1(\register_file_i/_1358_ ),
    .B2(net1847),
    .A2(\register_file_i/_1357_ ),
    .A1(net1830));
 sg13g2_o21ai_1 \register_file_i/_4413_  (.B1(\register_file_i/_1359_ ),
    .Y(\register_file_i/_1360_ ),
    .A1(net528),
    .A2(\register_file_i/_1356_ ));
 sg13g2_nand2_1 \register_file_i/_4414_  (.Y(\register_file_i/_1361_ ),
    .A(net1920),
    .B(\register_file_i/_1360_ ));
 sg13g2_mux4_1 \register_file_i/_4415_  (.S0(net2015),
    .A0(\register_file_i/rf_reg_524_ ),
    .A1(\register_file_i/rf_reg_556_ ),
    .A2(\register_file_i/rf_reg_588_ ),
    .A3(\register_file_i/rf_reg_620_ ),
    .S1(net541),
    .X(\register_file_i/_1362_ ));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(net1615));
 sg13g2_mux4_1 \register_file_i/_4417_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_652_ ),
    .A1(\register_file_i/rf_reg_684_ ),
    .A2(\register_file_i/rf_reg_716_ ),
    .A3(\register_file_i/rf_reg_748_ ),
    .S1(net543),
    .X(\register_file_i/_1364_ ));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net1615));
 sg13g2_mux2_1 \register_file_i/_4419_  (.A0(\register_file_i/rf_reg_396_ ),
    .A1(\register_file_i/rf_reg_428_ ),
    .S(net2010),
    .X(\register_file_i/_1366_ ));
 sg13g2_mux2_1 \register_file_i/_4420_  (.A0(\register_file_i/rf_reg_460_ ),
    .A1(\register_file_i/rf_reg_492_ ),
    .S(net2010),
    .X(\register_file_i/_1367_ ));
 sg13g2_a22oi_1 \register_file_i/_4421_  (.Y(\register_file_i/_1368_ ),
    .B1(\register_file_i/_1367_ ),
    .B2(net1820),
    .A2(\register_file_i/_1366_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4422_  (.A0(\register_file_i/rf_reg_332_ ),
    .A1(\register_file_i/rf_reg_364_ ),
    .S(net2011),
    .X(\register_file_i/_1369_ ));
 sg13g2_mux2_1 \register_file_i/_4423_  (.A0(\register_file_i/rf_reg_268_ ),
    .A1(\register_file_i/rf_reg_300_ ),
    .S(net2010),
    .X(\register_file_i/_1370_ ));
 sg13g2_a22oi_1 \register_file_i/_4424_  (.Y(\register_file_i/_1371_ ),
    .B1(\register_file_i/_1370_ ),
    .B2(net1798),
    .A2(\register_file_i/_1369_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4425_  (.A1(\register_file_i/_1368_ ),
    .A2(\register_file_i/_1371_ ),
    .Y(\register_file_i/_1372_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4426_  (.B2(net1693),
    .C1(\register_file_i/_1372_ ),
    .B1(\register_file_i/_1364_ ),
    .A1(net1792),
    .Y(\register_file_i/_1373_ ),
    .A2(\register_file_i/_1362_ ));
 sg13g2_nand3_1 \register_file_i/_4427_  (.B(\register_file_i/_1361_ ),
    .C(\register_file_i/_1373_ ),
    .A(\register_file_i/_1353_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_12_ ));
 sg13g2_mux2_1 \register_file_i/_4428_  (.A0(\register_file_i/rf_reg_925_ ),
    .A1(\register_file_i/rf_reg_957_ ),
    .S(net2072),
    .X(\register_file_i/_1374_ ));
 sg13g2_mux2_1 \register_file_i/_4429_  (.A0(\register_file_i/rf_reg_989_ ),
    .A1(\register_file_i/rf_reg_1021_ ),
    .S(net2072),
    .X(\register_file_i/_1375_ ));
 sg13g2_a22oi_1 \register_file_i/_4430_  (.Y(\register_file_i/_1376_ ),
    .B1(\register_file_i/_1375_ ),
    .B2(net1833),
    .A2(\register_file_i/_1374_ ),
    .A1(net1849));
 sg13g2_mux2_1 \register_file_i/_4431_  (.A0(\register_file_i/rf_reg_861_ ),
    .A1(\register_file_i/rf_reg_893_ ),
    .S(net2072),
    .X(\register_file_i/_1377_ ));
 sg13g2_mux2_1 \register_file_i/_4432_  (.A0(\register_file_i/rf_reg_797_ ),
    .A1(\register_file_i/rf_reg_829_ ),
    .S(net2072),
    .X(\register_file_i/_1378_ ));
 sg13g2_a22oi_1 \register_file_i/_4433_  (.Y(\register_file_i/_1379_ ),
    .B1(\register_file_i/_1378_ ),
    .B2(net1805),
    .A2(\register_file_i/_1377_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4434_  (.A2(\register_file_i/_1379_ ),
    .A1(\register_file_i/_1376_ ),
    .B1(net1926),
    .X(\register_file_i/_1380_ ));
 sg13g2_mux2_1 \register_file_i/_4435_  (.A0(\register_file_i/rf_reg_61_ ),
    .A1(\register_file_i/rf_reg_125_ ),
    .S(net534),
    .X(\register_file_i/_1381_ ));
 sg13g2_a22oi_1 \register_file_i/_4436_  (.Y(\register_file_i/_1382_ ),
    .B1(\register_file_i/_1381_ ),
    .B2(net2064),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_93_ ));
 sg13g2_mux2_1 \register_file_i/_4437_  (.A0(\register_file_i/rf_reg_221_ ),
    .A1(\register_file_i/rf_reg_253_ ),
    .S(net2062),
    .X(\register_file_i/_1383_ ));
 sg13g2_mux2_1 \register_file_i/_4438_  (.A0(\register_file_i/rf_reg_157_ ),
    .A1(\register_file_i/rf_reg_189_ ),
    .S(net2062),
    .X(\register_file_i/_1384_ ));
 sg13g2_a22oi_1 \register_file_i/_4439_  (.Y(\register_file_i/_1385_ ),
    .B1(\register_file_i/_1384_ ),
    .B2(net1846),
    .A2(\register_file_i/_1383_ ),
    .A1(net1830));
 sg13g2_o21ai_1 \register_file_i/_4440_  (.B1(\register_file_i/_1385_ ),
    .Y(\register_file_i/_1386_ ),
    .A1(net528),
    .A2(\register_file_i/_1382_ ));
 sg13g2_nand2_1 \register_file_i/_4441_  (.Y(\register_file_i/_1387_ ),
    .A(net1919),
    .B(\register_file_i/_1386_ ));
 sg13g2_mux4_1 \register_file_i/_4442_  (.S0(net2015),
    .A0(\register_file_i/rf_reg_541_ ),
    .A1(\register_file_i/rf_reg_573_ ),
    .A2(\register_file_i/rf_reg_605_ ),
    .A3(\register_file_i/rf_reg_637_ ),
    .S1(net541),
    .X(\register_file_i/_1388_ ));
 sg13g2_mux4_1 \register_file_i/_4443_  (.S0(net2015),
    .A0(\register_file_i/rf_reg_669_ ),
    .A1(\register_file_i/rf_reg_701_ ),
    .A2(\register_file_i/rf_reg_733_ ),
    .A3(\register_file_i/rf_reg_765_ ),
    .S1(net543),
    .X(\register_file_i/_1389_ ));
 sg13g2_buf_2 fanout351 (.A(net1615),
    .X(net351));
 sg13g2_mux2_1 \register_file_i/_4445_  (.A0(\register_file_i/rf_reg_413_ ),
    .A1(\register_file_i/rf_reg_445_ ),
    .S(net2011),
    .X(\register_file_i/_1391_ ));
 sg13g2_mux2_1 \register_file_i/_4446_  (.A0(\register_file_i/rf_reg_477_ ),
    .A1(\register_file_i/rf_reg_509_ ),
    .S(net2011),
    .X(\register_file_i/_1392_ ));
 sg13g2_a22oi_1 \register_file_i/_4447_  (.Y(\register_file_i/_1393_ ),
    .B1(\register_file_i/_1392_ ),
    .B2(net1820),
    .A2(\register_file_i/_1391_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4448_  (.A0(\register_file_i/rf_reg_349_ ),
    .A1(\register_file_i/rf_reg_381_ ),
    .S(net2011),
    .X(\register_file_i/_1394_ ));
 sg13g2_mux2_1 \register_file_i/_4449_  (.A0(\register_file_i/rf_reg_285_ ),
    .A1(\register_file_i/rf_reg_317_ ),
    .S(net2015),
    .X(\register_file_i/_1395_ ));
 sg13g2_a22oi_1 \register_file_i/_4450_  (.Y(\register_file_i/_1396_ ),
    .B1(\register_file_i/_1395_ ),
    .B2(net1798),
    .A2(\register_file_i/_1394_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4451_  (.A1(\register_file_i/_1393_ ),
    .A2(\register_file_i/_1396_ ),
    .Y(\register_file_i/_1397_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4452_  (.B2(net1693),
    .C1(\register_file_i/_1397_ ),
    .B1(\register_file_i/_1389_ ),
    .A1(net1792),
    .Y(\register_file_i/_1398_ ),
    .A2(\register_file_i/_1388_ ));
 sg13g2_nand3_1 \register_file_i/_4453_  (.B(\register_file_i/_1387_ ),
    .C(\register_file_i/_1398_ ),
    .A(\register_file_i/_1380_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net1616));
 sg13g2_mux2_1 \register_file_i/_4455_  (.A0(\register_file_i/rf_reg_907_ ),
    .A1(\register_file_i/rf_reg_939_ ),
    .S(net2057),
    .X(\register_file_i/_1400_ ));
 sg13g2_mux2_1 \register_file_i/_4456_  (.A0(\register_file_i/rf_reg_971_ ),
    .A1(\register_file_i/rf_reg_1003_ ),
    .S(net2056),
    .X(\register_file_i/_1401_ ));
 sg13g2_a22oi_1 \register_file_i/_4457_  (.Y(\register_file_i/_1402_ ),
    .B1(\register_file_i/_1401_ ),
    .B2(net1829),
    .A2(\register_file_i/_1400_ ),
    .A1(net1846));
 sg13g2_mux2_1 \register_file_i/_4458_  (.A0(\register_file_i/rf_reg_843_ ),
    .A1(\register_file_i/rf_reg_875_ ),
    .S(net2057),
    .X(\register_file_i/_1403_ ));
 sg13g2_mux2_1 \register_file_i/_4459_  (.A0(\register_file_i/rf_reg_779_ ),
    .A1(\register_file_i/rf_reg_811_ ),
    .S(net2056),
    .X(\register_file_i/_1404_ ));
 sg13g2_a22oi_1 \register_file_i/_4460_  (.Y(\register_file_i/_1405_ ),
    .B1(\register_file_i/_1404_ ),
    .B2(net1805),
    .A2(\register_file_i/_1403_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4461_  (.A2(\register_file_i/_1405_ ),
    .A1(\register_file_i/_1402_ ),
    .B1(net1925),
    .X(\register_file_i/_1406_ ));
 sg13g2_mux2_1 \register_file_i/_4462_  (.A0(\register_file_i/rf_reg_43_ ),
    .A1(\register_file_i/rf_reg_107_ ),
    .S(net533),
    .X(\register_file_i/_1407_ ));
 sg13g2_a22oi_1 \register_file_i/_4463_  (.Y(\register_file_i/_1408_ ),
    .B1(\register_file_i/_1407_ ),
    .B2(net2059),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_75_ ));
 sg13g2_mux2_1 \register_file_i/_4464_  (.A0(\register_file_i/rf_reg_203_ ),
    .A1(\register_file_i/rf_reg_235_ ),
    .S(net2062),
    .X(\register_file_i/_1409_ ));
 sg13g2_mux2_1 \register_file_i/_4465_  (.A0(\register_file_i/rf_reg_139_ ),
    .A1(\register_file_i/rf_reg_171_ ),
    .S(net2058),
    .X(\register_file_i/_1410_ ));
 sg13g2_a22oi_1 \register_file_i/_4466_  (.Y(\register_file_i/_1411_ ),
    .B1(\register_file_i/_1410_ ),
    .B2(net1845),
    .A2(\register_file_i/_1409_ ),
    .A1(net1828));
 sg13g2_o21ai_1 \register_file_i/_4467_  (.B1(\register_file_i/_1411_ ),
    .Y(\register_file_i/_1412_ ),
    .A1(net528),
    .A2(\register_file_i/_1408_ ));
 sg13g2_nand2_1 \register_file_i/_4468_  (.Y(\register_file_i/_1413_ ),
    .A(net1919),
    .B(\register_file_i/_1412_ ));
 sg13g2_mux4_1 \register_file_i/_4469_  (.S0(net2011),
    .A0(\register_file_i/rf_reg_523_ ),
    .A1(\register_file_i/rf_reg_555_ ),
    .A2(\register_file_i/rf_reg_587_ ),
    .A3(\register_file_i/rf_reg_619_ ),
    .S1(net541),
    .X(\register_file_i/_1414_ ));
 sg13g2_mux4_1 \register_file_i/_4470_  (.S0(net2010),
    .A0(\register_file_i/rf_reg_651_ ),
    .A1(\register_file_i/rf_reg_683_ ),
    .A2(\register_file_i/rf_reg_715_ ),
    .A3(\register_file_i/rf_reg_747_ ),
    .S1(net543),
    .X(\register_file_i/_1415_ ));
 sg13g2_mux2_1 \register_file_i/_4471_  (.A0(\register_file_i/rf_reg_395_ ),
    .A1(\register_file_i/rf_reg_427_ ),
    .S(net2010),
    .X(\register_file_i/_1416_ ));
 sg13g2_mux2_1 \register_file_i/_4472_  (.A0(\register_file_i/rf_reg_459_ ),
    .A1(\register_file_i/rf_reg_491_ ),
    .S(net2010),
    .X(\register_file_i/_1417_ ));
 sg13g2_a22oi_1 \register_file_i/_4473_  (.Y(\register_file_i/_1418_ ),
    .B1(\register_file_i/_1417_ ),
    .B2(net1820),
    .A2(\register_file_i/_1416_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4474_  (.A0(\register_file_i/rf_reg_331_ ),
    .A1(\register_file_i/rf_reg_363_ ),
    .S(net2010),
    .X(\register_file_i/_1419_ ));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net1616));
 sg13g2_mux2_1 \register_file_i/_4476_  (.A0(\register_file_i/rf_reg_267_ ),
    .A1(\register_file_i/rf_reg_299_ ),
    .S(net2010),
    .X(\register_file_i/_1421_ ));
 sg13g2_a22oi_1 \register_file_i/_4477_  (.Y(\register_file_i/_1422_ ),
    .B1(\register_file_i/_1421_ ),
    .B2(net1798),
    .A2(\register_file_i/_1419_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4478_  (.A1(\register_file_i/_1418_ ),
    .A2(\register_file_i/_1422_ ),
    .Y(\register_file_i/_1423_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4479_  (.B2(net1693),
    .C1(\register_file_i/_1423_ ),
    .B1(\register_file_i/_1415_ ),
    .A1(net1792),
    .Y(\register_file_i/_1424_ ),
    .A2(\register_file_i/_1414_ ));
 sg13g2_nand3_1 \register_file_i/_4480_  (.B(\register_file_i/_1413_ ),
    .C(\register_file_i/_1424_ ),
    .A(\register_file_i/_1406_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_mux2_1 \register_file_i/_4481_  (.A0(\register_file_i/rf_reg_906_ ),
    .A1(\register_file_i/rf_reg_938_ ),
    .S(net2056),
    .X(\register_file_i/_1425_ ));
 sg13g2_mux2_1 \register_file_i/_4482_  (.A0(\register_file_i/rf_reg_970_ ),
    .A1(\register_file_i/rf_reg_1002_ ),
    .S(net2056),
    .X(\register_file_i/_1426_ ));
 sg13g2_a22oi_1 \register_file_i/_4483_  (.Y(\register_file_i/_1427_ ),
    .B1(\register_file_i/_1426_ ),
    .B2(net1828),
    .A2(\register_file_i/_1425_ ),
    .A1(net1846));
 sg13g2_mux2_1 \register_file_i/_4484_  (.A0(\register_file_i/rf_reg_842_ ),
    .A1(\register_file_i/rf_reg_874_ ),
    .S(net2056),
    .X(\register_file_i/_1428_ ));
 sg13g2_mux2_1 \register_file_i/_4485_  (.A0(\register_file_i/rf_reg_778_ ),
    .A1(\register_file_i/rf_reg_810_ ),
    .S(net2056),
    .X(\register_file_i/_1429_ ));
 sg13g2_a22oi_1 \register_file_i/_4486_  (.Y(\register_file_i/_1430_ ),
    .B1(\register_file_i/_1429_ ),
    .B2(net1804),
    .A2(\register_file_i/_1428_ ),
    .A1(net1815));
 sg13g2_a21o_1 \register_file_i/_4487_  (.A2(\register_file_i/_1430_ ),
    .A1(\register_file_i/_1427_ ),
    .B1(net1925),
    .X(\register_file_i/_1431_ ));
 sg13g2_mux2_1 \register_file_i/_4488_  (.A0(\register_file_i/rf_reg_42_ ),
    .A1(\register_file_i/rf_reg_106_ ),
    .S(net533),
    .X(\register_file_i/_1432_ ));
 sg13g2_a22oi_1 \register_file_i/_4489_  (.Y(\register_file_i/_1433_ ),
    .B1(\register_file_i/_1432_ ),
    .B2(net2059),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_74_ ));
 sg13g2_buf_2 fanout348 (.A(_01801_),
    .X(net348));
 sg13g2_mux2_1 \register_file_i/_4491_  (.A0(\register_file_i/rf_reg_202_ ),
    .A1(\register_file_i/rf_reg_234_ ),
    .S(net2058),
    .X(\register_file_i/_1435_ ));
 sg13g2_mux2_1 \register_file_i/_4492_  (.A0(\register_file_i/rf_reg_138_ ),
    .A1(\register_file_i/rf_reg_170_ ),
    .S(net2058),
    .X(\register_file_i/_1436_ ));
 sg13g2_a22oi_1 \register_file_i/_4493_  (.Y(\register_file_i/_1437_ ),
    .B1(\register_file_i/_1436_ ),
    .B2(net1845),
    .A2(\register_file_i/_1435_ ),
    .A1(net1829));
 sg13g2_o21ai_1 \register_file_i/_4494_  (.B1(\register_file_i/_1437_ ),
    .Y(\register_file_i/_1438_ ),
    .A1(net527),
    .A2(\register_file_i/_1433_ ));
 sg13g2_nand2_1 \register_file_i/_4495_  (.Y(\register_file_i/_1439_ ),
    .A(net1920),
    .B(\register_file_i/_1438_ ));
 sg13g2_buf_2 fanout347 (.A(_01801_),
    .X(net347));
 sg13g2_mux4_1 \register_file_i/_4497_  (.S0(net2013),
    .A0(\register_file_i/rf_reg_522_ ),
    .A1(\register_file_i/rf_reg_554_ ),
    .A2(\register_file_i/rf_reg_586_ ),
    .A3(\register_file_i/rf_reg_618_ ),
    .S1(net544),
    .X(\register_file_i/_1441_ ));
 sg13g2_mux4_1 \register_file_i/_4498_  (.S0(net2013),
    .A0(\register_file_i/rf_reg_650_ ),
    .A1(\register_file_i/rf_reg_682_ ),
    .A2(\register_file_i/rf_reg_714_ ),
    .A3(\register_file_i/rf_reg_746_ ),
    .S1(net543),
    .X(\register_file_i/_1442_ ));
 sg13g2_mux2_1 \register_file_i/_4499_  (.A0(\register_file_i/rf_reg_394_ ),
    .A1(\register_file_i/rf_reg_426_ ),
    .S(net2012),
    .X(\register_file_i/_1443_ ));
 sg13g2_mux2_1 \register_file_i/_4500_  (.A0(\register_file_i/rf_reg_458_ ),
    .A1(\register_file_i/rf_reg_490_ ),
    .S(net2012),
    .X(\register_file_i/_1444_ ));
 sg13g2_a22oi_1 \register_file_i/_4501_  (.Y(\register_file_i/_1445_ ),
    .B1(\register_file_i/_1444_ ),
    .B2(net1820),
    .A2(\register_file_i/_1443_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4502_  (.A0(\register_file_i/rf_reg_330_ ),
    .A1(\register_file_i/rf_reg_362_ ),
    .S(net2012),
    .X(\register_file_i/_1446_ ));
 sg13g2_mux2_1 \register_file_i/_4503_  (.A0(\register_file_i/rf_reg_266_ ),
    .A1(\register_file_i/rf_reg_298_ ),
    .S(net2012),
    .X(\register_file_i/_1447_ ));
 sg13g2_a22oi_1 \register_file_i/_4504_  (.Y(\register_file_i/_1448_ ),
    .B1(\register_file_i/_1447_ ),
    .B2(net1798),
    .A2(\register_file_i/_1446_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4505_  (.A1(\register_file_i/_1445_ ),
    .A2(\register_file_i/_1448_ ),
    .Y(\register_file_i/_1449_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4506_  (.B2(net1693),
    .C1(\register_file_i/_1449_ ),
    .B1(\register_file_i/_1442_ ),
    .A1(net1792),
    .Y(\register_file_i/_1450_ ),
    .A2(\register_file_i/_1441_ ));
 sg13g2_nand3_1 \register_file_i/_4507_  (.B(\register_file_i/_1439_ ),
    .C(\register_file_i/_1450_ ),
    .A(\register_file_i/_1431_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_mux2_1 \register_file_i/_4508_  (.A0(\register_file_i/rf_reg_905_ ),
    .A1(\register_file_i/rf_reg_937_ ),
    .S(net2057),
    .X(\register_file_i/_1451_ ));
 sg13g2_mux2_1 \register_file_i/_4509_  (.A0(\register_file_i/rf_reg_969_ ),
    .A1(\register_file_i/rf_reg_1001_ ),
    .S(net2056),
    .X(\register_file_i/_1452_ ));
 sg13g2_a22oi_1 \register_file_i/_4510_  (.Y(\register_file_i/_1453_ ),
    .B1(\register_file_i/_1452_ ),
    .B2(net1828),
    .A2(\register_file_i/_1451_ ),
    .A1(net1846));
 sg13g2_mux2_1 \register_file_i/_4511_  (.A0(\register_file_i/rf_reg_841_ ),
    .A1(\register_file_i/rf_reg_873_ ),
    .S(net2057),
    .X(\register_file_i/_1454_ ));
 sg13g2_buf_1 fanout346 (.A(csr_restore_mret_id),
    .X(net346));
 sg13g2_mux2_1 \register_file_i/_4513_  (.A0(\register_file_i/rf_reg_777_ ),
    .A1(\register_file_i/rf_reg_809_ ),
    .S(net2056),
    .X(\register_file_i/_1456_ ));
 sg13g2_a22oi_1 \register_file_i/_4514_  (.Y(\register_file_i/_1457_ ),
    .B1(\register_file_i/_1456_ ),
    .B2(net1805),
    .A2(\register_file_i/_1454_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4515_  (.A2(\register_file_i/_1457_ ),
    .A1(\register_file_i/_1453_ ),
    .B1(net1925),
    .X(\register_file_i/_1458_ ));
 sg13g2_mux2_1 \register_file_i/_4516_  (.A0(\register_file_i/rf_reg_41_ ),
    .A1(\register_file_i/rf_reg_105_ ),
    .S(net533),
    .X(\register_file_i/_1459_ ));
 sg13g2_a22oi_1 \register_file_i/_4517_  (.Y(\register_file_i/_1460_ ),
    .B1(\register_file_i/_1459_ ),
    .B2(net2058),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_73_ ));
 sg13g2_mux2_1 \register_file_i/_4518_  (.A0(\register_file_i/rf_reg_201_ ),
    .A1(\register_file_i/rf_reg_233_ ),
    .S(net2058),
    .X(\register_file_i/_1461_ ));
 sg13g2_mux2_1 \register_file_i/_4519_  (.A0(\register_file_i/rf_reg_137_ ),
    .A1(\register_file_i/rf_reg_169_ ),
    .S(net2058),
    .X(\register_file_i/_1462_ ));
 sg13g2_a22oi_1 \register_file_i/_4520_  (.Y(\register_file_i/_1463_ ),
    .B1(\register_file_i/_1462_ ),
    .B2(net1845),
    .A2(\register_file_i/_1461_ ),
    .A1(net1829));
 sg13g2_o21ai_1 \register_file_i/_4521_  (.B1(\register_file_i/_1463_ ),
    .Y(\register_file_i/_1464_ ),
    .A1(net527),
    .A2(\register_file_i/_1460_ ));
 sg13g2_nand2_1 \register_file_i/_4522_  (.Y(\register_file_i/_1465_ ),
    .A(net1920),
    .B(\register_file_i/_1464_ ));
 sg13g2_mux4_1 \register_file_i/_4523_  (.S0(net2013),
    .A0(\register_file_i/rf_reg_521_ ),
    .A1(\register_file_i/rf_reg_553_ ),
    .A2(\register_file_i/rf_reg_585_ ),
    .A3(\register_file_i/rf_reg_617_ ),
    .S1(net544),
    .X(\register_file_i/_1466_ ));
 sg13g2_buf_2 fanout345 (.A(net346),
    .X(net345));
 sg13g2_mux4_1 \register_file_i/_4525_  (.S0(net2013),
    .A0(\register_file_i/rf_reg_649_ ),
    .A1(\register_file_i/rf_reg_681_ ),
    .A2(\register_file_i/rf_reg_713_ ),
    .A3(\register_file_i/rf_reg_745_ ),
    .S1(net542),
    .X(\register_file_i/_1468_ ));
 sg13g2_mux2_1 \register_file_i/_4526_  (.A0(\register_file_i/rf_reg_393_ ),
    .A1(\register_file_i/rf_reg_425_ ),
    .S(net2012),
    .X(\register_file_i/_1469_ ));
 sg13g2_buf_2 fanout344 (.A(net346),
    .X(net344));
 sg13g2_mux2_1 \register_file_i/_4528_  (.A0(\register_file_i/rf_reg_457_ ),
    .A1(\register_file_i/rf_reg_489_ ),
    .S(net2013),
    .X(\register_file_i/_1471_ ));
 sg13g2_a22oi_1 \register_file_i/_4529_  (.Y(\register_file_i/_1472_ ),
    .B1(\register_file_i/_1471_ ),
    .B2(net1820),
    .A2(\register_file_i/_1469_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4530_  (.A0(\register_file_i/rf_reg_329_ ),
    .A1(\register_file_i/rf_reg_361_ ),
    .S(net2012),
    .X(\register_file_i/_1473_ ));
 sg13g2_mux2_1 \register_file_i/_4531_  (.A0(\register_file_i/rf_reg_265_ ),
    .A1(\register_file_i/rf_reg_297_ ),
    .S(net2012),
    .X(\register_file_i/_1474_ ));
 sg13g2_a22oi_1 \register_file_i/_4532_  (.Y(\register_file_i/_1475_ ),
    .B1(\register_file_i/_1474_ ),
    .B2(net1798),
    .A2(\register_file_i/_1473_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4533_  (.A1(\register_file_i/_1472_ ),
    .A2(\register_file_i/_1475_ ),
    .Y(\register_file_i/_1476_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4534_  (.B2(net1693),
    .C1(\register_file_i/_1476_ ),
    .B1(\register_file_i/_1468_ ),
    .A1(net1792),
    .Y(\register_file_i/_1477_ ),
    .A2(\register_file_i/_1466_ ));
 sg13g2_nand3_1 \register_file_i/_4535_  (.B(\register_file_i/_1465_ ),
    .C(\register_file_i/_1477_ ),
    .A(\register_file_i/_1458_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_mux2_1 \register_file_i/_4536_  (.A0(\register_file_i/rf_reg_904_ ),
    .A1(\register_file_i/rf_reg_936_ ),
    .S(net2068),
    .X(\register_file_i/_1478_ ));
 sg13g2_mux2_1 \register_file_i/_4537_  (.A0(\register_file_i/rf_reg_968_ ),
    .A1(\register_file_i/rf_reg_1000_ ),
    .S(net2068),
    .X(\register_file_i/_1479_ ));
 sg13g2_a22oi_1 \register_file_i/_4538_  (.Y(\register_file_i/_1480_ ),
    .B1(\register_file_i/_1479_ ),
    .B2(net1831),
    .A2(\register_file_i/_1478_ ),
    .A1(net1848));
 sg13g2_mux2_1 \register_file_i/_4539_  (.A0(\register_file_i/rf_reg_840_ ),
    .A1(\register_file_i/rf_reg_872_ ),
    .S(net2066),
    .X(\register_file_i/_1481_ ));
 sg13g2_mux2_1 \register_file_i/_4540_  (.A0(\register_file_i/rf_reg_776_ ),
    .A1(\register_file_i/rf_reg_808_ ),
    .S(net2066),
    .X(\register_file_i/_1482_ ));
 sg13g2_a22oi_1 \register_file_i/_4541_  (.Y(\register_file_i/_1483_ ),
    .B1(\register_file_i/_1482_ ),
    .B2(net1805),
    .A2(\register_file_i/_1481_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4542_  (.A2(\register_file_i/_1483_ ),
    .A1(\register_file_i/_1480_ ),
    .B1(net1925),
    .X(\register_file_i/_1484_ ));
 sg13g2_mux2_1 \register_file_i/_4543_  (.A0(\register_file_i/rf_reg_40_ ),
    .A1(\register_file_i/rf_reg_104_ ),
    .S(net533),
    .X(\register_file_i/_1485_ ));
 sg13g2_a22oi_1 \register_file_i/_4544_  (.Y(\register_file_i/_1486_ ),
    .B1(\register_file_i/_1485_ ),
    .B2(net2067),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_72_ ));
 sg13g2_mux2_1 \register_file_i/_4545_  (.A0(\register_file_i/rf_reg_200_ ),
    .A1(\register_file_i/rf_reg_232_ ),
    .S(net2067),
    .X(\register_file_i/_1487_ ));
 sg13g2_mux2_1 \register_file_i/_4546_  (.A0(\register_file_i/rf_reg_136_ ),
    .A1(\register_file_i/rf_reg_168_ ),
    .S(net2067),
    .X(\register_file_i/_1488_ ));
 sg13g2_a22oi_1 \register_file_i/_4547_  (.Y(\register_file_i/_1489_ ),
    .B1(\register_file_i/_1488_ ),
    .B2(net1848),
    .A2(\register_file_i/_1487_ ),
    .A1(net1832));
 sg13g2_o21ai_1 \register_file_i/_4548_  (.B1(\register_file_i/_1489_ ),
    .Y(\register_file_i/_1490_ ),
    .A1(net527),
    .A2(\register_file_i/_1486_ ));
 sg13g2_nand2_1 \register_file_i/_4549_  (.Y(\register_file_i/_1491_ ),
    .A(net1919),
    .B(\register_file_i/_1490_ ));
 sg13g2_buf_2 fanout343 (.A(_03956_),
    .X(net343));
 sg13g2_mux4_1 \register_file_i/_4551_  (.S0(net2021),
    .A0(\register_file_i/rf_reg_520_ ),
    .A1(\register_file_i/rf_reg_552_ ),
    .A2(\register_file_i/rf_reg_584_ ),
    .A3(\register_file_i/rf_reg_616_ ),
    .S1(net544),
    .X(\register_file_i/_1493_ ));
 sg13g2_mux4_1 \register_file_i/_4552_  (.S0(net2021),
    .A0(\register_file_i/rf_reg_648_ ),
    .A1(\register_file_i/rf_reg_680_ ),
    .A2(\register_file_i/rf_reg_712_ ),
    .A3(\register_file_i/rf_reg_744_ ),
    .S1(net542),
    .X(\register_file_i/_1494_ ));
 sg13g2_mux2_1 \register_file_i/_4553_  (.A0(\register_file_i/rf_reg_392_ ),
    .A1(\register_file_i/rf_reg_424_ ),
    .S(net2020),
    .X(\register_file_i/_1495_ ));
 sg13g2_mux2_1 \register_file_i/_4554_  (.A0(\register_file_i/rf_reg_456_ ),
    .A1(\register_file_i/rf_reg_488_ ),
    .S(net2020),
    .X(\register_file_i/_1496_ ));
 sg13g2_a22oi_1 \register_file_i/_4555_  (.Y(\register_file_i/_1497_ ),
    .B1(\register_file_i/_1496_ ),
    .B2(net1821),
    .A2(\register_file_i/_1495_ ),
    .A1(net1838));
 sg13g2_mux2_1 \register_file_i/_4556_  (.A0(\register_file_i/rf_reg_328_ ),
    .A1(\register_file_i/rf_reg_360_ ),
    .S(net2020),
    .X(\register_file_i/_1498_ ));
 sg13g2_mux2_1 \register_file_i/_4557_  (.A0(\register_file_i/rf_reg_264_ ),
    .A1(\register_file_i/rf_reg_296_ ),
    .S(net2020),
    .X(\register_file_i/_1499_ ));
 sg13g2_a22oi_1 \register_file_i/_4558_  (.Y(\register_file_i/_1500_ ),
    .B1(\register_file_i/_1499_ ),
    .B2(net1799),
    .A2(\register_file_i/_1498_ ),
    .A1(net1810));
 sg13g2_buf_4 fanout342 (.X(net342),
    .A(net343));
 sg13g2_a21oi_1 \register_file_i/_4560_  (.A1(\register_file_i/_1497_ ),
    .A2(\register_file_i/_1500_ ),
    .Y(\register_file_i/_1502_ ),
    .B1(net1788));
 sg13g2_a221oi_1 \register_file_i/_4561_  (.B2(net1693),
    .C1(\register_file_i/_1502_ ),
    .B1(\register_file_i/_1494_ ),
    .A1(net1792),
    .Y(\register_file_i/_1503_ ),
    .A2(\register_file_i/_1493_ ));
 sg13g2_nand3_1 \register_file_i/_4562_  (.B(\register_file_i/_1491_ ),
    .C(\register_file_i/_1503_ ),
    .A(\register_file_i/_1484_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_mux2_1 \register_file_i/_4563_  (.A0(\register_file_i/rf_reg_903_ ),
    .A1(\register_file_i/rf_reg_935_ ),
    .S(net2068),
    .X(\register_file_i/_1504_ ));
 sg13g2_mux2_1 \register_file_i/_4564_  (.A0(\register_file_i/rf_reg_967_ ),
    .A1(\register_file_i/rf_reg_999_ ),
    .S(net2068),
    .X(\register_file_i/_1505_ ));
 sg13g2_a22oi_1 \register_file_i/_4565_  (.Y(\register_file_i/_1506_ ),
    .B1(\register_file_i/_1505_ ),
    .B2(net1831),
    .A2(\register_file_i/_1504_ ),
    .A1(net1848));
 sg13g2_mux2_1 \register_file_i/_4566_  (.A0(\register_file_i/rf_reg_839_ ),
    .A1(\register_file_i/rf_reg_871_ ),
    .S(net2066),
    .X(\register_file_i/_1507_ ));
 sg13g2_mux2_1 \register_file_i/_4567_  (.A0(\register_file_i/rf_reg_775_ ),
    .A1(\register_file_i/rf_reg_807_ ),
    .S(net2067),
    .X(\register_file_i/_1508_ ));
 sg13g2_a22oi_1 \register_file_i/_4568_  (.Y(\register_file_i/_1509_ ),
    .B1(\register_file_i/_1508_ ),
    .B2(net1805),
    .A2(\register_file_i/_1507_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4569_  (.A2(\register_file_i/_1509_ ),
    .A1(\register_file_i/_1506_ ),
    .B1(net1925),
    .X(\register_file_i/_1510_ ));
 sg13g2_buf_4 fanout341 (.X(net341),
    .A(net343));
 sg13g2_mux2_1 \register_file_i/_4571_  (.A0(\register_file_i/rf_reg_39_ ),
    .A1(\register_file_i/rf_reg_103_ ),
    .S(net535),
    .X(\register_file_i/_1512_ ));
 sg13g2_a22oi_1 \register_file_i/_4572_  (.Y(\register_file_i/_1513_ ),
    .B1(\register_file_i/_1512_ ),
    .B2(net2067),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_71_ ));
 sg13g2_buf_2 fanout340 (.A(net343),
    .X(net340));
 sg13g2_mux2_1 \register_file_i/_4574_  (.A0(\register_file_i/rf_reg_199_ ),
    .A1(\register_file_i/rf_reg_231_ ),
    .S(net2069),
    .X(\register_file_i/_1515_ ));
 sg13g2_mux2_1 \register_file_i/_4575_  (.A0(\register_file_i/rf_reg_135_ ),
    .A1(\register_file_i/rf_reg_167_ ),
    .S(net2070),
    .X(\register_file_i/_1516_ ));
 sg13g2_a22oi_1 \register_file_i/_4576_  (.Y(\register_file_i/_1517_ ),
    .B1(\register_file_i/_1516_ ),
    .B2(net1848),
    .A2(\register_file_i/_1515_ ),
    .A1(net1831));
 sg13g2_o21ai_1 \register_file_i/_4577_  (.B1(\register_file_i/_1517_ ),
    .Y(\register_file_i/_1518_ ),
    .A1(net527),
    .A2(\register_file_i/_1513_ ));
 sg13g2_nand2_1 \register_file_i/_4578_  (.Y(\register_file_i/_1519_ ),
    .A(net1919),
    .B(\register_file_i/_1518_ ));
 sg13g2_mux4_1 \register_file_i/_4579_  (.S0(net2021),
    .A0(\register_file_i/rf_reg_519_ ),
    .A1(\register_file_i/rf_reg_551_ ),
    .A2(\register_file_i/rf_reg_583_ ),
    .A3(\register_file_i/rf_reg_615_ ),
    .S1(net544),
    .X(\register_file_i/_1520_ ));
 sg13g2_mux4_1 \register_file_i/_4580_  (.S0(net2021),
    .A0(\register_file_i/rf_reg_647_ ),
    .A1(\register_file_i/rf_reg_679_ ),
    .A2(\register_file_i/rf_reg_711_ ),
    .A3(\register_file_i/rf_reg_743_ ),
    .S1(net542),
    .X(\register_file_i/_1521_ ));
 sg13g2_mux2_1 \register_file_i/_4581_  (.A0(\register_file_i/rf_reg_391_ ),
    .A1(\register_file_i/rf_reg_423_ ),
    .S(net2021),
    .X(\register_file_i/_1522_ ));
 sg13g2_mux2_1 \register_file_i/_4582_  (.A0(\register_file_i/rf_reg_455_ ),
    .A1(\register_file_i/rf_reg_487_ ),
    .S(net2021),
    .X(\register_file_i/_1523_ ));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(net343));
 sg13g2_a22oi_1 \register_file_i/_4584_  (.Y(\register_file_i/_1525_ ),
    .B1(\register_file_i/_1523_ ),
    .B2(net1821),
    .A2(\register_file_i/_1522_ ),
    .A1(net1838));
 sg13g2_mux2_1 \register_file_i/_4585_  (.A0(\register_file_i/rf_reg_327_ ),
    .A1(\register_file_i/rf_reg_359_ ),
    .S(net2020),
    .X(\register_file_i/_1526_ ));
 sg13g2_mux2_1 \register_file_i/_4586_  (.A0(\register_file_i/rf_reg_263_ ),
    .A1(\register_file_i/rf_reg_295_ ),
    .S(net2021),
    .X(\register_file_i/_1527_ ));
 sg13g2_a22oi_1 \register_file_i/_4587_  (.Y(\register_file_i/_1528_ ),
    .B1(\register_file_i/_1527_ ),
    .B2(net1799),
    .A2(\register_file_i/_1526_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4588_  (.A1(\register_file_i/_1525_ ),
    .A2(\register_file_i/_1528_ ),
    .Y(\register_file_i/_1529_ ),
    .B1(net1788));
 sg13g2_a221oi_1 \register_file_i/_4589_  (.B2(net1694),
    .C1(\register_file_i/_1529_ ),
    .B1(\register_file_i/_1521_ ),
    .A1(net1794),
    .Y(\register_file_i/_1530_ ),
    .A2(\register_file_i/_1520_ ));
 sg13g2_nand3_1 \register_file_i/_4590_  (.B(\register_file_i/_1519_ ),
    .C(\register_file_i/_1530_ ),
    .A(\register_file_i/_1510_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_mux2_1 \register_file_i/_4591_  (.A0(\register_file_i/rf_reg_902_ ),
    .A1(\register_file_i/rf_reg_934_ ),
    .S(net2070),
    .X(\register_file_i/_1531_ ));
 sg13g2_buf_2 fanout338 (.A(net343),
    .X(net338));
 sg13g2_mux2_1 \register_file_i/_4593_  (.A0(\register_file_i/rf_reg_966_ ),
    .A1(\register_file_i/rf_reg_998_ ),
    .S(net2068),
    .X(\register_file_i/_1533_ ));
 sg13g2_a22oi_1 \register_file_i/_4594_  (.Y(\register_file_i/_1534_ ),
    .B1(\register_file_i/_1533_ ),
    .B2(net1831),
    .A2(\register_file_i/_1531_ ),
    .A1(net1848));
 sg13g2_mux2_1 \register_file_i/_4595_  (.A0(\register_file_i/rf_reg_838_ ),
    .A1(\register_file_i/rf_reg_870_ ),
    .S(net2066),
    .X(\register_file_i/_1535_ ));
 sg13g2_mux2_1 \register_file_i/_4596_  (.A0(\register_file_i/rf_reg_774_ ),
    .A1(\register_file_i/rf_reg_806_ ),
    .S(net2066),
    .X(\register_file_i/_1536_ ));
 sg13g2_a22oi_1 \register_file_i/_4597_  (.Y(\register_file_i/_1537_ ),
    .B1(\register_file_i/_1536_ ),
    .B2(net1805),
    .A2(\register_file_i/_1535_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4598_  (.A2(\register_file_i/_1537_ ),
    .A1(\register_file_i/_1534_ ),
    .B1(net1925),
    .X(\register_file_i/_1538_ ));
 sg13g2_mux2_1 \register_file_i/_4599_  (.A0(\register_file_i/rf_reg_38_ ),
    .A1(\register_file_i/rf_reg_102_ ),
    .S(net535),
    .X(\register_file_i/_1539_ ));
 sg13g2_a22oi_1 \register_file_i/_4600_  (.Y(\register_file_i/_1540_ ),
    .B1(\register_file_i/_1539_ ),
    .B2(net2069),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_70_ ));
 sg13g2_mux2_1 \register_file_i/_4601_  (.A0(\register_file_i/rf_reg_198_ ),
    .A1(\register_file_i/rf_reg_230_ ),
    .S(net2069),
    .X(\register_file_i/_1541_ ));
 sg13g2_mux2_1 \register_file_i/_4602_  (.A0(\register_file_i/rf_reg_134_ ),
    .A1(\register_file_i/rf_reg_166_ ),
    .S(net2068),
    .X(\register_file_i/_1542_ ));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(net343));
 sg13g2_a22oi_1 \register_file_i/_4604_  (.Y(\register_file_i/_1544_ ),
    .B1(\register_file_i/_1542_ ),
    .B2(net1849),
    .A2(\register_file_i/_1541_ ),
    .A1(net1832));
 sg13g2_o21ai_1 \register_file_i/_4605_  (.B1(\register_file_i/_1544_ ),
    .Y(\register_file_i/_1545_ ),
    .A1(net527),
    .A2(\register_file_i/_1540_ ));
 sg13g2_nand2_1 \register_file_i/_4606_  (.Y(\register_file_i/_1546_ ),
    .A(net1919),
    .B(\register_file_i/_1545_ ));
 sg13g2_mux4_1 \register_file_i/_4607_  (.S0(net2024),
    .A0(\register_file_i/rf_reg_518_ ),
    .A1(\register_file_i/rf_reg_550_ ),
    .A2(\register_file_i/rf_reg_582_ ),
    .A3(\register_file_i/rf_reg_614_ ),
    .S1(net544),
    .X(\register_file_i/_1547_ ));
 sg13g2_mux4_1 \register_file_i/_4608_  (.S0(net2024),
    .A0(\register_file_i/rf_reg_646_ ),
    .A1(\register_file_i/rf_reg_678_ ),
    .A2(\register_file_i/rf_reg_710_ ),
    .A3(\register_file_i/rf_reg_742_ ),
    .S1(net542),
    .X(\register_file_i/_1548_ ));
 sg13g2_mux2_1 \register_file_i/_4609_  (.A0(\register_file_i/rf_reg_390_ ),
    .A1(\register_file_i/rf_reg_422_ ),
    .S(net2022),
    .X(\register_file_i/_1549_ ));
 sg13g2_mux2_1 \register_file_i/_4610_  (.A0(\register_file_i/rf_reg_454_ ),
    .A1(\register_file_i/rf_reg_486_ ),
    .S(net2022),
    .X(\register_file_i/_1550_ ));
 sg13g2_a22oi_1 \register_file_i/_4611_  (.Y(\register_file_i/_1551_ ),
    .B1(\register_file_i/_1550_ ),
    .B2(net1821),
    .A2(\register_file_i/_1549_ ),
    .A1(net1838));
 sg13g2_mux2_1 \register_file_i/_4612_  (.A0(\register_file_i/rf_reg_326_ ),
    .A1(\register_file_i/rf_reg_358_ ),
    .S(net2022),
    .X(\register_file_i/_1552_ ));
 sg13g2_mux2_1 \register_file_i/_4613_  (.A0(\register_file_i/rf_reg_262_ ),
    .A1(\register_file_i/rf_reg_294_ ),
    .S(net2022),
    .X(\register_file_i/_1553_ ));
 sg13g2_buf_2 fanout336 (.A(_07486_),
    .X(net336));
 sg13g2_a22oi_1 \register_file_i/_4615_  (.Y(\register_file_i/_1555_ ),
    .B1(\register_file_i/_1553_ ),
    .B2(net1799),
    .A2(\register_file_i/_1552_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4616_  (.A1(\register_file_i/_1551_ ),
    .A2(\register_file_i/_1555_ ),
    .Y(\register_file_i/_1556_ ),
    .B1(net1788));
 sg13g2_a221oi_1 \register_file_i/_4617_  (.B2(net1694),
    .C1(\register_file_i/_1556_ ),
    .B1(\register_file_i/_1548_ ),
    .A1(net1794),
    .Y(\register_file_i/_1557_ ),
    .A2(\register_file_i/_1547_ ));
 sg13g2_nand3_1 \register_file_i/_4618_  (.B(\register_file_i/_1546_ ),
    .C(\register_file_i/_1557_ ),
    .A(\register_file_i/_1538_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_mux2_1 \register_file_i/_4619_  (.A0(\register_file_i/rf_reg_901_ ),
    .A1(\register_file_i/rf_reg_933_ ),
    .S(net2068),
    .X(\register_file_i/_1558_ ));
 sg13g2_mux2_1 \register_file_i/_4620_  (.A0(\register_file_i/rf_reg_965_ ),
    .A1(\register_file_i/rf_reg_997_ ),
    .S(net2068),
    .X(\register_file_i/_1559_ ));
 sg13g2_a22oi_1 \register_file_i/_4621_  (.Y(\register_file_i/_1560_ ),
    .B1(\register_file_i/_1559_ ),
    .B2(net1831),
    .A2(\register_file_i/_1558_ ),
    .A1(net1848));
 sg13g2_mux2_1 \register_file_i/_4622_  (.A0(\register_file_i/rf_reg_837_ ),
    .A1(\register_file_i/rf_reg_869_ ),
    .S(net2067),
    .X(\register_file_i/_1561_ ));
 sg13g2_mux2_1 \register_file_i/_4623_  (.A0(\register_file_i/rf_reg_773_ ),
    .A1(\register_file_i/rf_reg_805_ ),
    .S(net2071),
    .X(\register_file_i/_1562_ ));
 sg13g2_a22oi_1 \register_file_i/_4624_  (.Y(\register_file_i/_1563_ ),
    .B1(\register_file_i/_1562_ ),
    .B2(net1805),
    .A2(\register_file_i/_1561_ ),
    .A1(net1816));
 sg13g2_a21o_1 \register_file_i/_4625_  (.A2(\register_file_i/_1563_ ),
    .A1(\register_file_i/_1560_ ),
    .B1(net1925),
    .X(\register_file_i/_1564_ ));
 sg13g2_mux2_1 \register_file_i/_4626_  (.A0(\register_file_i/rf_reg_37_ ),
    .A1(\register_file_i/rf_reg_101_ ),
    .S(net535),
    .X(\register_file_i/_1565_ ));
 sg13g2_a22oi_1 \register_file_i/_4627_  (.Y(\register_file_i/_1566_ ),
    .B1(\register_file_i/_1565_ ),
    .B2(net2069),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_69_ ));
 sg13g2_mux2_1 \register_file_i/_4628_  (.A0(\register_file_i/rf_reg_197_ ),
    .A1(\register_file_i/rf_reg_229_ ),
    .S(net2069),
    .X(\register_file_i/_1567_ ));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_07486_));
 sg13g2_mux2_1 \register_file_i/_4630_  (.A0(\register_file_i/rf_reg_133_ ),
    .A1(\register_file_i/rf_reg_165_ ),
    .S(net2070),
    .X(\register_file_i/_1569_ ));
 sg13g2_a22oi_1 \register_file_i/_4631_  (.Y(\register_file_i/_1570_ ),
    .B1(\register_file_i/_1569_ ),
    .B2(net1849),
    .A2(\register_file_i/_1567_ ),
    .A1(net1831));
 sg13g2_o21ai_1 \register_file_i/_4632_  (.B1(\register_file_i/_1570_ ),
    .Y(\register_file_i/_1571_ ),
    .A1(net527),
    .A2(\register_file_i/_1566_ ));
 sg13g2_nand2_1 \register_file_i/_4633_  (.Y(\register_file_i/_1572_ ),
    .A(net1919),
    .B(\register_file_i/_1571_ ));
 sg13g2_mux4_1 \register_file_i/_4634_  (.S0(net2025),
    .A0(\register_file_i/rf_reg_517_ ),
    .A1(\register_file_i/rf_reg_549_ ),
    .A2(\register_file_i/rf_reg_581_ ),
    .A3(\register_file_i/rf_reg_613_ ),
    .S1(net544),
    .X(\register_file_i/_1573_ ));
 sg13g2_mux4_1 \register_file_i/_4635_  (.S0(net2013),
    .A0(\register_file_i/rf_reg_645_ ),
    .A1(\register_file_i/rf_reg_677_ ),
    .A2(\register_file_i/rf_reg_709_ ),
    .A3(\register_file_i/rf_reg_741_ ),
    .S1(net542),
    .X(\register_file_i/_1574_ ));
 sg13g2_mux2_1 \register_file_i/_4636_  (.A0(\register_file_i/rf_reg_389_ ),
    .A1(\register_file_i/rf_reg_421_ ),
    .S(net2020),
    .X(\register_file_i/_1575_ ));
 sg13g2_mux2_1 \register_file_i/_4637_  (.A0(\register_file_i/rf_reg_453_ ),
    .A1(\register_file_i/rf_reg_485_ ),
    .S(net2012),
    .X(\register_file_i/_1576_ ));
 sg13g2_a22oi_1 \register_file_i/_4638_  (.Y(\register_file_i/_1577_ ),
    .B1(\register_file_i/_1576_ ),
    .B2(net1820),
    .A2(\register_file_i/_1575_ ),
    .A1(net1837));
 sg13g2_buf_2 fanout334 (.A(_07486_),
    .X(net334));
 sg13g2_buf_2 fanout333 (.A(_07619_),
    .X(net333));
 sg13g2_mux2_1 \register_file_i/_4641_  (.A0(\register_file_i/rf_reg_325_ ),
    .A1(\register_file_i/rf_reg_357_ ),
    .S(net2020),
    .X(\register_file_i/_1580_ ));
 sg13g2_mux2_1 \register_file_i/_4642_  (.A0(\register_file_i/rf_reg_261_ ),
    .A1(\register_file_i/rf_reg_293_ ),
    .S(net2020),
    .X(\register_file_i/_1581_ ));
 sg13g2_a22oi_1 \register_file_i/_4643_  (.Y(\register_file_i/_1582_ ),
    .B1(\register_file_i/_1581_ ),
    .B2(net1799),
    .A2(\register_file_i/_1580_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4644_  (.A1(\register_file_i/_1577_ ),
    .A2(\register_file_i/_1582_ ),
    .Y(\register_file_i/_1583_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4645_  (.B2(net1693),
    .C1(\register_file_i/_1583_ ),
    .B1(\register_file_i/_1574_ ),
    .A1(net1792),
    .Y(\register_file_i/_1584_ ),
    .A2(\register_file_i/_1573_ ));
 sg13g2_nand3_1 \register_file_i/_4646_  (.B(\register_file_i/_1572_ ),
    .C(\register_file_i/_1584_ ),
    .A(\register_file_i/_1564_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_5_ ));
 sg13g2_buf_2 fanout332 (.A(_01779_),
    .X(net332));
 sg13g2_mux2_1 \register_file_i/_4648_  (.A0(\register_file_i/rf_reg_900_ ),
    .A1(\register_file_i/rf_reg_932_ ),
    .S(net2066),
    .X(\register_file_i/_1586_ ));
 sg13g2_mux2_1 \register_file_i/_4649_  (.A0(\register_file_i/rf_reg_964_ ),
    .A1(\register_file_i/rf_reg_996_ ),
    .S(net2066),
    .X(\register_file_i/_1587_ ));
 sg13g2_buf_2 fanout331 (.A(net332),
    .X(net331));
 sg13g2_a22oi_1 \register_file_i/_4651_  (.Y(\register_file_i/_1589_ ),
    .B1(\register_file_i/_1587_ ),
    .B2(net1832),
    .A2(\register_file_i/_1586_ ),
    .A1(net1848));
 sg13g2_buf_2 fanout330 (.A(net332),
    .X(net330));
 sg13g2_mux2_1 \register_file_i/_4653_  (.A0(\register_file_i/rf_reg_836_ ),
    .A1(\register_file_i/rf_reg_868_ ),
    .S(net2067),
    .X(\register_file_i/_1591_ ));
 sg13g2_mux2_1 \register_file_i/_4654_  (.A0(\register_file_i/rf_reg_772_ ),
    .A1(\register_file_i/rf_reg_804_ ),
    .S(net2066),
    .X(\register_file_i/_1592_ ));
 sg13g2_buf_2 fanout329 (.A(net332),
    .X(net329));
 sg13g2_a22oi_1 \register_file_i/_4656_  (.Y(\register_file_i/_1594_ ),
    .B1(\register_file_i/_1592_ ),
    .B2(net1805),
    .A2(\register_file_i/_1591_ ),
    .A1(net1816));
 sg13g2_buf_2 fanout328 (.A(_03332_),
    .X(net328));
 sg13g2_a21o_1 \register_file_i/_4658_  (.A2(\register_file_i/_1594_ ),
    .A1(\register_file_i/_1589_ ),
    .B1(net1925),
    .X(\register_file_i/_1596_ ));
 sg13g2_buf_2 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_2 fanout326 (.A(net328),
    .X(net326));
 sg13g2_mux2_1 \register_file_i/_4661_  (.A0(\register_file_i/rf_reg_36_ ),
    .A1(\register_file_i/rf_reg_100_ ),
    .S(net535),
    .X(\register_file_i/_1599_ ));
 sg13g2_a22oi_1 \register_file_i/_4662_  (.Y(\register_file_i/_1600_ ),
    .B1(\register_file_i/_1599_ ),
    .B2(net2069),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_68_ ));
 sg13g2_mux2_1 \register_file_i/_4663_  (.A0(\register_file_i/rf_reg_196_ ),
    .A1(\register_file_i/rf_reg_228_ ),
    .S(net2069),
    .X(\register_file_i/_1601_ ));
 sg13g2_mux2_1 \register_file_i/_4664_  (.A0(\register_file_i/rf_reg_132_ ),
    .A1(\register_file_i/rf_reg_164_ ),
    .S(net2070),
    .X(\register_file_i/_1602_ ));
 sg13g2_a22oi_1 \register_file_i/_4665_  (.Y(\register_file_i/_1603_ ),
    .B1(\register_file_i/_1602_ ),
    .B2(net1848),
    .A2(\register_file_i/_1601_ ),
    .A1(net1831));
 sg13g2_o21ai_1 \register_file_i/_4666_  (.B1(\register_file_i/_1603_ ),
    .Y(\register_file_i/_1604_ ),
    .A1(net529),
    .A2(\register_file_i/_1600_ ));
 sg13g2_nand2_1 \register_file_i/_4667_  (.Y(\register_file_i/_1605_ ),
    .A(net1919),
    .B(\register_file_i/_1604_ ));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(net328));
 sg13g2_mux4_1 \register_file_i/_4669_  (.S0(net2024),
    .A0(\register_file_i/rf_reg_516_ ),
    .A1(\register_file_i/rf_reg_548_ ),
    .A2(\register_file_i/rf_reg_580_ ),
    .A3(\register_file_i/rf_reg_612_ ),
    .S1(net543),
    .X(\register_file_i/_1607_ ));
 sg13g2_mux4_1 \register_file_i/_4670_  (.S0(net2024),
    .A0(\register_file_i/rf_reg_644_ ),
    .A1(\register_file_i/rf_reg_676_ ),
    .A2(\register_file_i/rf_reg_708_ ),
    .A3(\register_file_i/rf_reg_740_ ),
    .S1(net542),
    .X(\register_file_i/_1608_ ));
 sg13g2_buf_2 fanout324 (.A(_03332_),
    .X(net324));
 sg13g2_mux2_1 \register_file_i/_4672_  (.A0(\register_file_i/rf_reg_388_ ),
    .A1(\register_file_i/rf_reg_420_ ),
    .S(net2022),
    .X(\register_file_i/_1610_ ));
 sg13g2_mux2_1 \register_file_i/_4673_  (.A0(\register_file_i/rf_reg_452_ ),
    .A1(\register_file_i/rf_reg_484_ ),
    .S(net2022),
    .X(\register_file_i/_1611_ ));
 sg13g2_a22oi_1 \register_file_i/_4674_  (.Y(\register_file_i/_1612_ ),
    .B1(\register_file_i/_1611_ ),
    .B2(net1821),
    .A2(\register_file_i/_1610_ ),
    .A1(net1838));
 sg13g2_mux2_1 \register_file_i/_4675_  (.A0(\register_file_i/rf_reg_324_ ),
    .A1(\register_file_i/rf_reg_356_ ),
    .S(net2023),
    .X(\register_file_i/_1613_ ));
 sg13g2_mux2_1 \register_file_i/_4676_  (.A0(\register_file_i/rf_reg_260_ ),
    .A1(\register_file_i/rf_reg_292_ ),
    .S(net2022),
    .X(\register_file_i/_1614_ ));
 sg13g2_a22oi_1 \register_file_i/_4677_  (.Y(\register_file_i/_1615_ ),
    .B1(\register_file_i/_1614_ ),
    .B2(net1804),
    .A2(\register_file_i/_1613_ ),
    .A1(net1815));
 sg13g2_a21oi_1 \register_file_i/_4678_  (.A1(\register_file_i/_1612_ ),
    .A2(\register_file_i/_1615_ ),
    .Y(\register_file_i/_1616_ ),
    .B1(net1788));
 sg13g2_a221oi_1 \register_file_i/_4679_  (.B2(net1695),
    .C1(\register_file_i/_1616_ ),
    .B1(\register_file_i/_1608_ ),
    .A1(net1794),
    .Y(\register_file_i/_1617_ ),
    .A2(\register_file_i/_1607_ ));
 sg13g2_nand3_1 \register_file_i/_4680_  (.B(\register_file_i/_1605_ ),
    .C(\register_file_i/_1617_ ),
    .A(\register_file_i/_1596_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_mux2_1 \register_file_i/_4681_  (.A0(\register_file_i/rf_reg_387_ ),
    .A1(\register_file_i/rf_reg_419_ ),
    .S(net2053),
    .X(\register_file_i/_1618_ ));
 sg13g2_mux2_1 \register_file_i/_4682_  (.A0(\register_file_i/rf_reg_451_ ),
    .A1(\register_file_i/rf_reg_483_ ),
    .S(net2054),
    .X(\register_file_i/_1619_ ));
 sg13g2_a22oi_1 \register_file_i/_4683_  (.Y(\register_file_i/_1620_ ),
    .B1(\register_file_i/_1619_ ),
    .B2(net1828),
    .A2(\register_file_i/_1618_ ),
    .A1(net1845));
 sg13g2_buf_2 fanout323 (.A(_04062_),
    .X(net323));
 sg13g2_mux2_1 \register_file_i/_4685_  (.A0(\register_file_i/rf_reg_323_ ),
    .A1(\register_file_i/rf_reg_355_ ),
    .S(net2055),
    .X(\register_file_i/_1622_ ));
 sg13g2_mux2_1 \register_file_i/_4686_  (.A0(\register_file_i/rf_reg_259_ ),
    .A1(\register_file_i/rf_reg_291_ ),
    .S(net2054),
    .X(\register_file_i/_1623_ ));
 sg13g2_a22oi_1 \register_file_i/_4687_  (.Y(\register_file_i/_1624_ ),
    .B1(\register_file_i/_1623_ ),
    .B2(net1804),
    .A2(\register_file_i/_1622_ ),
    .A1(net1815));
 sg13g2_a21o_1 \register_file_i/_4688_  (.A2(\register_file_i/_1624_ ),
    .A1(\register_file_i/_1620_ ),
    .B1(net1788),
    .X(\register_file_i/_1625_ ));
 sg13g2_buf_2 fanout322 (.A(net323),
    .X(net322));
 sg13g2_mux2_1 \register_file_i/_4690_  (.A0(\register_file_i/rf_reg_35_ ),
    .A1(\register_file_i/rf_reg_99_ ),
    .S(net532),
    .X(\register_file_i/_1627_ ));
 sg13g2_nand2_1 \register_file_i/_4691_  (.Y(\register_file_i/_1628_ ),
    .A(net2062),
    .B(\register_file_i/_1627_ ));
 sg13g2_nand3b_1 \register_file_i/_4692_  (.B(net537),
    .C(\register_file_i/rf_reg_67_ ),
    .Y(\register_file_i/_1629_ ),
    .A_N(net2063));
 sg13g2_a21oi_1 \register_file_i/_4693_  (.A1(\register_file_i/_1628_ ),
    .A2(\register_file_i/_1629_ ),
    .Y(\register_file_i/_1630_ ),
    .B1(net529));
 sg13g2_mux2_1 \register_file_i/_4694_  (.A0(\register_file_i/rf_reg_131_ ),
    .A1(\register_file_i/rf_reg_163_ ),
    .S(net2054),
    .X(\register_file_i/_1631_ ));
 sg13g2_mux2_1 \register_file_i/_4695_  (.A0(\register_file_i/rf_reg_195_ ),
    .A1(\register_file_i/rf_reg_227_ ),
    .S(net2054),
    .X(\register_file_i/_1632_ ));
 sg13g2_a22oi_1 \register_file_i/_4696_  (.Y(\register_file_i/_1633_ ),
    .B1(\register_file_i/_1632_ ),
    .B2(net1828),
    .A2(\register_file_i/_1631_ ),
    .A1(net1845));
 sg13g2_inv_1 \register_file_i/_4697_  (.Y(\register_file_i/_1634_ ),
    .A(\register_file_i/_1633_ ));
 sg13g2_o21ai_1 \register_file_i/_4698_  (.B1(net1920),
    .Y(\register_file_i/_1635_ ),
    .A1(\register_file_i/_1630_ ),
    .A2(\register_file_i/_1634_ ));
 sg13g2_mux4_1 \register_file_i/_4699_  (.S0(net2024),
    .A0(\register_file_i/rf_reg_643_ ),
    .A1(\register_file_i/rf_reg_675_ ),
    .A2(\register_file_i/rf_reg_707_ ),
    .A3(\register_file_i/rf_reg_739_ ),
    .S1(net543),
    .X(\register_file_i/_1636_ ));
 sg13g2_buf_2 fanout321 (.A(net323),
    .X(net321));
 sg13g2_mux4_1 \register_file_i/_4701_  (.S0(net2028),
    .A0(\register_file_i/rf_reg_515_ ),
    .A1(\register_file_i/rf_reg_547_ ),
    .A2(\register_file_i/rf_reg_579_ ),
    .A3(\register_file_i/rf_reg_611_ ),
    .S1(net545),
    .X(\register_file_i/_1638_ ));
 sg13g2_buf_2 fanout320 (.A(net323),
    .X(net320));
 sg13g2_mux2_1 \register_file_i/_4703_  (.A0(\register_file_i/rf_reg_771_ ),
    .A1(\register_file_i/rf_reg_803_ ),
    .S(net2023),
    .X(\register_file_i/_1640_ ));
 sg13g2_mux2_1 \register_file_i/_4704_  (.A0(\register_file_i/rf_reg_899_ ),
    .A1(\register_file_i/rf_reg_931_ ),
    .S(net2023),
    .X(\register_file_i/_1641_ ));
 sg13g2_a22oi_1 \register_file_i/_4705_  (.Y(\register_file_i/_1642_ ),
    .B1(\register_file_i/_1641_ ),
    .B2(net1838),
    .A2(\register_file_i/_1640_ ),
    .A1(net1804));
 sg13g2_mux2_1 \register_file_i/_4706_  (.A0(\register_file_i/rf_reg_835_ ),
    .A1(\register_file_i/rf_reg_867_ ),
    .S(net2023),
    .X(\register_file_i/_1643_ ));
 sg13g2_mux2_1 \register_file_i/_4707_  (.A0(\register_file_i/rf_reg_963_ ),
    .A1(\register_file_i/rf_reg_995_ ),
    .S(net2022),
    .X(\register_file_i/_1644_ ));
 sg13g2_a22oi_1 \register_file_i/_4708_  (.Y(\register_file_i/_1645_ ),
    .B1(\register_file_i/_1644_ ),
    .B2(net1821),
    .A2(\register_file_i/_1643_ ),
    .A1(net1815));
 sg13g2_a21oi_1 \register_file_i/_4709_  (.A1(\register_file_i/_1642_ ),
    .A2(\register_file_i/_1645_ ),
    .Y(\register_file_i/_1646_ ),
    .B1(net1927));
 sg13g2_a221oi_1 \register_file_i/_4710_  (.B2(net1793),
    .C1(\register_file_i/_1646_ ),
    .B1(\register_file_i/_1638_ ),
    .A1(net1695),
    .Y(\register_file_i/_1647_ ),
    .A2(\register_file_i/_1636_ ));
 sg13g2_nand3_1 \register_file_i/_4711_  (.B(\register_file_i/_1635_ ),
    .C(\register_file_i/_1647_ ),
    .A(\register_file_i/_1625_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_mux2_1 \register_file_i/_4712_  (.A0(\register_file_i/rf_reg_386_ ),
    .A1(\register_file_i/rf_reg_418_ ),
    .S(net2054),
    .X(\register_file_i/_1648_ ));
 sg13g2_mux2_1 \register_file_i/_4713_  (.A0(\register_file_i/rf_reg_450_ ),
    .A1(\register_file_i/rf_reg_482_ ),
    .S(net2054),
    .X(\register_file_i/_1649_ ));
 sg13g2_a22oi_1 \register_file_i/_4714_  (.Y(\register_file_i/_1650_ ),
    .B1(\register_file_i/_1649_ ),
    .B2(net1828),
    .A2(\register_file_i/_1648_ ),
    .A1(net1845));
 sg13g2_mux2_1 \register_file_i/_4715_  (.A0(\register_file_i/rf_reg_322_ ),
    .A1(\register_file_i/rf_reg_354_ ),
    .S(net2054),
    .X(\register_file_i/_1651_ ));
 sg13g2_mux2_1 \register_file_i/_4716_  (.A0(\register_file_i/rf_reg_258_ ),
    .A1(\register_file_i/rf_reg_290_ ),
    .S(net2054),
    .X(\register_file_i/_1652_ ));
 sg13g2_a22oi_1 \register_file_i/_4717_  (.Y(\register_file_i/_1653_ ),
    .B1(\register_file_i/_1652_ ),
    .B2(net1804),
    .A2(\register_file_i/_1651_ ),
    .A1(net1815));
 sg13g2_a21o_1 \register_file_i/_4718_  (.A2(\register_file_i/_1653_ ),
    .A1(\register_file_i/_1650_ ),
    .B1(net1788),
    .X(\register_file_i/_1654_ ));
 sg13g2_mux2_1 \register_file_i/_4719_  (.A0(\register_file_i/rf_reg_34_ ),
    .A1(\register_file_i/rf_reg_98_ ),
    .S(net532),
    .X(\register_file_i/_1655_ ));
 sg13g2_nand2_1 \register_file_i/_4720_  (.Y(\register_file_i/_1656_ ),
    .A(net2062),
    .B(\register_file_i/_1655_ ));
 sg13g2_nand3b_1 \register_file_i/_4721_  (.B(net537),
    .C(\register_file_i/rf_reg_66_ ),
    .Y(\register_file_i/_1657_ ),
    .A_N(net2063));
 sg13g2_a21oi_1 \register_file_i/_4722_  (.A1(\register_file_i/_1656_ ),
    .A2(\register_file_i/_1657_ ),
    .Y(\register_file_i/_1658_ ),
    .B1(net529));
 sg13g2_mux2_1 \register_file_i/_4723_  (.A0(\register_file_i/rf_reg_130_ ),
    .A1(\register_file_i/rf_reg_162_ ),
    .S(net2060),
    .X(\register_file_i/_1659_ ));
 sg13g2_mux2_1 \register_file_i/_4724_  (.A0(\register_file_i/rf_reg_194_ ),
    .A1(\register_file_i/rf_reg_226_ ),
    .S(net2060),
    .X(\register_file_i/_1660_ ));
 sg13g2_a22oi_1 \register_file_i/_4725_  (.Y(\register_file_i/_1661_ ),
    .B1(\register_file_i/_1660_ ),
    .B2(net1829),
    .A2(\register_file_i/_1659_ ),
    .A1(net1846));
 sg13g2_inv_1 \register_file_i/_4726_  (.Y(\register_file_i/_1662_ ),
    .A(\register_file_i/_1661_ ));
 sg13g2_o21ai_1 \register_file_i/_4727_  (.B1(net1920),
    .Y(\register_file_i/_1663_ ),
    .A1(\register_file_i/_1658_ ),
    .A2(\register_file_i/_1662_ ));
 sg13g2_mux4_1 \register_file_i/_4728_  (.S0(net2028),
    .A0(\register_file_i/rf_reg_642_ ),
    .A1(\register_file_i/rf_reg_674_ ),
    .A2(\register_file_i/rf_reg_706_ ),
    .A3(\register_file_i/rf_reg_738_ ),
    .S1(net543),
    .X(\register_file_i/_1664_ ));
 sg13g2_mux4_1 \register_file_i/_4729_  (.S0(net2028),
    .A0(\register_file_i/rf_reg_514_ ),
    .A1(\register_file_i/rf_reg_546_ ),
    .A2(\register_file_i/rf_reg_578_ ),
    .A3(\register_file_i/rf_reg_610_ ),
    .S1(net545),
    .X(\register_file_i/_1665_ ));
 sg13g2_mux2_1 \register_file_i/_4730_  (.A0(\register_file_i/rf_reg_770_ ),
    .A1(\register_file_i/rf_reg_802_ ),
    .S(net2053),
    .X(\register_file_i/_1666_ ));
 sg13g2_mux2_1 \register_file_i/_4731_  (.A0(\register_file_i/rf_reg_898_ ),
    .A1(\register_file_i/rf_reg_930_ ),
    .S(net2053),
    .X(\register_file_i/_1667_ ));
 sg13g2_a22oi_1 \register_file_i/_4732_  (.Y(\register_file_i/_1668_ ),
    .B1(\register_file_i/_1667_ ),
    .B2(net1845),
    .A2(\register_file_i/_1666_ ),
    .A1(net1804));
 sg13g2_mux2_1 \register_file_i/_4733_  (.A0(\register_file_i/rf_reg_834_ ),
    .A1(\register_file_i/rf_reg_866_ ),
    .S(net2053),
    .X(\register_file_i/_1669_ ));
 sg13g2_mux2_1 \register_file_i/_4734_  (.A0(\register_file_i/rf_reg_962_ ),
    .A1(\register_file_i/rf_reg_994_ ),
    .S(net2053),
    .X(\register_file_i/_1670_ ));
 sg13g2_a22oi_1 \register_file_i/_4735_  (.Y(\register_file_i/_1671_ ),
    .B1(\register_file_i/_1670_ ),
    .B2(net1828),
    .A2(\register_file_i/_1669_ ),
    .A1(net1815));
 sg13g2_a21oi_2 \register_file_i/_4736_  (.B1(net1927),
    .Y(\register_file_i/_1672_ ),
    .A2(\register_file_i/_1671_ ),
    .A1(\register_file_i/_1668_ ));
 sg13g2_a221oi_1 \register_file_i/_4737_  (.B2(net1793),
    .C1(\register_file_i/_1672_ ),
    .B1(\register_file_i/_1665_ ),
    .A1(net1695),
    .Y(\register_file_i/_1673_ ),
    .A2(\register_file_i/_1664_ ));
 sg13g2_nand3_1 \register_file_i/_4738_  (.B(\register_file_i/_1663_ ),
    .C(\register_file_i/_1673_ ),
    .A(\register_file_i/_1654_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_mux2_1 \register_file_i/_4739_  (.A0(\register_file_i/rf_reg_924_ ),
    .A1(\register_file_i/rf_reg_956_ ),
    .S(net2072),
    .X(\register_file_i/_1674_ ));
 sg13g2_mux2_1 \register_file_i/_4740_  (.A0(\register_file_i/rf_reg_988_ ),
    .A1(\register_file_i/rf_reg_1020_ ),
    .S(net2072),
    .X(\register_file_i/_1675_ ));
 sg13g2_a22oi_1 \register_file_i/_4741_  (.Y(\register_file_i/_1676_ ),
    .B1(\register_file_i/_1675_ ),
    .B2(net1833),
    .A2(\register_file_i/_1674_ ),
    .A1(net1850));
 sg13g2_mux2_1 \register_file_i/_4742_  (.A0(\register_file_i/rf_reg_860_ ),
    .A1(\register_file_i/rf_reg_892_ ),
    .S(net2073),
    .X(\register_file_i/_1677_ ));
 sg13g2_mux2_1 \register_file_i/_4743_  (.A0(\register_file_i/rf_reg_796_ ),
    .A1(\register_file_i/rf_reg_828_ ),
    .S(net2071),
    .X(\register_file_i/_1678_ ));
 sg13g2_a22oi_1 \register_file_i/_4744_  (.Y(\register_file_i/_1679_ ),
    .B1(\register_file_i/_1678_ ),
    .B2(net1806),
    .A2(\register_file_i/_1677_ ),
    .A1(net1817));
 sg13g2_a21o_1 \register_file_i/_4745_  (.A2(\register_file_i/_1679_ ),
    .A1(\register_file_i/_1676_ ),
    .B1(net1926),
    .X(\register_file_i/_1680_ ));
 sg13g2_mux2_1 \register_file_i/_4746_  (.A0(\register_file_i/rf_reg_60_ ),
    .A1(\register_file_i/rf_reg_124_ ),
    .S(net535),
    .X(\register_file_i/_1681_ ));
 sg13g2_a22oi_1 \register_file_i/_4747_  (.Y(\register_file_i/_1682_ ),
    .B1(\register_file_i/_1681_ ),
    .B2(net2074),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_92_ ));
 sg13g2_mux2_1 \register_file_i/_4748_  (.A0(\register_file_i/rf_reg_220_ ),
    .A1(\register_file_i/rf_reg_252_ ),
    .S(net2069),
    .X(\register_file_i/_1683_ ));
 sg13g2_mux2_1 \register_file_i/_4749_  (.A0(\register_file_i/rf_reg_156_ ),
    .A1(\register_file_i/rf_reg_188_ ),
    .S(net2074),
    .X(\register_file_i/_1684_ ));
 sg13g2_a22oi_1 \register_file_i/_4750_  (.Y(\register_file_i/_1685_ ),
    .B1(\register_file_i/_1684_ ),
    .B2(net1849),
    .A2(\register_file_i/_1683_ ),
    .A1(net1831));
 sg13g2_o21ai_1 \register_file_i/_4751_  (.B1(\register_file_i/_1685_ ),
    .Y(\register_file_i/_1686_ ),
    .A1(net529),
    .A2(\register_file_i/_1682_ ));
 sg13g2_nand2_1 \register_file_i/_4752_  (.Y(\register_file_i/_1687_ ),
    .A(net1919),
    .B(\register_file_i/_1686_ ));
 sg13g2_mux4_1 \register_file_i/_4753_  (.S0(net2028),
    .A0(\register_file_i/rf_reg_540_ ),
    .A1(\register_file_i/rf_reg_572_ ),
    .A2(\register_file_i/rf_reg_604_ ),
    .A3(\register_file_i/rf_reg_636_ ),
    .S1(net543),
    .X(\register_file_i/_1688_ ));
 sg13g2_mux4_1 \register_file_i/_4754_  (.S0(net2027),
    .A0(\register_file_i/rf_reg_668_ ),
    .A1(\register_file_i/rf_reg_700_ ),
    .A2(\register_file_i/rf_reg_732_ ),
    .A3(\register_file_i/rf_reg_764_ ),
    .S1(net545),
    .X(\register_file_i/_1689_ ));
 sg13g2_mux2_1 \register_file_i/_4755_  (.A0(\register_file_i/rf_reg_412_ ),
    .A1(\register_file_i/rf_reg_444_ ),
    .S(net2028),
    .X(\register_file_i/_1690_ ));
 sg13g2_mux2_1 \register_file_i/_4756_  (.A0(\register_file_i/rf_reg_476_ ),
    .A1(\register_file_i/rf_reg_508_ ),
    .S(net2028),
    .X(\register_file_i/_1691_ ));
 sg13g2_a22oi_1 \register_file_i/_4757_  (.Y(\register_file_i/_1692_ ),
    .B1(\register_file_i/_1691_ ),
    .B2(net1822),
    .A2(\register_file_i/_1690_ ),
    .A1(net1839));
 sg13g2_mux2_1 \register_file_i/_4758_  (.A0(\register_file_i/rf_reg_348_ ),
    .A1(\register_file_i/rf_reg_380_ ),
    .S(net2028),
    .X(\register_file_i/_1693_ ));
 sg13g2_mux2_1 \register_file_i/_4759_  (.A0(\register_file_i/rf_reg_284_ ),
    .A1(\register_file_i/rf_reg_316_ ),
    .S(net2028),
    .X(\register_file_i/_1694_ ));
 sg13g2_a22oi_1 \register_file_i/_4760_  (.Y(\register_file_i/_1695_ ),
    .B1(\register_file_i/_1694_ ),
    .B2(net1799),
    .A2(\register_file_i/_1693_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4761_  (.A1(\register_file_i/_1692_ ),
    .A2(\register_file_i/_1695_ ),
    .Y(\register_file_i/_1696_ ),
    .B1(net1789));
 sg13g2_a221oi_1 \register_file_i/_4762_  (.B2(net1695),
    .C1(\register_file_i/_1696_ ),
    .B1(\register_file_i/_1689_ ),
    .A1(net1794),
    .Y(\register_file_i/_1697_ ),
    .A2(\register_file_i/_1688_ ));
 sg13g2_nand3_1 \register_file_i/_4763_  (.B(\register_file_i/_1687_ ),
    .C(\register_file_i/_1697_ ),
    .A(\register_file_i/_1680_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_28_ ));
 sg13g2_mux2_1 \register_file_i/_4764_  (.A0(\register_file_i/rf_reg_385_ ),
    .A1(\register_file_i/rf_reg_417_ ),
    .S(net2060),
    .X(\register_file_i/_1698_ ));
 sg13g2_mux2_1 \register_file_i/_4765_  (.A0(\register_file_i/rf_reg_449_ ),
    .A1(\register_file_i/rf_reg_481_ ),
    .S(net2060),
    .X(\register_file_i/_1699_ ));
 sg13g2_a22oi_1 \register_file_i/_4766_  (.Y(\register_file_i/_1700_ ),
    .B1(\register_file_i/_1699_ ),
    .B2(net1830),
    .A2(\register_file_i/_1698_ ),
    .A1(net1847));
 sg13g2_mux2_1 \register_file_i/_4767_  (.A0(\register_file_i/rf_reg_321_ ),
    .A1(\register_file_i/rf_reg_353_ ),
    .S(net2060),
    .X(\register_file_i/_1701_ ));
 sg13g2_mux2_1 \register_file_i/_4768_  (.A0(\register_file_i/rf_reg_257_ ),
    .A1(\register_file_i/rf_reg_289_ ),
    .S(net2060),
    .X(\register_file_i/_1702_ ));
 sg13g2_a22oi_1 \register_file_i/_4769_  (.Y(\register_file_i/_1703_ ),
    .B1(\register_file_i/_1702_ ),
    .B2(net1806),
    .A2(\register_file_i/_1701_ ),
    .A1(net1817));
 sg13g2_a21o_1 \register_file_i/_4770_  (.A2(\register_file_i/_1703_ ),
    .A1(\register_file_i/_1700_ ),
    .B1(net1788),
    .X(\register_file_i/_1704_ ));
 sg13g2_mux2_1 \register_file_i/_4771_  (.A0(\register_file_i/rf_reg_33_ ),
    .A1(\register_file_i/rf_reg_97_ ),
    .S(net532),
    .X(\register_file_i/_1705_ ));
 sg13g2_nand2_1 \register_file_i/_4772_  (.Y(\register_file_i/_1706_ ),
    .A(net2061),
    .B(\register_file_i/_1705_ ));
 sg13g2_nand3b_1 \register_file_i/_4773_  (.B(net537),
    .C(\register_file_i/rf_reg_65_ ),
    .Y(\register_file_i/_1707_ ),
    .A_N(net2061));
 sg13g2_a21oi_1 \register_file_i/_4774_  (.A1(\register_file_i/_1706_ ),
    .A2(\register_file_i/_1707_ ),
    .Y(\register_file_i/_1708_ ),
    .B1(net525));
 sg13g2_mux2_1 \register_file_i/_4775_  (.A0(\register_file_i/rf_reg_129_ ),
    .A1(\register_file_i/rf_reg_161_ ),
    .S(net2061),
    .X(\register_file_i/_1709_ ));
 sg13g2_mux2_1 \register_file_i/_4776_  (.A0(\register_file_i/rf_reg_193_ ),
    .A1(\register_file_i/rf_reg_225_ ),
    .S(net2061),
    .X(\register_file_i/_1710_ ));
 sg13g2_a22oi_1 \register_file_i/_4777_  (.Y(\register_file_i/_1711_ ),
    .B1(\register_file_i/_1710_ ),
    .B2(net1829),
    .A2(\register_file_i/_1709_ ),
    .A1(net1846));
 sg13g2_inv_1 \register_file_i/_4778_  (.Y(\register_file_i/_1712_ ),
    .A(\register_file_i/_1711_ ));
 sg13g2_o21ai_1 \register_file_i/_4779_  (.B1(net1920),
    .Y(\register_file_i/_1713_ ),
    .A1(\register_file_i/_1708_ ),
    .A2(\register_file_i/_1712_ ));
 sg13g2_mux4_1 \register_file_i/_4780_  (.S0(net2025),
    .A0(\register_file_i/rf_reg_641_ ),
    .A1(\register_file_i/rf_reg_673_ ),
    .A2(\register_file_i/rf_reg_705_ ),
    .A3(\register_file_i/rf_reg_737_ ),
    .S1(net539),
    .X(\register_file_i/_1714_ ));
 sg13g2_mux4_1 \register_file_i/_4781_  (.S0(net2025),
    .A0(\register_file_i/rf_reg_513_ ),
    .A1(\register_file_i/rf_reg_545_ ),
    .A2(\register_file_i/rf_reg_577_ ),
    .A3(\register_file_i/rf_reg_609_ ),
    .S1(net545),
    .X(\register_file_i/_1715_ ));
 sg13g2_mux2_1 \register_file_i/_4782_  (.A0(\register_file_i/rf_reg_769_ ),
    .A1(\register_file_i/rf_reg_801_ ),
    .S(net2025),
    .X(\register_file_i/_1716_ ));
 sg13g2_mux2_1 \register_file_i/_4783_  (.A0(\register_file_i/rf_reg_897_ ),
    .A1(\register_file_i/rf_reg_929_ ),
    .S(net2025),
    .X(\register_file_i/_1717_ ));
 sg13g2_a22oi_1 \register_file_i/_4784_  (.Y(\register_file_i/_1718_ ),
    .B1(\register_file_i/_1717_ ),
    .B2(net1838),
    .A2(\register_file_i/_1716_ ),
    .A1(net1799));
 sg13g2_mux2_1 \register_file_i/_4785_  (.A0(\register_file_i/rf_reg_833_ ),
    .A1(\register_file_i/rf_reg_865_ ),
    .S(net2026),
    .X(\register_file_i/_1719_ ));
 sg13g2_mux2_1 \register_file_i/_4786_  (.A0(\register_file_i/rf_reg_961_ ),
    .A1(\register_file_i/rf_reg_993_ ),
    .S(net2025),
    .X(\register_file_i/_1720_ ));
 sg13g2_a22oi_1 \register_file_i/_4787_  (.Y(\register_file_i/_1721_ ),
    .B1(\register_file_i/_1720_ ),
    .B2(net1821),
    .A2(\register_file_i/_1719_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4788_  (.A1(\register_file_i/_1718_ ),
    .A2(\register_file_i/_1721_ ),
    .Y(\register_file_i/_1722_ ),
    .B1(net1927));
 sg13g2_a221oi_1 \register_file_i/_4789_  (.B2(net1793),
    .C1(\register_file_i/_1722_ ),
    .B1(\register_file_i/_1715_ ),
    .A1(net1694),
    .Y(\register_file_i/_1723_ ),
    .A2(\register_file_i/_1714_ ));
 sg13g2_nand3_1 \register_file_i/_4790_  (.B(\register_file_i/_1713_ ),
    .C(\register_file_i/_1723_ ),
    .A(\register_file_i/_1704_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_mux2_1 \register_file_i/_4791_  (.A0(\register_file_i/rf_reg_384_ ),
    .A1(\register_file_i/rf_reg_416_ ),
    .S(net2060),
    .X(\register_file_i/_1724_ ));
 sg13g2_mux2_1 \register_file_i/_4792_  (.A0(\register_file_i/rf_reg_448_ ),
    .A1(\register_file_i/rf_reg_480_ ),
    .S(net2061),
    .X(\register_file_i/_1725_ ));
 sg13g2_a22oi_1 \register_file_i/_4793_  (.Y(\register_file_i/_1726_ ),
    .B1(\register_file_i/_1725_ ),
    .B2(net1830),
    .A2(\register_file_i/_1724_ ),
    .A1(net1847));
 sg13g2_mux2_1 \register_file_i/_4794_  (.A0(\register_file_i/rf_reg_320_ ),
    .A1(\register_file_i/rf_reg_352_ ),
    .S(net2061),
    .X(\register_file_i/_1727_ ));
 sg13g2_mux2_1 \register_file_i/_4795_  (.A0(\register_file_i/rf_reg_256_ ),
    .A1(\register_file_i/rf_reg_288_ ),
    .S(net2060),
    .X(\register_file_i/_1728_ ));
 sg13g2_a22oi_1 \register_file_i/_4796_  (.Y(\register_file_i/_1729_ ),
    .B1(\register_file_i/_1728_ ),
    .B2(net1806),
    .A2(\register_file_i/_1727_ ),
    .A1(net1817));
 sg13g2_a21o_1 \register_file_i/_4797_  (.A2(\register_file_i/_1729_ ),
    .A1(\register_file_i/_1726_ ),
    .B1(net1788),
    .X(\register_file_i/_1730_ ));
 sg13g2_mux2_1 \register_file_i/_4798_  (.A0(\register_file_i/rf_reg_32_ ),
    .A1(\register_file_i/rf_reg_96_ ),
    .S(net532),
    .X(\register_file_i/_1731_ ));
 sg13g2_nand2_1 \register_file_i/_4799_  (.Y(\register_file_i/_1732_ ),
    .A(net2063),
    .B(\register_file_i/_1731_ ));
 sg13g2_nand3b_1 \register_file_i/_4800_  (.B(net537),
    .C(\register_file_i/rf_reg_64_ ),
    .Y(\register_file_i/_1733_ ),
    .A_N(net2063));
 sg13g2_a21oi_1 \register_file_i/_4801_  (.A1(\register_file_i/_1732_ ),
    .A2(\register_file_i/_1733_ ),
    .Y(\register_file_i/_1734_ ),
    .B1(net525));
 sg13g2_mux2_1 \register_file_i/_4802_  (.A0(\register_file_i/rf_reg_128_ ),
    .A1(\register_file_i/rf_reg_160_ ),
    .S(net2063),
    .X(\register_file_i/_1735_ ));
 sg13g2_mux2_1 \register_file_i/_4803_  (.A0(\register_file_i/rf_reg_192_ ),
    .A1(\register_file_i/rf_reg_224_ ),
    .S(net2063),
    .X(\register_file_i/_1736_ ));
 sg13g2_a22oi_1 \register_file_i/_4804_  (.Y(\register_file_i/_1737_ ),
    .B1(\register_file_i/_1736_ ),
    .B2(net1829),
    .A2(\register_file_i/_1735_ ),
    .A1(net1846));
 sg13g2_inv_1 \register_file_i/_4805_  (.Y(\register_file_i/_1738_ ),
    .A(\register_file_i/_1737_ ));
 sg13g2_o21ai_1 \register_file_i/_4806_  (.B1(net1920),
    .Y(\register_file_i/_1739_ ),
    .A1(\register_file_i/_1734_ ),
    .A2(\register_file_i/_1738_ ));
 sg13g2_mux4_1 \register_file_i/_4807_  (.S0(net2026),
    .A0(\register_file_i/rf_reg_640_ ),
    .A1(\register_file_i/rf_reg_672_ ),
    .A2(\register_file_i/rf_reg_704_ ),
    .A3(\register_file_i/rf_reg_736_ ),
    .S1(net539),
    .X(\register_file_i/_1740_ ));
 sg13g2_mux4_1 \register_file_i/_4808_  (.S0(net2025),
    .A0(\register_file_i/rf_reg_512_ ),
    .A1(\register_file_i/rf_reg_544_ ),
    .A2(\register_file_i/rf_reg_576_ ),
    .A3(\register_file_i/rf_reg_608_ ),
    .S1(net545),
    .X(\register_file_i/_1741_ ));
 sg13g2_mux2_1 \register_file_i/_4809_  (.A0(\register_file_i/rf_reg_768_ ),
    .A1(\register_file_i/rf_reg_800_ ),
    .S(net2042),
    .X(\register_file_i/_1742_ ));
 sg13g2_mux2_1 \register_file_i/_4810_  (.A0(\register_file_i/rf_reg_896_ ),
    .A1(\register_file_i/rf_reg_928_ ),
    .S(net2026),
    .X(\register_file_i/_1743_ ));
 sg13g2_a22oi_1 \register_file_i/_4811_  (.Y(\register_file_i/_1744_ ),
    .B1(\register_file_i/_1743_ ),
    .B2(net1842),
    .A2(\register_file_i/_1742_ ),
    .A1(net1801));
 sg13g2_mux2_1 \register_file_i/_4812_  (.A0(\register_file_i/rf_reg_832_ ),
    .A1(\register_file_i/rf_reg_864_ ),
    .S(net2026),
    .X(\register_file_i/_1745_ ));
 sg13g2_mux2_1 \register_file_i/_4813_  (.A0(\register_file_i/rf_reg_960_ ),
    .A1(\register_file_i/rf_reg_992_ ),
    .S(net2025),
    .X(\register_file_i/_1746_ ));
 sg13g2_a22oi_1 \register_file_i/_4814_  (.Y(\register_file_i/_1747_ ),
    .B1(\register_file_i/_1746_ ),
    .B2(net1821),
    .A2(\register_file_i/_1745_ ),
    .A1(net1810));
 sg13g2_a21oi_1 \register_file_i/_4815_  (.A1(\register_file_i/_1744_ ),
    .A2(\register_file_i/_1747_ ),
    .Y(\register_file_i/_1748_ ),
    .B1(net1927));
 sg13g2_a221oi_1 \register_file_i/_4816_  (.B2(net1793),
    .C1(\register_file_i/_1748_ ),
    .B1(\register_file_i/_1741_ ),
    .A1(net1694),
    .Y(\register_file_i/_1749_ ),
    .A2(\register_file_i/_1740_ ));
 sg13g2_nand3_1 \register_file_i/_4817_  (.B(\register_file_i/_1739_ ),
    .C(\register_file_i/_1749_ ),
    .A(\register_file_i/_1730_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_0_ ));
 sg13g2_mux2_1 \register_file_i/_4818_  (.A0(\register_file_i/rf_reg_923_ ),
    .A1(\register_file_i/rf_reg_955_ ),
    .S(net2074),
    .X(\register_file_i/_1750_ ));
 sg13g2_mux2_1 \register_file_i/_4819_  (.A0(\register_file_i/rf_reg_987_ ),
    .A1(\register_file_i/rf_reg_1019_ ),
    .S(net2073),
    .X(\register_file_i/_1751_ ));
 sg13g2_a22oi_1 \register_file_i/_4820_  (.Y(\register_file_i/_1752_ ),
    .B1(\register_file_i/_1751_ ),
    .B2(net1833),
    .A2(\register_file_i/_1750_ ),
    .A1(net1850));
 sg13g2_mux2_1 \register_file_i/_4821_  (.A0(\register_file_i/rf_reg_859_ ),
    .A1(\register_file_i/rf_reg_891_ ),
    .S(net2072),
    .X(\register_file_i/_1753_ ));
 sg13g2_mux2_1 \register_file_i/_4822_  (.A0(\register_file_i/rf_reg_795_ ),
    .A1(\register_file_i/rf_reg_827_ ),
    .S(net2072),
    .X(\register_file_i/_1754_ ));
 sg13g2_a22oi_1 \register_file_i/_4823_  (.Y(\register_file_i/_1755_ ),
    .B1(\register_file_i/_1754_ ),
    .B2(net1806),
    .A2(\register_file_i/_1753_ ),
    .A1(net1817));
 sg13g2_a21o_1 \register_file_i/_4824_  (.A2(\register_file_i/_1755_ ),
    .A1(\register_file_i/_1752_ ),
    .B1(net1926),
    .X(\register_file_i/_1756_ ));
 sg13g2_mux2_1 \register_file_i/_4825_  (.A0(\register_file_i/rf_reg_59_ ),
    .A1(\register_file_i/rf_reg_123_ ),
    .S(net535),
    .X(\register_file_i/_1757_ ));
 sg13g2_a22oi_1 \register_file_i/_4826_  (.Y(\register_file_i/_1758_ ),
    .B1(\register_file_i/_1757_ ),
    .B2(net2074),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_91_ ));
 sg13g2_mux2_1 \register_file_i/_4827_  (.A0(\register_file_i/rf_reg_219_ ),
    .A1(\register_file_i/rf_reg_251_ ),
    .S(net2074),
    .X(\register_file_i/_1759_ ));
 sg13g2_mux2_1 \register_file_i/_4828_  (.A0(\register_file_i/rf_reg_155_ ),
    .A1(\register_file_i/rf_reg_187_ ),
    .S(net2074),
    .X(\register_file_i/_1760_ ));
 sg13g2_a22oi_1 \register_file_i/_4829_  (.Y(\register_file_i/_1761_ ),
    .B1(\register_file_i/_1760_ ),
    .B2(net1849),
    .A2(\register_file_i/_1759_ ),
    .A1(net1833));
 sg13g2_o21ai_1 \register_file_i/_4830_  (.B1(\register_file_i/_1761_ ),
    .Y(\register_file_i/_1762_ ),
    .A1(net529),
    .A2(\register_file_i/_1758_ ));
 sg13g2_nand2_1 \register_file_i/_4831_  (.Y(\register_file_i/_1763_ ),
    .A(net1921),
    .B(\register_file_i/_1762_ ));
 sg13g2_mux4_1 \register_file_i/_4832_  (.S0(net2018),
    .A0(\register_file_i/rf_reg_539_ ),
    .A1(\register_file_i/rf_reg_571_ ),
    .A2(\register_file_i/rf_reg_603_ ),
    .A3(\register_file_i/rf_reg_635_ ),
    .S1(net539),
    .X(\register_file_i/_1764_ ));
 sg13g2_mux4_1 \register_file_i/_4833_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_667_ ),
    .A1(\register_file_i/rf_reg_699_ ),
    .A2(\register_file_i/rf_reg_731_ ),
    .A3(\register_file_i/rf_reg_763_ ),
    .S1(net545),
    .X(\register_file_i/_1765_ ));
 sg13g2_mux2_1 \register_file_i/_4834_  (.A0(\register_file_i/rf_reg_411_ ),
    .A1(\register_file_i/rf_reg_443_ ),
    .S(net2014),
    .X(\register_file_i/_1766_ ));
 sg13g2_mux2_1 \register_file_i/_4835_  (.A0(\register_file_i/rf_reg_475_ ),
    .A1(\register_file_i/rf_reg_507_ ),
    .S(net2014),
    .X(\register_file_i/_1767_ ));
 sg13g2_a22oi_1 \register_file_i/_4836_  (.Y(\register_file_i/_1768_ ),
    .B1(\register_file_i/_1767_ ),
    .B2(net1822),
    .A2(\register_file_i/_1766_ ),
    .A1(net1839));
 sg13g2_mux2_1 \register_file_i/_4837_  (.A0(\register_file_i/rf_reg_347_ ),
    .A1(\register_file_i/rf_reg_379_ ),
    .S(net2014),
    .X(\register_file_i/_1769_ ));
 sg13g2_mux2_1 \register_file_i/_4838_  (.A0(\register_file_i/rf_reg_283_ ),
    .A1(\register_file_i/rf_reg_315_ ),
    .S(net2014),
    .X(\register_file_i/_1770_ ));
 sg13g2_a22oi_1 \register_file_i/_4839_  (.Y(\register_file_i/_1771_ ),
    .B1(\register_file_i/_1770_ ),
    .B2(net1798),
    .A2(\register_file_i/_1769_ ),
    .A1(net1809));
 sg13g2_a21oi_2 \register_file_i/_4840_  (.B1(net1789),
    .Y(\register_file_i/_1772_ ),
    .A2(\register_file_i/_1771_ ),
    .A1(\register_file_i/_1768_ ));
 sg13g2_a221oi_1 \register_file_i/_4841_  (.B2(net1694),
    .C1(\register_file_i/_1772_ ),
    .B1(\register_file_i/_1765_ ),
    .A1(net1793),
    .Y(\register_file_i/_1773_ ),
    .A2(\register_file_i/_1764_ ));
 sg13g2_nand3_1 \register_file_i/_4842_  (.B(\register_file_i/_1763_ ),
    .C(\register_file_i/_1773_ ),
    .A(\register_file_i/_1756_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_mux2_1 \register_file_i/_4843_  (.A0(\register_file_i/rf_reg_922_ ),
    .A1(\register_file_i/rf_reg_954_ ),
    .S(net2075),
    .X(\register_file_i/_1774_ ));
 sg13g2_mux2_1 \register_file_i/_4844_  (.A0(\register_file_i/rf_reg_986_ ),
    .A1(\register_file_i/rf_reg_1018_ ),
    .S(net2075),
    .X(\register_file_i/_1775_ ));
 sg13g2_a22oi_1 \register_file_i/_4845_  (.Y(\register_file_i/_1776_ ),
    .B1(\register_file_i/_1775_ ),
    .B2(net1833),
    .A2(\register_file_i/_1774_ ),
    .A1(net1850));
 sg13g2_mux2_1 \register_file_i/_4846_  (.A0(\register_file_i/rf_reg_858_ ),
    .A1(\register_file_i/rf_reg_890_ ),
    .S(net2073),
    .X(\register_file_i/_1777_ ));
 sg13g2_mux2_1 \register_file_i/_4847_  (.A0(\register_file_i/rf_reg_794_ ),
    .A1(\register_file_i/rf_reg_826_ ),
    .S(net2073),
    .X(\register_file_i/_1778_ ));
 sg13g2_a22oi_1 \register_file_i/_4848_  (.Y(\register_file_i/_1779_ ),
    .B1(\register_file_i/_1778_ ),
    .B2(net1806),
    .A2(\register_file_i/_1777_ ),
    .A1(net1817));
 sg13g2_a21o_1 \register_file_i/_4849_  (.A2(\register_file_i/_1779_ ),
    .A1(\register_file_i/_1776_ ),
    .B1(net1926),
    .X(\register_file_i/_1780_ ));
 sg13g2_mux2_1 \register_file_i/_4850_  (.A0(\register_file_i/rf_reg_58_ ),
    .A1(\register_file_i/rf_reg_122_ ),
    .S(net535),
    .X(\register_file_i/_1781_ ));
 sg13g2_a22oi_1 \register_file_i/_4851_  (.Y(\register_file_i/_1782_ ),
    .B1(\register_file_i/_1781_ ),
    .B2(net2075),
    .A2(net1699),
    .A1(\register_file_i/rf_reg_90_ ));
 sg13g2_mux2_1 \register_file_i/_4852_  (.A0(\register_file_i/rf_reg_218_ ),
    .A1(\register_file_i/rf_reg_250_ ),
    .S(net2074),
    .X(\register_file_i/_1783_ ));
 sg13g2_mux2_1 \register_file_i/_4853_  (.A0(\register_file_i/rf_reg_154_ ),
    .A1(\register_file_i/rf_reg_186_ ),
    .S(net2074),
    .X(\register_file_i/_1784_ ));
 sg13g2_a22oi_1 \register_file_i/_4854_  (.Y(\register_file_i/_1785_ ),
    .B1(\register_file_i/_1784_ ),
    .B2(net1849),
    .A2(\register_file_i/_1783_ ),
    .A1(net1833));
 sg13g2_o21ai_1 \register_file_i/_4855_  (.B1(\register_file_i/_1785_ ),
    .Y(\register_file_i/_1786_ ),
    .A1(net529),
    .A2(\register_file_i/_1782_ ));
 sg13g2_nand2_1 \register_file_i/_4856_  (.Y(\register_file_i/_1787_ ),
    .A(net1921),
    .B(\register_file_i/_1786_ ));
 sg13g2_mux4_1 \register_file_i/_4857_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_538_ ),
    .A1(\register_file_i/rf_reg_570_ ),
    .A2(\register_file_i/rf_reg_602_ ),
    .A3(\register_file_i/rf_reg_634_ ),
    .S1(net539),
    .X(\register_file_i/_1788_ ));
 sg13g2_mux4_1 \register_file_i/_4858_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_666_ ),
    .A1(\register_file_i/rf_reg_698_ ),
    .A2(\register_file_i/rf_reg_730_ ),
    .A3(\register_file_i/rf_reg_762_ ),
    .S1(net545),
    .X(\register_file_i/_1789_ ));
 sg13g2_mux2_1 \register_file_i/_4859_  (.A0(\register_file_i/rf_reg_410_ ),
    .A1(\register_file_i/rf_reg_442_ ),
    .S(net2015),
    .X(\register_file_i/_1790_ ));
 sg13g2_mux2_1 \register_file_i/_4860_  (.A0(\register_file_i/rf_reg_474_ ),
    .A1(\register_file_i/rf_reg_506_ ),
    .S(net2015),
    .X(\register_file_i/_1791_ ));
 sg13g2_a22oi_1 \register_file_i/_4861_  (.Y(\register_file_i/_1792_ ),
    .B1(\register_file_i/_1791_ ),
    .B2(net1820),
    .A2(\register_file_i/_1790_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4862_  (.A0(\register_file_i/rf_reg_346_ ),
    .A1(\register_file_i/rf_reg_378_ ),
    .S(net2015),
    .X(\register_file_i/_1793_ ));
 sg13g2_mux2_1 \register_file_i/_4863_  (.A0(\register_file_i/rf_reg_282_ ),
    .A1(\register_file_i/rf_reg_314_ ),
    .S(net2015),
    .X(\register_file_i/_1794_ ));
 sg13g2_a22oi_1 \register_file_i/_4864_  (.Y(\register_file_i/_1795_ ),
    .B1(\register_file_i/_1794_ ),
    .B2(net1798),
    .A2(\register_file_i/_1793_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4865_  (.A1(\register_file_i/_1792_ ),
    .A2(\register_file_i/_1795_ ),
    .Y(\register_file_i/_1796_ ),
    .B1(net1789));
 sg13g2_a221oi_1 \register_file_i/_4866_  (.B2(net1694),
    .C1(\register_file_i/_1796_ ),
    .B1(\register_file_i/_1789_ ),
    .A1(net1793),
    .Y(\register_file_i/_1797_ ),
    .A2(\register_file_i/_1788_ ));
 sg13g2_nand3_1 \register_file_i/_4867_  (.B(\register_file_i/_1787_ ),
    .C(\register_file_i/_1797_ ),
    .A(\register_file_i/_1780_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_mux2_1 \register_file_i/_4868_  (.A0(\register_file_i/rf_reg_921_ ),
    .A1(\register_file_i/rf_reg_953_ ),
    .S(net2082),
    .X(\register_file_i/_1798_ ));
 sg13g2_mux2_1 \register_file_i/_4869_  (.A0(\register_file_i/rf_reg_985_ ),
    .A1(\register_file_i/rf_reg_1017_ ),
    .S(net2082),
    .X(\register_file_i/_1799_ ));
 sg13g2_a22oi_1 \register_file_i/_4870_  (.Y(\register_file_i/_1800_ ),
    .B1(\register_file_i/_1799_ ),
    .B2(net1835),
    .A2(\register_file_i/_1798_ ),
    .A1(net1853));
 sg13g2_mux2_1 \register_file_i/_4871_  (.A0(\register_file_i/rf_reg_857_ ),
    .A1(\register_file_i/rf_reg_889_ ),
    .S(net2083),
    .X(\register_file_i/_1801_ ));
 sg13g2_mux2_1 \register_file_i/_4872_  (.A0(\register_file_i/rf_reg_793_ ),
    .A1(\register_file_i/rf_reg_825_ ),
    .S(net2073),
    .X(\register_file_i/_1802_ ));
 sg13g2_a22oi_1 \register_file_i/_4873_  (.Y(\register_file_i/_1803_ ),
    .B1(\register_file_i/_1802_ ),
    .B2(net1807),
    .A2(\register_file_i/_1801_ ),
    .A1(net1818));
 sg13g2_a21o_1 \register_file_i/_4874_  (.A2(\register_file_i/_1803_ ),
    .A1(\register_file_i/_1800_ ),
    .B1(net1930),
    .X(\register_file_i/_1804_ ));
 sg13g2_mux2_1 \register_file_i/_4875_  (.A0(\register_file_i/rf_reg_57_ ),
    .A1(\register_file_i/rf_reg_121_ ),
    .S(net535),
    .X(\register_file_i/_1805_ ));
 sg13g2_a22oi_1 \register_file_i/_4876_  (.Y(\register_file_i/_1806_ ),
    .B1(\register_file_i/_1805_ ),
    .B2(net2075),
    .A2(net1700),
    .A1(\register_file_i/rf_reg_89_ ));
 sg13g2_mux2_1 \register_file_i/_4877_  (.A0(\register_file_i/rf_reg_217_ ),
    .A1(\register_file_i/rf_reg_249_ ),
    .S(net2073),
    .X(\register_file_i/_1807_ ));
 sg13g2_mux2_1 \register_file_i/_4878_  (.A0(\register_file_i/rf_reg_153_ ),
    .A1(\register_file_i/rf_reg_185_ ),
    .S(net2073),
    .X(\register_file_i/_1808_ ));
 sg13g2_a22oi_1 \register_file_i/_4879_  (.Y(\register_file_i/_1809_ ),
    .B1(\register_file_i/_1808_ ),
    .B2(net1849),
    .A2(\register_file_i/_1807_ ),
    .A1(net1833));
 sg13g2_o21ai_1 \register_file_i/_4880_  (.B1(\register_file_i/_1809_ ),
    .Y(\register_file_i/_1810_ ),
    .A1(net528),
    .A2(\register_file_i/_1806_ ));
 sg13g2_nand2_1 \register_file_i/_4881_  (.Y(\register_file_i/_1811_ ),
    .A(net1921),
    .B(\register_file_i/_1810_ ));
 sg13g2_mux4_1 \register_file_i/_4882_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_537_ ),
    .A1(\register_file_i/rf_reg_569_ ),
    .A2(\register_file_i/rf_reg_601_ ),
    .A3(\register_file_i/rf_reg_633_ ),
    .S1(net539),
    .X(\register_file_i/_1812_ ));
 sg13g2_mux4_1 \register_file_i/_4883_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_665_ ),
    .A1(\register_file_i/rf_reg_697_ ),
    .A2(\register_file_i/rf_reg_729_ ),
    .A3(\register_file_i/rf_reg_761_ ),
    .S1(net545),
    .X(\register_file_i/_1813_ ));
 sg13g2_mux2_1 \register_file_i/_4884_  (.A0(\register_file_i/rf_reg_409_ ),
    .A1(\register_file_i/rf_reg_441_ ),
    .S(net2016),
    .X(\register_file_i/_1814_ ));
 sg13g2_mux2_1 \register_file_i/_4885_  (.A0(\register_file_i/rf_reg_473_ ),
    .A1(\register_file_i/rf_reg_505_ ),
    .S(net2014),
    .X(\register_file_i/_1815_ ));
 sg13g2_a22oi_1 \register_file_i/_4886_  (.Y(\register_file_i/_1816_ ),
    .B1(\register_file_i/_1815_ ),
    .B2(net1820),
    .A2(\register_file_i/_1814_ ),
    .A1(net1837));
 sg13g2_mux2_1 \register_file_i/_4887_  (.A0(\register_file_i/rf_reg_345_ ),
    .A1(\register_file_i/rf_reg_377_ ),
    .S(net2016),
    .X(\register_file_i/_1817_ ));
 sg13g2_mux2_1 \register_file_i/_4888_  (.A0(\register_file_i/rf_reg_281_ ),
    .A1(\register_file_i/rf_reg_313_ ),
    .S(net2014),
    .X(\register_file_i/_1818_ ));
 sg13g2_a22oi_1 \register_file_i/_4889_  (.Y(\register_file_i/_1819_ ),
    .B1(\register_file_i/_1818_ ),
    .B2(net1798),
    .A2(\register_file_i/_1817_ ),
    .A1(net1809));
 sg13g2_a21oi_1 \register_file_i/_4890_  (.A1(\register_file_i/_1816_ ),
    .A2(\register_file_i/_1819_ ),
    .Y(\register_file_i/_1820_ ),
    .B1(net1787));
 sg13g2_a221oi_1 \register_file_i/_4891_  (.B2(net1694),
    .C1(\register_file_i/_1820_ ),
    .B1(\register_file_i/_1813_ ),
    .A1(net1793),
    .Y(\register_file_i/_1821_ ),
    .A2(\register_file_i/_1812_ ));
 sg13g2_nand3_1 \register_file_i/_4892_  (.B(\register_file_i/_1811_ ),
    .C(\register_file_i/_1821_ ),
    .A(\register_file_i/_1804_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_mux2_1 \register_file_i/_4893_  (.A0(\register_file_i/rf_reg_920_ ),
    .A1(\register_file_i/rf_reg_952_ ),
    .S(net2083),
    .X(\register_file_i/_1822_ ));
 sg13g2_mux2_1 \register_file_i/_4894_  (.A0(\register_file_i/rf_reg_984_ ),
    .A1(\register_file_i/rf_reg_1016_ ),
    .S(net2082),
    .X(\register_file_i/_1823_ ));
 sg13g2_a22oi_1 \register_file_i/_4895_  (.Y(\register_file_i/_1824_ ),
    .B1(\register_file_i/_1823_ ),
    .B2(net1835),
    .A2(\register_file_i/_1822_ ),
    .A1(net1853));
 sg13g2_mux2_1 \register_file_i/_4896_  (.A0(\register_file_i/rf_reg_856_ ),
    .A1(\register_file_i/rf_reg_888_ ),
    .S(net2082),
    .X(\register_file_i/_1825_ ));
 sg13g2_mux2_1 \register_file_i/_4897_  (.A0(\register_file_i/rf_reg_792_ ),
    .A1(\register_file_i/rf_reg_824_ ),
    .S(net2082),
    .X(\register_file_i/_1826_ ));
 sg13g2_a22oi_1 \register_file_i/_4898_  (.Y(\register_file_i/_1827_ ),
    .B1(\register_file_i/_1826_ ),
    .B2(net1807),
    .A2(\register_file_i/_1825_ ),
    .A1(net1818));
 sg13g2_a21o_1 \register_file_i/_4899_  (.A2(\register_file_i/_1827_ ),
    .A1(\register_file_i/_1824_ ),
    .B1(net1930),
    .X(\register_file_i/_1828_ ));
 sg13g2_mux2_1 \register_file_i/_4900_  (.A0(\register_file_i/rf_reg_56_ ),
    .A1(\register_file_i/rf_reg_120_ ),
    .S(net534),
    .X(\register_file_i/_1829_ ));
 sg13g2_a22oi_1 \register_file_i/_4901_  (.Y(\register_file_i/_1830_ ),
    .B1(\register_file_i/_1829_ ),
    .B2(net2075),
    .A2(net1703),
    .A1(\register_file_i/rf_reg_88_ ));
 sg13g2_mux2_1 \register_file_i/_4902_  (.A0(\register_file_i/rf_reg_216_ ),
    .A1(\register_file_i/rf_reg_248_ ),
    .S(net2082),
    .X(\register_file_i/_1831_ ));
 sg13g2_mux2_1 \register_file_i/_4903_  (.A0(\register_file_i/rf_reg_152_ ),
    .A1(\register_file_i/rf_reg_184_ ),
    .S(net2082),
    .X(\register_file_i/_1832_ ));
 sg13g2_a22oi_1 \register_file_i/_4904_  (.Y(\register_file_i/_1833_ ),
    .B1(\register_file_i/_1832_ ),
    .B2(net1853),
    .A2(\register_file_i/_1831_ ),
    .A1(net1835));
 sg13g2_o21ai_1 \register_file_i/_4905_  (.B1(\register_file_i/_1833_ ),
    .Y(\register_file_i/_1834_ ),
    .A1(net528),
    .A2(\register_file_i/_1830_ ));
 sg13g2_nand2_1 \register_file_i/_4906_  (.Y(\register_file_i/_1835_ ),
    .A(net1924),
    .B(\register_file_i/_1834_ ));
 sg13g2_mux4_1 \register_file_i/_4907_  (.S0(net2017),
    .A0(\register_file_i/rf_reg_536_ ),
    .A1(\register_file_i/rf_reg_568_ ),
    .A2(\register_file_i/rf_reg_600_ ),
    .A3(\register_file_i/rf_reg_632_ ),
    .S1(net539),
    .X(\register_file_i/_1836_ ));
 sg13g2_mux4_1 \register_file_i/_4908_  (.S0(net2034),
    .A0(\register_file_i/rf_reg_664_ ),
    .A1(\register_file_i/rf_reg_696_ ),
    .A2(\register_file_i/rf_reg_728_ ),
    .A3(\register_file_i/rf_reg_760_ ),
    .S1(net544),
    .X(\register_file_i/_1837_ ));
 sg13g2_mux2_1 \register_file_i/_4909_  (.A0(\register_file_i/rf_reg_408_ ),
    .A1(\register_file_i/rf_reg_440_ ),
    .S(net2034),
    .X(\register_file_i/_1838_ ));
 sg13g2_mux2_1 \register_file_i/_4910_  (.A0(\register_file_i/rf_reg_472_ ),
    .A1(\register_file_i/rf_reg_504_ ),
    .S(net2034),
    .X(\register_file_i/_1839_ ));
 sg13g2_a22oi_1 \register_file_i/_4911_  (.Y(\register_file_i/_1840_ ),
    .B1(\register_file_i/_1839_ ),
    .B2(net1823),
    .A2(\register_file_i/_1838_ ),
    .A1(net1840));
 sg13g2_mux2_1 \register_file_i/_4912_  (.A0(\register_file_i/rf_reg_344_ ),
    .A1(\register_file_i/rf_reg_376_ ),
    .S(net2034),
    .X(\register_file_i/_1841_ ));
 sg13g2_mux2_1 \register_file_i/_4913_  (.A0(\register_file_i/rf_reg_280_ ),
    .A1(\register_file_i/rf_reg_312_ ),
    .S(net2034),
    .X(\register_file_i/_1842_ ));
 sg13g2_a22oi_1 \register_file_i/_4914_  (.Y(\register_file_i/_1843_ ),
    .B1(\register_file_i/_1842_ ),
    .B2(net1801),
    .A2(\register_file_i/_1841_ ),
    .A1(net1812));
 sg13g2_a21oi_1 \register_file_i/_4915_  (.A1(\register_file_i/_1840_ ),
    .A2(\register_file_i/_1843_ ),
    .Y(\register_file_i/_1844_ ),
    .B1(net1790));
 sg13g2_a221oi_1 \register_file_i/_4916_  (.B2(net1696),
    .C1(\register_file_i/_1844_ ),
    .B1(\register_file_i/_1837_ ),
    .A1(net1795),
    .Y(\register_file_i/_1845_ ),
    .A2(\register_file_i/_1836_ ));
 sg13g2_nand3_1 \register_file_i/_4917_  (.B(\register_file_i/_1835_ ),
    .C(\register_file_i/_1845_ ),
    .A(\register_file_i/_1828_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_24_ ));
 sg13g2_mux2_1 \register_file_i/_4918_  (.A0(\register_file_i/rf_reg_919_ ),
    .A1(\register_file_i/rf_reg_951_ ),
    .S(net2027),
    .X(\register_file_i/_1846_ ));
 sg13g2_mux2_1 \register_file_i/_4919_  (.A0(\register_file_i/rf_reg_983_ ),
    .A1(\register_file_i/rf_reg_1015_ ),
    .S(net2027),
    .X(\register_file_i/_1847_ ));
 sg13g2_a22oi_1 \register_file_i/_4920_  (.Y(\register_file_i/_1848_ ),
    .B1(\register_file_i/_1847_ ),
    .B2(net1821),
    .A2(\register_file_i/_1846_ ),
    .A1(net1838));
 sg13g2_mux2_1 \register_file_i/_4921_  (.A0(\register_file_i/rf_reg_855_ ),
    .A1(\register_file_i/rf_reg_887_ ),
    .S(net2029),
    .X(\register_file_i/_1849_ ));
 sg13g2_mux2_1 \register_file_i/_4922_  (.A0(\register_file_i/rf_reg_791_ ),
    .A1(\register_file_i/rf_reg_823_ ),
    .S(net2027),
    .X(\register_file_i/_1850_ ));
 sg13g2_a22oi_1 \register_file_i/_4923_  (.Y(\register_file_i/_1851_ ),
    .B1(\register_file_i/_1850_ ),
    .B2(net1804),
    .A2(\register_file_i/_1849_ ),
    .A1(net1815));
 sg13g2_a21o_1 \register_file_i/_4924_  (.A2(\register_file_i/_1851_ ),
    .A1(\register_file_i/_1848_ ),
    .B1(net1928),
    .X(\register_file_i/_1852_ ));
 sg13g2_mux2_1 \register_file_i/_4925_  (.A0(\register_file_i/rf_reg_55_ ),
    .A1(\register_file_i/rf_reg_119_ ),
    .S(net534),
    .X(\register_file_i/_1853_ ));
 sg13g2_a22oi_1 \register_file_i/_4926_  (.Y(\register_file_i/_1854_ ),
    .B1(\register_file_i/_1853_ ),
    .B2(net2064),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_87_ ));
 sg13g2_mux2_1 \register_file_i/_4927_  (.A0(\register_file_i/rf_reg_215_ ),
    .A1(\register_file_i/rf_reg_247_ ),
    .S(net2063),
    .X(\register_file_i/_1855_ ));
 sg13g2_mux2_1 \register_file_i/_4928_  (.A0(\register_file_i/rf_reg_151_ ),
    .A1(\register_file_i/rf_reg_183_ ),
    .S(net2063),
    .X(\register_file_i/_1856_ ));
 sg13g2_a22oi_1 \register_file_i/_4929_  (.Y(\register_file_i/_1857_ ),
    .B1(\register_file_i/_1856_ ),
    .B2(net1847),
    .A2(\register_file_i/_1855_ ),
    .A1(net1829));
 sg13g2_o21ai_1 \register_file_i/_4930_  (.B1(\register_file_i/_1857_ ),
    .Y(\register_file_i/_1858_ ),
    .A1(net528),
    .A2(\register_file_i/_1854_ ));
 sg13g2_nand2_1 \register_file_i/_4931_  (.Y(\register_file_i/_1859_ ),
    .A(net1920),
    .B(\register_file_i/_1858_ ));
 sg13g2_mux4_1 \register_file_i/_4932_  (.S0(net2042),
    .A0(\register_file_i/rf_reg_535_ ),
    .A1(\register_file_i/rf_reg_567_ ),
    .A2(\register_file_i/rf_reg_599_ ),
    .A3(\register_file_i/rf_reg_631_ ),
    .S1(net538),
    .X(\register_file_i/_1860_ ));
 sg13g2_mux4_1 \register_file_i/_4933_  (.S0(net2042),
    .A0(\register_file_i/rf_reg_663_ ),
    .A1(\register_file_i/rf_reg_695_ ),
    .A2(\register_file_i/rf_reg_727_ ),
    .A3(\register_file_i/rf_reg_759_ ),
    .S1(net544),
    .X(\register_file_i/_1861_ ));
 sg13g2_mux2_1 \register_file_i/_4934_  (.A0(\register_file_i/rf_reg_407_ ),
    .A1(\register_file_i/rf_reg_439_ ),
    .S(net2042),
    .X(\register_file_i/_1862_ ));
 sg13g2_mux2_1 \register_file_i/_4935_  (.A0(\register_file_i/rf_reg_471_ ),
    .A1(\register_file_i/rf_reg_503_ ),
    .S(net2042),
    .X(\register_file_i/_1863_ ));
 sg13g2_a22oi_1 \register_file_i/_4936_  (.Y(\register_file_i/_1864_ ),
    .B1(\register_file_i/_1863_ ),
    .B2(net1825),
    .A2(\register_file_i/_1862_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4937_  (.A0(\register_file_i/rf_reg_343_ ),
    .A1(\register_file_i/rf_reg_375_ ),
    .S(net2042),
    .X(\register_file_i/_1865_ ));
 sg13g2_mux2_1 \register_file_i/_4938_  (.A0(\register_file_i/rf_reg_279_ ),
    .A1(\register_file_i/rf_reg_311_ ),
    .S(net2042),
    .X(\register_file_i/_1866_ ));
 sg13g2_a22oi_1 \register_file_i/_4939_  (.Y(\register_file_i/_1867_ ),
    .B1(\register_file_i/_1866_ ),
    .B2(net1801),
    .A2(\register_file_i/_1865_ ),
    .A1(net1812));
 sg13g2_a21oi_1 \register_file_i/_4940_  (.A1(\register_file_i/_1864_ ),
    .A2(\register_file_i/_1867_ ),
    .Y(\register_file_i/_1868_ ),
    .B1(net1791));
 sg13g2_a221oi_1 \register_file_i/_4941_  (.B2(net1696),
    .C1(\register_file_i/_1868_ ),
    .B1(\register_file_i/_1861_ ),
    .A1(net1795),
    .Y(\register_file_i/_1869_ ),
    .A2(\register_file_i/_1860_ ));
 sg13g2_nand3_1 \register_file_i/_4942_  (.B(\register_file_i/_1859_ ),
    .C(\register_file_i/_1869_ ),
    .A(\register_file_i/_1852_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_23_ ));
 sg13g2_mux2_1 \register_file_i/_4943_  (.A0(\register_file_i/rf_reg_918_ ),
    .A1(\register_file_i/rf_reg_950_ ),
    .S(net2082),
    .X(\register_file_i/_1870_ ));
 sg13g2_mux2_1 \register_file_i/_4944_  (.A0(\register_file_i/rf_reg_982_ ),
    .A1(\register_file_i/rf_reg_1014_ ),
    .S(net2083),
    .X(\register_file_i/_1871_ ));
 sg13g2_a22oi_1 \register_file_i/_4945_  (.Y(\register_file_i/_1872_ ),
    .B1(\register_file_i/_1871_ ),
    .B2(net1835),
    .A2(\register_file_i/_1870_ ),
    .A1(net1853));
 sg13g2_mux2_1 \register_file_i/_4946_  (.A0(\register_file_i/rf_reg_854_ ),
    .A1(\register_file_i/rf_reg_886_ ),
    .S(net2078),
    .X(\register_file_i/_1873_ ));
 sg13g2_mux2_1 \register_file_i/_4947_  (.A0(\register_file_i/rf_reg_790_ ),
    .A1(\register_file_i/rf_reg_822_ ),
    .S(net2078),
    .X(\register_file_i/_1874_ ));
 sg13g2_a22oi_1 \register_file_i/_4948_  (.Y(\register_file_i/_1875_ ),
    .B1(\register_file_i/_1874_ ),
    .B2(net1807),
    .A2(\register_file_i/_1873_ ),
    .A1(net1818));
 sg13g2_a21o_1 \register_file_i/_4949_  (.A2(\register_file_i/_1875_ ),
    .A1(\register_file_i/_1872_ ),
    .B1(net1930),
    .X(\register_file_i/_1876_ ));
 sg13g2_mux2_1 \register_file_i/_4950_  (.A0(\register_file_i/rf_reg_54_ ),
    .A1(\register_file_i/rf_reg_118_ ),
    .S(net532),
    .X(\register_file_i/_1877_ ));
 sg13g2_a22oi_1 \register_file_i/_4951_  (.Y(\register_file_i/_1878_ ),
    .B1(\register_file_i/_1877_ ),
    .B2(net2078),
    .A2(net1701),
    .A1(\register_file_i/rf_reg_86_ ));
 sg13g2_mux2_1 \register_file_i/_4952_  (.A0(\register_file_i/rf_reg_214_ ),
    .A1(\register_file_i/rf_reg_246_ ),
    .S(net2078),
    .X(\register_file_i/_1879_ ));
 sg13g2_mux2_1 \register_file_i/_4953_  (.A0(\register_file_i/rf_reg_150_ ),
    .A1(\register_file_i/rf_reg_182_ ),
    .S(net2078),
    .X(\register_file_i/_1880_ ));
 sg13g2_a22oi_1 \register_file_i/_4954_  (.Y(\register_file_i/_1881_ ),
    .B1(\register_file_i/_1880_ ),
    .B2(net1851),
    .A2(\register_file_i/_1879_ ),
    .A1(net1834));
 sg13g2_o21ai_1 \register_file_i/_4955_  (.B1(\register_file_i/_1881_ ),
    .Y(\register_file_i/_1882_ ),
    .A1(net528),
    .A2(\register_file_i/_1878_ ));
 sg13g2_nand2_1 \register_file_i/_4956_  (.Y(\register_file_i/_1883_ ),
    .A(net1924),
    .B(\register_file_i/_1882_ ));
 sg13g2_mux4_1 \register_file_i/_4957_  (.S0(net2048),
    .A0(\register_file_i/rf_reg_534_ ),
    .A1(\register_file_i/rf_reg_566_ ),
    .A2(\register_file_i/rf_reg_598_ ),
    .A3(\register_file_i/rf_reg_630_ ),
    .S1(net538),
    .X(\register_file_i/_1884_ ));
 sg13g2_mux4_1 \register_file_i/_4958_  (.S0(net2048),
    .A0(\register_file_i/rf_reg_662_ ),
    .A1(\register_file_i/rf_reg_694_ ),
    .A2(\register_file_i/rf_reg_726_ ),
    .A3(\register_file_i/rf_reg_758_ ),
    .S1(net538),
    .X(\register_file_i/_1885_ ));
 sg13g2_mux2_1 \register_file_i/_4959_  (.A0(\register_file_i/rf_reg_406_ ),
    .A1(\register_file_i/rf_reg_438_ ),
    .S(net2047),
    .X(\register_file_i/_1886_ ));
 sg13g2_mux2_1 \register_file_i/_4960_  (.A0(\register_file_i/rf_reg_470_ ),
    .A1(\register_file_i/rf_reg_502_ ),
    .S(net2047),
    .X(\register_file_i/_1887_ ));
 sg13g2_a22oi_1 \register_file_i/_4961_  (.Y(\register_file_i/_1888_ ),
    .B1(\register_file_i/_1887_ ),
    .B2(net1825),
    .A2(\register_file_i/_1886_ ),
    .A1(net1842));
 sg13g2_mux2_1 \register_file_i/_4962_  (.A0(\register_file_i/rf_reg_342_ ),
    .A1(\register_file_i/rf_reg_374_ ),
    .S(net2047),
    .X(\register_file_i/_1889_ ));
 sg13g2_mux2_1 \register_file_i/_4963_  (.A0(\register_file_i/rf_reg_278_ ),
    .A1(\register_file_i/rf_reg_310_ ),
    .S(net2047),
    .X(\register_file_i/_1890_ ));
 sg13g2_a22oi_1 \register_file_i/_4964_  (.Y(\register_file_i/_1891_ ),
    .B1(\register_file_i/_1890_ ),
    .B2(net1802),
    .A2(\register_file_i/_1889_ ),
    .A1(net1812));
 sg13g2_a21oi_1 \register_file_i/_4965_  (.A1(\register_file_i/_1888_ ),
    .A2(\register_file_i/_1891_ ),
    .Y(\register_file_i/_1892_ ),
    .B1(net1791));
 sg13g2_a221oi_1 \register_file_i/_4966_  (.B2(net1698),
    .C1(\register_file_i/_1892_ ),
    .B1(\register_file_i/_1885_ ),
    .A1(net1797),
    .Y(\register_file_i/_1893_ ),
    .A2(\register_file_i/_1884_ ));
 sg13g2_nand3_1 \register_file_i/_4967_  (.B(\register_file_i/_1883_ ),
    .C(\register_file_i/_1893_ ),
    .A(\register_file_i/_1876_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_22_ ));
 sg13g2_buf_2 fanout319 (.A(net323),
    .X(net319));
 sg13g2_buf_1 fanout318 (.A(_04077_),
    .X(net318));
 sg13g2_nor2b_2 \register_file_i/_4970_  (.A(net454),
    .B_N(net443),
    .Y(\register_file_i/_1896_ ));
 sg13g2_buf_2 fanout317 (.A(_04077_),
    .X(net317));
 sg13g2_buf_2 fanout316 (.A(net318),
    .X(net316));
 sg13g2_buf_2 fanout315 (.A(net318),
    .X(net315));
 sg13g2_buf_2 fanout314 (.A(net318),
    .X(net314));
 sg13g2_buf_4 fanout313 (.X(net313),
    .A(net318));
 sg13g2_mux2_1 \register_file_i/_4976_  (.A0(\register_file_i/rf_reg_927_ ),
    .A1(\register_file_i/rf_reg_959_ ),
    .S(net466),
    .X(\register_file_i/_1902_ ));
 sg13g2_buf_1 fanout312 (.A(net317),
    .X(net312));
 sg13g2_mux2_1 \register_file_i/_4978_  (.A0(\register_file_i/rf_reg_991_ ),
    .A1(\register_file_i/rf_reg_1023_ ),
    .S(net467),
    .X(\register_file_i/_1904_ ));
 sg13g2_and2_1 \register_file_i/_4979_  (.A(net442),
    .B(net449),
    .X(\register_file_i/_1905_ ));
 sg13g2_buf_2 fanout311 (.A(net317),
    .X(net311));
 sg13g2_buf_2 fanout310 (.A(net317),
    .X(net310));
 sg13g2_buf_2 fanout309 (.A(net317),
    .X(net309));
 sg13g2_a22oi_1 \register_file_i/_4983_  (.Y(\register_file_i/_1909_ ),
    .B1(\register_file_i/_1904_ ),
    .B2(net1758),
    .A2(\register_file_i/_1902_ ),
    .A1(net1775));
 sg13g2_nor2b_1 \register_file_i/_4984_  (.A(\id_stage_i.controller_i.instr_i_22_ ),
    .B_N(net449),
    .Y(\register_file_i/_1910_ ));
 sg13g2_buf_2 fanout308 (.A(net317),
    .X(net308));
 sg13g2_buf_2 fanout307 (.A(net317),
    .X(net307));
 sg13g2_mux2_1 \register_file_i/_4987_  (.A0(\register_file_i/rf_reg_863_ ),
    .A1(\register_file_i/rf_reg_895_ ),
    .S(net468),
    .X(\register_file_i/_1913_ ));
 sg13g2_buf_2 fanout306 (.A(net317),
    .X(net306));
 sg13g2_mux2_1 \register_file_i/_4989_  (.A0(\register_file_i/rf_reg_799_ ),
    .A1(\register_file_i/rf_reg_831_ ),
    .S(net469),
    .X(\register_file_i/_1915_ ));
 sg13g2_nor2_1 \register_file_i/_4990_  (.A(net443),
    .B(net448),
    .Y(\register_file_i/_1916_ ));
 sg13g2_buf_2 fanout305 (.A(net317),
    .X(net305));
 sg13g2_buf_4 fanout304 (.X(net304),
    .A(net318));
 sg13g2_a22oi_1 \register_file_i/_4993_  (.Y(\register_file_i/_1919_ ),
    .B1(\register_file_i/_1915_ ),
    .B2(net1739),
    .A2(\register_file_i/_1913_ ),
    .A1(net1750));
 sg13g2_nand2_2 \register_file_i/_4994_  (.Y(\register_file_i/_1920_ ),
    .A(\id_stage_i.controller_i.instr_i_24_ ),
    .B(net2007));
 sg13g2_buf_1 fanout303 (.A(_04061_),
    .X(net303));
 sg13g2_a21o_1 \register_file_i/_4996_  (.A2(\register_file_i/_1919_ ),
    .A1(\register_file_i/_1909_ ),
    .B1(net1917),
    .X(\register_file_i/_1922_ ));
 sg13g2_nor2_1 \register_file_i/_4997_  (.A(\id_stage_i.controller_i.instr_i_24_ ),
    .B(net2007),
    .Y(\register_file_i/_1923_ ));
 sg13g2_buf_1 fanout302 (.A(net303),
    .X(net302));
 sg13g2_buf_2 fanout301 (.A(net303),
    .X(net301));
 sg13g2_buf_2 fanout300 (.A(_04143_),
    .X(net300));
 sg13g2_buf_2 fanout299 (.A(net300),
    .X(net299));
 sg13g2_buf_2 fanout298 (.A(net300),
    .X(net298));
 sg13g2_mux2_1 \register_file_i/_5003_  (.A0(\register_file_i/rf_reg_63_ ),
    .A1(\register_file_i/rf_reg_127_ ),
    .S(net449),
    .X(\register_file_i/_1929_ ));
 sg13g2_buf_2 fanout297 (.A(net300),
    .X(net297));
 sg13g2_nor2b_1 \register_file_i/_5005_  (.A(net514),
    .B_N(net448),
    .Y(\register_file_i/_1931_ ));
 sg13g2_buf_2 fanout296 (.A(_07682_),
    .X(net296));
 sg13g2_a22oi_1 \register_file_i/_5007_  (.Y(\register_file_i/_1933_ ),
    .B1(net1691),
    .B2(\register_file_i/rf_reg_95_ ),
    .A2(\register_file_i/_1929_ ),
    .A1(net464));
 sg13g2_buf_2 fanout295 (.A(\cs_registers_i/_1404_ ),
    .X(net295));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(\cs_registers_i/_1404_ ));
 sg13g2_mux2_1 \register_file_i/_5010_  (.A0(\register_file_i/rf_reg_223_ ),
    .A1(\register_file_i/rf_reg_255_ ),
    .S(net472),
    .X(\register_file_i/_1936_ ));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(net294));
 sg13g2_mux2_1 \register_file_i/_5012_  (.A0(\register_file_i/rf_reg_159_ ),
    .A1(\register_file_i/rf_reg_191_ ),
    .S(net473),
    .X(\register_file_i/_1938_ ));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net294));
 sg13g2_a22oi_1 \register_file_i/_5014_  (.Y(\register_file_i/_1940_ ),
    .B1(\register_file_i/_1938_ ),
    .B2(net1784),
    .A2(\register_file_i/_1936_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5015_  (.B1(\register_file_i/_1940_ ),
    .Y(\register_file_i/_1941_ ),
    .A1(net444),
    .A2(\register_file_i/_1933_ ));
 sg13g2_nand2_1 \register_file_i/_5016_  (.Y(\register_file_i/_1942_ ),
    .A(net1910),
    .B(\register_file_i/_1941_ ));
 sg13g2_inv_1 \register_file_i/_5017_  (.Y(\register_file_i/_1943_ ),
    .A(\id_stage_i.controller_i.instr_i_24_ ));
 sg13g2_nor3_2 \register_file_i/_5018_  (.A(\register_file_i/_1943_ ),
    .B(net2007),
    .C(\id_stage_i.controller_i.instr_i_22_ ),
    .Y(\register_file_i/_1944_ ));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net294));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(net294));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_31_ ));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_31_ ));
 sg13g2_mux4_1 \register_file_i/_5023_  (.S0(net474),
    .A0(\register_file_i/rf_reg_543_ ),
    .A1(\register_file_i/rf_reg_575_ ),
    .A2(\register_file_i/rf_reg_607_ ),
    .A3(\register_file_i/rf_reg_639_ ),
    .S1(net455),
    .X(\register_file_i/_1949_ ));
 sg13g2_inv_1 \register_file_i/_5024_  (.Y(\register_file_i/_1950_ ),
    .A(net442));
 sg13g2_nor3_2 \register_file_i/_5025_  (.A(\register_file_i/_1943_ ),
    .B(net2007),
    .C(\register_file_i/_1950_ ),
    .Y(\register_file_i/_1951_ ));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ));
 sg13g2_mux4_1 \register_file_i/_5028_  (.S0(net475),
    .A0(\register_file_i/rf_reg_671_ ),
    .A1(\register_file_i/rf_reg_703_ ),
    .A2(\register_file_i/rf_reg_735_ ),
    .A3(\register_file_i/rf_reg_767_ ),
    .S1(net455),
    .X(\register_file_i/_1954_ ));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ));
 sg13g2_mux2_1 \register_file_i/_5031_  (.A0(\register_file_i/rf_reg_479_ ),
    .A1(\register_file_i/rf_reg_511_ ),
    .S(net477),
    .X(\register_file_i/_1957_ ));
 sg13g2_buf_2 fanout283 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_7_ ),
    .X(net283));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_7_ ));
 sg13g2_mux2_1 \register_file_i/_5034_  (.A0(\register_file_i/rf_reg_415_ ),
    .A1(\register_file_i/rf_reg_447_ ),
    .S(net478),
    .X(\register_file_i/_1960_ ));
 sg13g2_a22oi_1 \register_file_i/_5035_  (.Y(\register_file_i/_1961_ ),
    .B1(net1772),
    .B2(\register_file_i/_1960_ ),
    .A2(\register_file_i/_1957_ ),
    .A1(net1755));
 sg13g2_buf_2 fanout281 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_7_ ),
    .X(net281));
 sg13g2_mux2_1 \register_file_i/_5037_  (.A0(\register_file_i/rf_reg_351_ ),
    .A1(\register_file_i/rf_reg_383_ ),
    .S(net479),
    .X(\register_file_i/_1963_ ));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_0_ ));
 sg13g2_mux2_1 \register_file_i/_5039_  (.A0(\register_file_i/rf_reg_287_ ),
    .A1(\register_file_i/rf_reg_319_ ),
    .S(net480),
    .X(\register_file_i/_1965_ ));
 sg13g2_buf_2 fanout279 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_0_ ),
    .X(net279));
 sg13g2_a22oi_1 \register_file_i/_5041_  (.Y(\register_file_i/_1967_ ),
    .B1(\register_file_i/_1965_ ),
    .B2(net1735),
    .A2(net1743),
    .A1(\register_file_i/_1963_ ));
 sg13g2_nand2_2 \register_file_i/_5042_  (.Y(\register_file_i/_1968_ ),
    .A(\register_file_i/_1943_ ),
    .B(net2007));
 sg13g2_buf_2 fanout278 (.A(_04170_),
    .X(net278));
 sg13g2_a21oi_1 \register_file_i/_5044_  (.A1(\register_file_i/_1961_ ),
    .A2(\register_file_i/_1967_ ),
    .Y(\register_file_i/_1970_ ),
    .B1(net1723));
 sg13g2_a221oi_1 \register_file_i/_5045_  (.B2(\register_file_i/_1954_ ),
    .C1(\register_file_i/_1970_ ),
    .B1(net1686),
    .A1(net1728),
    .Y(\register_file_i/_1971_ ),
    .A2(\register_file_i/_1949_ ));
 sg13g2_nand3_1 \register_file_i/_5046_  (.B(\register_file_i/_1942_ ),
    .C(\register_file_i/_1971_ ),
    .A(\register_file_i/_1922_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_31_ ));
 sg13g2_mux2_1 \register_file_i/_5047_  (.A0(\register_file_i/rf_reg_926_ ),
    .A1(\register_file_i/rf_reg_958_ ),
    .S(net465),
    .X(\register_file_i/_1972_ ));
 sg13g2_mux2_1 \register_file_i/_5048_  (.A0(\register_file_i/rf_reg_990_ ),
    .A1(\register_file_i/rf_reg_1022_ ),
    .S(net467),
    .X(\register_file_i/_1973_ ));
 sg13g2_a22oi_1 \register_file_i/_5049_  (.Y(\register_file_i/_1974_ ),
    .B1(\register_file_i/_1973_ ),
    .B2(net1758),
    .A2(\register_file_i/_1972_ ),
    .A1(net1775));
 sg13g2_buf_2 fanout277 (.A(net278),
    .X(net277));
 sg13g2_mux2_1 \register_file_i/_5051_  (.A0(\register_file_i/rf_reg_862_ ),
    .A1(\register_file_i/rf_reg_894_ ),
    .S(net482),
    .X(\register_file_i/_1976_ ));
 sg13g2_mux2_1 \register_file_i/_5052_  (.A0(\register_file_i/rf_reg_798_ ),
    .A1(\register_file_i/rf_reg_830_ ),
    .S(net469),
    .X(\register_file_i/_1977_ ));
 sg13g2_a22oi_1 \register_file_i/_5053_  (.Y(\register_file_i/_1978_ ),
    .B1(\register_file_i/_1977_ ),
    .B2(net1734),
    .A2(\register_file_i/_1976_ ),
    .A1(net1745));
 sg13g2_a21o_1 \register_file_i/_5054_  (.A2(\register_file_i/_1978_ ),
    .A1(\register_file_i/_1974_ ),
    .B1(net1917),
    .X(\register_file_i/_1979_ ));
 sg13g2_mux2_1 \register_file_i/_5055_  (.A0(\register_file_i/rf_reg_62_ ),
    .A1(\register_file_i/rf_reg_126_ ),
    .S(net450),
    .X(\register_file_i/_1980_ ));
 sg13g2_buf_4 fanout276 (.X(net276),
    .A(net278));
 sg13g2_a22oi_1 \register_file_i/_5057_  (.Y(\register_file_i/_1982_ ),
    .B1(\register_file_i/_1980_ ),
    .B2(net515),
    .A2(net1691),
    .A1(\register_file_i/rf_reg_94_ ));
 sg13g2_mux2_1 \register_file_i/_5058_  (.A0(\register_file_i/rf_reg_222_ ),
    .A1(\register_file_i/rf_reg_254_ ),
    .S(net472),
    .X(\register_file_i/_1983_ ));
 sg13g2_mux2_1 \register_file_i/_5059_  (.A0(\register_file_i/rf_reg_158_ ),
    .A1(\register_file_i/rf_reg_190_ ),
    .S(net473),
    .X(\register_file_i/_1984_ ));
 sg13g2_a22oi_1 \register_file_i/_5060_  (.Y(\register_file_i/_1985_ ),
    .B1(\register_file_i/_1984_ ),
    .B2(net1784),
    .A2(\register_file_i/_1983_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5061_  (.B1(\register_file_i/_1985_ ),
    .Y(\register_file_i/_1986_ ),
    .A1(net444),
    .A2(\register_file_i/_1982_ ));
 sg13g2_nand2_1 \register_file_i/_5062_  (.Y(\register_file_i/_1987_ ),
    .A(net1910),
    .B(\register_file_i/_1986_ ));
 sg13g2_mux4_1 \register_file_i/_5063_  (.S0(net474),
    .A0(\register_file_i/rf_reg_542_ ),
    .A1(\register_file_i/rf_reg_574_ ),
    .A2(\register_file_i/rf_reg_606_ ),
    .A3(\register_file_i/rf_reg_638_ ),
    .S1(net455),
    .X(\register_file_i/_1988_ ));
 sg13g2_buf_2 fanout275 (.A(net278),
    .X(net275));
 sg13g2_buf_2 fanout274 (.A(_04218_),
    .X(net274));
 sg13g2_mux4_1 \register_file_i/_5066_  (.S0(net471),
    .A0(\register_file_i/rf_reg_670_ ),
    .A1(\register_file_i/rf_reg_702_ ),
    .A2(\register_file_i/rf_reg_734_ ),
    .A3(\register_file_i/rf_reg_766_ ),
    .S1(net457),
    .X(\register_file_i/_1991_ ));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_mux2_1 \register_file_i/_5068_  (.A0(\register_file_i/rf_reg_414_ ),
    .A1(\register_file_i/rf_reg_446_ ),
    .S(net483),
    .X(\register_file_i/_1993_ ));
 sg13g2_mux2_1 \register_file_i/_5069_  (.A0(\register_file_i/rf_reg_478_ ),
    .A1(\register_file_i/rf_reg_510_ ),
    .S(net478),
    .X(\register_file_i/_1994_ ));
 sg13g2_buf_2 fanout272 (.A(net274),
    .X(net272));
 sg13g2_a22oi_1 \register_file_i/_5071_  (.Y(\register_file_i/_1996_ ),
    .B1(\register_file_i/_1994_ ),
    .B2(net1756),
    .A2(\register_file_i/_1993_ ),
    .A1(net1772));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(_04306_));
 sg13g2_mux2_1 \register_file_i/_5073_  (.A0(\register_file_i/rf_reg_350_ ),
    .A1(\register_file_i/rf_reg_382_ ),
    .S(net479),
    .X(\register_file_i/_1998_ ));
 sg13g2_mux2_1 \register_file_i/_5074_  (.A0(\register_file_i/rf_reg_286_ ),
    .A1(\register_file_i/rf_reg_318_ ),
    .S(net480),
    .X(\register_file_i/_1999_ ));
 sg13g2_a22oi_1 \register_file_i/_5075_  (.Y(\register_file_i/_2000_ ),
    .B1(\register_file_i/_1999_ ),
    .B2(net1734),
    .A2(\register_file_i/_1998_ ),
    .A1(net1745));
 sg13g2_a21oi_1 \register_file_i/_5076_  (.A1(\register_file_i/_1996_ ),
    .A2(\register_file_i/_2000_ ),
    .Y(\register_file_i/_2001_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5077_  (.B2(net1686),
    .C1(\register_file_i/_2001_ ),
    .B1(\register_file_i/_1991_ ),
    .A1(net1728),
    .Y(\register_file_i/_2002_ ),
    .A2(\register_file_i/_1988_ ));
 sg13g2_nand3_1 \register_file_i/_5078_  (.B(\register_file_i/_1987_ ),
    .C(\register_file_i/_2002_ ),
    .A(\register_file_i/_1979_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_30_ ));
 sg13g2_mux2_1 \register_file_i/_5079_  (.A0(\register_file_i/rf_reg_917_ ),
    .A1(\register_file_i/rf_reg_949_ ),
    .S(net465),
    .X(\register_file_i/_2003_ ));
 sg13g2_mux2_1 \register_file_i/_5080_  (.A0(\register_file_i/rf_reg_981_ ),
    .A1(\register_file_i/rf_reg_1013_ ),
    .S(net467),
    .X(\register_file_i/_2004_ ));
 sg13g2_a22oi_1 \register_file_i/_5081_  (.Y(\register_file_i/_2005_ ),
    .B1(\register_file_i/_2004_ ),
    .B2(net1767),
    .A2(\register_file_i/_2003_ ),
    .A1(net1785));
 sg13g2_mux2_1 \register_file_i/_5082_  (.A0(\register_file_i/rf_reg_853_ ),
    .A1(\register_file_i/rf_reg_885_ ),
    .S(net481),
    .X(\register_file_i/_2006_ ));
 sg13g2_mux2_1 \register_file_i/_5083_  (.A0(\register_file_i/rf_reg_789_ ),
    .A1(\register_file_i/rf_reg_821_ ),
    .S(net469),
    .X(\register_file_i/_2007_ ));
 sg13g2_a22oi_1 \register_file_i/_5084_  (.Y(\register_file_i/_2008_ ),
    .B1(\register_file_i/_2007_ ),
    .B2(net1739),
    .A2(\register_file_i/_2006_ ),
    .A1(net1750));
 sg13g2_a21o_1 \register_file_i/_5085_  (.A2(\register_file_i/_2008_ ),
    .A1(\register_file_i/_2005_ ),
    .B1(net1917),
    .X(\register_file_i/_2009_ ));
 sg13g2_mux2_1 \register_file_i/_5086_  (.A0(\register_file_i/rf_reg_53_ ),
    .A1(\register_file_i/rf_reg_117_ ),
    .S(net450),
    .X(\register_file_i/_2010_ ));
 sg13g2_a22oi_1 \register_file_i/_5087_  (.Y(\register_file_i/_2011_ ),
    .B1(\register_file_i/_2010_ ),
    .B2(net515),
    .A2(net1691),
    .A1(\register_file_i/rf_reg_85_ ));
 sg13g2_mux2_1 \register_file_i/_5088_  (.A0(\register_file_i/rf_reg_213_ ),
    .A1(\register_file_i/rf_reg_245_ ),
    .S(net472),
    .X(\register_file_i/_2012_ ));
 sg13g2_mux2_1 \register_file_i/_5089_  (.A0(\register_file_i/rf_reg_149_ ),
    .A1(\register_file_i/rf_reg_181_ ),
    .S(net473),
    .X(\register_file_i/_2013_ ));
 sg13g2_a22oi_1 \register_file_i/_5090_  (.Y(\register_file_i/_2014_ ),
    .B1(\register_file_i/_2013_ ),
    .B2(net1785),
    .A2(\register_file_i/_2012_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5091_  (.B1(\register_file_i/_2014_ ),
    .Y(\register_file_i/_2015_ ),
    .A1(net444),
    .A2(\register_file_i/_2011_ ));
 sg13g2_nand2_1 \register_file_i/_5092_  (.Y(\register_file_i/_2016_ ),
    .A(net1910),
    .B(\register_file_i/_2015_ ));
 sg13g2_mux4_1 \register_file_i/_5093_  (.S0(net474),
    .A0(\register_file_i/rf_reg_533_ ),
    .A1(\register_file_i/rf_reg_565_ ),
    .A2(\register_file_i/rf_reg_597_ ),
    .A3(\register_file_i/rf_reg_629_ ),
    .S1(net455),
    .X(\register_file_i/_2017_ ));
 sg13g2_mux4_1 \register_file_i/_5094_  (.S0(net470),
    .A0(\register_file_i/rf_reg_661_ ),
    .A1(\register_file_i/rf_reg_693_ ),
    .A2(\register_file_i/rf_reg_725_ ),
    .A3(\register_file_i/rf_reg_757_ ),
    .S1(net457),
    .X(\register_file_i/_2018_ ));
 sg13g2_buf_2 fanout270 (.A(_04306_),
    .X(net270));
 sg13g2_mux2_1 \register_file_i/_5096_  (.A0(\register_file_i/rf_reg_405_ ),
    .A1(\register_file_i/rf_reg_437_ ),
    .S(net483),
    .X(\register_file_i/_2020_ ));
 sg13g2_mux2_1 \register_file_i/_5097_  (.A0(\register_file_i/rf_reg_469_ ),
    .A1(\register_file_i/rf_reg_501_ ),
    .S(net478),
    .X(\register_file_i/_2021_ ));
 sg13g2_a22oi_1 \register_file_i/_5098_  (.Y(\register_file_i/_2022_ ),
    .B1(\register_file_i/_2021_ ),
    .B2(net1756),
    .A2(\register_file_i/_2020_ ),
    .A1(net1773));
 sg13g2_mux2_1 \register_file_i/_5099_  (.A0(\register_file_i/rf_reg_341_ ),
    .A1(\register_file_i/rf_reg_373_ ),
    .S(net479),
    .X(\register_file_i/_2023_ ));
 sg13g2_mux2_1 \register_file_i/_5100_  (.A0(\register_file_i/rf_reg_277_ ),
    .A1(\register_file_i/rf_reg_309_ ),
    .S(net480),
    .X(\register_file_i/_2024_ ));
 sg13g2_a22oi_1 \register_file_i/_5101_  (.Y(\register_file_i/_2025_ ),
    .B1(\register_file_i/_2024_ ),
    .B2(net1735),
    .A2(\register_file_i/_2023_ ),
    .A1(net1746));
 sg13g2_a21oi_1 \register_file_i/_5102_  (.A1(\register_file_i/_2022_ ),
    .A2(\register_file_i/_2025_ ),
    .Y(\register_file_i/_2026_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5103_  (.B2(net1686),
    .C1(\register_file_i/_2026_ ),
    .B1(\register_file_i/_2018_ ),
    .A1(net1728),
    .Y(\register_file_i/_2027_ ),
    .A2(\register_file_i/_2017_ ));
 sg13g2_nand3_1 \register_file_i/_5104_  (.B(\register_file_i/_2016_ ),
    .C(\register_file_i/_2027_ ),
    .A(\register_file_i/_2009_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_21_ ));
 sg13g2_buf_2 fanout269 (.A(_04369_),
    .X(net269));
 sg13g2_mux2_1 \register_file_i/_5106_  (.A0(\register_file_i/rf_reg_916_ ),
    .A1(\register_file_i/rf_reg_948_ ),
    .S(net484),
    .X(\register_file_i/_2029_ ));
 sg13g2_mux2_1 \register_file_i/_5107_  (.A0(\register_file_i/rf_reg_980_ ),
    .A1(\register_file_i/rf_reg_1012_ ),
    .S(net466),
    .X(\register_file_i/_2030_ ));
 sg13g2_a22oi_1 \register_file_i/_5108_  (.Y(\register_file_i/_2031_ ),
    .B1(\register_file_i/_2030_ ),
    .B2(net1758),
    .A2(\register_file_i/_2029_ ),
    .A1(net1775));
 sg13g2_mux2_1 \register_file_i/_5109_  (.A0(\register_file_i/rf_reg_852_ ),
    .A1(\register_file_i/rf_reg_884_ ),
    .S(net481),
    .X(\register_file_i/_2032_ ));
 sg13g2_mux2_1 \register_file_i/_5110_  (.A0(\register_file_i/rf_reg_788_ ),
    .A1(\register_file_i/rf_reg_820_ ),
    .S(net469),
    .X(\register_file_i/_2033_ ));
 sg13g2_a22oi_1 \register_file_i/_5111_  (.Y(\register_file_i/_2034_ ),
    .B1(\register_file_i/_2033_ ),
    .B2(net1734),
    .A2(\register_file_i/_2032_ ),
    .A1(net1745));
 sg13g2_a21o_1 \register_file_i/_5112_  (.A2(\register_file_i/_2034_ ),
    .A1(\register_file_i/_2031_ ),
    .B1(net1917),
    .X(\register_file_i/_2035_ ));
 sg13g2_mux2_1 \register_file_i/_5113_  (.A0(\register_file_i/rf_reg_52_ ),
    .A1(\register_file_i/rf_reg_116_ ),
    .S(net450),
    .X(\register_file_i/_2036_ ));
 sg13g2_a22oi_1 \register_file_i/_5114_  (.Y(\register_file_i/_2037_ ),
    .B1(\register_file_i/_2036_ ),
    .B2(net515),
    .A2(net1691),
    .A1(\register_file_i/rf_reg_84_ ));
 sg13g2_mux2_1 \register_file_i/_5115_  (.A0(\register_file_i/rf_reg_212_ ),
    .A1(\register_file_i/rf_reg_244_ ),
    .S(net471),
    .X(\register_file_i/_2038_ ));
 sg13g2_mux2_1 \register_file_i/_5116_  (.A0(\register_file_i/rf_reg_148_ ),
    .A1(\register_file_i/rf_reg_180_ ),
    .S(net473),
    .X(\register_file_i/_2039_ ));
 sg13g2_a22oi_1 \register_file_i/_5117_  (.Y(\register_file_i/_2040_ ),
    .B1(\register_file_i/_2039_ ),
    .B2(net1785),
    .A2(\register_file_i/_2038_ ),
    .A1(net1767));
 sg13g2_o21ai_1 \register_file_i/_5118_  (.B1(\register_file_i/_2040_ ),
    .Y(\register_file_i/_2041_ ),
    .A1(net444),
    .A2(\register_file_i/_2037_ ));
 sg13g2_nand2_1 \register_file_i/_5119_  (.Y(\register_file_i/_2042_ ),
    .A(net1911),
    .B(\register_file_i/_2041_ ));
 sg13g2_mux4_1 \register_file_i/_5120_  (.S0(net474),
    .A0(\register_file_i/rf_reg_532_ ),
    .A1(\register_file_i/rf_reg_564_ ),
    .A2(\register_file_i/rf_reg_596_ ),
    .A3(\register_file_i/rf_reg_628_ ),
    .S1(net455),
    .X(\register_file_i/_2043_ ));
 sg13g2_mux4_1 \register_file_i/_5121_  (.S0(net470),
    .A0(\register_file_i/rf_reg_660_ ),
    .A1(\register_file_i/rf_reg_692_ ),
    .A2(\register_file_i/rf_reg_724_ ),
    .A3(\register_file_i/rf_reg_756_ ),
    .S1(net457),
    .X(\register_file_i/_2044_ ));
 sg13g2_mux2_1 \register_file_i/_5122_  (.A0(\register_file_i/rf_reg_404_ ),
    .A1(\register_file_i/rf_reg_436_ ),
    .S(net483),
    .X(\register_file_i/_2045_ ));
 sg13g2_mux2_1 \register_file_i/_5123_  (.A0(\register_file_i/rf_reg_468_ ),
    .A1(\register_file_i/rf_reg_500_ ),
    .S(net477),
    .X(\register_file_i/_2046_ ));
 sg13g2_a22oi_1 \register_file_i/_5124_  (.Y(\register_file_i/_2047_ ),
    .B1(\register_file_i/_2046_ ),
    .B2(net1756),
    .A2(\register_file_i/_2045_ ),
    .A1(net1773));
 sg13g2_mux2_1 \register_file_i/_5125_  (.A0(\register_file_i/rf_reg_340_ ),
    .A1(\register_file_i/rf_reg_372_ ),
    .S(net479),
    .X(\register_file_i/_2048_ ));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(net269));
 sg13g2_mux2_1 \register_file_i/_5127_  (.A0(\register_file_i/rf_reg_276_ ),
    .A1(\register_file_i/rf_reg_308_ ),
    .S(net485),
    .X(\register_file_i/_2050_ ));
 sg13g2_a22oi_1 \register_file_i/_5128_  (.Y(\register_file_i/_2051_ ),
    .B1(\register_file_i/_2050_ ),
    .B2(net1732),
    .A2(\register_file_i/_2048_ ),
    .A1(net1746));
 sg13g2_a21oi_1 \register_file_i/_5129_  (.A1(\register_file_i/_2047_ ),
    .A2(\register_file_i/_2051_ ),
    .Y(\register_file_i/_2052_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5130_  (.B2(net1686),
    .C1(\register_file_i/_2052_ ),
    .B1(\register_file_i/_2044_ ),
    .A1(net1727),
    .Y(\register_file_i/_2053_ ),
    .A2(\register_file_i/_2043_ ));
 sg13g2_nand3_1 \register_file_i/_5131_  (.B(\register_file_i/_2042_ ),
    .C(\register_file_i/_2053_ ),
    .A(\register_file_i/_2035_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_mux2_1 \register_file_i/_5132_  (.A0(\register_file_i/rf_reg_915_ ),
    .A1(\register_file_i/rf_reg_947_ ),
    .S(net484),
    .X(\register_file_i/_2054_ ));
 sg13g2_mux2_1 \register_file_i/_5133_  (.A0(\register_file_i/rf_reg_979_ ),
    .A1(\register_file_i/rf_reg_1011_ ),
    .S(net466),
    .X(\register_file_i/_2055_ ));
 sg13g2_a22oi_1 \register_file_i/_5134_  (.Y(\register_file_i/_2056_ ),
    .B1(\register_file_i/_2055_ ),
    .B2(net1758),
    .A2(\register_file_i/_2054_ ),
    .A1(net1775));
 sg13g2_mux2_1 \register_file_i/_5135_  (.A0(\register_file_i/rf_reg_851_ ),
    .A1(\register_file_i/rf_reg_883_ ),
    .S(net481),
    .X(\register_file_i/_2057_ ));
 sg13g2_mux2_1 \register_file_i/_5136_  (.A0(\register_file_i/rf_reg_787_ ),
    .A1(\register_file_i/rf_reg_819_ ),
    .S(net469),
    .X(\register_file_i/_2058_ ));
 sg13g2_a22oi_1 \register_file_i/_5137_  (.Y(\register_file_i/_2059_ ),
    .B1(\register_file_i/_2058_ ),
    .B2(net1734),
    .A2(\register_file_i/_2057_ ),
    .A1(net1745));
 sg13g2_a21o_1 \register_file_i/_5138_  (.A2(\register_file_i/_2059_ ),
    .A1(\register_file_i/_2056_ ),
    .B1(net1916),
    .X(\register_file_i/_2060_ ));
 sg13g2_mux2_1 \register_file_i/_5139_  (.A0(\register_file_i/rf_reg_51_ ),
    .A1(\register_file_i/rf_reg_115_ ),
    .S(net450),
    .X(\register_file_i/_2061_ ));
 sg13g2_a22oi_1 \register_file_i/_5140_  (.Y(\register_file_i/_2062_ ),
    .B1(\register_file_i/_2061_ ),
    .B2(net514),
    .A2(net1691),
    .A1(\register_file_i/rf_reg_83_ ));
 sg13g2_buf_2 fanout267 (.A(net269),
    .X(net267));
 sg13g2_mux2_1 \register_file_i/_5142_  (.A0(\register_file_i/rf_reg_211_ ),
    .A1(\register_file_i/rf_reg_243_ ),
    .S(net471),
    .X(\register_file_i/_2064_ ));
 sg13g2_mux2_1 \register_file_i/_5143_  (.A0(\register_file_i/rf_reg_147_ ),
    .A1(\register_file_i/rf_reg_179_ ),
    .S(net473),
    .X(\register_file_i/_2065_ ));
 sg13g2_a22oi_1 \register_file_i/_5144_  (.Y(\register_file_i/_2066_ ),
    .B1(\register_file_i/_2065_ ),
    .B2(net1785),
    .A2(\register_file_i/_2064_ ),
    .A1(net1767));
 sg13g2_o21ai_1 \register_file_i/_5145_  (.B1(\register_file_i/_2066_ ),
    .Y(\register_file_i/_2067_ ),
    .A1(net443),
    .A2(\register_file_i/_2062_ ));
 sg13g2_nand2_1 \register_file_i/_5146_  (.Y(\register_file_i/_2068_ ),
    .A(net1910),
    .B(\register_file_i/_2067_ ));
 sg13g2_buf_4 fanout266 (.X(net266),
    .A(_04608_));
 sg13g2_mux4_1 \register_file_i/_5148_  (.S0(net474),
    .A0(\register_file_i/rf_reg_531_ ),
    .A1(\register_file_i/rf_reg_563_ ),
    .A2(\register_file_i/rf_reg_595_ ),
    .A3(\register_file_i/rf_reg_627_ ),
    .S1(net459),
    .X(\register_file_i/_2070_ ));
 sg13g2_mux4_1 \register_file_i/_5149_  (.S0(net470),
    .A0(\register_file_i/rf_reg_659_ ),
    .A1(\register_file_i/rf_reg_691_ ),
    .A2(\register_file_i/rf_reg_723_ ),
    .A3(\register_file_i/rf_reg_755_ ),
    .S1(net457),
    .X(\register_file_i/_2071_ ));
 sg13g2_mux2_1 \register_file_i/_5150_  (.A0(\register_file_i/rf_reg_403_ ),
    .A1(\register_file_i/rf_reg_435_ ),
    .S(net482),
    .X(\register_file_i/_2072_ ));
 sg13g2_mux2_1 \register_file_i/_5151_  (.A0(\register_file_i/rf_reg_467_ ),
    .A1(\register_file_i/rf_reg_499_ ),
    .S(net477),
    .X(\register_file_i/_2073_ ));
 sg13g2_a22oi_1 \register_file_i/_5152_  (.Y(\register_file_i/_2074_ ),
    .B1(\register_file_i/_2073_ ),
    .B2(net1755),
    .A2(\register_file_i/_2072_ ),
    .A1(net1773));
 sg13g2_mux2_1 \register_file_i/_5153_  (.A0(\register_file_i/rf_reg_339_ ),
    .A1(\register_file_i/rf_reg_371_ ),
    .S(net479),
    .X(\register_file_i/_2075_ ));
 sg13g2_mux2_1 \register_file_i/_5154_  (.A0(\register_file_i/rf_reg_275_ ),
    .A1(\register_file_i/rf_reg_307_ ),
    .S(net485),
    .X(\register_file_i/_2076_ ));
 sg13g2_a22oi_1 \register_file_i/_5155_  (.Y(\register_file_i/_2077_ ),
    .B1(\register_file_i/_2076_ ),
    .B2(net1732),
    .A2(\register_file_i/_2075_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5156_  (.A1(\register_file_i/_2074_ ),
    .A2(\register_file_i/_2077_ ),
    .Y(\register_file_i/_2078_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5157_  (.B2(net1685),
    .C1(\register_file_i/_2078_ ),
    .B1(\register_file_i/_2071_ ),
    .A1(net1727),
    .Y(\register_file_i/_2079_ ),
    .A2(\register_file_i/_2070_ ));
 sg13g2_nand3_1 \register_file_i/_5158_  (.B(\register_file_i/_2068_ ),
    .C(\register_file_i/_2079_ ),
    .A(\register_file_i/_2060_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_mux2_1 \register_file_i/_5159_  (.A0(\register_file_i/rf_reg_914_ ),
    .A1(\register_file_i/rf_reg_946_ ),
    .S(net484),
    .X(\register_file_i/_2080_ ));
 sg13g2_mux2_1 \register_file_i/_5160_  (.A0(\register_file_i/rf_reg_978_ ),
    .A1(\register_file_i/rf_reg_1010_ ),
    .S(net466),
    .X(\register_file_i/_2081_ ));
 sg13g2_a22oi_1 \register_file_i/_5161_  (.Y(\register_file_i/_2082_ ),
    .B1(\register_file_i/_2081_ ),
    .B2(net1757),
    .A2(\register_file_i/_2080_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5162_  (.A0(\register_file_i/rf_reg_850_ ),
    .A1(\register_file_i/rf_reg_882_ ),
    .S(net481),
    .X(\register_file_i/_2083_ ));
 sg13g2_buf_1 fanout265 (.A(net266),
    .X(net265));
 sg13g2_mux2_1 \register_file_i/_5164_  (.A0(\register_file_i/rf_reg_786_ ),
    .A1(\register_file_i/rf_reg_818_ ),
    .S(net487),
    .X(\register_file_i/_2085_ ));
 sg13g2_a22oi_1 \register_file_i/_5165_  (.Y(\register_file_i/_2086_ ),
    .B1(\register_file_i/_2085_ ),
    .B2(net1733),
    .A2(\register_file_i/_2083_ ),
    .A1(net1744));
 sg13g2_a21o_1 \register_file_i/_5166_  (.A2(\register_file_i/_2086_ ),
    .A1(\register_file_i/_2082_ ),
    .B1(net1916),
    .X(\register_file_i/_2087_ ));
 sg13g2_mux2_1 \register_file_i/_5167_  (.A0(\register_file_i/rf_reg_50_ ),
    .A1(\register_file_i/rf_reg_114_ ),
    .S(net450),
    .X(\register_file_i/_2088_ ));
 sg13g2_a22oi_1 \register_file_i/_5168_  (.Y(\register_file_i/_2089_ ),
    .B1(\register_file_i/_2088_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_82_ ));
 sg13g2_mux2_1 \register_file_i/_5169_  (.A0(\register_file_i/rf_reg_210_ ),
    .A1(\register_file_i/rf_reg_242_ ),
    .S(net471),
    .X(\register_file_i/_2090_ ));
 sg13g2_mux2_1 \register_file_i/_5170_  (.A0(\register_file_i/rf_reg_146_ ),
    .A1(\register_file_i/rf_reg_178_ ),
    .S(net472),
    .X(\register_file_i/_2091_ ));
 sg13g2_a22oi_1 \register_file_i/_5171_  (.Y(\register_file_i/_2092_ ),
    .B1(\register_file_i/_2091_ ),
    .B2(net1784),
    .A2(\register_file_i/_2090_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5172_  (.B1(\register_file_i/_2092_ ),
    .Y(\register_file_i/_2093_ ),
    .A1(net443),
    .A2(\register_file_i/_2089_ ));
 sg13g2_nand2_1 \register_file_i/_5173_  (.Y(\register_file_i/_2094_ ),
    .A(net1910),
    .B(\register_file_i/_2093_ ));
 sg13g2_mux4_1 \register_file_i/_5174_  (.S0(net474),
    .A0(\register_file_i/rf_reg_530_ ),
    .A1(\register_file_i/rf_reg_562_ ),
    .A2(\register_file_i/rf_reg_594_ ),
    .A3(\register_file_i/rf_reg_626_ ),
    .S1(net459),
    .X(\register_file_i/_2095_ ));
 sg13g2_buf_4 fanout264 (.X(net264),
    .A(net266));
 sg13g2_mux4_1 \register_file_i/_5176_  (.S0(net488),
    .A0(\register_file_i/rf_reg_658_ ),
    .A1(\register_file_i/rf_reg_690_ ),
    .A2(\register_file_i/rf_reg_722_ ),
    .A3(\register_file_i/rf_reg_754_ ),
    .S1(net457),
    .X(\register_file_i/_2097_ ));
 sg13g2_mux2_1 \register_file_i/_5177_  (.A0(\register_file_i/rf_reg_402_ ),
    .A1(\register_file_i/rf_reg_434_ ),
    .S(net482),
    .X(\register_file_i/_2098_ ));
 sg13g2_buf_2 fanout263 (.A(\cs_registers_i/_0594_ ),
    .X(net263));
 sg13g2_mux2_1 \register_file_i/_5179_  (.A0(\register_file_i/rf_reg_466_ ),
    .A1(\register_file_i/rf_reg_498_ ),
    .S(net489),
    .X(\register_file_i/_2100_ ));
 sg13g2_a22oi_1 \register_file_i/_5180_  (.Y(\register_file_i/_2101_ ),
    .B1(\register_file_i/_2100_ ),
    .B2(net1755),
    .A2(\register_file_i/_2098_ ),
    .A1(net1772));
 sg13g2_mux2_1 \register_file_i/_5181_  (.A0(\register_file_i/rf_reg_338_ ),
    .A1(\register_file_i/rf_reg_370_ ),
    .S(net478),
    .X(\register_file_i/_2102_ ));
 sg13g2_mux2_1 \register_file_i/_5182_  (.A0(\register_file_i/rf_reg_274_ ),
    .A1(\register_file_i/rf_reg_306_ ),
    .S(net485),
    .X(\register_file_i/_2103_ ));
 sg13g2_a22oi_1 \register_file_i/_5183_  (.Y(\register_file_i/_2104_ ),
    .B1(\register_file_i/_2103_ ),
    .B2(net1732),
    .A2(\register_file_i/_2102_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5184_  (.A1(\register_file_i/_2101_ ),
    .A2(\register_file_i/_2104_ ),
    .Y(\register_file_i/_2105_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5185_  (.B2(net1685),
    .C1(\register_file_i/_2105_ ),
    .B1(\register_file_i/_2097_ ),
    .A1(net1727),
    .Y(\register_file_i/_2106_ ),
    .A2(\register_file_i/_2095_ ));
 sg13g2_nand3_1 \register_file_i/_5186_  (.B(\register_file_i/_2094_ ),
    .C(\register_file_i/_2106_ ),
    .A(\register_file_i/_2087_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_18_ ));
 sg13g2_mux2_1 \register_file_i/_5187_  (.A0(\register_file_i/rf_reg_913_ ),
    .A1(\register_file_i/rf_reg_945_ ),
    .S(net484),
    .X(\register_file_i/_2107_ ));
 sg13g2_mux2_1 \register_file_i/_5188_  (.A0(\register_file_i/rf_reg_977_ ),
    .A1(\register_file_i/rf_reg_1009_ ),
    .S(net466),
    .X(\register_file_i/_2108_ ));
 sg13g2_a22oi_1 \register_file_i/_5189_  (.Y(\register_file_i/_2109_ ),
    .B1(\register_file_i/_2108_ ),
    .B2(net1757),
    .A2(\register_file_i/_2107_ ),
    .A1(net1775));
 sg13g2_mux2_1 \register_file_i/_5190_  (.A0(\register_file_i/rf_reg_849_ ),
    .A1(\register_file_i/rf_reg_881_ ),
    .S(net481),
    .X(\register_file_i/_2110_ ));
 sg13g2_mux2_1 \register_file_i/_5191_  (.A0(\register_file_i/rf_reg_785_ ),
    .A1(\register_file_i/rf_reg_817_ ),
    .S(net486),
    .X(\register_file_i/_2111_ ));
 sg13g2_a22oi_1 \register_file_i/_5192_  (.Y(\register_file_i/_2112_ ),
    .B1(\register_file_i/_2111_ ),
    .B2(net1733),
    .A2(\register_file_i/_2110_ ),
    .A1(net1744));
 sg13g2_a21o_1 \register_file_i/_5193_  (.A2(\register_file_i/_2112_ ),
    .A1(\register_file_i/_2109_ ),
    .B1(net1916),
    .X(\register_file_i/_2113_ ));
 sg13g2_mux2_1 \register_file_i/_5194_  (.A0(\register_file_i/rf_reg_49_ ),
    .A1(\register_file_i/rf_reg_113_ ),
    .S(net450),
    .X(\register_file_i/_2114_ ));
 sg13g2_a22oi_1 \register_file_i/_5195_  (.Y(\register_file_i/_2115_ ),
    .B1(\register_file_i/_2114_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_81_ ));
 sg13g2_mux2_1 \register_file_i/_5196_  (.A0(\register_file_i/rf_reg_209_ ),
    .A1(\register_file_i/rf_reg_241_ ),
    .S(net471),
    .X(\register_file_i/_2116_ ));
 sg13g2_mux2_1 \register_file_i/_5197_  (.A0(\register_file_i/rf_reg_145_ ),
    .A1(\register_file_i/rf_reg_177_ ),
    .S(net472),
    .X(\register_file_i/_2117_ ));
 sg13g2_a22oi_1 \register_file_i/_5198_  (.Y(\register_file_i/_2118_ ),
    .B1(\register_file_i/_2117_ ),
    .B2(net1785),
    .A2(\register_file_i/_2116_ ),
    .A1(net1767));
 sg13g2_o21ai_1 \register_file_i/_5199_  (.B1(\register_file_i/_2118_ ),
    .Y(\register_file_i/_2119_ ),
    .A1(net443),
    .A2(\register_file_i/_2115_ ));
 sg13g2_nand2_1 \register_file_i/_5200_  (.Y(\register_file_i/_2120_ ),
    .A(net1910),
    .B(\register_file_i/_2119_ ));
 sg13g2_buf_1 fanout262 (.A(net263),
    .X(net262));
 sg13g2_mux4_1 \register_file_i/_5202_  (.S0(net474),
    .A0(\register_file_i/rf_reg_529_ ),
    .A1(\register_file_i/rf_reg_561_ ),
    .A2(\register_file_i/rf_reg_593_ ),
    .A3(\register_file_i/rf_reg_625_ ),
    .S1(net458),
    .X(\register_file_i/_2122_ ));
 sg13g2_mux4_1 \register_file_i/_5203_  (.S0(net488),
    .A0(\register_file_i/rf_reg_657_ ),
    .A1(\register_file_i/rf_reg_689_ ),
    .A2(\register_file_i/rf_reg_721_ ),
    .A3(\register_file_i/rf_reg_753_ ),
    .S1(net457),
    .X(\register_file_i/_2123_ ));
 sg13g2_mux2_1 \register_file_i/_5204_  (.A0(\register_file_i/rf_reg_401_ ),
    .A1(\register_file_i/rf_reg_433_ ),
    .S(net482),
    .X(\register_file_i/_2124_ ));
 sg13g2_mux2_1 \register_file_i/_5205_  (.A0(\register_file_i/rf_reg_465_ ),
    .A1(\register_file_i/rf_reg_497_ ),
    .S(net489),
    .X(\register_file_i/_2125_ ));
 sg13g2_a22oi_1 \register_file_i/_5206_  (.Y(\register_file_i/_2126_ ),
    .B1(\register_file_i/_2125_ ),
    .B2(net1755),
    .A2(\register_file_i/_2124_ ),
    .A1(net1773));
 sg13g2_mux2_1 \register_file_i/_5207_  (.A0(\register_file_i/rf_reg_337_ ),
    .A1(\register_file_i/rf_reg_369_ ),
    .S(net478),
    .X(\register_file_i/_2127_ ));
 sg13g2_mux2_1 \register_file_i/_5208_  (.A0(\register_file_i/rf_reg_273_ ),
    .A1(\register_file_i/rf_reg_305_ ),
    .S(net485),
    .X(\register_file_i/_2128_ ));
 sg13g2_a22oi_1 \register_file_i/_5209_  (.Y(\register_file_i/_2129_ ),
    .B1(\register_file_i/_2128_ ),
    .B2(net1732),
    .A2(\register_file_i/_2127_ ),
    .A1(net1743));
 sg13g2_buf_2 fanout261 (.A(net263),
    .X(net261));
 sg13g2_a21oi_1 \register_file_i/_5211_  (.A1(\register_file_i/_2126_ ),
    .A2(\register_file_i/_2129_ ),
    .Y(\register_file_i/_2131_ ),
    .B1(net1723));
 sg13g2_a221oi_1 \register_file_i/_5212_  (.B2(net1685),
    .C1(\register_file_i/_2131_ ),
    .B1(\register_file_i/_2123_ ),
    .A1(net1728),
    .Y(\register_file_i/_2132_ ),
    .A2(\register_file_i/_2122_ ));
 sg13g2_nand3_1 \register_file_i/_5213_  (.B(\register_file_i/_2120_ ),
    .C(\register_file_i/_2132_ ),
    .A(\register_file_i/_2113_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_17_ ));
 sg13g2_mux2_1 \register_file_i/_5214_  (.A0(\register_file_i/rf_reg_912_ ),
    .A1(\register_file_i/rf_reg_944_ ),
    .S(net484),
    .X(\register_file_i/_2133_ ));
 sg13g2_mux2_1 \register_file_i/_5215_  (.A0(\register_file_i/rf_reg_976_ ),
    .A1(\register_file_i/rf_reg_1008_ ),
    .S(net466),
    .X(\register_file_i/_2134_ ));
 sg13g2_a22oi_1 \register_file_i/_5216_  (.Y(\register_file_i/_2135_ ),
    .B1(\register_file_i/_2134_ ),
    .B2(net1757),
    .A2(\register_file_i/_2133_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5217_  (.A0(\register_file_i/rf_reg_848_ ),
    .A1(\register_file_i/rf_reg_880_ ),
    .S(net481),
    .X(\register_file_i/_2136_ ));
 sg13g2_mux2_1 \register_file_i/_5218_  (.A0(\register_file_i/rf_reg_784_ ),
    .A1(\register_file_i/rf_reg_816_ ),
    .S(net486),
    .X(\register_file_i/_2137_ ));
 sg13g2_a22oi_1 \register_file_i/_5219_  (.Y(\register_file_i/_2138_ ),
    .B1(\register_file_i/_2137_ ),
    .B2(net1733),
    .A2(\register_file_i/_2136_ ),
    .A1(net1744));
 sg13g2_a21o_1 \register_file_i/_5220_  (.A2(\register_file_i/_2138_ ),
    .A1(\register_file_i/_2135_ ),
    .B1(net1916),
    .X(\register_file_i/_2139_ ));
 sg13g2_buf_2 fanout260 (.A(\cs_registers_i/_0594_ ),
    .X(net260));
 sg13g2_mux2_1 \register_file_i/_5222_  (.A0(\register_file_i/rf_reg_48_ ),
    .A1(\register_file_i/rf_reg_112_ ),
    .S(net451),
    .X(\register_file_i/_2141_ ));
 sg13g2_a22oi_1 \register_file_i/_5223_  (.Y(\register_file_i/_2142_ ),
    .B1(\register_file_i/_2141_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_80_ ));
 sg13g2_buf_4 fanout259 (.X(net259),
    .A(\cs_registers_i/_0594_ ));
 sg13g2_mux2_1 \register_file_i/_5225_  (.A0(\register_file_i/rf_reg_208_ ),
    .A1(\register_file_i/rf_reg_240_ ),
    .S(net490),
    .X(\register_file_i/_2144_ ));
 sg13g2_mux2_1 \register_file_i/_5226_  (.A0(\register_file_i/rf_reg_144_ ),
    .A1(\register_file_i/rf_reg_176_ ),
    .S(net472),
    .X(\register_file_i/_2145_ ));
 sg13g2_a22oi_1 \register_file_i/_5227_  (.Y(\register_file_i/_2146_ ),
    .B1(\register_file_i/_2145_ ),
    .B2(net1784),
    .A2(\register_file_i/_2144_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5228_  (.B1(\register_file_i/_2146_ ),
    .Y(\register_file_i/_2147_ ),
    .A1(net443),
    .A2(\register_file_i/_2142_ ));
 sg13g2_nand2_1 \register_file_i/_5229_  (.Y(\register_file_i/_2148_ ),
    .A(net1910),
    .B(\register_file_i/_2147_ ));
 sg13g2_mux4_1 \register_file_i/_5230_  (.S0(net473),
    .A0(\register_file_i/rf_reg_528_ ),
    .A1(\register_file_i/rf_reg_560_ ),
    .A2(\register_file_i/rf_reg_592_ ),
    .A3(\register_file_i/rf_reg_624_ ),
    .S1(net458),
    .X(\register_file_i/_2149_ ));
 sg13g2_mux4_1 \register_file_i/_5231_  (.S0(net488),
    .A0(\register_file_i/rf_reg_656_ ),
    .A1(\register_file_i/rf_reg_688_ ),
    .A2(\register_file_i/rf_reg_720_ ),
    .A3(\register_file_i/rf_reg_752_ ),
    .S1(net457),
    .X(\register_file_i/_2150_ ));
 sg13g2_mux2_1 \register_file_i/_5232_  (.A0(\register_file_i/rf_reg_400_ ),
    .A1(\register_file_i/rf_reg_432_ ),
    .S(net482),
    .X(\register_file_i/_2151_ ));
 sg13g2_mux2_1 \register_file_i/_5233_  (.A0(\register_file_i/rf_reg_464_ ),
    .A1(\register_file_i/rf_reg_496_ ),
    .S(net489),
    .X(\register_file_i/_2152_ ));
 sg13g2_buf_4 fanout258 (.X(net258),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_10_ ));
 sg13g2_a22oi_1 \register_file_i/_5235_  (.Y(\register_file_i/_2154_ ),
    .B1(\register_file_i/_2152_ ),
    .B2(net1756),
    .A2(\register_file_i/_2151_ ),
    .A1(net1772));
 sg13g2_mux2_1 \register_file_i/_5236_  (.A0(\register_file_i/rf_reg_336_ ),
    .A1(\register_file_i/rf_reg_368_ ),
    .S(net478),
    .X(\register_file_i/_2155_ ));
 sg13g2_mux2_1 \register_file_i/_5237_  (.A0(\register_file_i/rf_reg_272_ ),
    .A1(\register_file_i/rf_reg_304_ ),
    .S(net485),
    .X(\register_file_i/_2156_ ));
 sg13g2_a22oi_1 \register_file_i/_5238_  (.Y(\register_file_i/_2157_ ),
    .B1(\register_file_i/_2156_ ),
    .B2(net1732),
    .A2(\register_file_i/_2155_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5239_  (.A1(\register_file_i/_2154_ ),
    .A2(\register_file_i/_2157_ ),
    .Y(\register_file_i/_2158_ ),
    .B1(net1723));
 sg13g2_a221oi_1 \register_file_i/_5240_  (.B2(net1685),
    .C1(\register_file_i/_2158_ ),
    .B1(\register_file_i/_2150_ ),
    .A1(net1728),
    .Y(\register_file_i/_2159_ ),
    .A2(\register_file_i/_2149_ ));
 sg13g2_nand3_1 \register_file_i/_5241_  (.B(\register_file_i/_2148_ ),
    .C(\register_file_i/_2159_ ),
    .A(\register_file_i/_2139_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_16_ ));
 sg13g2_mux2_1 \register_file_i/_5242_  (.A0(\register_file_i/rf_reg_911_ ),
    .A1(\register_file_i/rf_reg_943_ ),
    .S(net483),
    .X(\register_file_i/_2160_ ));
 sg13g2_buf_2 fanout257 (.A(csr_save_cause),
    .X(net257));
 sg13g2_mux2_1 \register_file_i/_5244_  (.A0(\register_file_i/rf_reg_975_ ),
    .A1(\register_file_i/rf_reg_1007_ ),
    .S(net492),
    .X(\register_file_i/_2162_ ));
 sg13g2_a22oi_1 \register_file_i/_5245_  (.Y(\register_file_i/_2163_ ),
    .B1(\register_file_i/_2162_ ),
    .B2(net1757),
    .A2(\register_file_i/_2160_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5246_  (.A0(\register_file_i/rf_reg_847_ ),
    .A1(\register_file_i/rf_reg_879_ ),
    .S(net481),
    .X(\register_file_i/_2164_ ));
 sg13g2_mux2_1 \register_file_i/_5247_  (.A0(\register_file_i/rf_reg_783_ ),
    .A1(\register_file_i/rf_reg_815_ ),
    .S(net486),
    .X(\register_file_i/_2165_ ));
 sg13g2_a22oi_1 \register_file_i/_5248_  (.Y(\register_file_i/_2166_ ),
    .B1(\register_file_i/_2165_ ),
    .B2(net1739),
    .A2(\register_file_i/_2164_ ),
    .A1(net1750));
 sg13g2_a21o_1 \register_file_i/_5249_  (.A2(\register_file_i/_2166_ ),
    .A1(\register_file_i/_2163_ ),
    .B1(net1916),
    .X(\register_file_i/_2167_ ));
 sg13g2_mux2_1 \register_file_i/_5250_  (.A0(\register_file_i/rf_reg_47_ ),
    .A1(\register_file_i/rf_reg_111_ ),
    .S(net451),
    .X(\register_file_i/_2168_ ));
 sg13g2_a22oi_1 \register_file_i/_5251_  (.Y(\register_file_i/_2169_ ),
    .B1(\register_file_i/_2168_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_79_ ));
 sg13g2_mux2_1 \register_file_i/_5252_  (.A0(\register_file_i/rf_reg_207_ ),
    .A1(\register_file_i/rf_reg_239_ ),
    .S(net490),
    .X(\register_file_i/_2170_ ));
 sg13g2_mux2_1 \register_file_i/_5253_  (.A0(\register_file_i/rf_reg_143_ ),
    .A1(\register_file_i/rf_reg_175_ ),
    .S(net472),
    .X(\register_file_i/_2171_ ));
 sg13g2_buf_4 fanout256 (.X(net256),
    .A(csr_save_cause));
 sg13g2_a22oi_1 \register_file_i/_5255_  (.Y(\register_file_i/_2173_ ),
    .B1(\register_file_i/_2171_ ),
    .B2(net1784),
    .A2(\register_file_i/_2170_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5256_  (.B1(\register_file_i/_2173_ ),
    .Y(\register_file_i/_2174_ ),
    .A1(net443),
    .A2(\register_file_i/_2169_ ));
 sg13g2_nand2_1 \register_file_i/_5257_  (.Y(\register_file_i/_2175_ ),
    .A(net1910),
    .B(\register_file_i/_2174_ ));
 sg13g2_mux4_1 \register_file_i/_5258_  (.S0(net473),
    .A0(\register_file_i/rf_reg_527_ ),
    .A1(\register_file_i/rf_reg_559_ ),
    .A2(\register_file_i/rf_reg_591_ ),
    .A3(\register_file_i/rf_reg_623_ ),
    .S1(net458),
    .X(\register_file_i/_2176_ ));
 sg13g2_mux4_1 \register_file_i/_5259_  (.S0(net487),
    .A0(\register_file_i/rf_reg_655_ ),
    .A1(\register_file_i/rf_reg_687_ ),
    .A2(\register_file_i/rf_reg_719_ ),
    .A3(\register_file_i/rf_reg_751_ ),
    .S1(net457),
    .X(\register_file_i/_2177_ ));
 sg13g2_mux2_1 \register_file_i/_5260_  (.A0(\register_file_i/rf_reg_399_ ),
    .A1(\register_file_i/rf_reg_431_ ),
    .S(net482),
    .X(\register_file_i/_2178_ ));
 sg13g2_mux2_1 \register_file_i/_5261_  (.A0(\register_file_i/rf_reg_463_ ),
    .A1(\register_file_i/rf_reg_495_ ),
    .S(net489),
    .X(\register_file_i/_2179_ ));
 sg13g2_a22oi_1 \register_file_i/_5262_  (.Y(\register_file_i/_2180_ ),
    .B1(\register_file_i/_2179_ ),
    .B2(net1755),
    .A2(\register_file_i/_2178_ ),
    .A1(net1772));
 sg13g2_mux2_1 \register_file_i/_5263_  (.A0(\register_file_i/rf_reg_335_ ),
    .A1(\register_file_i/rf_reg_367_ ),
    .S(net478),
    .X(\register_file_i/_2181_ ));
 sg13g2_mux2_1 \register_file_i/_5264_  (.A0(\register_file_i/rf_reg_271_ ),
    .A1(\register_file_i/rf_reg_303_ ),
    .S(net485),
    .X(\register_file_i/_2182_ ));
 sg13g2_buf_2 fanout255 (.A(csr_save_cause),
    .X(net255));
 sg13g2_a22oi_1 \register_file_i/_5266_  (.Y(\register_file_i/_2184_ ),
    .B1(\register_file_i/_2182_ ),
    .B2(net1732),
    .A2(\register_file_i/_2181_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5267_  (.A1(\register_file_i/_2180_ ),
    .A2(\register_file_i/_2184_ ),
    .Y(\register_file_i/_2185_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5268_  (.B2(net1685),
    .C1(\register_file_i/_2185_ ),
    .B1(\register_file_i/_2177_ ),
    .A1(net1727),
    .Y(\register_file_i/_2186_ ),
    .A2(\register_file_i/_2176_ ));
 sg13g2_nand3_1 \register_file_i/_5269_  (.B(\register_file_i/_2175_ ),
    .C(\register_file_i/_2186_ ),
    .A(\register_file_i/_2167_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_15_ ));
 sg13g2_mux2_1 \register_file_i/_5270_  (.A0(\register_file_i/rf_reg_910_ ),
    .A1(\register_file_i/rf_reg_942_ ),
    .S(net483),
    .X(\register_file_i/_2187_ ));
 sg13g2_mux2_1 \register_file_i/_5271_  (.A0(\register_file_i/rf_reg_974_ ),
    .A1(\register_file_i/rf_reg_1006_ ),
    .S(net491),
    .X(\register_file_i/_2188_ ));
 sg13g2_a22oi_1 \register_file_i/_5272_  (.Y(\register_file_i/_2189_ ),
    .B1(\register_file_i/_2188_ ),
    .B2(net1757),
    .A2(\register_file_i/_2187_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5273_  (.A0(\register_file_i/rf_reg_846_ ),
    .A1(\register_file_i/rf_reg_878_ ),
    .S(net481),
    .X(\register_file_i/_2190_ ));
 sg13g2_mux2_1 \register_file_i/_5274_  (.A0(\register_file_i/rf_reg_782_ ),
    .A1(\register_file_i/rf_reg_814_ ),
    .S(net486),
    .X(\register_file_i/_2191_ ));
 sg13g2_a22oi_1 \register_file_i/_5275_  (.Y(\register_file_i/_2192_ ),
    .B1(\register_file_i/_2191_ ),
    .B2(net1733),
    .A2(\register_file_i/_2190_ ),
    .A1(net1744));
 sg13g2_a21o_1 \register_file_i/_5276_  (.A2(\register_file_i/_2192_ ),
    .A1(\register_file_i/_2189_ ),
    .B1(net1916),
    .X(\register_file_i/_2193_ ));
 sg13g2_mux2_1 \register_file_i/_5277_  (.A0(\register_file_i/rf_reg_46_ ),
    .A1(\register_file_i/rf_reg_110_ ),
    .S(net451),
    .X(\register_file_i/_2194_ ));
 sg13g2_a22oi_1 \register_file_i/_5278_  (.Y(\register_file_i/_2195_ ),
    .B1(\register_file_i/_2194_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_78_ ));
 sg13g2_mux2_1 \register_file_i/_5279_  (.A0(\register_file_i/rf_reg_206_ ),
    .A1(\register_file_i/rf_reg_238_ ),
    .S(net490),
    .X(\register_file_i/_2196_ ));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_04618_));
 sg13g2_mux2_1 \register_file_i/_5281_  (.A0(\register_file_i/rf_reg_142_ ),
    .A1(\register_file_i/rf_reg_174_ ),
    .S(net493),
    .X(\register_file_i/_2198_ ));
 sg13g2_a22oi_1 \register_file_i/_5282_  (.Y(\register_file_i/_2199_ ),
    .B1(\register_file_i/_2198_ ),
    .B2(net1784),
    .A2(\register_file_i/_2196_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5283_  (.B1(\register_file_i/_2199_ ),
    .Y(\register_file_i/_2200_ ),
    .A1(net443),
    .A2(\register_file_i/_2195_ ));
 sg13g2_nand2_1 \register_file_i/_5284_  (.Y(\register_file_i/_2201_ ),
    .A(net1911),
    .B(\register_file_i/_2200_ ));
 sg13g2_mux4_1 \register_file_i/_5285_  (.S0(net473),
    .A0(\register_file_i/rf_reg_526_ ),
    .A1(\register_file_i/rf_reg_558_ ),
    .A2(\register_file_i/rf_reg_590_ ),
    .A3(\register_file_i/rf_reg_622_ ),
    .S1(net458),
    .X(\register_file_i/_2202_ ));
 sg13g2_mux4_1 \register_file_i/_5286_  (.S0(net487),
    .A0(\register_file_i/rf_reg_654_ ),
    .A1(\register_file_i/rf_reg_686_ ),
    .A2(\register_file_i/rf_reg_718_ ),
    .A3(\register_file_i/rf_reg_750_ ),
    .S1(net456),
    .X(\register_file_i/_2203_ ));
 sg13g2_mux2_1 \register_file_i/_5287_  (.A0(\register_file_i/rf_reg_398_ ),
    .A1(\register_file_i/rf_reg_430_ ),
    .S(net482),
    .X(\register_file_i/_2204_ ));
 sg13g2_mux2_1 \register_file_i/_5288_  (.A0(\register_file_i/rf_reg_462_ ),
    .A1(\register_file_i/rf_reg_494_ ),
    .S(net489),
    .X(\register_file_i/_2205_ ));
 sg13g2_a22oi_1 \register_file_i/_5289_  (.Y(\register_file_i/_2206_ ),
    .B1(\register_file_i/_2205_ ),
    .B2(net1755),
    .A2(\register_file_i/_2204_ ),
    .A1(net1772));
 sg13g2_buf_2 fanout253 (.A(_04618_),
    .X(net253));
 sg13g2_buf_2 fanout252 (.A(_04704_),
    .X(net252));
 sg13g2_mux2_1 \register_file_i/_5292_  (.A0(\register_file_i/rf_reg_334_ ),
    .A1(\register_file_i/rf_reg_366_ ),
    .S(net494),
    .X(\register_file_i/_2209_ ));
 sg13g2_mux2_1 \register_file_i/_5293_  (.A0(\register_file_i/rf_reg_270_ ),
    .A1(\register_file_i/rf_reg_302_ ),
    .S(net485),
    .X(\register_file_i/_2210_ ));
 sg13g2_a22oi_1 \register_file_i/_5294_  (.Y(\register_file_i/_2211_ ),
    .B1(\register_file_i/_2210_ ),
    .B2(net1732),
    .A2(\register_file_i/_2209_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5295_  (.A1(\register_file_i/_2206_ ),
    .A2(\register_file_i/_2211_ ),
    .Y(\register_file_i/_2212_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5296_  (.B2(net1685),
    .C1(\register_file_i/_2212_ ),
    .B1(\register_file_i/_2203_ ),
    .A1(net1727),
    .Y(\register_file_i/_2213_ ),
    .A2(\register_file_i/_2202_ ));
 sg13g2_nand3_1 \register_file_i/_5297_  (.B(\register_file_i/_2201_ ),
    .C(\register_file_i/_2213_ ),
    .A(\register_file_i/_2193_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_14_ ));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(net252));
 sg13g2_mux2_1 \register_file_i/_5299_  (.A0(\register_file_i/rf_reg_909_ ),
    .A1(\register_file_i/rf_reg_941_ ),
    .S(net483),
    .X(\register_file_i/_2215_ ));
 sg13g2_mux2_1 \register_file_i/_5300_  (.A0(\register_file_i/rf_reg_973_ ),
    .A1(\register_file_i/rf_reg_1005_ ),
    .S(net491),
    .X(\register_file_i/_2216_ ));
 sg13g2_buf_1 fanout250 (.A(_04946_),
    .X(net250));
 sg13g2_a22oi_1 \register_file_i/_5302_  (.Y(\register_file_i/_2218_ ),
    .B1(\register_file_i/_2216_ ),
    .B2(net1757),
    .A2(\register_file_i/_2215_ ),
    .A1(net1774));
 sg13g2_buf_2 fanout249 (.A(_04946_),
    .X(net249));
 sg13g2_mux2_1 \register_file_i/_5304_  (.A0(\register_file_i/rf_reg_845_ ),
    .A1(\register_file_i/rf_reg_877_ ),
    .S(net480),
    .X(\register_file_i/_2220_ ));
 sg13g2_mux2_1 \register_file_i/_5305_  (.A0(\register_file_i/rf_reg_781_ ),
    .A1(\register_file_i/rf_reg_813_ ),
    .S(net486),
    .X(\register_file_i/_2221_ ));
 sg13g2_buf_4 fanout248 (.X(net248),
    .A(net249));
 sg13g2_a22oi_1 \register_file_i/_5307_  (.Y(\register_file_i/_2223_ ),
    .B1(\register_file_i/_2221_ ),
    .B2(net1733),
    .A2(\register_file_i/_2220_ ),
    .A1(net1744));
 sg13g2_buf_2 fanout247 (.A(_05079_),
    .X(net247));
 sg13g2_a21o_1 \register_file_i/_5309_  (.A2(\register_file_i/_2223_ ),
    .A1(\register_file_i/_2218_ ),
    .B1(net1916),
    .X(\register_file_i/_2225_ ));
 sg13g2_buf_2 fanout246 (.A(_05079_),
    .X(net246));
 sg13g2_buf_1 fanout245 (.A(_05556_),
    .X(net245));
 sg13g2_buf_4 fanout244 (.X(net244),
    .A(net245));
 sg13g2_mux2_1 \register_file_i/_5313_  (.A0(\register_file_i/rf_reg_45_ ),
    .A1(\register_file_i/rf_reg_109_ ),
    .S(net451),
    .X(\register_file_i/_2229_ ));
 sg13g2_a22oi_1 \register_file_i/_5314_  (.Y(\register_file_i/_2230_ ),
    .B1(\register_file_i/_2229_ ),
    .B2(net514),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_77_ ));
 sg13g2_mux2_1 \register_file_i/_5315_  (.A0(\register_file_i/rf_reg_205_ ),
    .A1(\register_file_i/rf_reg_237_ ),
    .S(net490),
    .X(\register_file_i/_2231_ ));
 sg13g2_mux2_1 \register_file_i/_5316_  (.A0(\register_file_i/rf_reg_141_ ),
    .A1(\register_file_i/rf_reg_173_ ),
    .S(net493),
    .X(\register_file_i/_2232_ ));
 sg13g2_a22oi_1 \register_file_i/_5317_  (.Y(\register_file_i/_2233_ ),
    .B1(\register_file_i/_2232_ ),
    .B2(net1784),
    .A2(\register_file_i/_2231_ ),
    .A1(net1767));
 sg13g2_o21ai_1 \register_file_i/_5318_  (.B1(\register_file_i/_2233_ ),
    .Y(\register_file_i/_2234_ ),
    .A1(net445),
    .A2(\register_file_i/_2230_ ));
 sg13g2_nand2_1 \register_file_i/_5319_  (.Y(\register_file_i/_2235_ ),
    .A(net1911),
    .B(\register_file_i/_2234_ ));
 sg13g2_buf_2 fanout243 (.A(net245),
    .X(net243));
 sg13g2_mux4_1 \register_file_i/_5321_  (.S0(net495),
    .A0(\register_file_i/rf_reg_525_ ),
    .A1(\register_file_i/rf_reg_557_ ),
    .A2(\register_file_i/rf_reg_589_ ),
    .A3(\register_file_i/rf_reg_621_ ),
    .S1(net458),
    .X(\register_file_i/_2237_ ));
 sg13g2_mux4_1 \register_file_i/_5322_  (.S0(net487),
    .A0(\register_file_i/rf_reg_653_ ),
    .A1(\register_file_i/rf_reg_685_ ),
    .A2(\register_file_i/rf_reg_717_ ),
    .A3(\register_file_i/rf_reg_749_ ),
    .S1(net456),
    .X(\register_file_i/_2238_ ));
 sg13g2_buf_4 fanout242 (.X(net242),
    .A(net245));
 sg13g2_mux2_1 \register_file_i/_5324_  (.A0(\register_file_i/rf_reg_397_ ),
    .A1(\register_file_i/rf_reg_429_ ),
    .S(net482),
    .X(\register_file_i/_2240_ ));
 sg13g2_mux2_1 \register_file_i/_5325_  (.A0(\register_file_i/rf_reg_461_ ),
    .A1(\register_file_i/rf_reg_493_ ),
    .S(net488),
    .X(\register_file_i/_2241_ ));
 sg13g2_a22oi_1 \register_file_i/_5326_  (.Y(\register_file_i/_2242_ ),
    .B1(\register_file_i/_2241_ ),
    .B2(net1755),
    .A2(\register_file_i/_2240_ ),
    .A1(net1772));
 sg13g2_mux2_1 \register_file_i/_5327_  (.A0(\register_file_i/rf_reg_333_ ),
    .A1(\register_file_i/rf_reg_365_ ),
    .S(net494),
    .X(\register_file_i/_2243_ ));
 sg13g2_mux2_1 \register_file_i/_5328_  (.A0(\register_file_i/rf_reg_269_ ),
    .A1(\register_file_i/rf_reg_301_ ),
    .S(net484),
    .X(\register_file_i/_2244_ ));
 sg13g2_a22oi_1 \register_file_i/_5329_  (.Y(\register_file_i/_2245_ ),
    .B1(\register_file_i/_2244_ ),
    .B2(net1732),
    .A2(\register_file_i/_2243_ ),
    .A1(net1743));
 sg13g2_a21oi_1 \register_file_i/_5330_  (.A1(\register_file_i/_2242_ ),
    .A2(\register_file_i/_2245_ ),
    .Y(\register_file_i/_2246_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5331_  (.B2(net1682),
    .C1(\register_file_i/_2246_ ),
    .B1(\register_file_i/_2238_ ),
    .A1(net1724),
    .Y(\register_file_i/_2247_ ),
    .A2(\register_file_i/_2237_ ));
 sg13g2_nand3_1 \register_file_i/_5332_  (.B(\register_file_i/_2235_ ),
    .C(\register_file_i/_2247_ ),
    .A(\register_file_i/_2225_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_13_ ));
 sg13g2_mux2_1 \register_file_i/_5333_  (.A0(\register_file_i/rf_reg_908_ ),
    .A1(\register_file_i/rf_reg_940_ ),
    .S(net483),
    .X(\register_file_i/_2248_ ));
 sg13g2_mux2_1 \register_file_i/_5334_  (.A0(\register_file_i/rf_reg_972_ ),
    .A1(\register_file_i/rf_reg_1004_ ),
    .S(net491),
    .X(\register_file_i/_2249_ ));
 sg13g2_a22oi_1 \register_file_i/_5335_  (.Y(\register_file_i/_2250_ ),
    .B1(\register_file_i/_2249_ ),
    .B2(net1760),
    .A2(\register_file_i/_2248_ ),
    .A1(net1778));
 sg13g2_buf_2 fanout241 (.A(_02086_),
    .X(net241));
 sg13g2_mux2_1 \register_file_i/_5337_  (.A0(\register_file_i/rf_reg_844_ ),
    .A1(\register_file_i/rf_reg_876_ ),
    .S(net497),
    .X(\register_file_i/_2252_ ));
 sg13g2_mux2_1 \register_file_i/_5338_  (.A0(\register_file_i/rf_reg_780_ ),
    .A1(\register_file_i/rf_reg_812_ ),
    .S(net486),
    .X(\register_file_i/_2253_ ));
 sg13g2_a22oi_1 \register_file_i/_5339_  (.Y(\register_file_i/_2254_ ),
    .B1(\register_file_i/_2253_ ),
    .B2(net1736),
    .A2(\register_file_i/_2252_ ),
    .A1(net1747));
 sg13g2_a21o_1 \register_file_i/_5340_  (.A2(\register_file_i/_2254_ ),
    .A1(\register_file_i/_2250_ ),
    .B1(net1915),
    .X(\register_file_i/_2255_ ));
 sg13g2_mux2_1 \register_file_i/_5341_  (.A0(\register_file_i/rf_reg_44_ ),
    .A1(\register_file_i/rf_reg_108_ ),
    .S(net451),
    .X(\register_file_i/_2256_ ));
 sg13g2_buf_2 fanout240 (.A(_02638_),
    .X(net240));
 sg13g2_a22oi_1 \register_file_i/_5343_  (.Y(\register_file_i/_2258_ ),
    .B1(\register_file_i/_2256_ ),
    .B2(net516),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_76_ ));
 sg13g2_mux2_1 \register_file_i/_5344_  (.A0(\register_file_i/rf_reg_204_ ),
    .A1(\register_file_i/rf_reg_236_ ),
    .S(net490),
    .X(\register_file_i/_2259_ ));
 sg13g2_mux2_1 \register_file_i/_5345_  (.A0(\register_file_i/rf_reg_140_ ),
    .A1(\register_file_i/rf_reg_172_ ),
    .S(net493),
    .X(\register_file_i/_2260_ ));
 sg13g2_a22oi_1 \register_file_i/_5346_  (.Y(\register_file_i/_2261_ ),
    .B1(\register_file_i/_2260_ ),
    .B2(net1779),
    .A2(\register_file_i/_2259_ ),
    .A1(net1765));
 sg13g2_o21ai_1 \register_file_i/_5347_  (.B1(\register_file_i/_2261_ ),
    .Y(\register_file_i/_2262_ ),
    .A1(net445),
    .A2(\register_file_i/_2258_ ));
 sg13g2_nand2_1 \register_file_i/_5348_  (.Y(\register_file_i/_2263_ ),
    .A(net1908),
    .B(\register_file_i/_2262_ ));
 sg13g2_mux4_1 \register_file_i/_5349_  (.S0(net495),
    .A0(\register_file_i/rf_reg_524_ ),
    .A1(\register_file_i/rf_reg_556_ ),
    .A2(\register_file_i/rf_reg_588_ ),
    .A3(\register_file_i/rf_reg_620_ ),
    .S1(net458),
    .X(\register_file_i/_2264_ ));
 sg13g2_buf_1 fanout239 (.A(_03323_),
    .X(net239));
 sg13g2_mux4_1 \register_file_i/_5351_  (.S0(net487),
    .A0(\register_file_i/rf_reg_652_ ),
    .A1(\register_file_i/rf_reg_684_ ),
    .A2(\register_file_i/rf_reg_716_ ),
    .A3(\register_file_i/rf_reg_748_ ),
    .S1(net460),
    .X(\register_file_i/_2266_ ));
 sg13g2_buf_2 fanout238 (.A(_03323_),
    .X(net238));
 sg13g2_mux2_1 \register_file_i/_5353_  (.A0(\register_file_i/rf_reg_396_ ),
    .A1(\register_file_i/rf_reg_428_ ),
    .S(net498),
    .X(\register_file_i/_2268_ ));
 sg13g2_mux2_1 \register_file_i/_5354_  (.A0(\register_file_i/rf_reg_460_ ),
    .A1(\register_file_i/rf_reg_492_ ),
    .S(net488),
    .X(\register_file_i/_2269_ ));
 sg13g2_a22oi_1 \register_file_i/_5355_  (.Y(\register_file_i/_2270_ ),
    .B1(\register_file_i/_2269_ ),
    .B2(net1752),
    .A2(\register_file_i/_2268_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5356_  (.A0(\register_file_i/rf_reg_332_ ),
    .A1(\register_file_i/rf_reg_364_ ),
    .S(net494),
    .X(\register_file_i/_2271_ ));
 sg13g2_mux2_1 \register_file_i/_5357_  (.A0(\register_file_i/rf_reg_268_ ),
    .A1(\register_file_i/rf_reg_300_ ),
    .S(net484),
    .X(\register_file_i/_2272_ ));
 sg13g2_a22oi_1 \register_file_i/_5358_  (.Y(\register_file_i/_2273_ ),
    .B1(\register_file_i/_2272_ ),
    .B2(net1730),
    .A2(\register_file_i/_2271_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5359_  (.A1(\register_file_i/_2270_ ),
    .A2(\register_file_i/_2273_ ),
    .Y(\register_file_i/_2274_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5360_  (.B2(net1682),
    .C1(\register_file_i/_2274_ ),
    .B1(\register_file_i/_2266_ ),
    .A1(net1724),
    .Y(\register_file_i/_2275_ ),
    .A2(\register_file_i/_2264_ ));
 sg13g2_nand3_1 \register_file_i/_5361_  (.B(\register_file_i/_2263_ ),
    .C(\register_file_i/_2275_ ),
    .A(\register_file_i/_2255_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_12_ ));
 sg13g2_mux2_1 \register_file_i/_5362_  (.A0(\register_file_i/rf_reg_925_ ),
    .A1(\register_file_i/rf_reg_957_ ),
    .S(net483),
    .X(\register_file_i/_2276_ ));
 sg13g2_mux2_1 \register_file_i/_5363_  (.A0(\register_file_i/rf_reg_989_ ),
    .A1(\register_file_i/rf_reg_1021_ ),
    .S(net491),
    .X(\register_file_i/_2277_ ));
 sg13g2_a22oi_1 \register_file_i/_5364_  (.Y(\register_file_i/_2278_ ),
    .B1(\register_file_i/_2277_ ),
    .B2(net1764),
    .A2(\register_file_i/_2276_ ),
    .A1(net1782));
 sg13g2_mux2_1 \register_file_i/_5365_  (.A0(\register_file_i/rf_reg_861_ ),
    .A1(\register_file_i/rf_reg_893_ ),
    .S(net496),
    .X(\register_file_i/_2279_ ));
 sg13g2_mux2_1 \register_file_i/_5366_  (.A0(\register_file_i/rf_reg_797_ ),
    .A1(\register_file_i/rf_reg_829_ ),
    .S(net486),
    .X(\register_file_i/_2280_ ));
 sg13g2_a22oi_1 \register_file_i/_5367_  (.Y(\register_file_i/_2281_ ),
    .B1(\register_file_i/_2280_ ),
    .B2(net1737),
    .A2(\register_file_i/_2279_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5368_  (.A2(\register_file_i/_2281_ ),
    .A1(\register_file_i/_2278_ ),
    .B1(net1914),
    .X(\register_file_i/_2282_ ));
 sg13g2_mux2_1 \register_file_i/_5369_  (.A0(\register_file_i/rf_reg_61_ ),
    .A1(\register_file_i/rf_reg_125_ ),
    .S(net451),
    .X(\register_file_i/_2283_ ));
 sg13g2_a22oi_1 \register_file_i/_5370_  (.Y(\register_file_i/_2284_ ),
    .B1(\register_file_i/_2283_ ),
    .B2(net516),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_93_ ));
 sg13g2_mux2_1 \register_file_i/_5371_  (.A0(\register_file_i/rf_reg_221_ ),
    .A1(\register_file_i/rf_reg_253_ ),
    .S(net490),
    .X(\register_file_i/_2285_ ));
 sg13g2_mux2_1 \register_file_i/_5372_  (.A0(\register_file_i/rf_reg_157_ ),
    .A1(\register_file_i/rf_reg_189_ ),
    .S(net492),
    .X(\register_file_i/_2286_ ));
 sg13g2_a22oi_1 \register_file_i/_5373_  (.Y(\register_file_i/_2287_ ),
    .B1(\register_file_i/_2286_ ),
    .B2(net1779),
    .A2(\register_file_i/_2285_ ),
    .A1(net1761));
 sg13g2_o21ai_1 \register_file_i/_5374_  (.B1(\register_file_i/_2287_ ),
    .Y(\register_file_i/_2288_ ),
    .A1(net445),
    .A2(\register_file_i/_2284_ ));
 sg13g2_nand2_1 \register_file_i/_5375_  (.Y(\register_file_i/_2289_ ),
    .A(net1907),
    .B(\register_file_i/_2288_ ));
 sg13g2_mux4_1 \register_file_i/_5376_  (.S0(net495),
    .A0(\register_file_i/rf_reg_541_ ),
    .A1(\register_file_i/rf_reg_573_ ),
    .A2(\register_file_i/rf_reg_605_ ),
    .A3(\register_file_i/rf_reg_637_ ),
    .S1(net458),
    .X(\register_file_i/_2290_ ));
 sg13g2_mux4_1 \register_file_i/_5377_  (.S0(net487),
    .A0(\register_file_i/rf_reg_669_ ),
    .A1(\register_file_i/rf_reg_701_ ),
    .A2(\register_file_i/rf_reg_733_ ),
    .A3(\register_file_i/rf_reg_765_ ),
    .S1(net460),
    .X(\register_file_i/_2291_ ));
 sg13g2_buf_2 fanout237 (.A(_03323_),
    .X(net237));
 sg13g2_mux2_1 \register_file_i/_5379_  (.A0(\register_file_i/rf_reg_413_ ),
    .A1(\register_file_i/rf_reg_445_ ),
    .S(net498),
    .X(\register_file_i/_2293_ ));
 sg13g2_mux2_1 \register_file_i/_5380_  (.A0(\register_file_i/rf_reg_477_ ),
    .A1(\register_file_i/rf_reg_509_ ),
    .S(net488),
    .X(\register_file_i/_2294_ ));
 sg13g2_a22oi_1 \register_file_i/_5381_  (.Y(\register_file_i/_2295_ ),
    .B1(\register_file_i/_2294_ ),
    .B2(net1752),
    .A2(\register_file_i/_2293_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5382_  (.A0(\register_file_i/rf_reg_349_ ),
    .A1(\register_file_i/rf_reg_381_ ),
    .S(net494),
    .X(\register_file_i/_2296_ ));
 sg13g2_mux2_1 \register_file_i/_5383_  (.A0(\register_file_i/rf_reg_285_ ),
    .A1(\register_file_i/rf_reg_317_ ),
    .S(net484),
    .X(\register_file_i/_2297_ ));
 sg13g2_a22oi_1 \register_file_i/_5384_  (.Y(\register_file_i/_2298_ ),
    .B1(\register_file_i/_2297_ ),
    .B2(net1730),
    .A2(\register_file_i/_2296_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5385_  (.A1(\register_file_i/_2295_ ),
    .A2(\register_file_i/_2298_ ),
    .Y(\register_file_i/_2299_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5386_  (.B2(net1682),
    .C1(\register_file_i/_2299_ ),
    .B1(\register_file_i/_2291_ ),
    .A1(net1724),
    .Y(\register_file_i/_2300_ ),
    .A2(\register_file_i/_2290_ ));
 sg13g2_nand3_1 \register_file_i/_5387_  (.B(\register_file_i/_2289_ ),
    .C(\register_file_i/_2300_ ),
    .A(\register_file_i/_2282_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_29_ ));
 sg13g2_buf_4 fanout236 (.X(net236),
    .A(_03323_));
 sg13g2_mux2_1 \register_file_i/_5389_  (.A0(\register_file_i/rf_reg_907_ ),
    .A1(\register_file_i/rf_reg_939_ ),
    .S(net499),
    .X(\register_file_i/_2302_ ));
 sg13g2_mux2_1 \register_file_i/_5390_  (.A0(\register_file_i/rf_reg_971_ ),
    .A1(\register_file_i/rf_reg_1003_ ),
    .S(net491),
    .X(\register_file_i/_2303_ ));
 sg13g2_a22oi_1 \register_file_i/_5391_  (.Y(\register_file_i/_2304_ ),
    .B1(\register_file_i/_2303_ ),
    .B2(net1763),
    .A2(\register_file_i/_2302_ ),
    .A1(net1780));
 sg13g2_mux2_1 \register_file_i/_5392_  (.A0(\register_file_i/rf_reg_843_ ),
    .A1(\register_file_i/rf_reg_875_ ),
    .S(net496),
    .X(\register_file_i/_2305_ ));
 sg13g2_mux2_1 \register_file_i/_5393_  (.A0(\register_file_i/rf_reg_779_ ),
    .A1(\register_file_i/rf_reg_811_ ),
    .S(net486),
    .X(\register_file_i/_2306_ ));
 sg13g2_a22oi_1 \register_file_i/_5394_  (.Y(\register_file_i/_2307_ ),
    .B1(\register_file_i/_2306_ ),
    .B2(net1737),
    .A2(\register_file_i/_2305_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5395_  (.A2(\register_file_i/_2307_ ),
    .A1(\register_file_i/_2304_ ),
    .B1(net1913),
    .X(\register_file_i/_2308_ ));
 sg13g2_mux2_1 \register_file_i/_5396_  (.A0(\register_file_i/rf_reg_43_ ),
    .A1(\register_file_i/rf_reg_107_ ),
    .S(net451),
    .X(\register_file_i/_2309_ ));
 sg13g2_a22oi_1 \register_file_i/_5397_  (.Y(\register_file_i/_2310_ ),
    .B1(\register_file_i/_2309_ ),
    .B2(net516),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_75_ ));
 sg13g2_mux2_1 \register_file_i/_5398_  (.A0(\register_file_i/rf_reg_203_ ),
    .A1(\register_file_i/rf_reg_235_ ),
    .S(net490),
    .X(\register_file_i/_2311_ ));
 sg13g2_mux2_1 \register_file_i/_5399_  (.A0(\register_file_i/rf_reg_139_ ),
    .A1(\register_file_i/rf_reg_171_ ),
    .S(net492),
    .X(\register_file_i/_2312_ ));
 sg13g2_a22oi_1 \register_file_i/_5400_  (.Y(\register_file_i/_2313_ ),
    .B1(\register_file_i/_2312_ ),
    .B2(net1780),
    .A2(\register_file_i/_2311_ ),
    .A1(net1760));
 sg13g2_o21ai_1 \register_file_i/_5401_  (.B1(\register_file_i/_2313_ ),
    .Y(\register_file_i/_2314_ ),
    .A1(net445),
    .A2(\register_file_i/_2310_ ));
 sg13g2_nand2_1 \register_file_i/_5402_  (.Y(\register_file_i/_2315_ ),
    .A(net1907),
    .B(\register_file_i/_2314_ ));
 sg13g2_mux4_1 \register_file_i/_5403_  (.S0(net495),
    .A0(\register_file_i/rf_reg_523_ ),
    .A1(\register_file_i/rf_reg_555_ ),
    .A2(\register_file_i/rf_reg_587_ ),
    .A3(\register_file_i/rf_reg_619_ ),
    .S1(net458),
    .X(\register_file_i/_2316_ ));
 sg13g2_mux4_1 \register_file_i/_5404_  (.S0(net487),
    .A0(\register_file_i/rf_reg_651_ ),
    .A1(\register_file_i/rf_reg_683_ ),
    .A2(\register_file_i/rf_reg_715_ ),
    .A3(\register_file_i/rf_reg_747_ ),
    .S1(net460),
    .X(\register_file_i/_2317_ ));
 sg13g2_mux2_1 \register_file_i/_5405_  (.A0(\register_file_i/rf_reg_395_ ),
    .A1(\register_file_i/rf_reg_427_ ),
    .S(net498),
    .X(\register_file_i/_2318_ ));
 sg13g2_mux2_1 \register_file_i/_5406_  (.A0(\register_file_i/rf_reg_459_ ),
    .A1(\register_file_i/rf_reg_491_ ),
    .S(net488),
    .X(\register_file_i/_2319_ ));
 sg13g2_a22oi_1 \register_file_i/_5407_  (.Y(\register_file_i/_2320_ ),
    .B1(\register_file_i/_2319_ ),
    .B2(net1752),
    .A2(\register_file_i/_2318_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5408_  (.A0(\register_file_i/rf_reg_331_ ),
    .A1(\register_file_i/rf_reg_363_ ),
    .S(net494),
    .X(\register_file_i/_2321_ ));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(_03323_));
 sg13g2_mux2_1 \register_file_i/_5410_  (.A0(\register_file_i/rf_reg_267_ ),
    .A1(\register_file_i/rf_reg_299_ ),
    .S(net500),
    .X(\register_file_i/_2323_ ));
 sg13g2_a22oi_1 \register_file_i/_5411_  (.Y(\register_file_i/_2324_ ),
    .B1(\register_file_i/_2323_ ),
    .B2(net1730),
    .A2(\register_file_i/_2321_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5412_  (.A1(\register_file_i/_2320_ ),
    .A2(\register_file_i/_2324_ ),
    .Y(\register_file_i/_2325_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5413_  (.B2(net1682),
    .C1(\register_file_i/_2325_ ),
    .B1(\register_file_i/_2317_ ),
    .A1(net1724),
    .Y(\register_file_i/_2326_ ),
    .A2(\register_file_i/_2316_ ));
 sg13g2_nand3_1 \register_file_i/_5414_  (.B(\register_file_i/_2315_ ),
    .C(\register_file_i/_2326_ ),
    .A(\register_file_i/_2308_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ));
 sg13g2_mux2_1 \register_file_i/_5415_  (.A0(\register_file_i/rf_reg_906_ ),
    .A1(\register_file_i/rf_reg_938_ ),
    .S(net499),
    .X(\register_file_i/_2327_ ));
 sg13g2_mux2_1 \register_file_i/_5416_  (.A0(\register_file_i/rf_reg_970_ ),
    .A1(\register_file_i/rf_reg_1002_ ),
    .S(net491),
    .X(\register_file_i/_2328_ ));
 sg13g2_a22oi_1 \register_file_i/_5417_  (.Y(\register_file_i/_2329_ ),
    .B1(\register_file_i/_2328_ ),
    .B2(net1760),
    .A2(\register_file_i/_2327_ ),
    .A1(net1779));
 sg13g2_mux2_1 \register_file_i/_5418_  (.A0(\register_file_i/rf_reg_842_ ),
    .A1(\register_file_i/rf_reg_874_ ),
    .S(net496),
    .X(\register_file_i/_2330_ ));
 sg13g2_mux2_1 \register_file_i/_5419_  (.A0(\register_file_i/rf_reg_778_ ),
    .A1(\register_file_i/rf_reg_810_ ),
    .S(net485),
    .X(\register_file_i/_2331_ ));
 sg13g2_a22oi_1 \register_file_i/_5420_  (.Y(\register_file_i/_2332_ ),
    .B1(\register_file_i/_2331_ ),
    .B2(net1736),
    .A2(\register_file_i/_2330_ ),
    .A1(net1747));
 sg13g2_a21o_1 \register_file_i/_5421_  (.A2(\register_file_i/_2332_ ),
    .A1(\register_file_i/_2329_ ),
    .B1(net1913),
    .X(\register_file_i/_2333_ ));
 sg13g2_mux2_1 \register_file_i/_5422_  (.A0(\register_file_i/rf_reg_42_ ),
    .A1(\register_file_i/rf_reg_106_ ),
    .S(net451),
    .X(\register_file_i/_2334_ ));
 sg13g2_a22oi_1 \register_file_i/_5423_  (.Y(\register_file_i/_2335_ ),
    .B1(\register_file_i/_2334_ ),
    .B2(net516),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_74_ ));
 sg13g2_buf_4 fanout234 (.X(net234),
    .A(_03905_));
 sg13g2_mux2_1 \register_file_i/_5425_  (.A0(\register_file_i/rf_reg_202_ ),
    .A1(\register_file_i/rf_reg_234_ ),
    .S(net489),
    .X(\register_file_i/_2337_ ));
 sg13g2_mux2_1 \register_file_i/_5426_  (.A0(\register_file_i/rf_reg_138_ ),
    .A1(\register_file_i/rf_reg_170_ ),
    .S(net492),
    .X(\register_file_i/_2338_ ));
 sg13g2_a22oi_1 \register_file_i/_5427_  (.Y(\register_file_i/_2339_ ),
    .B1(\register_file_i/_2338_ ),
    .B2(net1778),
    .A2(\register_file_i/_2337_ ),
    .A1(net1761));
 sg13g2_o21ai_1 \register_file_i/_5428_  (.B1(\register_file_i/_2339_ ),
    .Y(\register_file_i/_2340_ ),
    .A1(net445),
    .A2(\register_file_i/_2335_ ));
 sg13g2_nand2_1 \register_file_i/_5429_  (.Y(\register_file_i/_2341_ ),
    .A(net1908),
    .B(\register_file_i/_2340_ ));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(_04046_));
 sg13g2_mux4_1 \register_file_i/_5431_  (.S0(net495),
    .A0(\register_file_i/rf_reg_522_ ),
    .A1(\register_file_i/rf_reg_554_ ),
    .A2(\register_file_i/rf_reg_586_ ),
    .A3(\register_file_i/rf_reg_618_ ),
    .S1(net461),
    .X(\register_file_i/_2343_ ));
 sg13g2_mux4_1 \register_file_i/_5432_  (.S0(net487),
    .A0(\register_file_i/rf_reg_650_ ),
    .A1(\register_file_i/rf_reg_682_ ),
    .A2(\register_file_i/rf_reg_714_ ),
    .A3(\register_file_i/rf_reg_746_ ),
    .S1(net460),
    .X(\register_file_i/_2344_ ));
 sg13g2_mux2_1 \register_file_i/_5433_  (.A0(\register_file_i/rf_reg_394_ ),
    .A1(\register_file_i/rf_reg_426_ ),
    .S(net497),
    .X(\register_file_i/_2345_ ));
 sg13g2_mux2_1 \register_file_i/_5434_  (.A0(\register_file_i/rf_reg_458_ ),
    .A1(\register_file_i/rf_reg_490_ ),
    .S(net488),
    .X(\register_file_i/_2346_ ));
 sg13g2_a22oi_1 \register_file_i/_5435_  (.Y(\register_file_i/_2347_ ),
    .B1(\register_file_i/_2346_ ),
    .B2(net1752),
    .A2(\register_file_i/_2345_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5436_  (.A0(\register_file_i/rf_reg_330_ ),
    .A1(\register_file_i/rf_reg_362_ ),
    .S(net493),
    .X(\register_file_i/_2348_ ));
 sg13g2_mux2_1 \register_file_i/_5437_  (.A0(\register_file_i/rf_reg_266_ ),
    .A1(\register_file_i/rf_reg_298_ ),
    .S(net500),
    .X(\register_file_i/_2349_ ));
 sg13g2_a22oi_1 \register_file_i/_5438_  (.Y(\register_file_i/_2350_ ),
    .B1(\register_file_i/_2349_ ),
    .B2(net1730),
    .A2(\register_file_i/_2348_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5439_  (.A1(\register_file_i/_2347_ ),
    .A2(\register_file_i/_2350_ ),
    .Y(\register_file_i/_2351_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5440_  (.B2(net1682),
    .C1(\register_file_i/_2351_ ),
    .B1(\register_file_i/_2344_ ),
    .A1(net1724),
    .Y(\register_file_i/_2352_ ),
    .A2(\register_file_i/_2343_ ));
 sg13g2_nand3_1 \register_file_i/_5441_  (.B(\register_file_i/_2341_ ),
    .C(\register_file_i/_2352_ ),
    .A(\register_file_i/_2333_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_10_ ));
 sg13g2_mux2_1 \register_file_i/_5442_  (.A0(\register_file_i/rf_reg_905_ ),
    .A1(\register_file_i/rf_reg_937_ ),
    .S(net499),
    .X(\register_file_i/_2353_ ));
 sg13g2_mux2_1 \register_file_i/_5443_  (.A0(\register_file_i/rf_reg_969_ ),
    .A1(\register_file_i/rf_reg_1001_ ),
    .S(net491),
    .X(\register_file_i/_2354_ ));
 sg13g2_a22oi_1 \register_file_i/_5444_  (.Y(\register_file_i/_2355_ ),
    .B1(\register_file_i/_2354_ ),
    .B2(net1760),
    .A2(\register_file_i/_2353_ ),
    .A1(net1778));
 sg13g2_mux2_1 \register_file_i/_5445_  (.A0(\register_file_i/rf_reg_841_ ),
    .A1(\register_file_i/rf_reg_873_ ),
    .S(net496),
    .X(\register_file_i/_2356_ ));
 sg13g2_buf_2 fanout232 (.A(_04046_),
    .X(net232));
 sg13g2_mux2_1 \register_file_i/_5447_  (.A0(\register_file_i/rf_reg_777_ ),
    .A1(\register_file_i/rf_reg_809_ ),
    .S(net502),
    .X(\register_file_i/_2358_ ));
 sg13g2_a22oi_1 \register_file_i/_5448_  (.Y(\register_file_i/_2359_ ),
    .B1(\register_file_i/_2358_ ),
    .B2(net1737),
    .A2(\register_file_i/_2356_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5449_  (.A2(\register_file_i/_2359_ ),
    .A1(\register_file_i/_2355_ ),
    .B1(net1913),
    .X(\register_file_i/_2360_ ));
 sg13g2_mux2_1 \register_file_i/_5450_  (.A0(\register_file_i/rf_reg_41_ ),
    .A1(\register_file_i/rf_reg_105_ ),
    .S(net450),
    .X(\register_file_i/_2361_ ));
 sg13g2_a22oi_1 \register_file_i/_5451_  (.Y(\register_file_i/_2362_ ),
    .B1(\register_file_i/_2361_ ),
    .B2(net516),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_73_ ));
 sg13g2_mux2_1 \register_file_i/_5452_  (.A0(\register_file_i/rf_reg_201_ ),
    .A1(\register_file_i/rf_reg_233_ ),
    .S(net489),
    .X(\register_file_i/_2363_ ));
 sg13g2_mux2_1 \register_file_i/_5453_  (.A0(\register_file_i/rf_reg_137_ ),
    .A1(\register_file_i/rf_reg_169_ ),
    .S(net492),
    .X(\register_file_i/_2364_ ));
 sg13g2_a22oi_1 \register_file_i/_5454_  (.Y(\register_file_i/_2365_ ),
    .B1(\register_file_i/_2364_ ),
    .B2(net1778),
    .A2(\register_file_i/_2363_ ),
    .A1(net1761));
 sg13g2_o21ai_1 \register_file_i/_5455_  (.B1(\register_file_i/_2365_ ),
    .Y(\register_file_i/_2366_ ),
    .A1(net445),
    .A2(\register_file_i/_2362_ ));
 sg13g2_nand2_1 \register_file_i/_5456_  (.Y(\register_file_i/_2367_ ),
    .A(net1908),
    .B(\register_file_i/_2366_ ));
 sg13g2_mux4_1 \register_file_i/_5457_  (.S0(net495),
    .A0(\register_file_i/rf_reg_521_ ),
    .A1(\register_file_i/rf_reg_553_ ),
    .A2(\register_file_i/rf_reg_585_ ),
    .A3(\register_file_i/rf_reg_617_ ),
    .S1(net461),
    .X(\register_file_i/_2368_ ));
 sg13g2_buf_2 fanout231 (.A(_04046_),
    .X(net231));
 sg13g2_mux4_1 \register_file_i/_5459_  (.S0(net503),
    .A0(\register_file_i/rf_reg_649_ ),
    .A1(\register_file_i/rf_reg_681_ ),
    .A2(\register_file_i/rf_reg_713_ ),
    .A3(\register_file_i/rf_reg_745_ ),
    .S1(net459),
    .X(\register_file_i/_2370_ ));
 sg13g2_mux2_1 \register_file_i/_5460_  (.A0(\register_file_i/rf_reg_393_ ),
    .A1(\register_file_i/rf_reg_425_ ),
    .S(net497),
    .X(\register_file_i/_2371_ ));
 sg13g2_buf_4 fanout230 (.X(net230),
    .A(_04046_));
 sg13g2_mux2_1 \register_file_i/_5462_  (.A0(\register_file_i/rf_reg_457_ ),
    .A1(\register_file_i/rf_reg_489_ ),
    .S(net504),
    .X(\register_file_i/_2373_ ));
 sg13g2_a22oi_1 \register_file_i/_5463_  (.Y(\register_file_i/_2374_ ),
    .B1(\register_file_i/_2373_ ),
    .B2(net1752),
    .A2(\register_file_i/_2371_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5464_  (.A0(\register_file_i/rf_reg_329_ ),
    .A1(\register_file_i/rf_reg_361_ ),
    .S(net493),
    .X(\register_file_i/_2375_ ));
 sg13g2_mux2_1 \register_file_i/_5465_  (.A0(\register_file_i/rf_reg_265_ ),
    .A1(\register_file_i/rf_reg_297_ ),
    .S(net500),
    .X(\register_file_i/_2376_ ));
 sg13g2_a22oi_1 \register_file_i/_5466_  (.Y(\register_file_i/_2377_ ),
    .B1(\register_file_i/_2376_ ),
    .B2(net1730),
    .A2(\register_file_i/_2375_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5467_  (.A1(\register_file_i/_2374_ ),
    .A2(\register_file_i/_2377_ ),
    .Y(\register_file_i/_2378_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5468_  (.B2(net1682),
    .C1(\register_file_i/_2378_ ),
    .B1(\register_file_i/_2370_ ),
    .A1(net1724),
    .Y(\register_file_i/_2379_ ),
    .A2(\register_file_i/_2368_ ));
 sg13g2_nand3_1 \register_file_i/_5469_  (.B(\register_file_i/_2367_ ),
    .C(\register_file_i/_2379_ ),
    .A(\register_file_i/_2360_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_9_ ));
 sg13g2_mux2_1 \register_file_i/_5470_  (.A0(\register_file_i/rf_reg_904_ ),
    .A1(\register_file_i/rf_reg_936_ ),
    .S(net499),
    .X(\register_file_i/_2380_ ));
 sg13g2_mux2_1 \register_file_i/_5471_  (.A0(\register_file_i/rf_reg_968_ ),
    .A1(\register_file_i/rf_reg_1000_ ),
    .S(net491),
    .X(\register_file_i/_2381_ ));
 sg13g2_a22oi_1 \register_file_i/_5472_  (.Y(\register_file_i/_2382_ ),
    .B1(\register_file_i/_2381_ ),
    .B2(net1762),
    .A2(\register_file_i/_2380_ ),
    .A1(net1781));
 sg13g2_mux2_1 \register_file_i/_5473_  (.A0(\register_file_i/rf_reg_840_ ),
    .A1(\register_file_i/rf_reg_872_ ),
    .S(net496),
    .X(\register_file_i/_2383_ ));
 sg13g2_mux2_1 \register_file_i/_5474_  (.A0(\register_file_i/rf_reg_776_ ),
    .A1(\register_file_i/rf_reg_808_ ),
    .S(net501),
    .X(\register_file_i/_2384_ ));
 sg13g2_a22oi_1 \register_file_i/_5475_  (.Y(\register_file_i/_2385_ ),
    .B1(\register_file_i/_2384_ ),
    .B2(net1737),
    .A2(\register_file_i/_2383_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5476_  (.A2(\register_file_i/_2385_ ),
    .A1(\register_file_i/_2382_ ),
    .B1(net1913),
    .X(\register_file_i/_2386_ ));
 sg13g2_mux2_1 \register_file_i/_5477_  (.A0(\register_file_i/rf_reg_40_ ),
    .A1(\register_file_i/rf_reg_104_ ),
    .S(net450),
    .X(\register_file_i/_2387_ ));
 sg13g2_a22oi_1 \register_file_i/_5478_  (.Y(\register_file_i/_2388_ ),
    .B1(\register_file_i/_2387_ ),
    .B2(net515),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_72_ ));
 sg13g2_mux2_1 \register_file_i/_5479_  (.A0(\register_file_i/rf_reg_200_ ),
    .A1(\register_file_i/rf_reg_232_ ),
    .S(net489),
    .X(\register_file_i/_2389_ ));
 sg13g2_mux2_1 \register_file_i/_5480_  (.A0(\register_file_i/rf_reg_136_ ),
    .A1(\register_file_i/rf_reg_168_ ),
    .S(net492),
    .X(\register_file_i/_2390_ ));
 sg13g2_a22oi_1 \register_file_i/_5481_  (.Y(\register_file_i/_2391_ ),
    .B1(\register_file_i/_2390_ ),
    .B2(net1780),
    .A2(\register_file_i/_2389_ ),
    .A1(net1763));
 sg13g2_o21ai_1 \register_file_i/_5482_  (.B1(\register_file_i/_2391_ ),
    .Y(\register_file_i/_2392_ ),
    .A1(net444),
    .A2(\register_file_i/_2388_ ));
 sg13g2_nand2_1 \register_file_i/_5483_  (.Y(\register_file_i/_2393_ ),
    .A(net1907),
    .B(\register_file_i/_2392_ ));
 sg13g2_buf_1 fanout229 (.A(_04242_),
    .X(net229));
 sg13g2_mux4_1 \register_file_i/_5485_  (.S0(net495),
    .A0(\register_file_i/rf_reg_520_ ),
    .A1(\register_file_i/rf_reg_552_ ),
    .A2(\register_file_i/rf_reg_584_ ),
    .A3(\register_file_i/rf_reg_616_ ),
    .S1(net461),
    .X(\register_file_i/_2395_ ));
 sg13g2_mux4_1 \register_file_i/_5486_  (.S0(net503),
    .A0(\register_file_i/rf_reg_648_ ),
    .A1(\register_file_i/rf_reg_680_ ),
    .A2(\register_file_i/rf_reg_712_ ),
    .A3(\register_file_i/rf_reg_744_ ),
    .S1(net459),
    .X(\register_file_i/_2396_ ));
 sg13g2_mux2_1 \register_file_i/_5487_  (.A0(\register_file_i/rf_reg_392_ ),
    .A1(\register_file_i/rf_reg_424_ ),
    .S(net497),
    .X(\register_file_i/_2397_ ));
 sg13g2_mux2_1 \register_file_i/_5488_  (.A0(\register_file_i/rf_reg_456_ ),
    .A1(\register_file_i/rf_reg_488_ ),
    .S(net504),
    .X(\register_file_i/_2398_ ));
 sg13g2_a22oi_1 \register_file_i/_5489_  (.Y(\register_file_i/_2399_ ),
    .B1(\register_file_i/_2398_ ),
    .B2(net1753),
    .A2(\register_file_i/_2397_ ),
    .A1(net1777));
 sg13g2_mux2_1 \register_file_i/_5490_  (.A0(\register_file_i/rf_reg_328_ ),
    .A1(\register_file_i/rf_reg_360_ ),
    .S(net493),
    .X(\register_file_i/_2400_ ));
 sg13g2_mux2_1 \register_file_i/_5491_  (.A0(\register_file_i/rf_reg_264_ ),
    .A1(\register_file_i/rf_reg_296_ ),
    .S(net500),
    .X(\register_file_i/_2401_ ));
 sg13g2_a22oi_1 \register_file_i/_5492_  (.Y(\register_file_i/_2402_ ),
    .B1(\register_file_i/_2401_ ),
    .B2(net1731),
    .A2(\register_file_i/_2400_ ),
    .A1(net1742));
 sg13g2_buf_2 fanout228 (.A(net229),
    .X(net228));
 sg13g2_a21oi_1 \register_file_i/_5494_  (.A1(\register_file_i/_2399_ ),
    .A2(\register_file_i/_2402_ ),
    .Y(\register_file_i/_2404_ ),
    .B1(net1720));
 sg13g2_a221oi_1 \register_file_i/_5495_  (.B2(net1682),
    .C1(\register_file_i/_2404_ ),
    .B1(\register_file_i/_2396_ ),
    .A1(net1724),
    .Y(\register_file_i/_2405_ ),
    .A2(\register_file_i/_2395_ ));
 sg13g2_nand3_1 \register_file_i/_5496_  (.B(\register_file_i/_2393_ ),
    .C(\register_file_i/_2405_ ),
    .A(\register_file_i/_2386_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ));
 sg13g2_mux2_1 \register_file_i/_5497_  (.A0(\register_file_i/rf_reg_903_ ),
    .A1(\register_file_i/rf_reg_935_ ),
    .S(net499),
    .X(\register_file_i/_2406_ ));
 sg13g2_mux2_1 \register_file_i/_5498_  (.A0(\register_file_i/rf_reg_967_ ),
    .A1(\register_file_i/rf_reg_999_ ),
    .S(net490),
    .X(\register_file_i/_2407_ ));
 sg13g2_a22oi_1 \register_file_i/_5499_  (.Y(\register_file_i/_2408_ ),
    .B1(\register_file_i/_2407_ ),
    .B2(net1762),
    .A2(\register_file_i/_2406_ ),
    .A1(net1780));
 sg13g2_mux2_1 \register_file_i/_5500_  (.A0(\register_file_i/rf_reg_839_ ),
    .A1(\register_file_i/rf_reg_871_ ),
    .S(net496),
    .X(\register_file_i/_2409_ ));
 sg13g2_mux2_1 \register_file_i/_5501_  (.A0(\register_file_i/rf_reg_775_ ),
    .A1(\register_file_i/rf_reg_807_ ),
    .S(net501),
    .X(\register_file_i/_2410_ ));
 sg13g2_a22oi_1 \register_file_i/_5502_  (.Y(\register_file_i/_2411_ ),
    .B1(\register_file_i/_2410_ ),
    .B2(net1737),
    .A2(\register_file_i/_2409_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5503_  (.A2(\register_file_i/_2411_ ),
    .A1(\register_file_i/_2408_ ),
    .B1(net1913),
    .X(\register_file_i/_2412_ ));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(net229));
 sg13g2_mux2_1 \register_file_i/_5505_  (.A0(\register_file_i/rf_reg_39_ ),
    .A1(\register_file_i/rf_reg_103_ ),
    .S(net453),
    .X(\register_file_i/_2414_ ));
 sg13g2_a22oi_1 \register_file_i/_5506_  (.Y(\register_file_i/_2415_ ),
    .B1(\register_file_i/_2414_ ),
    .B2(net515),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_71_ ));
 sg13g2_buf_2 fanout226 (.A(net229),
    .X(net226));
 sg13g2_mux2_1 \register_file_i/_5508_  (.A0(\register_file_i/rf_reg_199_ ),
    .A1(\register_file_i/rf_reg_231_ ),
    .S(net505),
    .X(\register_file_i/_2417_ ));
 sg13g2_mux2_1 \register_file_i/_5509_  (.A0(\register_file_i/rf_reg_135_ ),
    .A1(\register_file_i/rf_reg_167_ ),
    .S(net492),
    .X(\register_file_i/_2418_ ));
 sg13g2_a22oi_1 \register_file_i/_5510_  (.Y(\register_file_i/_2419_ ),
    .B1(\register_file_i/_2418_ ),
    .B2(net1780),
    .A2(\register_file_i/_2417_ ),
    .A1(net1762));
 sg13g2_o21ai_1 \register_file_i/_5511_  (.B1(\register_file_i/_2419_ ),
    .Y(\register_file_i/_2420_ ),
    .A1(net444),
    .A2(\register_file_i/_2415_ ));
 sg13g2_nand2_1 \register_file_i/_5512_  (.Y(\register_file_i/_2421_ ),
    .A(net1907),
    .B(\register_file_i/_2420_ ));
 sg13g2_mux4_1 \register_file_i/_5513_  (.S0(net494),
    .A0(\register_file_i/rf_reg_519_ ),
    .A1(\register_file_i/rf_reg_551_ ),
    .A2(\register_file_i/rf_reg_583_ ),
    .A3(\register_file_i/rf_reg_615_ ),
    .S1(net461),
    .X(\register_file_i/_2422_ ));
 sg13g2_mux4_1 \register_file_i/_5514_  (.S0(net503),
    .A0(\register_file_i/rf_reg_647_ ),
    .A1(\register_file_i/rf_reg_679_ ),
    .A2(\register_file_i/rf_reg_711_ ),
    .A3(\register_file_i/rf_reg_743_ ),
    .S1(net459),
    .X(\register_file_i/_2423_ ));
 sg13g2_mux2_1 \register_file_i/_5515_  (.A0(\register_file_i/rf_reg_391_ ),
    .A1(\register_file_i/rf_reg_423_ ),
    .S(net497),
    .X(\register_file_i/_2424_ ));
 sg13g2_mux2_1 \register_file_i/_5516_  (.A0(\register_file_i/rf_reg_455_ ),
    .A1(\register_file_i/rf_reg_487_ ),
    .S(net504),
    .X(\register_file_i/_2425_ ));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_04361_));
 sg13g2_a22oi_1 \register_file_i/_5518_  (.Y(\register_file_i/_2427_ ),
    .B1(\register_file_i/_2425_ ),
    .B2(net1753),
    .A2(\register_file_i/_2424_ ),
    .A1(net1777));
 sg13g2_mux2_1 \register_file_i/_5519_  (.A0(\register_file_i/rf_reg_327_ ),
    .A1(\register_file_i/rf_reg_359_ ),
    .S(net493),
    .X(\register_file_i/_2428_ ));
 sg13g2_mux2_1 \register_file_i/_5520_  (.A0(\register_file_i/rf_reg_263_ ),
    .A1(\register_file_i/rf_reg_295_ ),
    .S(net500),
    .X(\register_file_i/_2429_ ));
 sg13g2_a22oi_1 \register_file_i/_5521_  (.Y(\register_file_i/_2430_ ),
    .B1(\register_file_i/_2429_ ),
    .B2(net1731),
    .A2(\register_file_i/_2428_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5522_  (.A1(\register_file_i/_2427_ ),
    .A2(\register_file_i/_2430_ ),
    .Y(\register_file_i/_2431_ ),
    .B1(net1720));
 sg13g2_a221oi_1 \register_file_i/_5523_  (.B2(net1683),
    .C1(\register_file_i/_2431_ ),
    .B1(\register_file_i/_2423_ ),
    .A1(net1726),
    .Y(\register_file_i/_2432_ ),
    .A2(\register_file_i/_2422_ ));
 sg13g2_nand3_1 \register_file_i/_5524_  (.B(\register_file_i/_2421_ ),
    .C(\register_file_i/_2432_ ),
    .A(\register_file_i/_2412_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_7_ ));
 sg13g2_mux2_1 \register_file_i/_5525_  (.A0(\register_file_i/rf_reg_902_ ),
    .A1(\register_file_i/rf_reg_934_ ),
    .S(net498),
    .X(\register_file_i/_2433_ ));
 sg13g2_buf_4 fanout224 (.X(net224),
    .A(_04361_));
 sg13g2_mux2_1 \register_file_i/_5527_  (.A0(\register_file_i/rf_reg_966_ ),
    .A1(\register_file_i/rf_reg_998_ ),
    .S(net507),
    .X(\register_file_i/_2435_ ));
 sg13g2_a22oi_1 \register_file_i/_5528_  (.Y(\register_file_i/_2436_ ),
    .B1(\register_file_i/_2435_ ),
    .B2(net1762),
    .A2(\register_file_i/_2433_ ),
    .A1(net1780));
 sg13g2_mux2_1 \register_file_i/_5529_  (.A0(\register_file_i/rf_reg_838_ ),
    .A1(\register_file_i/rf_reg_870_ ),
    .S(net496),
    .X(\register_file_i/_2437_ ));
 sg13g2_mux2_1 \register_file_i/_5530_  (.A0(\register_file_i/rf_reg_774_ ),
    .A1(\register_file_i/rf_reg_806_ ),
    .S(net501),
    .X(\register_file_i/_2438_ ));
 sg13g2_a22oi_1 \register_file_i/_5531_  (.Y(\register_file_i/_2439_ ),
    .B1(\register_file_i/_2438_ ),
    .B2(net1737),
    .A2(\register_file_i/_2437_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5532_  (.A2(\register_file_i/_2439_ ),
    .A1(\register_file_i/_2436_ ),
    .B1(net1913),
    .X(\register_file_i/_2440_ ));
 sg13g2_mux2_1 \register_file_i/_5533_  (.A0(\register_file_i/rf_reg_38_ ),
    .A1(\register_file_i/rf_reg_102_ ),
    .S(net453),
    .X(\register_file_i/_2441_ ));
 sg13g2_a22oi_1 \register_file_i/_5534_  (.Y(\register_file_i/_2442_ ),
    .B1(\register_file_i/_2441_ ),
    .B2(net515),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_70_ ));
 sg13g2_mux2_1 \register_file_i/_5535_  (.A0(\register_file_i/rf_reg_198_ ),
    .A1(\register_file_i/rf_reg_230_ ),
    .S(net505),
    .X(\register_file_i/_2443_ ));
 sg13g2_mux2_1 \register_file_i/_5536_  (.A0(\register_file_i/rf_reg_134_ ),
    .A1(\register_file_i/rf_reg_166_ ),
    .S(net492),
    .X(\register_file_i/_2444_ ));
 sg13g2_buf_4 fanout223 (.X(net223),
    .A(_04361_));
 sg13g2_a22oi_1 \register_file_i/_5538_  (.Y(\register_file_i/_2446_ ),
    .B1(\register_file_i/_2444_ ),
    .B2(net1781),
    .A2(\register_file_i/_2443_ ),
    .A1(net1763));
 sg13g2_o21ai_1 \register_file_i/_5539_  (.B1(\register_file_i/_2446_ ),
    .Y(\register_file_i/_2447_ ),
    .A1(net444),
    .A2(\register_file_i/_2442_ ));
 sg13g2_nand2_1 \register_file_i/_5540_  (.Y(\register_file_i/_2448_ ),
    .A(net1907),
    .B(\register_file_i/_2447_ ));
 sg13g2_mux4_1 \register_file_i/_5541_  (.S0(net494),
    .A0(\register_file_i/rf_reg_518_ ),
    .A1(\register_file_i/rf_reg_550_ ),
    .A2(\register_file_i/rf_reg_582_ ),
    .A3(\register_file_i/rf_reg_614_ ),
    .S1(net461),
    .X(\register_file_i/_2449_ ));
 sg13g2_mux4_1 \register_file_i/_5542_  (.S0(net502),
    .A0(\register_file_i/rf_reg_646_ ),
    .A1(\register_file_i/rf_reg_678_ ),
    .A2(\register_file_i/rf_reg_710_ ),
    .A3(\register_file_i/rf_reg_742_ ),
    .S1(net459),
    .X(\register_file_i/_2450_ ));
 sg13g2_mux2_1 \register_file_i/_5543_  (.A0(\register_file_i/rf_reg_390_ ),
    .A1(\register_file_i/rf_reg_422_ ),
    .S(net497),
    .X(\register_file_i/_2451_ ));
 sg13g2_mux2_1 \register_file_i/_5544_  (.A0(\register_file_i/rf_reg_454_ ),
    .A1(\register_file_i/rf_reg_486_ ),
    .S(net504),
    .X(\register_file_i/_2452_ ));
 sg13g2_a22oi_1 \register_file_i/_5545_  (.Y(\register_file_i/_2453_ ),
    .B1(\register_file_i/_2452_ ),
    .B2(net1753),
    .A2(\register_file_i/_2451_ ),
    .A1(net1771));
 sg13g2_mux2_1 \register_file_i/_5546_  (.A0(\register_file_i/rf_reg_326_ ),
    .A1(\register_file_i/rf_reg_358_ ),
    .S(net493),
    .X(\register_file_i/_2454_ ));
 sg13g2_mux2_1 \register_file_i/_5547_  (.A0(\register_file_i/rf_reg_262_ ),
    .A1(\register_file_i/rf_reg_294_ ),
    .S(net500),
    .X(\register_file_i/_2455_ ));
 sg13g2_buf_2 fanout222 (.A(_04378_),
    .X(net222));
 sg13g2_a22oi_1 \register_file_i/_5549_  (.Y(\register_file_i/_2457_ ),
    .B1(\register_file_i/_2455_ ),
    .B2(net1731),
    .A2(\register_file_i/_2454_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5550_  (.A1(\register_file_i/_2453_ ),
    .A2(\register_file_i/_2457_ ),
    .Y(\register_file_i/_2458_ ),
    .B1(net1720));
 sg13g2_a221oi_1 \register_file_i/_5551_  (.B2(net1683),
    .C1(\register_file_i/_2458_ ),
    .B1(\register_file_i/_2450_ ),
    .A1(net1726),
    .Y(\register_file_i/_2459_ ),
    .A2(\register_file_i/_2449_ ));
 sg13g2_nand3_1 \register_file_i/_5552_  (.B(\register_file_i/_2448_ ),
    .C(\register_file_i/_2459_ ),
    .A(\register_file_i/_2440_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_6_ ));
 sg13g2_mux2_1 \register_file_i/_5553_  (.A0(\register_file_i/rf_reg_901_ ),
    .A1(\register_file_i/rf_reg_933_ ),
    .S(net498),
    .X(\register_file_i/_2460_ ));
 sg13g2_mux2_1 \register_file_i/_5554_  (.A0(\register_file_i/rf_reg_965_ ),
    .A1(\register_file_i/rf_reg_997_ ),
    .S(net506),
    .X(\register_file_i/_2461_ ));
 sg13g2_a22oi_1 \register_file_i/_5555_  (.Y(\register_file_i/_2462_ ),
    .B1(\register_file_i/_2461_ ),
    .B2(net1762),
    .A2(\register_file_i/_2460_ ),
    .A1(net1780));
 sg13g2_mux2_1 \register_file_i/_5556_  (.A0(\register_file_i/rf_reg_837_ ),
    .A1(\register_file_i/rf_reg_869_ ),
    .S(net496),
    .X(\register_file_i/_2463_ ));
 sg13g2_mux2_1 \register_file_i/_5557_  (.A0(\register_file_i/rf_reg_773_ ),
    .A1(\register_file_i/rf_reg_805_ ),
    .S(net501),
    .X(\register_file_i/_2464_ ));
 sg13g2_a22oi_1 \register_file_i/_5558_  (.Y(\register_file_i/_2465_ ),
    .B1(\register_file_i/_2464_ ),
    .B2(net1737),
    .A2(\register_file_i/_2463_ ),
    .A1(net1748));
 sg13g2_a21o_1 \register_file_i/_5559_  (.A2(\register_file_i/_2465_ ),
    .A1(\register_file_i/_2462_ ),
    .B1(net1913),
    .X(\register_file_i/_2466_ ));
 sg13g2_mux2_1 \register_file_i/_5560_  (.A0(\register_file_i/rf_reg_37_ ),
    .A1(\register_file_i/rf_reg_101_ ),
    .S(net452),
    .X(\register_file_i/_2467_ ));
 sg13g2_a22oi_1 \register_file_i/_5561_  (.Y(\register_file_i/_2468_ ),
    .B1(\register_file_i/_2467_ ),
    .B2(net515),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_69_ ));
 sg13g2_mux2_1 \register_file_i/_5562_  (.A0(\register_file_i/rf_reg_197_ ),
    .A1(\register_file_i/rf_reg_229_ ),
    .S(net505),
    .X(\register_file_i/_2469_ ));
 sg13g2_buf_1 fanout221 (.A(net222),
    .X(net221));
 sg13g2_mux2_1 \register_file_i/_5564_  (.A0(\register_file_i/rf_reg_133_ ),
    .A1(\register_file_i/rf_reg_165_ ),
    .S(net508),
    .X(\register_file_i/_2471_ ));
 sg13g2_a22oi_1 \register_file_i/_5565_  (.Y(\register_file_i/_2472_ ),
    .B1(\register_file_i/_2471_ ),
    .B2(net1781),
    .A2(\register_file_i/_2469_ ),
    .A1(net1762));
 sg13g2_o21ai_1 \register_file_i/_5566_  (.B1(\register_file_i/_2472_ ),
    .Y(\register_file_i/_2473_ ),
    .A1(net444),
    .A2(\register_file_i/_2468_ ));
 sg13g2_nand2_1 \register_file_i/_5567_  (.Y(\register_file_i/_2474_ ),
    .A(net1907),
    .B(\register_file_i/_2473_ ));
 sg13g2_mux4_1 \register_file_i/_5568_  (.S0(net494),
    .A0(\register_file_i/rf_reg_517_ ),
    .A1(\register_file_i/rf_reg_549_ ),
    .A2(\register_file_i/rf_reg_581_ ),
    .A3(\register_file_i/rf_reg_613_ ),
    .S1(net461),
    .X(\register_file_i/_2475_ ));
 sg13g2_mux4_1 \register_file_i/_5569_  (.S0(net502),
    .A0(\register_file_i/rf_reg_645_ ),
    .A1(\register_file_i/rf_reg_677_ ),
    .A2(\register_file_i/rf_reg_709_ ),
    .A3(\register_file_i/rf_reg_741_ ),
    .S1(net459),
    .X(\register_file_i/_2476_ ));
 sg13g2_mux2_1 \register_file_i/_5570_  (.A0(\register_file_i/rf_reg_389_ ),
    .A1(\register_file_i/rf_reg_421_ ),
    .S(net497),
    .X(\register_file_i/_2477_ ));
 sg13g2_mux2_1 \register_file_i/_5571_  (.A0(\register_file_i/rf_reg_453_ ),
    .A1(\register_file_i/rf_reg_485_ ),
    .S(net504),
    .X(\register_file_i/_2478_ ));
 sg13g2_a22oi_1 \register_file_i/_5572_  (.Y(\register_file_i/_2479_ ),
    .B1(\register_file_i/_2478_ ),
    .B2(net1752),
    .A2(\register_file_i/_2477_ ),
    .A1(net1770));
 sg13g2_buf_2 fanout220 (.A(net222),
    .X(net220));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(_04523_));
 sg13g2_mux2_1 \register_file_i/_5575_  (.A0(\register_file_i/rf_reg_325_ ),
    .A1(\register_file_i/rf_reg_357_ ),
    .S(net509),
    .X(\register_file_i/_2482_ ));
 sg13g2_mux2_1 \register_file_i/_5576_  (.A0(\register_file_i/rf_reg_261_ ),
    .A1(\register_file_i/rf_reg_293_ ),
    .S(net500),
    .X(\register_file_i/_2483_ ));
 sg13g2_a22oi_1 \register_file_i/_5577_  (.Y(\register_file_i/_2484_ ),
    .B1(\register_file_i/_2483_ ),
    .B2(net1731),
    .A2(\register_file_i/_2482_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5578_  (.A1(\register_file_i/_2479_ ),
    .A2(\register_file_i/_2484_ ),
    .Y(\register_file_i/_2485_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5579_  (.B2(net1682),
    .C1(\register_file_i/_2485_ ),
    .B1(\register_file_i/_2476_ ),
    .A1(net1724),
    .Y(\register_file_i/_2486_ ),
    .A2(\register_file_i/_2475_ ));
 sg13g2_nand3_1 \register_file_i/_5580_  (.B(\register_file_i/_2474_ ),
    .C(\register_file_i/_2486_ ),
    .A(\register_file_i/_2466_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_5_ ));
 sg13g2_buf_4 fanout218 (.X(net218),
    .A(net219));
 sg13g2_mux2_1 \register_file_i/_5582_  (.A0(\register_file_i/rf_reg_900_ ),
    .A1(\register_file_i/rf_reg_932_ ),
    .S(net498),
    .X(\register_file_i/_2488_ ));
 sg13g2_mux2_1 \register_file_i/_5583_  (.A0(\register_file_i/rf_reg_964_ ),
    .A1(\register_file_i/rf_reg_996_ ),
    .S(net506),
    .X(\register_file_i/_2489_ ));
 sg13g2_buf_2 fanout217 (.A(net219),
    .X(net217));
 sg13g2_a22oi_1 \register_file_i/_5585_  (.Y(\register_file_i/_2491_ ),
    .B1(\register_file_i/_2489_ ),
    .B2(net1763),
    .A2(\register_file_i/_2488_ ),
    .A1(net1780));
 sg13g2_buf_2 fanout216 (.A(_05684_),
    .X(net216));
 sg13g2_mux2_1 \register_file_i/_5587_  (.A0(\register_file_i/rf_reg_836_ ),
    .A1(\register_file_i/rf_reg_868_ ),
    .S(net495),
    .X(\register_file_i/_2493_ ));
 sg13g2_mux2_1 \register_file_i/_5588_  (.A0(\register_file_i/rf_reg_772_ ),
    .A1(\register_file_i/rf_reg_804_ ),
    .S(net501),
    .X(\register_file_i/_2494_ ));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(_05684_));
 sg13g2_a22oi_1 \register_file_i/_5590_  (.Y(\register_file_i/_2496_ ),
    .B1(\register_file_i/_2494_ ),
    .B2(net1737),
    .A2(\register_file_i/_2493_ ),
    .A1(net1748));
 sg13g2_buf_2 fanout214 (.A(_05804_),
    .X(net214));
 sg13g2_a21o_1 \register_file_i/_5592_  (.A2(\register_file_i/_2496_ ),
    .A1(\register_file_i/_2491_ ),
    .B1(net1913),
    .X(\register_file_i/_2498_ ));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(net214));
 sg13g2_buf_2 fanout212 (.A(_08439_),
    .X(net212));
 sg13g2_mux2_1 \register_file_i/_5595_  (.A0(\register_file_i/rf_reg_36_ ),
    .A1(\register_file_i/rf_reg_100_ ),
    .S(net452),
    .X(\register_file_i/_2501_ ));
 sg13g2_a22oi_1 \register_file_i/_5596_  (.Y(\register_file_i/_2502_ ),
    .B1(\register_file_i/_2501_ ),
    .B2(net515),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_68_ ));
 sg13g2_mux2_1 \register_file_i/_5597_  (.A0(\register_file_i/rf_reg_196_ ),
    .A1(\register_file_i/rf_reg_228_ ),
    .S(net505),
    .X(\register_file_i/_2503_ ));
 sg13g2_mux2_1 \register_file_i/_5598_  (.A0(\register_file_i/rf_reg_132_ ),
    .A1(\register_file_i/rf_reg_164_ ),
    .S(net508),
    .X(\register_file_i/_2504_ ));
 sg13g2_a22oi_1 \register_file_i/_5599_  (.Y(\register_file_i/_2505_ ),
    .B1(\register_file_i/_2504_ ),
    .B2(net1781),
    .A2(\register_file_i/_2503_ ),
    .A1(net1762));
 sg13g2_o21ai_1 \register_file_i/_5600_  (.B1(\register_file_i/_2505_ ),
    .Y(\register_file_i/_2506_ ),
    .A1(net446),
    .A2(\register_file_i/_2502_ ));
 sg13g2_nand2_1 \register_file_i/_5601_  (.Y(\register_file_i/_2507_ ),
    .A(net1907),
    .B(\register_file_i/_2506_ ));
 sg13g2_buf_2 fanout211 (.A(net212),
    .X(net211));
 sg13g2_mux4_1 \register_file_i/_5603_  (.S0(net510),
    .A0(\register_file_i/rf_reg_516_ ),
    .A1(\register_file_i/rf_reg_548_ ),
    .A2(\register_file_i/rf_reg_580_ ),
    .A3(\register_file_i/rf_reg_612_ ),
    .S1(net460),
    .X(\register_file_i/_2509_ ));
 sg13g2_mux4_1 \register_file_i/_5604_  (.S0(net502),
    .A0(\register_file_i/rf_reg_644_ ),
    .A1(\register_file_i/rf_reg_676_ ),
    .A2(\register_file_i/rf_reg_708_ ),
    .A3(\register_file_i/rf_reg_740_ ),
    .S1(net459),
    .X(\register_file_i/_2510_ ));
 sg13g2_buf_4 fanout210 (.X(net210),
    .A(net212));
 sg13g2_mux2_1 \register_file_i/_5606_  (.A0(\register_file_i/rf_reg_388_ ),
    .A1(\register_file_i/rf_reg_420_ ),
    .S(net497),
    .X(\register_file_i/_2512_ ));
 sg13g2_mux2_1 \register_file_i/_5607_  (.A0(\register_file_i/rf_reg_452_ ),
    .A1(\register_file_i/rf_reg_484_ ),
    .S(net503),
    .X(\register_file_i/_2513_ ));
 sg13g2_a22oi_1 \register_file_i/_5608_  (.Y(\register_file_i/_2514_ ),
    .B1(\register_file_i/_2513_ ),
    .B2(net1753),
    .A2(\register_file_i/_2512_ ),
    .A1(net1771));
 sg13g2_mux2_1 \register_file_i/_5609_  (.A0(\register_file_i/rf_reg_324_ ),
    .A1(\register_file_i/rf_reg_356_ ),
    .S(net509),
    .X(\register_file_i/_2515_ ));
 sg13g2_mux2_1 \register_file_i/_5610_  (.A0(\register_file_i/rf_reg_260_ ),
    .A1(\register_file_i/rf_reg_292_ ),
    .S(net499),
    .X(\register_file_i/_2516_ ));
 sg13g2_a22oi_1 \register_file_i/_5611_  (.Y(\register_file_i/_2517_ ),
    .B1(\register_file_i/_2516_ ),
    .B2(net1736),
    .A2(\register_file_i/_2515_ ),
    .A1(net1747));
 sg13g2_a21oi_1 \register_file_i/_5612_  (.A1(\register_file_i/_2514_ ),
    .A2(\register_file_i/_2517_ ),
    .Y(\register_file_i/_2518_ ),
    .B1(net1720));
 sg13g2_a221oi_1 \register_file_i/_5613_  (.B2(net1684),
    .C1(\register_file_i/_2518_ ),
    .B1(\register_file_i/_2510_ ),
    .A1(net1726),
    .Y(\register_file_i/_2519_ ),
    .A2(\register_file_i/_2509_ ));
 sg13g2_nand3_1 \register_file_i/_5614_  (.B(\register_file_i/_2507_ ),
    .C(\register_file_i/_2519_ ),
    .A(\register_file_i/_2498_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ));
 sg13g2_mux2_1 \register_file_i/_5615_  (.A0(\register_file_i/rf_reg_387_ ),
    .A1(\register_file_i/rf_reg_419_ ),
    .S(net498),
    .X(\register_file_i/_2520_ ));
 sg13g2_mux2_1 \register_file_i/_5616_  (.A0(\register_file_i/rf_reg_451_ ),
    .A1(\register_file_i/rf_reg_483_ ),
    .S(net506),
    .X(\register_file_i/_2521_ ));
 sg13g2_a22oi_1 \register_file_i/_5617_  (.Y(\register_file_i/_2522_ ),
    .B1(\register_file_i/_2521_ ),
    .B2(net1760),
    .A2(\register_file_i/_2520_ ),
    .A1(net1778));
 sg13g2_buf_2 fanout209 (.A(net212),
    .X(net209));
 sg13g2_mux2_1 \register_file_i/_5619_  (.A0(\register_file_i/rf_reg_323_ ),
    .A1(\register_file_i/rf_reg_355_ ),
    .S(net512),
    .X(\register_file_i/_2524_ ));
 sg13g2_mux2_1 \register_file_i/_5620_  (.A0(\register_file_i/rf_reg_259_ ),
    .A1(\register_file_i/rf_reg_291_ ),
    .S(net501),
    .X(\register_file_i/_2525_ ));
 sg13g2_a22oi_1 \register_file_i/_5621_  (.Y(\register_file_i/_2526_ ),
    .B1(\register_file_i/_2525_ ),
    .B2(net1736),
    .A2(\register_file_i/_2524_ ),
    .A1(net1747));
 sg13g2_a21o_1 \register_file_i/_5622_  (.A2(\register_file_i/_2526_ ),
    .A1(\register_file_i/_2522_ ),
    .B1(net1720),
    .X(\register_file_i/_2527_ ));
 sg13g2_buf_1 fanout208 (.A(net209),
    .X(net208));
 sg13g2_mux2_1 \register_file_i/_5624_  (.A0(\register_file_i/rf_reg_35_ ),
    .A1(\register_file_i/rf_reg_99_ ),
    .S(net449),
    .X(\register_file_i/_2529_ ));
 sg13g2_nand2_1 \register_file_i/_5625_  (.Y(\register_file_i/_2530_ ),
    .A(net517),
    .B(\register_file_i/_2529_ ));
 sg13g2_nand3b_1 \register_file_i/_5626_  (.B(net454),
    .C(\register_file_i/rf_reg_67_ ),
    .Y(\register_file_i/_2531_ ),
    .A_N(net470));
 sg13g2_a21oi_1 \register_file_i/_5627_  (.A1(\register_file_i/_2530_ ),
    .A2(\register_file_i/_2531_ ),
    .Y(\register_file_i/_2532_ ),
    .B1(net446));
 sg13g2_mux2_1 \register_file_i/_5628_  (.A0(\register_file_i/rf_reg_131_ ),
    .A1(\register_file_i/rf_reg_163_ ),
    .S(net477),
    .X(\register_file_i/_2533_ ));
 sg13g2_mux2_1 \register_file_i/_5629_  (.A0(\register_file_i/rf_reg_195_ ),
    .A1(\register_file_i/rf_reg_227_ ),
    .S(net508),
    .X(\register_file_i/_2534_ ));
 sg13g2_a22oi_1 \register_file_i/_5630_  (.Y(\register_file_i/_2535_ ),
    .B1(\register_file_i/_2534_ ),
    .B2(net1760),
    .A2(\register_file_i/_2533_ ),
    .A1(net1778));
 sg13g2_inv_1 \register_file_i/_5631_  (.Y(\register_file_i/_2536_ ),
    .A(\register_file_i/_2535_ ));
 sg13g2_o21ai_1 \register_file_i/_5632_  (.B1(net1908),
    .Y(\register_file_i/_2537_ ),
    .A1(\register_file_i/_2532_ ),
    .A2(\register_file_i/_2536_ ));
 sg13g2_mux4_1 \register_file_i/_5633_  (.S0(net510),
    .A0(\register_file_i/rf_reg_643_ ),
    .A1(\register_file_i/rf_reg_675_ ),
    .A2(\register_file_i/rf_reg_707_ ),
    .A3(\register_file_i/rf_reg_739_ ),
    .S1(net460),
    .X(\register_file_i/_2538_ ));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net209));
 sg13g2_mux4_1 \register_file_i/_5635_  (.S0(net502),
    .A0(\register_file_i/rf_reg_515_ ),
    .A1(\register_file_i/rf_reg_547_ ),
    .A2(\register_file_i/rf_reg_579_ ),
    .A3(\register_file_i/rf_reg_611_ ),
    .S1(net462),
    .X(\register_file_i/_2540_ ));
 sg13g2_buf_4 fanout206 (.X(net206),
    .A(net209));
 sg13g2_mux2_1 \register_file_i/_5637_  (.A0(\register_file_i/rf_reg_771_ ),
    .A1(\register_file_i/rf_reg_803_ ),
    .S(net524),
    .X(\register_file_i/_2542_ ));
 sg13g2_mux2_1 \register_file_i/_5638_  (.A0(\register_file_i/rf_reg_899_ ),
    .A1(\register_file_i/rf_reg_931_ ),
    .S(net503),
    .X(\register_file_i/_2543_ ));
 sg13g2_a22oi_1 \register_file_i/_5639_  (.Y(\register_file_i/_2544_ ),
    .B1(\register_file_i/_2543_ ),
    .B2(net1771),
    .A2(\register_file_i/_2542_ ),
    .A1(net1736));
 sg13g2_mux2_1 \register_file_i/_5640_  (.A0(\register_file_i/rf_reg_835_ ),
    .A1(\register_file_i/rf_reg_867_ ),
    .S(net509),
    .X(\register_file_i/_2545_ ));
 sg13g2_mux2_1 \register_file_i/_5641_  (.A0(\register_file_i/rf_reg_963_ ),
    .A1(\register_file_i/rf_reg_995_ ),
    .S(net499),
    .X(\register_file_i/_2546_ ));
 sg13g2_a22oi_1 \register_file_i/_5642_  (.Y(\register_file_i/_2547_ ),
    .B1(\register_file_i/_2546_ ),
    .B2(net1753),
    .A2(\register_file_i/_2545_ ),
    .A1(net1747));
 sg13g2_a21oi_1 \register_file_i/_5643_  (.A1(\register_file_i/_2544_ ),
    .A2(\register_file_i/_2547_ ),
    .Y(\register_file_i/_2548_ ),
    .B1(net1915));
 sg13g2_a221oi_1 \register_file_i/_5644_  (.B2(net1725),
    .C1(\register_file_i/_2548_ ),
    .B1(\register_file_i/_2540_ ),
    .A1(net1684),
    .Y(\register_file_i/_2549_ ),
    .A2(\register_file_i/_2538_ ));
 sg13g2_nand3_1 \register_file_i/_5645_  (.B(\register_file_i/_2537_ ),
    .C(\register_file_i/_2549_ ),
    .A(\register_file_i/_2527_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_3_ ));
 sg13g2_mux2_1 \register_file_i/_5646_  (.A0(\register_file_i/rf_reg_386_ ),
    .A1(\register_file_i/rf_reg_418_ ),
    .S(net498),
    .X(\register_file_i/_2550_ ));
 sg13g2_mux2_1 \register_file_i/_5647_  (.A0(\register_file_i/rf_reg_450_ ),
    .A1(\register_file_i/rf_reg_482_ ),
    .S(net506),
    .X(\register_file_i/_2551_ ));
 sg13g2_a22oi_1 \register_file_i/_5648_  (.Y(\register_file_i/_2552_ ),
    .B1(\register_file_i/_2551_ ),
    .B2(net1760),
    .A2(\register_file_i/_2550_ ),
    .A1(net1778));
 sg13g2_mux2_1 \register_file_i/_5649_  (.A0(\register_file_i/rf_reg_322_ ),
    .A1(\register_file_i/rf_reg_354_ ),
    .S(net511),
    .X(\register_file_i/_2553_ ));
 sg13g2_mux2_1 \register_file_i/_5650_  (.A0(\register_file_i/rf_reg_258_ ),
    .A1(\register_file_i/rf_reg_290_ ),
    .S(net501),
    .X(\register_file_i/_2554_ ));
 sg13g2_a22oi_1 \register_file_i/_5651_  (.Y(\register_file_i/_2555_ ),
    .B1(\register_file_i/_2554_ ),
    .B2(net1736),
    .A2(\register_file_i/_2553_ ),
    .A1(net1747));
 sg13g2_a21o_1 \register_file_i/_5652_  (.A2(\register_file_i/_2555_ ),
    .A1(\register_file_i/_2552_ ),
    .B1(net1720),
    .X(\register_file_i/_2556_ ));
 sg13g2_mux2_1 \register_file_i/_5653_  (.A0(\register_file_i/rf_reg_34_ ),
    .A1(\register_file_i/rf_reg_98_ ),
    .S(net449),
    .X(\register_file_i/_2557_ ));
 sg13g2_nand2_1 \register_file_i/_5654_  (.Y(\register_file_i/_2558_ ),
    .A(net517),
    .B(\register_file_i/_2557_ ));
 sg13g2_nand3b_1 \register_file_i/_5655_  (.B(net454),
    .C(\register_file_i/rf_reg_66_ ),
    .Y(\register_file_i/_2559_ ),
    .A_N(net470));
 sg13g2_a21oi_1 \register_file_i/_5656_  (.A1(\register_file_i/_2558_ ),
    .A2(\register_file_i/_2559_ ),
    .Y(\register_file_i/_2560_ ),
    .B1(net446));
 sg13g2_mux2_1 \register_file_i/_5657_  (.A0(\register_file_i/rf_reg_130_ ),
    .A1(\register_file_i/rf_reg_162_ ),
    .S(net477),
    .X(\register_file_i/_2561_ ));
 sg13g2_mux2_1 \register_file_i/_5658_  (.A0(\register_file_i/rf_reg_194_ ),
    .A1(\register_file_i/rf_reg_226_ ),
    .S(net471),
    .X(\register_file_i/_2562_ ));
 sg13g2_a22oi_1 \register_file_i/_5659_  (.Y(\register_file_i/_2563_ ),
    .B1(\register_file_i/_2562_ ),
    .B2(net1761),
    .A2(\register_file_i/_2561_ ),
    .A1(net1779));
 sg13g2_inv_1 \register_file_i/_5660_  (.Y(\register_file_i/_2564_ ),
    .A(\register_file_i/_2563_ ));
 sg13g2_o21ai_1 \register_file_i/_5661_  (.B1(net1908),
    .Y(\register_file_i/_2565_ ),
    .A1(\register_file_i/_2560_ ),
    .A2(\register_file_i/_2564_ ));
 sg13g2_mux4_1 \register_file_i/_5662_  (.S0(net510),
    .A0(\register_file_i/rf_reg_642_ ),
    .A1(\register_file_i/rf_reg_674_ ),
    .A2(\register_file_i/rf_reg_706_ ),
    .A3(\register_file_i/rf_reg_738_ ),
    .S1(net460),
    .X(\register_file_i/_2566_ ));
 sg13g2_mux4_1 \register_file_i/_5663_  (.S0(net502),
    .A0(\register_file_i/rf_reg_514_ ),
    .A1(\register_file_i/rf_reg_546_ ),
    .A2(\register_file_i/rf_reg_578_ ),
    .A3(\register_file_i/rf_reg_610_ ),
    .S1(net462),
    .X(\register_file_i/_2567_ ));
 sg13g2_mux2_1 \register_file_i/_5664_  (.A0(\register_file_i/rf_reg_770_ ),
    .A1(\register_file_i/rf_reg_802_ ),
    .S(net524),
    .X(\register_file_i/_2568_ ));
 sg13g2_mux2_1 \register_file_i/_5665_  (.A0(\register_file_i/rf_reg_898_ ),
    .A1(\register_file_i/rf_reg_930_ ),
    .S(net503),
    .X(\register_file_i/_2569_ ));
 sg13g2_a22oi_1 \register_file_i/_5666_  (.Y(\register_file_i/_2570_ ),
    .B1(\register_file_i/_2569_ ),
    .B2(net1778),
    .A2(\register_file_i/_2568_ ),
    .A1(net1736));
 sg13g2_mux2_1 \register_file_i/_5667_  (.A0(\register_file_i/rf_reg_834_ ),
    .A1(\register_file_i/rf_reg_866_ ),
    .S(net509),
    .X(\register_file_i/_2571_ ));
 sg13g2_mux2_1 \register_file_i/_5668_  (.A0(\register_file_i/rf_reg_962_ ),
    .A1(\register_file_i/rf_reg_994_ ),
    .S(net499),
    .X(\register_file_i/_2572_ ));
 sg13g2_a22oi_1 \register_file_i/_5669_  (.Y(\register_file_i/_2573_ ),
    .B1(\register_file_i/_2572_ ),
    .B2(net1760),
    .A2(\register_file_i/_2571_ ),
    .A1(net1747));
 sg13g2_a21oi_2 \register_file_i/_5670_  (.B1(net1915),
    .Y(\register_file_i/_2574_ ),
    .A2(\register_file_i/_2573_ ),
    .A1(\register_file_i/_2570_ ));
 sg13g2_a221oi_1 \register_file_i/_5671_  (.B2(net1725),
    .C1(\register_file_i/_2574_ ),
    .B1(\register_file_i/_2567_ ),
    .A1(net1684),
    .Y(\register_file_i/_2575_ ),
    .A2(\register_file_i/_2566_ ));
 sg13g2_nand3_1 \register_file_i/_5672_  (.B(\register_file_i/_2565_ ),
    .C(\register_file_i/_2575_ ),
    .A(\register_file_i/_2556_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_mux2_1 \register_file_i/_5673_  (.A0(\register_file_i/rf_reg_924_ ),
    .A1(\register_file_i/rf_reg_956_ ),
    .S(net468),
    .X(\register_file_i/_2576_ ));
 sg13g2_mux2_1 \register_file_i/_5674_  (.A0(\register_file_i/rf_reg_988_ ),
    .A1(\register_file_i/rf_reg_1020_ ),
    .S(net506),
    .X(\register_file_i/_2577_ ));
 sg13g2_a22oi_1 \register_file_i/_5675_  (.Y(\register_file_i/_2578_ ),
    .B1(\register_file_i/_2577_ ),
    .B2(net1764),
    .A2(\register_file_i/_2576_ ),
    .A1(net1783));
 sg13g2_mux2_1 \register_file_i/_5676_  (.A0(\register_file_i/rf_reg_860_ ),
    .A1(\register_file_i/rf_reg_892_ ),
    .S(net511),
    .X(\register_file_i/_2579_ ));
 sg13g2_mux2_1 \register_file_i/_5677_  (.A0(\register_file_i/rf_reg_796_ ),
    .A1(\register_file_i/rf_reg_828_ ),
    .S(net501),
    .X(\register_file_i/_2580_ ));
 sg13g2_a22oi_1 \register_file_i/_5678_  (.Y(\register_file_i/_2581_ ),
    .B1(\register_file_i/_2580_ ),
    .B2(net1738),
    .A2(\register_file_i/_2579_ ),
    .A1(net1749));
 sg13g2_a21o_1 \register_file_i/_5679_  (.A2(\register_file_i/_2581_ ),
    .A1(\register_file_i/_2578_ ),
    .B1(net1914),
    .X(\register_file_i/_2582_ ));
 sg13g2_mux2_1 \register_file_i/_5680_  (.A0(\register_file_i/rf_reg_60_ ),
    .A1(\register_file_i/rf_reg_124_ ),
    .S(net452),
    .X(\register_file_i/_2583_ ));
 sg13g2_a22oi_1 \register_file_i/_5681_  (.Y(\register_file_i/_2584_ ),
    .B1(\register_file_i/_2583_ ),
    .B2(net517),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_92_ ));
 sg13g2_mux2_1 \register_file_i/_5682_  (.A0(\register_file_i/rf_reg_220_ ),
    .A1(\register_file_i/rf_reg_252_ ),
    .S(net505),
    .X(\register_file_i/_2585_ ));
 sg13g2_mux2_1 \register_file_i/_5683_  (.A0(\register_file_i/rf_reg_156_ ),
    .A1(\register_file_i/rf_reg_188_ ),
    .S(net507),
    .X(\register_file_i/_2586_ ));
 sg13g2_a22oi_1 \register_file_i/_5684_  (.Y(\register_file_i/_2587_ ),
    .B1(\register_file_i/_2586_ ),
    .B2(net1782),
    .A2(\register_file_i/_2585_ ),
    .A1(net1762));
 sg13g2_o21ai_1 \register_file_i/_5685_  (.B1(\register_file_i/_2587_ ),
    .Y(\register_file_i/_2588_ ),
    .A1(net446),
    .A2(\register_file_i/_2584_ ));
 sg13g2_nand2_1 \register_file_i/_5686_  (.Y(\register_file_i/_2589_ ),
    .A(net1907),
    .B(\register_file_i/_2588_ ));
 sg13g2_mux4_1 \register_file_i/_5687_  (.S0(net510),
    .A0(\register_file_i/rf_reg_540_ ),
    .A1(\register_file_i/rf_reg_572_ ),
    .A2(\register_file_i/rf_reg_604_ ),
    .A3(\register_file_i/rf_reg_636_ ),
    .S1(net460),
    .X(\register_file_i/_2590_ ));
 sg13g2_mux4_1 \register_file_i/_5688_  (.S0(net502),
    .A0(\register_file_i/rf_reg_668_ ),
    .A1(\register_file_i/rf_reg_700_ ),
    .A2(\register_file_i/rf_reg_732_ ),
    .A3(\register_file_i/rf_reg_764_ ),
    .S1(net462),
    .X(\register_file_i/_2591_ ));
 sg13g2_mux2_1 \register_file_i/_5689_  (.A0(\register_file_i/rf_reg_412_ ),
    .A1(\register_file_i/rf_reg_444_ ),
    .S(net524),
    .X(\register_file_i/_2592_ ));
 sg13g2_mux2_1 \register_file_i/_5690_  (.A0(\register_file_i/rf_reg_476_ ),
    .A1(\register_file_i/rf_reg_508_ ),
    .S(net503),
    .X(\register_file_i/_2593_ ));
 sg13g2_a22oi_1 \register_file_i/_5691_  (.Y(\register_file_i/_2594_ ),
    .B1(\register_file_i/_2593_ ),
    .B2(net1754),
    .A2(\register_file_i/_2592_ ),
    .A1(net1771));
 sg13g2_mux2_1 \register_file_i/_5692_  (.A0(\register_file_i/rf_reg_348_ ),
    .A1(\register_file_i/rf_reg_380_ ),
    .S(net509),
    .X(\register_file_i/_2595_ ));
 sg13g2_mux2_1 \register_file_i/_5693_  (.A0(\register_file_i/rf_reg_284_ ),
    .A1(\register_file_i/rf_reg_316_ ),
    .S(net476),
    .X(\register_file_i/_2596_ ));
 sg13g2_a22oi_1 \register_file_i/_5694_  (.Y(\register_file_i/_2597_ ),
    .B1(\register_file_i/_2596_ ),
    .B2(net1731),
    .A2(\register_file_i/_2595_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5695_  (.A1(\register_file_i/_2594_ ),
    .A2(\register_file_i/_2597_ ),
    .Y(\register_file_i/_2598_ ),
    .B1(net1721));
 sg13g2_a221oi_1 \register_file_i/_5696_  (.B2(net1684),
    .C1(\register_file_i/_2598_ ),
    .B1(\register_file_i/_2591_ ),
    .A1(net1726),
    .Y(\register_file_i/_2599_ ),
    .A2(\register_file_i/_2590_ ));
 sg13g2_nand3_1 \register_file_i/_5697_  (.B(\register_file_i/_2589_ ),
    .C(\register_file_i/_2599_ ),
    .A(\register_file_i/_2582_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_28_ ));
 sg13g2_mux2_1 \register_file_i/_5698_  (.A0(\register_file_i/rf_reg_385_ ),
    .A1(\register_file_i/rf_reg_417_ ),
    .S(net468),
    .X(\register_file_i/_2600_ ));
 sg13g2_mux2_1 \register_file_i/_5699_  (.A0(\register_file_i/rf_reg_449_ ),
    .A1(\register_file_i/rf_reg_481_ ),
    .S(net506),
    .X(\register_file_i/_2601_ ));
 sg13g2_a22oi_1 \register_file_i/_5700_  (.Y(\register_file_i/_2602_ ),
    .B1(\register_file_i/_2601_ ),
    .B2(net1765),
    .A2(\register_file_i/_2600_ ),
    .A1(net1783));
 sg13g2_mux2_1 \register_file_i/_5701_  (.A0(\register_file_i/rf_reg_321_ ),
    .A1(\register_file_i/rf_reg_353_ ),
    .S(net511),
    .X(\register_file_i/_2603_ ));
 sg13g2_mux2_1 \register_file_i/_5702_  (.A0(\register_file_i/rf_reg_257_ ),
    .A1(\register_file_i/rf_reg_289_ ),
    .S(net500),
    .X(\register_file_i/_2604_ ));
 sg13g2_a22oi_1 \register_file_i/_5703_  (.Y(\register_file_i/_2605_ ),
    .B1(\register_file_i/_2604_ ),
    .B2(net1738),
    .A2(\register_file_i/_2603_ ),
    .A1(net1749));
 sg13g2_a21o_1 \register_file_i/_5704_  (.A2(\register_file_i/_2605_ ),
    .A1(\register_file_i/_2602_ ),
    .B1(net1720),
    .X(\register_file_i/_2606_ ));
 sg13g2_mux2_1 \register_file_i/_5705_  (.A0(\register_file_i/rf_reg_33_ ),
    .A1(\register_file_i/rf_reg_97_ ),
    .S(net449),
    .X(\register_file_i/_2607_ ));
 sg13g2_nand2_1 \register_file_i/_5706_  (.Y(\register_file_i/_2608_ ),
    .A(net517),
    .B(\register_file_i/_2607_ ));
 sg13g2_nand3b_1 \register_file_i/_5707_  (.B(net454),
    .C(\register_file_i/rf_reg_65_ ),
    .Y(\register_file_i/_2609_ ),
    .A_N(net470));
 sg13g2_a21oi_1 \register_file_i/_5708_  (.A1(\register_file_i/_2608_ ),
    .A2(\register_file_i/_2609_ ),
    .Y(\register_file_i/_2610_ ),
    .B1(net442));
 sg13g2_mux2_1 \register_file_i/_5709_  (.A0(\register_file_i/rf_reg_129_ ),
    .A1(\register_file_i/rf_reg_161_ ),
    .S(net477),
    .X(\register_file_i/_2611_ ));
 sg13g2_mux2_1 \register_file_i/_5710_  (.A0(\register_file_i/rf_reg_193_ ),
    .A1(\register_file_i/rf_reg_225_ ),
    .S(net471),
    .X(\register_file_i/_2612_ ));
 sg13g2_a22oi_1 \register_file_i/_5711_  (.Y(\register_file_i/_2613_ ),
    .B1(\register_file_i/_2612_ ),
    .B2(net1761),
    .A2(\register_file_i/_2611_ ),
    .A1(net1779));
 sg13g2_inv_1 \register_file_i/_5712_  (.Y(\register_file_i/_2614_ ),
    .A(\register_file_i/_2613_ ));
 sg13g2_o21ai_1 \register_file_i/_5713_  (.B1(net1908),
    .Y(\register_file_i/_2615_ ),
    .A1(\register_file_i/_2610_ ),
    .A2(\register_file_i/_2614_ ));
 sg13g2_mux4_1 \register_file_i/_5714_  (.S0(net510),
    .A0(\register_file_i/rf_reg_641_ ),
    .A1(\register_file_i/rf_reg_673_ ),
    .A2(\register_file_i/rf_reg_705_ ),
    .A3(\register_file_i/rf_reg_737_ ),
    .S1(net456),
    .X(\register_file_i/_2616_ ));
 sg13g2_mux4_1 \register_file_i/_5715_  (.S0(net502),
    .A0(\register_file_i/rf_reg_513_ ),
    .A1(\register_file_i/rf_reg_545_ ),
    .A2(\register_file_i/rf_reg_577_ ),
    .A3(\register_file_i/rf_reg_609_ ),
    .S1(net462),
    .X(\register_file_i/_2617_ ));
 sg13g2_mux2_1 \register_file_i/_5716_  (.A0(\register_file_i/rf_reg_769_ ),
    .A1(\register_file_i/rf_reg_801_ ),
    .S(net512),
    .X(\register_file_i/_2618_ ));
 sg13g2_mux2_1 \register_file_i/_5717_  (.A0(\register_file_i/rf_reg_897_ ),
    .A1(\register_file_i/rf_reg_929_ ),
    .S(net503),
    .X(\register_file_i/_2619_ ));
 sg13g2_a22oi_1 \register_file_i/_5718_  (.Y(\register_file_i/_2620_ ),
    .B1(\register_file_i/_2619_ ),
    .B2(net1771),
    .A2(\register_file_i/_2618_ ),
    .A1(net1731));
 sg13g2_mux2_1 \register_file_i/_5719_  (.A0(\register_file_i/rf_reg_833_ ),
    .A1(\register_file_i/rf_reg_865_ ),
    .S(net508),
    .X(\register_file_i/_2621_ ));
 sg13g2_mux2_1 \register_file_i/_5720_  (.A0(\register_file_i/rf_reg_961_ ),
    .A1(\register_file_i/rf_reg_993_ ),
    .S(net476),
    .X(\register_file_i/_2622_ ));
 sg13g2_a22oi_1 \register_file_i/_5721_  (.Y(\register_file_i/_2623_ ),
    .B1(\register_file_i/_2622_ ),
    .B2(net1753),
    .A2(\register_file_i/_2621_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5722_  (.A1(\register_file_i/_2620_ ),
    .A2(\register_file_i/_2623_ ),
    .Y(\register_file_i/_2624_ ),
    .B1(net1915));
 sg13g2_a221oi_1 \register_file_i/_5723_  (.B2(net1725),
    .C1(\register_file_i/_2624_ ),
    .B1(\register_file_i/_2617_ ),
    .A1(net1683),
    .Y(\register_file_i/_2625_ ),
    .A2(\register_file_i/_2616_ ));
 sg13g2_nand3_1 \register_file_i/_5724_  (.B(\register_file_i/_2615_ ),
    .C(\register_file_i/_2625_ ),
    .A(\register_file_i/_2606_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_1_ ));
 sg13g2_mux2_1 \register_file_i/_5725_  (.A0(\register_file_i/rf_reg_384_ ),
    .A1(\register_file_i/rf_reg_416_ ),
    .S(net468),
    .X(\register_file_i/_2626_ ));
 sg13g2_mux2_1 \register_file_i/_5726_  (.A0(\register_file_i/rf_reg_448_ ),
    .A1(\register_file_i/rf_reg_480_ ),
    .S(net506),
    .X(\register_file_i/_2627_ ));
 sg13g2_a22oi_1 \register_file_i/_5727_  (.Y(\register_file_i/_2628_ ),
    .B1(\register_file_i/_2627_ ),
    .B2(net1765),
    .A2(\register_file_i/_2626_ ),
    .A1(net1783));
 sg13g2_mux2_1 \register_file_i/_5728_  (.A0(\register_file_i/rf_reg_320_ ),
    .A1(\register_file_i/rf_reg_352_ ),
    .S(net511),
    .X(\register_file_i/_2629_ ));
 sg13g2_mux2_1 \register_file_i/_5729_  (.A0(\register_file_i/rf_reg_256_ ),
    .A1(\register_file_i/rf_reg_288_ ),
    .S(net465),
    .X(\register_file_i/_2630_ ));
 sg13g2_a22oi_1 \register_file_i/_5730_  (.Y(\register_file_i/_2631_ ),
    .B1(\register_file_i/_2630_ ),
    .B2(net1738),
    .A2(\register_file_i/_2629_ ),
    .A1(net1749));
 sg13g2_a21o_1 \register_file_i/_5731_  (.A2(\register_file_i/_2631_ ),
    .A1(\register_file_i/_2628_ ),
    .B1(net1720),
    .X(\register_file_i/_2632_ ));
 sg13g2_mux2_1 \register_file_i/_5732_  (.A0(\register_file_i/rf_reg_32_ ),
    .A1(\register_file_i/rf_reg_96_ ),
    .S(net449),
    .X(\register_file_i/_2633_ ));
 sg13g2_nand2_1 \register_file_i/_5733_  (.Y(\register_file_i/_2634_ ),
    .A(net513),
    .B(\register_file_i/_2633_ ));
 sg13g2_nand3b_1 \register_file_i/_5734_  (.B(net454),
    .C(\register_file_i/rf_reg_64_ ),
    .Y(\register_file_i/_2635_ ),
    .A_N(net470));
 sg13g2_a21oi_1 \register_file_i/_5735_  (.A1(\register_file_i/_2634_ ),
    .A2(\register_file_i/_2635_ ),
    .Y(\register_file_i/_2636_ ),
    .B1(net442));
 sg13g2_mux2_1 \register_file_i/_5736_  (.A0(\register_file_i/rf_reg_128_ ),
    .A1(\register_file_i/rf_reg_160_ ),
    .S(net477),
    .X(\register_file_i/_2637_ ));
 sg13g2_mux2_1 \register_file_i/_5737_  (.A0(\register_file_i/rf_reg_192_ ),
    .A1(\register_file_i/rf_reg_224_ ),
    .S(net471),
    .X(\register_file_i/_2638_ ));
 sg13g2_a22oi_1 \register_file_i/_5738_  (.Y(\register_file_i/_2639_ ),
    .B1(\register_file_i/_2638_ ),
    .B2(net1761),
    .A2(\register_file_i/_2637_ ),
    .A1(net1779));
 sg13g2_inv_1 \register_file_i/_5739_  (.Y(\register_file_i/_2640_ ),
    .A(\register_file_i/_2639_ ));
 sg13g2_o21ai_1 \register_file_i/_5740_  (.B1(net1908),
    .Y(\register_file_i/_2641_ ),
    .A1(\register_file_i/_2636_ ),
    .A2(\register_file_i/_2640_ ));
 sg13g2_mux4_1 \register_file_i/_5741_  (.S0(net510),
    .A0(\register_file_i/rf_reg_640_ ),
    .A1(\register_file_i/rf_reg_672_ ),
    .A2(\register_file_i/rf_reg_704_ ),
    .A3(\register_file_i/rf_reg_736_ ),
    .S1(net456),
    .X(\register_file_i/_2642_ ));
 sg13g2_mux4_1 \register_file_i/_5742_  (.S0(net475),
    .A0(\register_file_i/rf_reg_512_ ),
    .A1(\register_file_i/rf_reg_544_ ),
    .A2(\register_file_i/rf_reg_576_ ),
    .A3(\register_file_i/rf_reg_608_ ),
    .S1(net462),
    .X(\register_file_i/_2643_ ));
 sg13g2_mux2_1 \register_file_i/_5743_  (.A0(\register_file_i/rf_reg_768_ ),
    .A1(\register_file_i/rf_reg_800_ ),
    .S(net512),
    .X(\register_file_i/_2644_ ));
 sg13g2_mux2_1 \register_file_i/_5744_  (.A0(\register_file_i/rf_reg_896_ ),
    .A1(\register_file_i/rf_reg_928_ ),
    .S(net480),
    .X(\register_file_i/_2645_ ));
 sg13g2_a22oi_1 \register_file_i/_5745_  (.Y(\register_file_i/_2646_ ),
    .B1(\register_file_i/_2645_ ),
    .B2(net1774),
    .A2(\register_file_i/_2644_ ),
    .A1(net1733));
 sg13g2_mux2_1 \register_file_i/_5746_  (.A0(\register_file_i/rf_reg_832_ ),
    .A1(\register_file_i/rf_reg_864_ ),
    .S(net508),
    .X(\register_file_i/_2647_ ));
 sg13g2_mux2_1 \register_file_i/_5747_  (.A0(\register_file_i/rf_reg_960_ ),
    .A1(\register_file_i/rf_reg_992_ ),
    .S(net476),
    .X(\register_file_i/_2648_ ));
 sg13g2_a22oi_1 \register_file_i/_5748_  (.Y(\register_file_i/_2649_ ),
    .B1(\register_file_i/_2648_ ),
    .B2(net1753),
    .A2(\register_file_i/_2647_ ),
    .A1(net1742));
 sg13g2_a21oi_1 \register_file_i/_5749_  (.A1(\register_file_i/_2646_ ),
    .A2(\register_file_i/_2649_ ),
    .Y(\register_file_i/_2650_ ),
    .B1(net1915));
 sg13g2_a221oi_1 \register_file_i/_5750_  (.B2(net1725),
    .C1(\register_file_i/_2650_ ),
    .B1(\register_file_i/_2643_ ),
    .A1(net1683),
    .Y(\register_file_i/_2651_ ),
    .A2(\register_file_i/_2642_ ));
 sg13g2_nand3_1 \register_file_i/_5751_  (.B(\register_file_i/_2641_ ),
    .C(\register_file_i/_2651_ ),
    .A(\register_file_i/_2632_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_0_ ));
 sg13g2_mux2_1 \register_file_i/_5752_  (.A0(\register_file_i/rf_reg_923_ ),
    .A1(\register_file_i/rf_reg_955_ ),
    .S(net468),
    .X(\register_file_i/_2652_ ));
 sg13g2_mux2_1 \register_file_i/_5753_  (.A0(\register_file_i/rf_reg_987_ ),
    .A1(\register_file_i/rf_reg_1019_ ),
    .S(net506),
    .X(\register_file_i/_2653_ ));
 sg13g2_a22oi_1 \register_file_i/_5754_  (.Y(\register_file_i/_2654_ ),
    .B1(\register_file_i/_2653_ ),
    .B2(net1764),
    .A2(\register_file_i/_2652_ ),
    .A1(net1783));
 sg13g2_mux2_1 \register_file_i/_5755_  (.A0(\register_file_i/rf_reg_859_ ),
    .A1(\register_file_i/rf_reg_891_ ),
    .S(net511),
    .X(\register_file_i/_2655_ ));
 sg13g2_mux2_1 \register_file_i/_5756_  (.A0(\register_file_i/rf_reg_795_ ),
    .A1(\register_file_i/rf_reg_827_ ),
    .S(net465),
    .X(\register_file_i/_2656_ ));
 sg13g2_a22oi_1 \register_file_i/_5757_  (.Y(\register_file_i/_2657_ ),
    .B1(\register_file_i/_2656_ ),
    .B2(net1738),
    .A2(\register_file_i/_2655_ ),
    .A1(net1749));
 sg13g2_a21o_1 \register_file_i/_5758_  (.A2(\register_file_i/_2657_ ),
    .A1(\register_file_i/_2654_ ),
    .B1(net1914),
    .X(\register_file_i/_2658_ ));
 sg13g2_mux2_1 \register_file_i/_5759_  (.A0(\register_file_i/rf_reg_59_ ),
    .A1(\register_file_i/rf_reg_123_ ),
    .S(net452),
    .X(\register_file_i/_2659_ ));
 sg13g2_a22oi_1 \register_file_i/_5760_  (.Y(\register_file_i/_2660_ ),
    .B1(\register_file_i/_2659_ ),
    .B2(net517),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_91_ ));
 sg13g2_mux2_1 \register_file_i/_5761_  (.A0(\register_file_i/rf_reg_219_ ),
    .A1(\register_file_i/rf_reg_251_ ),
    .S(net505),
    .X(\register_file_i/_2661_ ));
 sg13g2_mux2_1 \register_file_i/_5762_  (.A0(\register_file_i/rf_reg_155_ ),
    .A1(\register_file_i/rf_reg_187_ ),
    .S(net507),
    .X(\register_file_i/_2662_ ));
 sg13g2_a22oi_1 \register_file_i/_5763_  (.Y(\register_file_i/_2663_ ),
    .B1(\register_file_i/_2662_ ),
    .B2(net1782),
    .A2(\register_file_i/_2661_ ),
    .A1(net1764));
 sg13g2_o21ai_1 \register_file_i/_5764_  (.B1(\register_file_i/_2663_ ),
    .Y(\register_file_i/_2664_ ),
    .A1(net446),
    .A2(\register_file_i/_2660_ ));
 sg13g2_nand2_1 \register_file_i/_5765_  (.Y(\register_file_i/_2665_ ),
    .A(net1909),
    .B(\register_file_i/_2664_ ));
 sg13g2_mux4_1 \register_file_i/_5766_  (.S0(net510),
    .A0(\register_file_i/rf_reg_539_ ),
    .A1(\register_file_i/rf_reg_571_ ),
    .A2(\register_file_i/rf_reg_603_ ),
    .A3(\register_file_i/rf_reg_635_ ),
    .S1(net456),
    .X(\register_file_i/_2666_ ));
 sg13g2_mux4_1 \register_file_i/_5767_  (.S0(net475),
    .A0(\register_file_i/rf_reg_667_ ),
    .A1(\register_file_i/rf_reg_699_ ),
    .A2(\register_file_i/rf_reg_731_ ),
    .A3(\register_file_i/rf_reg_763_ ),
    .S1(net462),
    .X(\register_file_i/_2667_ ));
 sg13g2_mux2_1 \register_file_i/_5768_  (.A0(\register_file_i/rf_reg_411_ ),
    .A1(\register_file_i/rf_reg_443_ ),
    .S(net512),
    .X(\register_file_i/_2668_ ));
 sg13g2_mux2_1 \register_file_i/_5769_  (.A0(\register_file_i/rf_reg_475_ ),
    .A1(\register_file_i/rf_reg_507_ ),
    .S(net480),
    .X(\register_file_i/_2669_ ));
 sg13g2_a22oi_1 \register_file_i/_5770_  (.Y(\register_file_i/_2670_ ),
    .B1(\register_file_i/_2669_ ),
    .B2(net1754),
    .A2(\register_file_i/_2668_ ),
    .A1(net1771));
 sg13g2_mux2_1 \register_file_i/_5771_  (.A0(\register_file_i/rf_reg_347_ ),
    .A1(\register_file_i/rf_reg_379_ ),
    .S(net508),
    .X(\register_file_i/_2671_ ));
 sg13g2_mux2_1 \register_file_i/_5772_  (.A0(\register_file_i/rf_reg_283_ ),
    .A1(\register_file_i/rf_reg_315_ ),
    .S(net476),
    .X(\register_file_i/_2672_ ));
 sg13g2_a22oi_1 \register_file_i/_5773_  (.Y(\register_file_i/_2673_ ),
    .B1(\register_file_i/_2672_ ),
    .B2(net1730),
    .A2(\register_file_i/_2671_ ),
    .A1(net1741));
 sg13g2_a21oi_2 \register_file_i/_5774_  (.B1(net1721),
    .Y(\register_file_i/_2674_ ),
    .A2(\register_file_i/_2673_ ),
    .A1(\register_file_i/_2670_ ));
 sg13g2_a221oi_1 \register_file_i/_5775_  (.B2(net1683),
    .C1(\register_file_i/_2674_ ),
    .B1(\register_file_i/_2667_ ),
    .A1(net1725),
    .Y(\register_file_i/_2675_ ),
    .A2(\register_file_i/_2666_ ));
 sg13g2_nand3_1 \register_file_i/_5776_  (.B(\register_file_i/_2665_ ),
    .C(\register_file_i/_2675_ ),
    .A(\register_file_i/_2658_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_27_ ));
 sg13g2_mux2_1 \register_file_i/_5777_  (.A0(\register_file_i/rf_reg_922_ ),
    .A1(\register_file_i/rf_reg_954_ ),
    .S(net467),
    .X(\register_file_i/_2676_ ));
 sg13g2_mux2_1 \register_file_i/_5778_  (.A0(\register_file_i/rf_reg_986_ ),
    .A1(\register_file_i/rf_reg_1018_ ),
    .S(net505),
    .X(\register_file_i/_2677_ ));
 sg13g2_a22oi_1 \register_file_i/_5779_  (.Y(\register_file_i/_2678_ ),
    .B1(\register_file_i/_2677_ ),
    .B2(net1764),
    .A2(\register_file_i/_2676_ ),
    .A1(net1782));
 sg13g2_mux2_1 \register_file_i/_5780_  (.A0(\register_file_i/rf_reg_858_ ),
    .A1(\register_file_i/rf_reg_890_ ),
    .S(net511),
    .X(\register_file_i/_2679_ ));
 sg13g2_mux2_1 \register_file_i/_5781_  (.A0(\register_file_i/rf_reg_794_ ),
    .A1(\register_file_i/rf_reg_826_ ),
    .S(net465),
    .X(\register_file_i/_2680_ ));
 sg13g2_a22oi_1 \register_file_i/_5782_  (.Y(\register_file_i/_2681_ ),
    .B1(\register_file_i/_2680_ ),
    .B2(net1738),
    .A2(\register_file_i/_2679_ ),
    .A1(net1749));
 sg13g2_a21o_1 \register_file_i/_5783_  (.A2(\register_file_i/_2681_ ),
    .A1(\register_file_i/_2678_ ),
    .B1(net1914),
    .X(\register_file_i/_2682_ ));
 sg13g2_mux2_1 \register_file_i/_5784_  (.A0(\register_file_i/rf_reg_58_ ),
    .A1(\register_file_i/rf_reg_122_ ),
    .S(net452),
    .X(\register_file_i/_2683_ ));
 sg13g2_a22oi_1 \register_file_i/_5785_  (.Y(\register_file_i/_2684_ ),
    .B1(\register_file_i/_2683_ ),
    .B2(net517),
    .A2(net1688),
    .A1(\register_file_i/rf_reg_90_ ));
 sg13g2_mux2_1 \register_file_i/_5786_  (.A0(\register_file_i/rf_reg_218_ ),
    .A1(\register_file_i/rf_reg_250_ ),
    .S(net505),
    .X(\register_file_i/_2685_ ));
 sg13g2_mux2_1 \register_file_i/_5787_  (.A0(\register_file_i/rf_reg_154_ ),
    .A1(\register_file_i/rf_reg_186_ ),
    .S(net507),
    .X(\register_file_i/_2686_ ));
 sg13g2_a22oi_1 \register_file_i/_5788_  (.Y(\register_file_i/_2687_ ),
    .B1(\register_file_i/_2686_ ),
    .B2(net1782),
    .A2(\register_file_i/_2685_ ),
    .A1(net1764));
 sg13g2_o21ai_1 \register_file_i/_5789_  (.B1(\register_file_i/_2687_ ),
    .Y(\register_file_i/_2688_ ),
    .A1(net446),
    .A2(\register_file_i/_2684_ ));
 sg13g2_nand2_1 \register_file_i/_5790_  (.Y(\register_file_i/_2689_ ),
    .A(net1909),
    .B(\register_file_i/_2688_ ));
 sg13g2_mux4_1 \register_file_i/_5791_  (.S0(net509),
    .A0(\register_file_i/rf_reg_538_ ),
    .A1(\register_file_i/rf_reg_570_ ),
    .A2(\register_file_i/rf_reg_602_ ),
    .A3(\register_file_i/rf_reg_634_ ),
    .S1(net456),
    .X(\register_file_i/_2690_ ));
 sg13g2_mux4_1 \register_file_i/_5792_  (.S0(net475),
    .A0(\register_file_i/rf_reg_666_ ),
    .A1(\register_file_i/rf_reg_698_ ),
    .A2(\register_file_i/rf_reg_730_ ),
    .A3(\register_file_i/rf_reg_762_ ),
    .S1(net462),
    .X(\register_file_i/_2691_ ));
 sg13g2_mux2_1 \register_file_i/_5793_  (.A0(\register_file_i/rf_reg_410_ ),
    .A1(\register_file_i/rf_reg_442_ ),
    .S(net512),
    .X(\register_file_i/_2692_ ));
 sg13g2_mux2_1 \register_file_i/_5794_  (.A0(\register_file_i/rf_reg_474_ ),
    .A1(\register_file_i/rf_reg_506_ ),
    .S(net480),
    .X(\register_file_i/_2693_ ));
 sg13g2_a22oi_1 \register_file_i/_5795_  (.Y(\register_file_i/_2694_ ),
    .B1(\register_file_i/_2693_ ),
    .B2(net1752),
    .A2(\register_file_i/_2692_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5796_  (.A0(\register_file_i/rf_reg_346_ ),
    .A1(\register_file_i/rf_reg_378_ ),
    .S(net508),
    .X(\register_file_i/_2695_ ));
 sg13g2_mux2_1 \register_file_i/_5797_  (.A0(\register_file_i/rf_reg_282_ ),
    .A1(\register_file_i/rf_reg_314_ ),
    .S(net476),
    .X(\register_file_i/_2696_ ));
 sg13g2_a22oi_1 \register_file_i/_5798_  (.Y(\register_file_i/_2697_ ),
    .B1(\register_file_i/_2696_ ),
    .B2(net1730),
    .A2(\register_file_i/_2695_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5799_  (.A1(\register_file_i/_2694_ ),
    .A2(\register_file_i/_2697_ ),
    .Y(\register_file_i/_2698_ ),
    .B1(net1721));
 sg13g2_a221oi_1 \register_file_i/_5800_  (.B2(net1683),
    .C1(\register_file_i/_2698_ ),
    .B1(\register_file_i/_2691_ ),
    .A1(net1725),
    .Y(\register_file_i/_2699_ ),
    .A2(\register_file_i/_2690_ ));
 sg13g2_nand3_1 \register_file_i/_5801_  (.B(\register_file_i/_2689_ ),
    .C(\register_file_i/_2699_ ),
    .A(\register_file_i/_2682_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_26_ ));
 sg13g2_mux2_1 \register_file_i/_5802_  (.A0(\register_file_i/rf_reg_921_ ),
    .A1(\register_file_i/rf_reg_953_ ),
    .S(net467),
    .X(\register_file_i/_2700_ ));
 sg13g2_mux2_1 \register_file_i/_5803_  (.A0(\register_file_i/rf_reg_985_ ),
    .A1(\register_file_i/rf_reg_1017_ ),
    .S(net469),
    .X(\register_file_i/_2701_ ));
 sg13g2_a22oi_1 \register_file_i/_5804_  (.Y(\register_file_i/_2702_ ),
    .B1(\register_file_i/_2701_ ),
    .B2(net1768),
    .A2(\register_file_i/_2700_ ),
    .A1(net1786));
 sg13g2_mux2_1 \register_file_i/_5805_  (.A0(\register_file_i/rf_reg_857_ ),
    .A1(\register_file_i/rf_reg_889_ ),
    .S(net511),
    .X(\register_file_i/_2703_ ));
 sg13g2_mux2_1 \register_file_i/_5806_  (.A0(\register_file_i/rf_reg_793_ ),
    .A1(\register_file_i/rf_reg_825_ ),
    .S(net465),
    .X(\register_file_i/_2704_ ));
 sg13g2_a22oi_1 \register_file_i/_5807_  (.Y(\register_file_i/_2705_ ),
    .B1(\register_file_i/_2704_ ),
    .B2(net1739),
    .A2(\register_file_i/_2703_ ),
    .A1(net1750));
 sg13g2_a21o_1 \register_file_i/_5808_  (.A2(\register_file_i/_2705_ ),
    .A1(\register_file_i/_2702_ ),
    .B1(net1918),
    .X(\register_file_i/_2706_ ));
 sg13g2_mux2_1 \register_file_i/_5809_  (.A0(\register_file_i/rf_reg_57_ ),
    .A1(\register_file_i/rf_reg_121_ ),
    .S(net452),
    .X(\register_file_i/_2707_ ));
 sg13g2_a22oi_1 \register_file_i/_5810_  (.Y(\register_file_i/_2708_ ),
    .B1(\register_file_i/_2707_ ),
    .B2(net517),
    .A2(net1689),
    .A1(\register_file_i/rf_reg_89_ ));
 sg13g2_mux2_1 \register_file_i/_5811_  (.A0(\register_file_i/rf_reg_217_ ),
    .A1(\register_file_i/rf_reg_249_ ),
    .S(net504),
    .X(\register_file_i/_2709_ ));
 sg13g2_mux2_1 \register_file_i/_5812_  (.A0(\register_file_i/rf_reg_153_ ),
    .A1(\register_file_i/rf_reg_185_ ),
    .S(net507),
    .X(\register_file_i/_2710_ ));
 sg13g2_a22oi_1 \register_file_i/_5813_  (.Y(\register_file_i/_2711_ ),
    .B1(\register_file_i/_2710_ ),
    .B2(net1782),
    .A2(\register_file_i/_2709_ ),
    .A1(net1764));
 sg13g2_o21ai_1 \register_file_i/_5814_  (.B1(\register_file_i/_2711_ ),
    .Y(\register_file_i/_2712_ ),
    .A1(net446),
    .A2(\register_file_i/_2708_ ));
 sg13g2_nand2_1 \register_file_i/_5815_  (.Y(\register_file_i/_2713_ ),
    .A(net1909),
    .B(\register_file_i/_2712_ ));
 sg13g2_mux4_1 \register_file_i/_5816_  (.S0(net509),
    .A0(\register_file_i/rf_reg_537_ ),
    .A1(\register_file_i/rf_reg_569_ ),
    .A2(\register_file_i/rf_reg_601_ ),
    .A3(\register_file_i/rf_reg_633_ ),
    .S1(net456),
    .X(\register_file_i/_2714_ ));
 sg13g2_mux4_1 \register_file_i/_5817_  (.S0(net475),
    .A0(\register_file_i/rf_reg_665_ ),
    .A1(\register_file_i/rf_reg_697_ ),
    .A2(\register_file_i/rf_reg_729_ ),
    .A3(\register_file_i/rf_reg_761_ ),
    .S1(net462),
    .X(\register_file_i/_2715_ ));
 sg13g2_mux2_1 \register_file_i/_5818_  (.A0(\register_file_i/rf_reg_409_ ),
    .A1(\register_file_i/rf_reg_441_ ),
    .S(net512),
    .X(\register_file_i/_2716_ ));
 sg13g2_mux2_1 \register_file_i/_5819_  (.A0(\register_file_i/rf_reg_473_ ),
    .A1(\register_file_i/rf_reg_505_ ),
    .S(net480),
    .X(\register_file_i/_2717_ ));
 sg13g2_a22oi_1 \register_file_i/_5820_  (.Y(\register_file_i/_2718_ ),
    .B1(\register_file_i/_2717_ ),
    .B2(net1752),
    .A2(\register_file_i/_2716_ ),
    .A1(net1770));
 sg13g2_mux2_1 \register_file_i/_5821_  (.A0(\register_file_i/rf_reg_345_ ),
    .A1(\register_file_i/rf_reg_377_ ),
    .S(net508),
    .X(\register_file_i/_2719_ ));
 sg13g2_mux2_1 \register_file_i/_5822_  (.A0(\register_file_i/rf_reg_281_ ),
    .A1(\register_file_i/rf_reg_313_ ),
    .S(net476),
    .X(\register_file_i/_2720_ ));
 sg13g2_a22oi_1 \register_file_i/_5823_  (.Y(\register_file_i/_2721_ ),
    .B1(\register_file_i/_2720_ ),
    .B2(net1730),
    .A2(\register_file_i/_2719_ ),
    .A1(net1741));
 sg13g2_a21oi_1 \register_file_i/_5824_  (.A1(\register_file_i/_2718_ ),
    .A2(\register_file_i/_2721_ ),
    .Y(\register_file_i/_2722_ ),
    .B1(net1719));
 sg13g2_a221oi_1 \register_file_i/_5825_  (.B2(net1683),
    .C1(\register_file_i/_2722_ ),
    .B1(\register_file_i/_2715_ ),
    .A1(net1725),
    .Y(\register_file_i/_2723_ ),
    .A2(\register_file_i/_2714_ ));
 sg13g2_nand3_1 \register_file_i/_5826_  (.B(\register_file_i/_2713_ ),
    .C(\register_file_i/_2723_ ),
    .A(\register_file_i/_2706_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_25_ ));
 sg13g2_mux2_1 \register_file_i/_5827_  (.A0(\register_file_i/rf_reg_920_ ),
    .A1(\register_file_i/rf_reg_952_ ),
    .S(net467),
    .X(\register_file_i/_2724_ ));
 sg13g2_mux2_1 \register_file_i/_5828_  (.A0(\register_file_i/rf_reg_984_ ),
    .A1(\register_file_i/rf_reg_1016_ ),
    .S(net468),
    .X(\register_file_i/_2725_ ));
 sg13g2_a22oi_1 \register_file_i/_5829_  (.Y(\register_file_i/_2726_ ),
    .B1(\register_file_i/_2725_ ),
    .B2(net1768),
    .A2(\register_file_i/_2724_ ),
    .A1(net1786));
 sg13g2_mux2_1 \register_file_i/_5830_  (.A0(\register_file_i/rf_reg_856_ ),
    .A1(\register_file_i/rf_reg_888_ ),
    .S(net511),
    .X(\register_file_i/_2727_ ));
 sg13g2_mux2_1 \register_file_i/_5831_  (.A0(\register_file_i/rf_reg_792_ ),
    .A1(\register_file_i/rf_reg_824_ ),
    .S(net465),
    .X(\register_file_i/_2728_ ));
 sg13g2_a22oi_1 \register_file_i/_5832_  (.Y(\register_file_i/_2729_ ),
    .B1(\register_file_i/_2728_ ),
    .B2(net1739),
    .A2(\register_file_i/_2727_ ),
    .A1(net1750));
 sg13g2_a21o_1 \register_file_i/_5833_  (.A2(\register_file_i/_2729_ ),
    .A1(\register_file_i/_2726_ ),
    .B1(net1918),
    .X(\register_file_i/_2730_ ));
 sg13g2_mux2_1 \register_file_i/_5834_  (.A0(\register_file_i/rf_reg_56_ ),
    .A1(\register_file_i/rf_reg_120_ ),
    .S(net452),
    .X(\register_file_i/_2731_ ));
 sg13g2_a22oi_1 \register_file_i/_5835_  (.Y(\register_file_i/_2732_ ),
    .B1(\register_file_i/_2731_ ),
    .B2(net516),
    .A2(net1692),
    .A1(\register_file_i/rf_reg_88_ ));
 sg13g2_mux2_1 \register_file_i/_5836_  (.A0(\register_file_i/rf_reg_216_ ),
    .A1(\register_file_i/rf_reg_248_ ),
    .S(net504),
    .X(\register_file_i/_2733_ ));
 sg13g2_mux2_1 \register_file_i/_5837_  (.A0(\register_file_i/rf_reg_152_ ),
    .A1(\register_file_i/rf_reg_184_ ),
    .S(net507),
    .X(\register_file_i/_2734_ ));
 sg13g2_a22oi_1 \register_file_i/_5838_  (.Y(\register_file_i/_2735_ ),
    .B1(\register_file_i/_2734_ ),
    .B2(net1786),
    .A2(\register_file_i/_2733_ ),
    .A1(net1768));
 sg13g2_o21ai_1 \register_file_i/_5839_  (.B1(\register_file_i/_2735_ ),
    .Y(\register_file_i/_2736_ ),
    .A1(net446),
    .A2(\register_file_i/_2732_ ));
 sg13g2_nand2_1 \register_file_i/_5840_  (.Y(\register_file_i/_2737_ ),
    .A(net1912),
    .B(\register_file_i/_2736_ ));
 sg13g2_mux4_1 \register_file_i/_5841_  (.S0(net509),
    .A0(\register_file_i/rf_reg_536_ ),
    .A1(\register_file_i/rf_reg_568_ ),
    .A2(\register_file_i/rf_reg_600_ ),
    .A3(\register_file_i/rf_reg_632_ ),
    .S1(net456),
    .X(\register_file_i/_2738_ ));
 sg13g2_mux4_1 \register_file_i/_5842_  (.S0(net475),
    .A0(\register_file_i/rf_reg_664_ ),
    .A1(\register_file_i/rf_reg_696_ ),
    .A2(\register_file_i/rf_reg_728_ ),
    .A3(\register_file_i/rf_reg_760_ ),
    .S1(net461),
    .X(\register_file_i/_2739_ ));
 sg13g2_mux2_1 \register_file_i/_5843_  (.A0(\register_file_i/rf_reg_408_ ),
    .A1(\register_file_i/rf_reg_440_ ),
    .S(net512),
    .X(\register_file_i/_2740_ ));
 sg13g2_mux2_1 \register_file_i/_5844_  (.A0(\register_file_i/rf_reg_472_ ),
    .A1(\register_file_i/rf_reg_504_ ),
    .S(net479),
    .X(\register_file_i/_2741_ ));
 sg13g2_a22oi_1 \register_file_i/_5845_  (.Y(\register_file_i/_2742_ ),
    .B1(\register_file_i/_2741_ ),
    .B2(net1755),
    .A2(\register_file_i/_2740_ ),
    .A1(net1772));
 sg13g2_mux2_1 \register_file_i/_5846_  (.A0(\register_file_i/rf_reg_344_ ),
    .A1(\register_file_i/rf_reg_376_ ),
    .S(net470),
    .X(\register_file_i/_2743_ ));
 sg13g2_mux2_1 \register_file_i/_5847_  (.A0(\register_file_i/rf_reg_280_ ),
    .A1(\register_file_i/rf_reg_312_ ),
    .S(net476),
    .X(\register_file_i/_2744_ ));
 sg13g2_a22oi_1 \register_file_i/_5848_  (.Y(\register_file_i/_2745_ ),
    .B1(\register_file_i/_2744_ ),
    .B2(net1733),
    .A2(\register_file_i/_2743_ ),
    .A1(net1744));
 sg13g2_a21oi_1 \register_file_i/_5849_  (.A1(\register_file_i/_2742_ ),
    .A2(\register_file_i/_2745_ ),
    .Y(\register_file_i/_2746_ ),
    .B1(net1722));
 sg13g2_a221oi_1 \register_file_i/_5850_  (.B2(net1685),
    .C1(\register_file_i/_2746_ ),
    .B1(\register_file_i/_2739_ ),
    .A1(net1727),
    .Y(\register_file_i/_2747_ ),
    .A2(\register_file_i/_2738_ ));
 sg13g2_nand3_1 \register_file_i/_5851_  (.B(\register_file_i/_2737_ ),
    .C(\register_file_i/_2747_ ),
    .A(\register_file_i/_2730_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_24_ ));
 sg13g2_mux2_1 \register_file_i/_5852_  (.A0(\register_file_i/rf_reg_919_ ),
    .A1(\register_file_i/rf_reg_951_ ),
    .S(net467),
    .X(\register_file_i/_2748_ ));
 sg13g2_mux2_1 \register_file_i/_5853_  (.A0(\register_file_i/rf_reg_983_ ),
    .A1(\register_file_i/rf_reg_1015_ ),
    .S(net468),
    .X(\register_file_i/_2749_ ));
 sg13g2_a22oi_1 \register_file_i/_5854_  (.Y(\register_file_i/_2750_ ),
    .B1(\register_file_i/_2749_ ),
    .B2(net1753),
    .A2(\register_file_i/_2748_ ),
    .A1(net1771));
 sg13g2_mux2_1 \register_file_i/_5855_  (.A0(\register_file_i/rf_reg_855_ ),
    .A1(\register_file_i/rf_reg_887_ ),
    .S(net510),
    .X(\register_file_i/_2751_ ));
 sg13g2_mux2_1 \register_file_i/_5856_  (.A0(\register_file_i/rf_reg_791_ ),
    .A1(\register_file_i/rf_reg_823_ ),
    .S(net465),
    .X(\register_file_i/_2752_ ));
 sg13g2_a22oi_1 \register_file_i/_5857_  (.Y(\register_file_i/_2753_ ),
    .B1(\register_file_i/_2752_ ),
    .B2(net1736),
    .A2(\register_file_i/_2751_ ),
    .A1(net1747));
 sg13g2_a21o_1 \register_file_i/_5858_  (.A2(\register_file_i/_2753_ ),
    .A1(\register_file_i/_2750_ ),
    .B1(net1916),
    .X(\register_file_i/_2754_ ));
 sg13g2_mux2_1 \register_file_i/_5859_  (.A0(\register_file_i/rf_reg_55_ ),
    .A1(\register_file_i/rf_reg_119_ ),
    .S(net452),
    .X(\register_file_i/_2755_ ));
 sg13g2_a22oi_1 \register_file_i/_5860_  (.Y(\register_file_i/_2756_ ),
    .B1(\register_file_i/_2755_ ),
    .B2(net516),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_87_ ));
 sg13g2_mux2_1 \register_file_i/_5861_  (.A0(\register_file_i/rf_reg_215_ ),
    .A1(\register_file_i/rf_reg_247_ ),
    .S(net504),
    .X(\register_file_i/_2757_ ));
 sg13g2_mux2_1 \register_file_i/_5862_  (.A0(\register_file_i/rf_reg_151_ ),
    .A1(\register_file_i/rf_reg_183_ ),
    .S(net507),
    .X(\register_file_i/_2758_ ));
 sg13g2_a22oi_1 \register_file_i/_5863_  (.Y(\register_file_i/_2759_ ),
    .B1(\register_file_i/_2758_ ),
    .B2(net1779),
    .A2(\register_file_i/_2757_ ),
    .A1(net1761));
 sg13g2_o21ai_1 \register_file_i/_5864_  (.B1(\register_file_i/_2759_ ),
    .Y(\register_file_i/_2760_ ),
    .A1(net445),
    .A2(\register_file_i/_2756_ ));
 sg13g2_nand2_1 \register_file_i/_5865_  (.Y(\register_file_i/_2761_ ),
    .A(net1908),
    .B(\register_file_i/_2760_ ));
 sg13g2_mux4_1 \register_file_i/_5866_  (.S0(net466),
    .A0(\register_file_i/rf_reg_535_ ),
    .A1(\register_file_i/rf_reg_567_ ),
    .A2(\register_file_i/rf_reg_599_ ),
    .A3(\register_file_i/rf_reg_631_ ),
    .S1(net455),
    .X(\register_file_i/_2762_ ));
 sg13g2_mux4_1 \register_file_i/_5867_  (.S0(net475),
    .A0(\register_file_i/rf_reg_663_ ),
    .A1(\register_file_i/rf_reg_695_ ),
    .A2(\register_file_i/rf_reg_727_ ),
    .A3(\register_file_i/rf_reg_759_ ),
    .S1(net461),
    .X(\register_file_i/_2763_ ));
 sg13g2_mux2_1 \register_file_i/_5868_  (.A0(\register_file_i/rf_reg_407_ ),
    .A1(\register_file_i/rf_reg_439_ ),
    .S(net512),
    .X(\register_file_i/_2764_ ));
 sg13g2_mux2_1 \register_file_i/_5869_  (.A0(\register_file_i/rf_reg_471_ ),
    .A1(\register_file_i/rf_reg_503_ ),
    .S(net479),
    .X(\register_file_i/_2765_ ));
 sg13g2_a22oi_1 \register_file_i/_5870_  (.Y(\register_file_i/_2766_ ),
    .B1(\register_file_i/_2765_ ),
    .B2(net1757),
    .A2(\register_file_i/_2764_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5871_  (.A0(\register_file_i/rf_reg_343_ ),
    .A1(\register_file_i/rf_reg_375_ ),
    .S(net469),
    .X(\register_file_i/_2767_ ));
 sg13g2_mux2_1 \register_file_i/_5872_  (.A0(\register_file_i/rf_reg_279_ ),
    .A1(\register_file_i/rf_reg_311_ ),
    .S(net476),
    .X(\register_file_i/_2768_ ));
 sg13g2_a22oi_1 \register_file_i/_5873_  (.Y(\register_file_i/_2769_ ),
    .B1(\register_file_i/_2768_ ),
    .B2(net1733),
    .A2(\register_file_i/_2767_ ),
    .A1(net1744));
 sg13g2_a21oi_1 \register_file_i/_5874_  (.A1(\register_file_i/_2766_ ),
    .A2(\register_file_i/_2769_ ),
    .Y(\register_file_i/_2770_ ),
    .B1(net1723));
 sg13g2_a221oi_1 \register_file_i/_5875_  (.B2(net1685),
    .C1(\register_file_i/_2770_ ),
    .B1(\register_file_i/_2763_ ),
    .A1(net1727),
    .Y(\register_file_i/_2771_ ),
    .A2(\register_file_i/_2762_ ));
 sg13g2_nand3_1 \register_file_i/_5876_  (.B(\register_file_i/_2761_ ),
    .C(\register_file_i/_2771_ ),
    .A(\register_file_i/_2754_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_23_ ));
 sg13g2_mux2_1 \register_file_i/_5877_  (.A0(\register_file_i/rf_reg_918_ ),
    .A1(\register_file_i/rf_reg_950_ ),
    .S(net467),
    .X(\register_file_i/_2772_ ));
 sg13g2_mux2_1 \register_file_i/_5878_  (.A0(\register_file_i/rf_reg_982_ ),
    .A1(\register_file_i/rf_reg_1014_ ),
    .S(net468),
    .X(\register_file_i/_2773_ ));
 sg13g2_a22oi_1 \register_file_i/_5879_  (.Y(\register_file_i/_2774_ ),
    .B1(\register_file_i/_2773_ ),
    .B2(net1768),
    .A2(\register_file_i/_2772_ ),
    .A1(net1786));
 sg13g2_mux2_1 \register_file_i/_5880_  (.A0(\register_file_i/rf_reg_854_ ),
    .A1(\register_file_i/rf_reg_886_ ),
    .S(net472),
    .X(\register_file_i/_2775_ ));
 sg13g2_mux2_1 \register_file_i/_5881_  (.A0(\register_file_i/rf_reg_790_ ),
    .A1(\register_file_i/rf_reg_822_ ),
    .S(net464),
    .X(\register_file_i/_2776_ ));
 sg13g2_a22oi_1 \register_file_i/_5882_  (.Y(\register_file_i/_2777_ ),
    .B1(\register_file_i/_2776_ ),
    .B2(net1739),
    .A2(\register_file_i/_2775_ ),
    .A1(net1750));
 sg13g2_a21o_1 \register_file_i/_5883_  (.A2(\register_file_i/_2777_ ),
    .A1(\register_file_i/_2774_ ),
    .B1(net1918),
    .X(\register_file_i/_2778_ ));
 sg13g2_mux2_1 \register_file_i/_5884_  (.A0(\register_file_i/rf_reg_54_ ),
    .A1(\register_file_i/rf_reg_118_ ),
    .S(net449),
    .X(\register_file_i/_2779_ ));
 sg13g2_a22oi_1 \register_file_i/_5885_  (.Y(\register_file_i/_2780_ ),
    .B1(\register_file_i/_2779_ ),
    .B2(net516),
    .A2(net1690),
    .A1(\register_file_i/rf_reg_86_ ));
 sg13g2_mux2_1 \register_file_i/_5886_  (.A0(\register_file_i/rf_reg_214_ ),
    .A1(\register_file_i/rf_reg_246_ ),
    .S(net477),
    .X(\register_file_i/_2781_ ));
 sg13g2_mux2_1 \register_file_i/_5887_  (.A0(\register_file_i/rf_reg_150_ ),
    .A1(\register_file_i/rf_reg_182_ ),
    .S(net507),
    .X(\register_file_i/_2782_ ));
 sg13g2_a22oi_1 \register_file_i/_5888_  (.Y(\register_file_i/_2783_ ),
    .B1(\register_file_i/_2782_ ),
    .B2(net1784),
    .A2(\register_file_i/_2781_ ),
    .A1(net1766));
 sg13g2_o21ai_1 \register_file_i/_5889_  (.B1(\register_file_i/_2783_ ),
    .Y(\register_file_i/_2784_ ),
    .A1(net445),
    .A2(\register_file_i/_2780_ ));
 sg13g2_nand2_1 \register_file_i/_5890_  (.Y(\register_file_i/_2785_ ),
    .A(net1912),
    .B(\register_file_i/_2784_ ));
 sg13g2_mux4_1 \register_file_i/_5891_  (.S0(net466),
    .A0(\register_file_i/rf_reg_534_ ),
    .A1(\register_file_i/rf_reg_566_ ),
    .A2(\register_file_i/rf_reg_598_ ),
    .A3(\register_file_i/rf_reg_630_ ),
    .S1(net455),
    .X(\register_file_i/_2786_ ));
 sg13g2_mux4_1 \register_file_i/_5892_  (.S0(net474),
    .A0(\register_file_i/rf_reg_662_ ),
    .A1(\register_file_i/rf_reg_694_ ),
    .A2(\register_file_i/rf_reg_726_ ),
    .A3(\register_file_i/rf_reg_758_ ),
    .S1(net455),
    .X(\register_file_i/_2787_ ));
 sg13g2_mux2_1 \register_file_i/_5893_  (.A0(\register_file_i/rf_reg_406_ ),
    .A1(\register_file_i/rf_reg_438_ ),
    .S(net478),
    .X(\register_file_i/_2788_ ));
 sg13g2_mux2_1 \register_file_i/_5894_  (.A0(\register_file_i/rf_reg_470_ ),
    .A1(\register_file_i/rf_reg_502_ ),
    .S(net479),
    .X(\register_file_i/_2789_ ));
 sg13g2_a22oi_1 \register_file_i/_5895_  (.Y(\register_file_i/_2790_ ),
    .B1(\register_file_i/_2789_ ),
    .B2(net1757),
    .A2(\register_file_i/_2788_ ),
    .A1(net1774));
 sg13g2_mux2_1 \register_file_i/_5896_  (.A0(\register_file_i/rf_reg_342_ ),
    .A1(\register_file_i/rf_reg_374_ ),
    .S(net469),
    .X(\register_file_i/_2791_ ));
 sg13g2_mux2_1 \register_file_i/_5897_  (.A0(\register_file_i/rf_reg_278_ ),
    .A1(\register_file_i/rf_reg_310_ ),
    .S(net475),
    .X(\register_file_i/_2792_ ));
 sg13g2_a22oi_1 \register_file_i/_5898_  (.Y(\register_file_i/_2793_ ),
    .B1(\register_file_i/_2792_ ),
    .B2(net1734),
    .A2(\register_file_i/_2791_ ),
    .A1(net1744));
 sg13g2_a21oi_1 \register_file_i/_5899_  (.A1(\register_file_i/_2790_ ),
    .A2(\register_file_i/_2793_ ),
    .Y(\register_file_i/_2794_ ),
    .B1(net1723));
 sg13g2_a221oi_1 \register_file_i/_5900_  (.B2(net1686),
    .C1(\register_file_i/_2794_ ),
    .B1(\register_file_i/_2787_ ),
    .A1(net1727),
    .Y(\register_file_i/_2795_ ),
    .A2(\register_file_i/_2786_ ));
 sg13g2_nand3_1 \register_file_i/_5901_  (.B(\register_file_i/_2785_ ),
    .C(\register_file_i/_2795_ ),
    .A(\register_file_i/_2778_ ),
    .Y(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_22_ ));
 sg13g2_buf_2 fanout205 (.A(_08443_),
    .X(net205));
 sg13g2_buf_2 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_2 fanout203 (.A(net204),
    .X(net203));
 sg13g2_nand2_2 \register_file_i/_5905_  (.Y(\register_file_i/_2799_ ),
    .A(net1991),
    .B(net2099));
 sg13g2_nand4_1 \register_file_i/_5906_  (.B(rf_we_wb),
    .C(\id_stage_i.controller_i.instr_i_8_ ),
    .A(net553),
    .Y(\register_file_i/_2800_ ),
    .D(net1993));
 sg13g2_nor2_1 \register_file_i/_5907_  (.A(\register_file_i/_2799_ ),
    .B(\register_file_i/_2800_ ),
    .Y(\register_file_i/_2801_ ));
 sg13g2_buf_2 fanout202 (.A(net204),
    .X(net202));
 sg13g2_mux2_1 \register_file_i/_5909_  (.A0(\register_file_i/rf_reg_1000_ ),
    .A1(net877),
    .S(net985),
    .X(\register_file_i/_0000_ ));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(net204));
 sg13g2_mux2_1 \register_file_i/_5911_  (.A0(\register_file_i/rf_reg_1001_ ),
    .A1(net806),
    .S(net985),
    .X(\register_file_i/_0001_ ));
 sg13g2_buf_8 fanout200 (.A(net204),
    .X(net200));
 sg13g2_mux2_1 \register_file_i/_5913_  (.A0(\register_file_i/rf_reg_1002_ ),
    .A1(net797),
    .S(net986),
    .X(\register_file_i/_0002_ ));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net204));
 sg13g2_mux2_1 \register_file_i/_5915_  (.A0(\register_file_i/rf_reg_1003_ ),
    .A1(net792),
    .S(net985),
    .X(\register_file_i/_0003_ ));
 sg13g2_buf_2 fanout198 (.A(alu_operand_a_ex_0_),
    .X(net198));
 sg13g2_mux2_1 \register_file_i/_5917_  (.A0(\register_file_i/rf_reg_1004_ ),
    .A1(net801),
    .S(net986),
    .X(\register_file_i/_0004_ ));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(alu_operand_a_ex_0_));
 sg13g2_mux2_1 \register_file_i/_5919_  (.A0(\register_file_i/rf_reg_1005_ ),
    .A1(net788),
    .S(net987),
    .X(\register_file_i/_0005_ ));
 sg13g2_buf_2 fanout196 (.A(alu_operand_a_ex_22_),
    .X(net196));
 sg13g2_mux2_1 \register_file_i/_5921_  (.A0(\register_file_i/rf_reg_1006_ ),
    .A1(net750),
    .S(net987),
    .X(\register_file_i/_0006_ ));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(net196));
 sg13g2_mux2_1 \register_file_i/_5923_  (.A0(\register_file_i/rf_reg_1007_ ),
    .A1(net782),
    .S(net987),
    .X(\register_file_i/_0007_ ));
 sg13g2_buf_2 fanout194 (.A(_01326_),
    .X(net194));
 sg13g2_mux2_1 \register_file_i/_5925_  (.A0(\register_file_i/rf_reg_1008_ ),
    .A1(net711),
    .S(net987),
    .X(\register_file_i/_0008_ ));
 sg13g2_buf_8 fanout193 (.A(net194),
    .X(net193));
 sg13g2_mux2_1 \register_file_i/_5927_  (.A0(\register_file_i/rf_reg_1009_ ),
    .A1(net725),
    .S(net987),
    .X(\register_file_i/_0009_ ));
 sg13g2_buf_16 fanout192 (.X(net192),
    .A(net193));
 sg13g2_nand2_2 \register_file_i/_5929_  (.Y(\register_file_i/_2813_ ),
    .A(\id_stage_i.controller_i.instr_i_8_ ),
    .B(net1993));
 sg13g2_nor2b_1 \register_file_i/_5930_  (.A(net553),
    .B_N(rf_we_wb),
    .Y(\register_file_i/_2814_ ));
 sg13g2_nor2_1 \register_file_i/_5931_  (.A(net1991),
    .B(net2099),
    .Y(\register_file_i/_2815_ ));
 sg13g2_and2_1 \register_file_i/_5932_  (.A(\register_file_i/_2814_ ),
    .B(\register_file_i/_2815_ ),
    .X(\register_file_i/_2816_ ));
 sg13g2_nand2b_2 \register_file_i/_5933_  (.Y(\register_file_i/_2817_ ),
    .B(\register_file_i/_2816_ ),
    .A_N(\register_file_i/_2813_ ));
 sg13g2_buf_2 fanout191 (.A(_01763_),
    .X(net191));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5936_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_100_ ),
    .S(net871),
    .X(\register_file_i/_0010_ ));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(net191));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5939_  (.A0(\register_file_i/rf_reg_1010_ ),
    .A1(net705),
    .S(net988),
    .X(\register_file_i/_0011_ ));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5941_  (.A0(\register_file_i/rf_reg_1011_ ),
    .A1(net700),
    .S(net988),
    .X(\register_file_i/_0012_ ));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5943_  (.A0(\register_file_i/rf_reg_1012_ ),
    .A1(net739),
    .S(net987),
    .X(\register_file_i/_0013_ ));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5945_  (.A0(\register_file_i/rf_reg_1013_ ),
    .A1(net674),
    .S(net987),
    .X(\register_file_i/_0014_ ));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5947_  (.A0(\register_file_i/rf_reg_1014_ ),
    .A1(net695),
    .S(net989),
    .X(\register_file_i/_0015_ ));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(net191));
 sg13g2_mux2_1 \register_file_i/_5949_  (.A0(\register_file_i/rf_reg_1015_ ),
    .A1(net687),
    .S(net987),
    .X(\register_file_i/_0016_ ));
 sg13g2_buf_2 fanout182 (.A(net1347),
    .X(net182));
 sg13g2_mux2_1 \register_file_i/_5951_  (.A0(\register_file_i/rf_reg_1016_ ),
    .A1(net685),
    .S(net989),
    .X(\register_file_i/_0017_ ));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(net1347));
 sg13g2_mux2_1 \register_file_i/_5953_  (.A0(\register_file_i/rf_reg_1017_ ),
    .A1(net603),
    .S(net989),
    .X(\register_file_i/_0018_ ));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net1348));
 sg13g2_mux2_1 \register_file_i/_5955_  (.A0(\register_file_i/rf_reg_1018_ ),
    .A1(net667),
    .S(net990),
    .X(\register_file_i/_0019_ ));
 sg13g2_buf_2 fanout179 (.A(net1347),
    .X(net179));
 sg13g2_mux2_1 \register_file_i/_5957_  (.A0(\register_file_i/rf_reg_1019_ ),
    .A1(net584),
    .S(net985),
    .X(\register_file_i/_0020_ ));
 sg13g2_buf_2 fanout178 (.A(_01814_),
    .X(net178));
 sg13g2_mux2_1 \register_file_i/_5959_  (.A0(net998),
    .A1(\register_file_i/rf_reg_101_ ),
    .S(net871),
    .X(\register_file_i/_0021_ ));
 sg13g2_buf_4 fanout177 (.X(net177),
    .A(net1347));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net1347));
 sg13g2_mux2_1 \register_file_i/_5962_  (.A0(\register_file_i/rf_reg_1020_ ),
    .A1(net579),
    .S(net986),
    .X(\register_file_i/_0022_ ));
 sg13g2_buf_2 fanout175 (.A(net1347),
    .X(net175));
 sg13g2_mux2_1 \register_file_i/_5964_  (.A0(\register_file_i/rf_reg_1021_ ),
    .A1(net570),
    .S(net990),
    .X(\register_file_i/_0023_ ));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net1348));
 sg13g2_mux2_1 \register_file_i/_5966_  (.A0(\register_file_i/rf_reg_1022_ ),
    .A1(net574),
    .S(net988),
    .X(\register_file_i/_0024_ ));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net1347));
 sg13g2_mux2_1 \register_file_i/_5968_  (.A0(\register_file_i/rf_reg_1023_ ),
    .A1(net564),
    .S(net988),
    .X(\register_file_i/_0025_ ));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net1347));
 sg13g2_mux2_1 \register_file_i/_5970_  (.A0(net883),
    .A1(\register_file_i/rf_reg_102_ ),
    .S(net871),
    .X(\register_file_i/_0026_ ));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net1348));
 sg13g2_mux2_1 \register_file_i/_5972_  (.A0(net994),
    .A1(\register_file_i/rf_reg_103_ ),
    .S(net871),
    .X(\register_file_i/_0027_ ));
 sg13g2_buf_1 fanout170 (.A(_02686_),
    .X(net170));
 sg13g2_mux2_1 \register_file_i/_5974_  (.A0(net878),
    .A1(\register_file_i/rf_reg_104_ ),
    .S(net871),
    .X(\register_file_i/_0028_ ));
 sg13g2_buf_2 fanout169 (.A(_02686_),
    .X(net169));
 sg13g2_mux2_1 \register_file_i/_5976_  (.A0(net807),
    .A1(\register_file_i/rf_reg_105_ ),
    .S(net869),
    .X(\register_file_i/_0029_ ));
 sg13g2_buf_4 fanout168 (.X(net168),
    .A(_04289_));
 sg13g2_mux2_1 \register_file_i/_5978_  (.A0(net798),
    .A1(\register_file_i/rf_reg_106_ ),
    .S(net869),
    .X(\register_file_i/_0030_ ));
 sg13g2_buf_4 fanout167 (.X(net167),
    .A(_04289_));
 sg13g2_mux2_1 \register_file_i/_5980_  (.A0(net793),
    .A1(\register_file_i/rf_reg_107_ ),
    .S(net869),
    .X(\register_file_i/_0031_ ));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(_04289_));
 sg13g2_mux2_1 \register_file_i/_5982_  (.A0(net802),
    .A1(\register_file_i/rf_reg_108_ ),
    .S(net869),
    .X(\register_file_i/_0032_ ));
 sg13g2_buf_2 fanout165 (.A(_04317_),
    .X(net165));
 sg13g2_mux2_1 \register_file_i/_5984_  (.A0(net789),
    .A1(\register_file_i/rf_reg_109_ ),
    .S(net869),
    .X(\register_file_i/_0033_ ));
 sg13g2_buf_2 fanout164 (.A(_04317_),
    .X(net164));
 sg13g2_buf_2 fanout163 (.A(_04438_),
    .X(net163));
 sg13g2_mux2_1 \register_file_i/_5987_  (.A0(net751),
    .A1(\register_file_i/rf_reg_110_ ),
    .S(net873),
    .X(\register_file_i/_0034_ ));
 sg13g2_buf_2 fanout162 (.A(_04438_),
    .X(net162));
 sg13g2_mux2_1 \register_file_i/_5989_  (.A0(net783),
    .A1(\register_file_i/rf_reg_111_ ),
    .S(net873),
    .X(\register_file_i/_0035_ ));
 sg13g2_buf_2 fanout161 (.A(_04589_),
    .X(net161));
 sg13g2_mux2_1 \register_file_i/_5991_  (.A0(net710),
    .A1(\register_file_i/rf_reg_112_ ),
    .S(net873),
    .X(\register_file_i/_0036_ ));
 sg13g2_buf_2 fanout160 (.A(_04589_),
    .X(net160));
 sg13g2_mux2_1 \register_file_i/_5993_  (.A0(net726),
    .A1(\register_file_i/rf_reg_113_ ),
    .S(net874),
    .X(\register_file_i/_0037_ ));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(_04593_));
 sg13g2_mux2_1 \register_file_i/_5995_  (.A0(net706),
    .A1(\register_file_i/rf_reg_114_ ),
    .S(net873),
    .X(\register_file_i/_0038_ ));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net159));
 sg13g2_mux2_1 \register_file_i/_5997_  (.A0(net701),
    .A1(\register_file_i/rf_reg_115_ ),
    .S(net874),
    .X(\register_file_i/_0039_ ));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net159));
 sg13g2_mux2_1 \register_file_i/_5999_  (.A0(rf_wdata_wb_20_),
    .A1(\register_file_i/rf_reg_116_ ),
    .S(net873),
    .X(\register_file_i/_0040_ ));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net159));
 sg13g2_mux2_1 \register_file_i/_6001_  (.A0(net673),
    .A1(\register_file_i/rf_reg_117_ ),
    .S(net873),
    .X(\register_file_i/_0041_ ));
 sg13g2_buf_2 fanout155 (.A(\cs_registers_i/_1421_ ),
    .X(net155));
 sg13g2_mux2_1 \register_file_i/_6003_  (.A0(net695),
    .A1(\register_file_i/rf_reg_118_ ),
    .S(net873),
    .X(\register_file_i/_0042_ ));
 sg13g2_buf_2 fanout154 (.A(net155),
    .X(net154));
 sg13g2_mux2_1 \register_file_i/_6005_  (.A0(net692),
    .A1(\register_file_i/rf_reg_119_ ),
    .S(net870),
    .X(\register_file_i/_0043_ ));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(net155));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_01210_));
 sg13g2_mux2_1 \register_file_i/_6008_  (.A0(net686),
    .A1(\register_file_i/rf_reg_120_ ),
    .S(net870),
    .X(\register_file_i/_0044_ ));
 sg13g2_buf_8 fanout151 (.A(net152),
    .X(net151));
 sg13g2_mux2_1 \register_file_i/_6010_  (.A0(net602),
    .A1(\register_file_i/rf_reg_121_ ),
    .S(net872),
    .X(\register_file_i/_0045_ ));
 sg13g2_buf_4 fanout150 (.X(net150),
    .A(alu_operand_a_ex_23_));
 sg13g2_mux2_1 \register_file_i/_6012_  (.A0(net668),
    .A1(\register_file_i/rf_reg_122_ ),
    .S(net871),
    .X(\register_file_i/_0046_ ));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_mux2_1 \register_file_i/_6014_  (.A0(net585),
    .A1(\register_file_i/rf_reg_123_ ),
    .S(net871),
    .X(\register_file_i/_0047_ ));
 sg13g2_buf_16 fanout148 (.X(net148),
    .A(alu_operand_a_ex_7_));
 sg13g2_mux2_1 \register_file_i/_6016_  (.A0(net580),
    .A1(\register_file_i/rf_reg_124_ ),
    .S(net871),
    .X(\register_file_i/_0048_ ));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(csr_addr_7_));
 sg13g2_mux2_1 \register_file_i/_6018_  (.A0(net572),
    .A1(\register_file_i/rf_reg_125_ ),
    .S(net869),
    .X(\register_file_i/_0049_ ));
 sg13g2_buf_2 fanout146 (.A(net147),
    .X(net146));
 sg13g2_mux2_1 \register_file_i/_6020_  (.A0(rf_wdata_wb_30_),
    .A1(\register_file_i/rf_reg_126_ ),
    .S(net874),
    .X(\register_file_i/_0050_ ));
 sg13g2_buf_4 fanout145 (.X(net145),
    .A(net146));
 sg13g2_mux2_1 \register_file_i/_6022_  (.A0(net565),
    .A1(\register_file_i/rf_reg_127_ ),
    .S(net873),
    .X(\register_file_i/_0051_ ));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net146));
 sg13g2_nor2_2 \register_file_i/_6024_  (.A(\id_stage_i.controller_i.instr_i_8_ ),
    .B(net1993),
    .Y(\register_file_i/_2866_ ));
 sg13g2_nand2b_2 \register_file_i/_6025_  (.Y(\register_file_i/_2867_ ),
    .B(rf_we_wb),
    .A_N(net553));
 sg13g2_nand2b_2 \register_file_i/_6026_  (.Y(\register_file_i/_2868_ ),
    .B(net1991),
    .A_N(net2099));
 sg13g2_nor2_1 \register_file_i/_6027_  (.A(\register_file_i/_2867_ ),
    .B(\register_file_i/_2868_ ),
    .Y(\register_file_i/_2869_ ));
 sg13g2_nand2_1 \register_file_i/_6028_  (.Y(\register_file_i/_2870_ ),
    .A(\register_file_i/_2866_ ),
    .B(\register_file_i/_2869_ ));
 sg13g2_buf_2 fanout143 (.A(_04032_),
    .X(net143));
 sg13g2_mux2_1 \register_file_i/_6030_  (.A0(net756),
    .A1(\register_file_i/rf_reg_128_ ),
    .S(net865),
    .X(\register_file_i/_0052_ ));
 sg13g2_buf_2 fanout142 (.A(_04032_),
    .X(net142));
 sg13g2_mux2_1 \register_file_i/_6032_  (.A0(net1003),
    .A1(\register_file_i/rf_reg_129_ ),
    .S(net864),
    .X(\register_file_i/_0053_ ));
 sg13g2_buf_2 fanout141 (.A(_04820_),
    .X(net141));
 sg13g2_mux2_1 \register_file_i/_6034_  (.A0(net886),
    .A1(\register_file_i/rf_reg_130_ ),
    .S(net864),
    .X(\register_file_i/_0054_ ));
 sg13g2_buf_1 fanout140 (.A(net141),
    .X(net140));
 sg13g2_mux2_1 \register_file_i/_6036_  (.A0(net1023),
    .A1(\register_file_i/rf_reg_131_ ),
    .S(net864),
    .X(\register_file_i/_0055_ ));
 sg13g2_mux2_1 \register_file_i/_6037_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_132_ ),
    .S(net863),
    .X(\register_file_i/_0056_ ));
 sg13g2_mux2_1 \register_file_i/_6038_  (.A0(net998),
    .A1(\register_file_i/rf_reg_133_ ),
    .S(net863),
    .X(\register_file_i/_0057_ ));
 sg13g2_mux2_1 \register_file_i/_6039_  (.A0(net882),
    .A1(\register_file_i/rf_reg_134_ ),
    .S(net863),
    .X(\register_file_i/_0058_ ));
 sg13g2_mux2_1 \register_file_i/_6040_  (.A0(net993),
    .A1(\register_file_i/rf_reg_135_ ),
    .S(net863),
    .X(\register_file_i/_0059_ ));
 sg13g2_mux2_1 \register_file_i/_6041_  (.A0(net878),
    .A1(\register_file_i/rf_reg_136_ ),
    .S(net863),
    .X(\register_file_i/_0060_ ));
 sg13g2_mux2_1 \register_file_i/_6042_  (.A0(net806),
    .A1(\register_file_i/rf_reg_137_ ),
    .S(net864),
    .X(\register_file_i/_0061_ ));
 sg13g2_buf_4 fanout139 (.X(net139),
    .A(net141));
 sg13g2_mux2_1 \register_file_i/_6044_  (.A0(net797),
    .A1(\register_file_i/rf_reg_138_ ),
    .S(net864),
    .X(\register_file_i/_0062_ ));
 sg13g2_mux2_1 \register_file_i/_6045_  (.A0(net793),
    .A1(\register_file_i/rf_reg_139_ ),
    .S(net863),
    .X(\register_file_i/_0063_ ));
 sg13g2_mux2_1 \register_file_i/_6046_  (.A0(net802),
    .A1(\register_file_i/rf_reg_140_ ),
    .S(net864),
    .X(\register_file_i/_0064_ ));
 sg13g2_mux2_1 \register_file_i/_6047_  (.A0(net789),
    .A1(\register_file_i/rf_reg_141_ ),
    .S(net865),
    .X(\register_file_i/_0065_ ));
 sg13g2_mux2_1 \register_file_i/_6048_  (.A0(net751),
    .A1(\register_file_i/rf_reg_142_ ),
    .S(net865),
    .X(\register_file_i/_0066_ ));
 sg13g2_mux2_1 \register_file_i/_6049_  (.A0(net783),
    .A1(\register_file_i/rf_reg_143_ ),
    .S(net866),
    .X(\register_file_i/_0067_ ));
 sg13g2_mux2_1 \register_file_i/_6050_  (.A0(net710),
    .A1(\register_file_i/rf_reg_144_ ),
    .S(net865),
    .X(\register_file_i/_0068_ ));
 sg13g2_mux2_1 \register_file_i/_6051_  (.A0(net726),
    .A1(\register_file_i/rf_reg_145_ ),
    .S(net866),
    .X(\register_file_i/_0069_ ));
 sg13g2_mux2_1 \register_file_i/_6052_  (.A0(net706),
    .A1(\register_file_i/rf_reg_146_ ),
    .S(net865),
    .X(\register_file_i/_0070_ ));
 sg13g2_mux2_1 \register_file_i/_6053_  (.A0(net701),
    .A1(\register_file_i/rf_reg_147_ ),
    .S(net865),
    .X(\register_file_i/_0071_ ));
 sg13g2_buf_2 fanout138 (.A(_05064_),
    .X(net138));
 sg13g2_mux2_1 \register_file_i/_6055_  (.A0(net740),
    .A1(\register_file_i/rf_reg_148_ ),
    .S(net866),
    .X(\register_file_i/_0072_ ));
 sg13g2_mux2_1 \register_file_i/_6056_  (.A0(net673),
    .A1(\register_file_i/rf_reg_149_ ),
    .S(net866),
    .X(\register_file_i/_0073_ ));
 sg13g2_mux2_1 \register_file_i/_6057_  (.A0(net696),
    .A1(\register_file_i/rf_reg_150_ ),
    .S(net867),
    .X(\register_file_i/_0074_ ));
 sg13g2_mux2_1 \register_file_i/_6058_  (.A0(net692),
    .A1(\register_file_i/rf_reg_151_ ),
    .S(net864),
    .X(\register_file_i/_0075_ ));
 sg13g2_mux2_1 \register_file_i/_6059_  (.A0(net686),
    .A1(\register_file_i/rf_reg_152_ ),
    .S(net867),
    .X(\register_file_i/_0076_ ));
 sg13g2_mux2_1 \register_file_i/_6060_  (.A0(net602),
    .A1(\register_file_i/rf_reg_153_ ),
    .S(net868),
    .X(\register_file_i/_0077_ ));
 sg13g2_mux2_1 \register_file_i/_6061_  (.A0(net667),
    .A1(\register_file_i/rf_reg_154_ ),
    .S(net868),
    .X(\register_file_i/_0078_ ));
 sg13g2_mux2_1 \register_file_i/_6062_  (.A0(net585),
    .A1(\register_file_i/rf_reg_155_ ),
    .S(net863),
    .X(\register_file_i/_0079_ ));
 sg13g2_mux2_1 \register_file_i/_6063_  (.A0(net580),
    .A1(\register_file_i/rf_reg_156_ ),
    .S(net863),
    .X(\register_file_i/_0080_ ));
 sg13g2_mux2_1 \register_file_i/_6064_  (.A0(net570),
    .A1(\register_file_i/rf_reg_157_ ),
    .S(net864),
    .X(\register_file_i/_0081_ ));
 sg13g2_mux2_1 \register_file_i/_6065_  (.A0(rf_wdata_wb_30_),
    .A1(\register_file_i/rf_reg_158_ ),
    .S(net865),
    .X(\register_file_i/_0082_ ));
 sg13g2_mux2_1 \register_file_i/_6066_  (.A0(net565),
    .A1(\register_file_i/rf_reg_159_ ),
    .S(net865),
    .X(\register_file_i/_0083_ ));
 sg13g2_inv_1 \register_file_i/_6067_  (.Y(\register_file_i/_2877_ ),
    .A(net1993));
 sg13g2_nor2_2 \register_file_i/_6068_  (.A(\id_stage_i.controller_i.instr_i_8_ ),
    .B(\register_file_i/_2877_ ),
    .Y(\register_file_i/_2878_ ));
 sg13g2_nand2_1 \register_file_i/_6069_  (.Y(\register_file_i/_2879_ ),
    .A(\register_file_i/_2869_ ),
    .B(\register_file_i/_2878_ ));
 sg13g2_buf_4 fanout137 (.X(net137),
    .A(net138));
 sg13g2_mux2_1 \register_file_i/_6071_  (.A0(net756),
    .A1(\register_file_i/rf_reg_160_ ),
    .S(net859),
    .X(\register_file_i/_0084_ ));
 sg13g2_mux2_1 \register_file_i/_6072_  (.A0(net1002),
    .A1(\register_file_i/rf_reg_161_ ),
    .S(net858),
    .X(\register_file_i/_0085_ ));
 sg13g2_mux2_1 \register_file_i/_6073_  (.A0(net886),
    .A1(\register_file_i/rf_reg_162_ ),
    .S(net858),
    .X(\register_file_i/_0086_ ));
 sg13g2_mux2_1 \register_file_i/_6074_  (.A0(net1023),
    .A1(\register_file_i/rf_reg_163_ ),
    .S(net858),
    .X(\register_file_i/_0087_ ));
 sg13g2_mux2_1 \register_file_i/_6075_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_164_ ),
    .S(net857),
    .X(\register_file_i/_0088_ ));
 sg13g2_mux2_1 \register_file_i/_6076_  (.A0(net997),
    .A1(\register_file_i/rf_reg_165_ ),
    .S(net857),
    .X(\register_file_i/_0089_ ));
 sg13g2_mux2_1 \register_file_i/_6077_  (.A0(net882),
    .A1(\register_file_i/rf_reg_166_ ),
    .S(net857),
    .X(\register_file_i/_0090_ ));
 sg13g2_mux2_1 \register_file_i/_6078_  (.A0(net993),
    .A1(\register_file_i/rf_reg_167_ ),
    .S(net857),
    .X(\register_file_i/_0091_ ));
 sg13g2_mux2_1 \register_file_i/_6079_  (.A0(net878),
    .A1(\register_file_i/rf_reg_168_ ),
    .S(net857),
    .X(\register_file_i/_0092_ ));
 sg13g2_mux2_1 \register_file_i/_6080_  (.A0(net807),
    .A1(\register_file_i/rf_reg_169_ ),
    .S(net858),
    .X(\register_file_i/_0093_ ));
 sg13g2_buf_2 fanout136 (.A(_05296_),
    .X(net136));
 sg13g2_mux2_1 \register_file_i/_6082_  (.A0(net798),
    .A1(\register_file_i/rf_reg_170_ ),
    .S(net858),
    .X(\register_file_i/_0094_ ));
 sg13g2_mux2_1 \register_file_i/_6083_  (.A0(net793),
    .A1(\register_file_i/rf_reg_171_ ),
    .S(net857),
    .X(\register_file_i/_0095_ ));
 sg13g2_mux2_1 \register_file_i/_6084_  (.A0(net802),
    .A1(\register_file_i/rf_reg_172_ ),
    .S(net858),
    .X(\register_file_i/_0096_ ));
 sg13g2_mux2_1 \register_file_i/_6085_  (.A0(net789),
    .A1(\register_file_i/rf_reg_173_ ),
    .S(net859),
    .X(\register_file_i/_0097_ ));
 sg13g2_mux2_1 \register_file_i/_6086_  (.A0(net751),
    .A1(\register_file_i/rf_reg_174_ ),
    .S(net859),
    .X(\register_file_i/_0098_ ));
 sg13g2_mux2_1 \register_file_i/_6087_  (.A0(net783),
    .A1(\register_file_i/rf_reg_175_ ),
    .S(net860),
    .X(\register_file_i/_0099_ ));
 sg13g2_mux2_1 \register_file_i/_6088_  (.A0(net710),
    .A1(\register_file_i/rf_reg_176_ ),
    .S(net859),
    .X(\register_file_i/_0100_ ));
 sg13g2_mux2_1 \register_file_i/_6089_  (.A0(net726),
    .A1(\register_file_i/rf_reg_177_ ),
    .S(net860),
    .X(\register_file_i/_0101_ ));
 sg13g2_mux2_1 \register_file_i/_6090_  (.A0(net706),
    .A1(\register_file_i/rf_reg_178_ ),
    .S(net860),
    .X(\register_file_i/_0102_ ));
 sg13g2_mux2_1 \register_file_i/_6091_  (.A0(net701),
    .A1(\register_file_i/rf_reg_179_ ),
    .S(net859),
    .X(\register_file_i/_0103_ ));
 sg13g2_buf_2 fanout135 (.A(net136),
    .X(net135));
 sg13g2_mux2_1 \register_file_i/_6093_  (.A0(net740),
    .A1(\register_file_i/rf_reg_180_ ),
    .S(net860),
    .X(\register_file_i/_0104_ ));
 sg13g2_mux2_1 \register_file_i/_6094_  (.A0(net673),
    .A1(\register_file_i/rf_reg_181_ ),
    .S(net860),
    .X(\register_file_i/_0105_ ));
 sg13g2_mux2_1 \register_file_i/_6095_  (.A0(net696),
    .A1(\register_file_i/rf_reg_182_ ),
    .S(net859),
    .X(\register_file_i/_0106_ ));
 sg13g2_mux2_1 \register_file_i/_6096_  (.A0(net692),
    .A1(\register_file_i/rf_reg_183_ ),
    .S(net858),
    .X(\register_file_i/_0107_ ));
 sg13g2_mux2_1 \register_file_i/_6097_  (.A0(net686),
    .A1(\register_file_i/rf_reg_184_ ),
    .S(net861),
    .X(\register_file_i/_0108_ ));
 sg13g2_mux2_1 \register_file_i/_6098_  (.A0(net602),
    .A1(\register_file_i/rf_reg_185_ ),
    .S(net861),
    .X(\register_file_i/_0109_ ));
 sg13g2_mux2_1 \register_file_i/_6099_  (.A0(net667),
    .A1(\register_file_i/rf_reg_186_ ),
    .S(net862),
    .X(\register_file_i/_0110_ ));
 sg13g2_mux2_1 \register_file_i/_6100_  (.A0(net585),
    .A1(\register_file_i/rf_reg_187_ ),
    .S(net857),
    .X(\register_file_i/_0111_ ));
 sg13g2_mux2_1 \register_file_i/_6101_  (.A0(net579),
    .A1(\register_file_i/rf_reg_188_ ),
    .S(net857),
    .X(\register_file_i/_0112_ ));
 sg13g2_mux2_1 \register_file_i/_6102_  (.A0(net572),
    .A1(\register_file_i/rf_reg_189_ ),
    .S(net858),
    .X(\register_file_i/_0113_ ));
 sg13g2_mux2_1 \register_file_i/_6103_  (.A0(net576),
    .A1(\register_file_i/rf_reg_190_ ),
    .S(net859),
    .X(\register_file_i/_0114_ ));
 sg13g2_mux2_1 \register_file_i/_6104_  (.A0(net565),
    .A1(\register_file_i/rf_reg_191_ ),
    .S(net859),
    .X(\register_file_i/_0115_ ));
 sg13g2_inv_1 \register_file_i/_6105_  (.Y(\register_file_i/_2883_ ),
    .A(\id_stage_i.controller_i.instr_i_8_ ));
 sg13g2_nor2_2 \register_file_i/_6106_  (.A(\register_file_i/_2883_ ),
    .B(net1993),
    .Y(\register_file_i/_2884_ ));
 sg13g2_nand2_1 \register_file_i/_6107_  (.Y(\register_file_i/_2885_ ),
    .A(\register_file_i/_2869_ ),
    .B(\register_file_i/_2884_ ));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net136));
 sg13g2_mux2_1 \register_file_i/_6109_  (.A0(net756),
    .A1(\register_file_i/rf_reg_192_ ),
    .S(net854),
    .X(\register_file_i/_0116_ ));
 sg13g2_mux2_1 \register_file_i/_6110_  (.A0(net1003),
    .A1(\register_file_i/rf_reg_193_ ),
    .S(net852),
    .X(\register_file_i/_0117_ ));
 sg13g2_mux2_1 \register_file_i/_6111_  (.A0(net886),
    .A1(\register_file_i/rf_reg_194_ ),
    .S(net852),
    .X(\register_file_i/_0118_ ));
 sg13g2_mux2_1 \register_file_i/_6112_  (.A0(net1024),
    .A1(\register_file_i/rf_reg_195_ ),
    .S(net852),
    .X(\register_file_i/_0119_ ));
 sg13g2_mux2_1 \register_file_i/_6113_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_196_ ),
    .S(net853),
    .X(\register_file_i/_0120_ ));
 sg13g2_mux2_1 \register_file_i/_6114_  (.A0(net998),
    .A1(\register_file_i/rf_reg_197_ ),
    .S(net853),
    .X(\register_file_i/_0121_ ));
 sg13g2_mux2_1 \register_file_i/_6115_  (.A0(net883),
    .A1(\register_file_i/rf_reg_198_ ),
    .S(net853),
    .X(\register_file_i/_0122_ ));
 sg13g2_mux2_1 \register_file_i/_6116_  (.A0(net994),
    .A1(\register_file_i/rf_reg_199_ ),
    .S(net853),
    .X(\register_file_i/_0123_ ));
 sg13g2_mux2_1 \register_file_i/_6117_  (.A0(net879),
    .A1(\register_file_i/rf_reg_200_ ),
    .S(net852),
    .X(\register_file_i/_0124_ ));
 sg13g2_mux2_1 \register_file_i/_6118_  (.A0(net807),
    .A1(\register_file_i/rf_reg_201_ ),
    .S(net852),
    .X(\register_file_i/_0125_ ));
 sg13g2_buf_1 fanout133 (.A(_08523_),
    .X(net133));
 sg13g2_mux2_1 \register_file_i/_6120_  (.A0(net798),
    .A1(\register_file_i/rf_reg_202_ ),
    .S(net852),
    .X(\register_file_i/_0126_ ));
 sg13g2_mux2_1 \register_file_i/_6121_  (.A0(net793),
    .A1(\register_file_i/rf_reg_203_ ),
    .S(net852),
    .X(\register_file_i/_0127_ ));
 sg13g2_mux2_1 \register_file_i/_6122_  (.A0(net802),
    .A1(\register_file_i/rf_reg_204_ ),
    .S(net852),
    .X(\register_file_i/_0128_ ));
 sg13g2_mux2_1 \register_file_i/_6123_  (.A0(net789),
    .A1(\register_file_i/rf_reg_205_ ),
    .S(net854),
    .X(\register_file_i/_0129_ ));
 sg13g2_mux2_1 \register_file_i/_6124_  (.A0(net751),
    .A1(\register_file_i/rf_reg_206_ ),
    .S(net854),
    .X(\register_file_i/_0130_ ));
 sg13g2_mux2_1 \register_file_i/_6125_  (.A0(net783),
    .A1(\register_file_i/rf_reg_207_ ),
    .S(net854),
    .X(\register_file_i/_0131_ ));
 sg13g2_mux2_1 \register_file_i/_6126_  (.A0(net710),
    .A1(\register_file_i/rf_reg_208_ ),
    .S(net854),
    .X(\register_file_i/_0132_ ));
 sg13g2_mux2_1 \register_file_i/_6127_  (.A0(net726),
    .A1(\register_file_i/rf_reg_209_ ),
    .S(net855),
    .X(\register_file_i/_0133_ ));
 sg13g2_mux2_1 \register_file_i/_6128_  (.A0(net706),
    .A1(\register_file_i/rf_reg_210_ ),
    .S(net854),
    .X(\register_file_i/_0134_ ));
 sg13g2_mux2_1 \register_file_i/_6129_  (.A0(net701),
    .A1(\register_file_i/rf_reg_211_ ),
    .S(net855),
    .X(\register_file_i/_0135_ ));
 sg13g2_buf_1 fanout132 (.A(net133),
    .X(net132));
 sg13g2_mux2_1 \register_file_i/_6131_  (.A0(net740),
    .A1(\register_file_i/rf_reg_212_ ),
    .S(net855),
    .X(\register_file_i/_0136_ ));
 sg13g2_mux2_1 \register_file_i/_6132_  (.A0(net673),
    .A1(\register_file_i/rf_reg_213_ ),
    .S(net855),
    .X(\register_file_i/_0137_ ));
 sg13g2_mux2_1 \register_file_i/_6133_  (.A0(net695),
    .A1(\register_file_i/rf_reg_214_ ),
    .S(net854),
    .X(\register_file_i/_0138_ ));
 sg13g2_mux2_1 \register_file_i/_6134_  (.A0(net692),
    .A1(\register_file_i/rf_reg_215_ ),
    .S(net853),
    .X(\register_file_i/_0139_ ));
 sg13g2_mux2_1 \register_file_i/_6135_  (.A0(net686),
    .A1(\register_file_i/rf_reg_216_ ),
    .S(net856),
    .X(\register_file_i/_0140_ ));
 sg13g2_mux2_1 \register_file_i/_6136_  (.A0(net602),
    .A1(\register_file_i/rf_reg_217_ ),
    .S(net853),
    .X(\register_file_i/_0141_ ));
 sg13g2_mux2_1 \register_file_i/_6137_  (.A0(net667),
    .A1(\register_file_i/rf_reg_218_ ),
    .S(net856),
    .X(\register_file_i/_0142_ ));
 sg13g2_mux2_1 \register_file_i/_6138_  (.A0(net585),
    .A1(\register_file_i/rf_reg_219_ ),
    .S(net856),
    .X(\register_file_i/_0143_ ));
 sg13g2_mux2_1 \register_file_i/_6139_  (.A0(net579),
    .A1(\register_file_i/rf_reg_220_ ),
    .S(net856),
    .X(\register_file_i/_0144_ ));
 sg13g2_mux2_1 \register_file_i/_6140_  (.A0(net570),
    .A1(\register_file_i/rf_reg_221_ ),
    .S(net853),
    .X(\register_file_i/_0145_ ));
 sg13g2_mux2_1 \register_file_i/_6141_  (.A0(net576),
    .A1(\register_file_i/rf_reg_222_ ),
    .S(net855),
    .X(\register_file_i/_0146_ ));
 sg13g2_mux2_1 \register_file_i/_6142_  (.A0(net565),
    .A1(\register_file_i/rf_reg_223_ ),
    .S(net854),
    .X(\register_file_i/_0147_ ));
 sg13g2_buf_2 fanout131 (.A(net133),
    .X(net131));
 sg13g2_nor3_1 \register_file_i/_6144_  (.A(\register_file_i/_2813_ ),
    .B(\register_file_i/_2867_ ),
    .C(\register_file_i/_2868_ ),
    .Y(\register_file_i/_2890_ ));
 sg13g2_buf_2 fanout130 (.A(net133),
    .X(net130));
 sg13g2_mux2_1 \register_file_i/_6146_  (.A0(\register_file_i/rf_reg_224_ ),
    .A1(net756),
    .S(net980),
    .X(\register_file_i/_0148_ ));
 sg13g2_buf_1 fanout129 (.A(net133),
    .X(net129));
 sg13g2_mux2_1 \register_file_i/_6148_  (.A0(\register_file_i/rf_reg_225_ ),
    .A1(net1003),
    .S(net979),
    .X(\register_file_i/_0149_ ));
 sg13g2_buf_2 fanout128 (.A(net133),
    .X(net128));
 sg13g2_mux2_1 \register_file_i/_6150_  (.A0(\register_file_i/rf_reg_226_ ),
    .A1(net887),
    .S(net979),
    .X(\register_file_i/_0150_ ));
 sg13g2_buf_2 fanout127 (.A(alu_operand_a_ex_21_),
    .X(net127));
 sg13g2_mux2_1 \register_file_i/_6152_  (.A0(\register_file_i/rf_reg_227_ ),
    .A1(net1024),
    .S(net979),
    .X(\register_file_i/_0151_ ));
 sg13g2_buf_4 fanout126 (.X(net126),
    .A(alu_operand_a_ex_21_));
 sg13g2_mux2_1 \register_file_i/_6154_  (.A0(\register_file_i/rf_reg_228_ ),
    .A1(net1018),
    .S(net981),
    .X(\register_file_i/_0152_ ));
 sg13g2_buf_4 fanout125 (.X(net125),
    .A(alu_operand_a_ex_24_));
 sg13g2_mux2_1 \register_file_i/_6156_  (.A0(\register_file_i/rf_reg_229_ ),
    .A1(net998),
    .S(net981),
    .X(\register_file_i/_0153_ ));
 sg13g2_buf_2 fanout124 (.A(_01280_),
    .X(net124));
 sg13g2_mux2_1 \register_file_i/_6158_  (.A0(\register_file_i/rf_reg_230_ ),
    .A1(net883),
    .S(net981),
    .X(\register_file_i/_0154_ ));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123));
 sg13g2_mux2_1 \register_file_i/_6160_  (.A0(\register_file_i/rf_reg_231_ ),
    .A1(net994),
    .S(net981),
    .X(\register_file_i/_0155_ ));
 sg13g2_mux2_1 \register_file_i/_6161_  (.A0(\register_file_i/rf_reg_232_ ),
    .A1(net879),
    .S(net979),
    .X(\register_file_i/_0156_ ));
 sg13g2_mux2_1 \register_file_i/_6162_  (.A0(\register_file_i/rf_reg_233_ ),
    .A1(net806),
    .S(net979),
    .X(\register_file_i/_0157_ ));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(net124));
 sg13g2_mux2_1 \register_file_i/_6164_  (.A0(\register_file_i/rf_reg_234_ ),
    .A1(net798),
    .S(net979),
    .X(\register_file_i/_0158_ ));
 sg13g2_mux2_1 \register_file_i/_6165_  (.A0(\register_file_i/rf_reg_235_ ),
    .A1(net793),
    .S(net979),
    .X(\register_file_i/_0159_ ));
 sg13g2_mux2_1 \register_file_i/_6166_  (.A0(\register_file_i/rf_reg_236_ ),
    .A1(net802),
    .S(net979),
    .X(\register_file_i/_0160_ ));
 sg13g2_mux2_1 \register_file_i/_6167_  (.A0(\register_file_i/rf_reg_237_ ),
    .A1(net789),
    .S(net982),
    .X(\register_file_i/_0161_ ));
 sg13g2_mux2_1 \register_file_i/_6168_  (.A0(\register_file_i/rf_reg_238_ ),
    .A1(net751),
    .S(net982),
    .X(\register_file_i/_0162_ ));
 sg13g2_mux2_1 \register_file_i/_6169_  (.A0(\register_file_i/rf_reg_239_ ),
    .A1(net783),
    .S(net982),
    .X(\register_file_i/_0163_ ));
 sg13g2_mux2_1 \register_file_i/_6170_  (.A0(\register_file_i/rf_reg_240_ ),
    .A1(net710),
    .S(net982),
    .X(\register_file_i/_0164_ ));
 sg13g2_mux2_1 \register_file_i/_6171_  (.A0(\register_file_i/rf_reg_241_ ),
    .A1(net726),
    .S(net983),
    .X(\register_file_i/_0165_ ));
 sg13g2_mux2_1 \register_file_i/_6172_  (.A0(\register_file_i/rf_reg_242_ ),
    .A1(net706),
    .S(net983),
    .X(\register_file_i/_0166_ ));
 sg13g2_mux2_1 \register_file_i/_6173_  (.A0(\register_file_i/rf_reg_243_ ),
    .A1(net701),
    .S(net982),
    .X(\register_file_i/_0167_ ));
 sg13g2_buf_8 fanout121 (.A(_01469_),
    .X(net121));
 sg13g2_mux2_1 \register_file_i/_6175_  (.A0(\register_file_i/rf_reg_244_ ),
    .A1(net740),
    .S(net983),
    .X(\register_file_i/_0168_ ));
 sg13g2_mux2_1 \register_file_i/_6176_  (.A0(\register_file_i/rf_reg_245_ ),
    .A1(net673),
    .S(net983),
    .X(\register_file_i/_0169_ ));
 sg13g2_mux2_1 \register_file_i/_6177_  (.A0(\register_file_i/rf_reg_246_ ),
    .A1(net695),
    .S(net982),
    .X(\register_file_i/_0170_ ));
 sg13g2_mux2_1 \register_file_i/_6178_  (.A0(\register_file_i/rf_reg_247_ ),
    .A1(net692),
    .S(net980),
    .X(\register_file_i/_0171_ ));
 sg13g2_mux2_1 \register_file_i/_6179_  (.A0(\register_file_i/rf_reg_248_ ),
    .A1(net686),
    .S(net984),
    .X(\register_file_i/_0172_ ));
 sg13g2_mux2_1 \register_file_i/_6180_  (.A0(\register_file_i/rf_reg_249_ ),
    .A1(net602),
    .S(net980),
    .X(\register_file_i/_0173_ ));
 sg13g2_mux2_1 \register_file_i/_6181_  (.A0(\register_file_i/rf_reg_250_ ),
    .A1(net667),
    .S(net984),
    .X(\register_file_i/_0174_ ));
 sg13g2_mux2_1 \register_file_i/_6182_  (.A0(\register_file_i/rf_reg_251_ ),
    .A1(net585),
    .S(net981),
    .X(\register_file_i/_0175_ ));
 sg13g2_mux2_1 \register_file_i/_6183_  (.A0(\register_file_i/rf_reg_252_ ),
    .A1(net579),
    .S(net981),
    .X(\register_file_i/_0176_ ));
 sg13g2_mux2_1 \register_file_i/_6184_  (.A0(\register_file_i/rf_reg_253_ ),
    .A1(net570),
    .S(net980),
    .X(\register_file_i/_0177_ ));
 sg13g2_mux2_1 \register_file_i/_6185_  (.A0(\register_file_i/rf_reg_254_ ),
    .A1(net576),
    .S(net982),
    .X(\register_file_i/_0178_ ));
 sg13g2_mux2_1 \register_file_i/_6186_  (.A0(\register_file_i/rf_reg_255_ ),
    .A1(net565),
    .S(net982),
    .X(\register_file_i/_0179_ ));
 sg13g2_nand2b_2 \register_file_i/_6187_  (.Y(\register_file_i/_2901_ ),
    .B(net2099),
    .A_N(net1991));
 sg13g2_nor2_2 \register_file_i/_6188_  (.A(\register_file_i/_2867_ ),
    .B(\register_file_i/_2901_ ),
    .Y(\register_file_i/_2902_ ));
 sg13g2_nand2_2 \register_file_i/_6189_  (.Y(\register_file_i/_2903_ ),
    .A(\register_file_i/_2866_ ),
    .B(\register_file_i/_2902_ ));
 sg13g2_buf_8 fanout120 (.A(_01469_),
    .X(net120));
 sg13g2_mux2_1 \register_file_i/_6191_  (.A0(net755),
    .A1(\register_file_i/rf_reg_256_ ),
    .S(net848),
    .X(\register_file_i/_0180_ ));
 sg13g2_mux2_1 \register_file_i/_6192_  (.A0(net1002),
    .A1(\register_file_i/rf_reg_257_ ),
    .S(net848),
    .X(\register_file_i/_0181_ ));
 sg13g2_mux2_1 \register_file_i/_6193_  (.A0(net886),
    .A1(\register_file_i/rf_reg_258_ ),
    .S(net848),
    .X(\register_file_i/_0182_ ));
 sg13g2_mux2_1 \register_file_i/_6194_  (.A0(net1021),
    .A1(\register_file_i/rf_reg_259_ ),
    .S(net848),
    .X(\register_file_i/_0183_ ));
 sg13g2_mux2_1 \register_file_i/_6195_  (.A0(net1015),
    .A1(\register_file_i/rf_reg_260_ ),
    .S(net848),
    .X(\register_file_i/_0184_ ));
 sg13g2_mux2_1 \register_file_i/_6196_  (.A0(net995),
    .A1(\register_file_i/rf_reg_261_ ),
    .S(net847),
    .X(\register_file_i/_0185_ ));
 sg13g2_mux2_1 \register_file_i/_6197_  (.A0(net880),
    .A1(\register_file_i/rf_reg_262_ ),
    .S(net848),
    .X(\register_file_i/_0186_ ));
 sg13g2_mux2_1 \register_file_i/_6198_  (.A0(net991),
    .A1(\register_file_i/rf_reg_263_ ),
    .S(net848),
    .X(\register_file_i/_0187_ ));
 sg13g2_mux2_1 \register_file_i/_6199_  (.A0(net875),
    .A1(\register_file_i/rf_reg_264_ ),
    .S(net848),
    .X(\register_file_i/_0188_ ));
 sg13g2_mux2_1 \register_file_i/_6200_  (.A0(net804),
    .A1(\register_file_i/rf_reg_265_ ),
    .S(net847),
    .X(\register_file_i/_0189_ ));
 sg13g2_buf_16 fanout119 (.X(net119),
    .A(net120));
 sg13g2_mux2_1 \register_file_i/_6202_  (.A0(net795),
    .A1(\register_file_i/rf_reg_266_ ),
    .S(net847),
    .X(\register_file_i/_0190_ ));
 sg13g2_mux2_1 \register_file_i/_6203_  (.A0(net790),
    .A1(\register_file_i/rf_reg_267_ ),
    .S(net847),
    .X(\register_file_i/_0191_ ));
 sg13g2_mux2_1 \register_file_i/_6204_  (.A0(net799),
    .A1(\register_file_i/rf_reg_268_ ),
    .S(net847),
    .X(\register_file_i/_0192_ ));
 sg13g2_mux2_1 \register_file_i/_6205_  (.A0(net785),
    .A1(\register_file_i/rf_reg_269_ ),
    .S(net847),
    .X(\register_file_i/_0193_ ));
 sg13g2_mux2_1 \register_file_i/_6206_  (.A0(net747),
    .A1(\register_file_i/rf_reg_270_ ),
    .S(net850),
    .X(\register_file_i/_0194_ ));
 sg13g2_mux2_1 \register_file_i/_6207_  (.A0(net780),
    .A1(\register_file_i/rf_reg_271_ ),
    .S(net850),
    .X(\register_file_i/_0195_ ));
 sg13g2_mux2_1 \register_file_i/_6208_  (.A0(net709),
    .A1(\register_file_i/rf_reg_272_ ),
    .S(net851),
    .X(\register_file_i/_0196_ ));
 sg13g2_mux2_1 \register_file_i/_6209_  (.A0(net724),
    .A1(\register_file_i/rf_reg_273_ ),
    .S(net850),
    .X(\register_file_i/_0197_ ));
 sg13g2_mux2_1 \register_file_i/_6210_  (.A0(net703),
    .A1(\register_file_i/rf_reg_274_ ),
    .S(net850),
    .X(\register_file_i/_0198_ ));
 sg13g2_mux2_1 \register_file_i/_6211_  (.A0(net699),
    .A1(\register_file_i/rf_reg_275_ ),
    .S(net850),
    .X(\register_file_i/_0199_ ));
 sg13g2_buf_2 fanout118 (.A(net120),
    .X(net118));
 sg13g2_mux2_1 \register_file_i/_6213_  (.A0(net737),
    .A1(\register_file_i/rf_reg_276_ ),
    .S(net851),
    .X(\register_file_i/_0200_ ));
 sg13g2_mux2_1 \register_file_i/_6214_  (.A0(net670),
    .A1(\register_file_i/rf_reg_277_ ),
    .S(net851),
    .X(\register_file_i/_0201_ ));
 sg13g2_mux2_1 \register_file_i/_6215_  (.A0(net694),
    .A1(\register_file_i/rf_reg_278_ ),
    .S(net851),
    .X(\register_file_i/_0202_ ));
 sg13g2_mux2_1 \register_file_i/_6216_  (.A0(net689),
    .A1(\register_file_i/rf_reg_279_ ),
    .S(net851),
    .X(\register_file_i/_0203_ ));
 sg13g2_mux2_1 \register_file_i/_6217_  (.A0(net684),
    .A1(\register_file_i/rf_reg_280_ ),
    .S(net850),
    .X(\register_file_i/_0204_ ));
 sg13g2_mux2_1 \register_file_i/_6218_  (.A0(net599),
    .A1(\register_file_i/rf_reg_281_ ),
    .S(net849),
    .X(\register_file_i/_0205_ ));
 sg13g2_mux2_1 \register_file_i/_6219_  (.A0(net665),
    .A1(\register_file_i/rf_reg_282_ ),
    .S(net849),
    .X(\register_file_i/_0206_ ));
 sg13g2_mux2_1 \register_file_i/_6220_  (.A0(net581),
    .A1(\register_file_i/rf_reg_283_ ),
    .S(net847),
    .X(\register_file_i/_0207_ ));
 sg13g2_mux2_1 \register_file_i/_6221_  (.A0(net577),
    .A1(\register_file_i/rf_reg_284_ ),
    .S(net849),
    .X(\register_file_i/_0208_ ));
 sg13g2_mux2_1 \register_file_i/_6222_  (.A0(net567),
    .A1(\register_file_i/rf_reg_285_ ),
    .S(net847),
    .X(\register_file_i/_0209_ ));
 sg13g2_mux2_1 \register_file_i/_6223_  (.A0(net576),
    .A1(\register_file_i/rf_reg_286_ ),
    .S(net850),
    .X(\register_file_i/_0210_ ));
 sg13g2_mux2_1 \register_file_i/_6224_  (.A0(net562),
    .A1(\register_file_i/rf_reg_287_ ),
    .S(net850),
    .X(\register_file_i/_0211_ ));
 sg13g2_nand2_2 \register_file_i/_6225_  (.Y(\register_file_i/_2907_ ),
    .A(\register_file_i/_2878_ ),
    .B(\register_file_i/_2902_ ));
 sg13g2_buf_16 fanout117 (.X(net117),
    .A(net121));
 sg13g2_mux2_1 \register_file_i/_6227_  (.A0(net755),
    .A1(\register_file_i/rf_reg_288_ ),
    .S(net843),
    .X(\register_file_i/_0212_ ));
 sg13g2_mux2_1 \register_file_i/_6228_  (.A0(net1002),
    .A1(\register_file_i/rf_reg_289_ ),
    .S(net843),
    .X(\register_file_i/_0213_ ));
 sg13g2_mux2_1 \register_file_i/_6229_  (.A0(net886),
    .A1(\register_file_i/rf_reg_290_ ),
    .S(net843),
    .X(\register_file_i/_0214_ ));
 sg13g2_mux2_1 \register_file_i/_6230_  (.A0(net1021),
    .A1(\register_file_i/rf_reg_291_ ),
    .S(net843),
    .X(\register_file_i/_0215_ ));
 sg13g2_mux2_1 \register_file_i/_6231_  (.A0(net1015),
    .A1(\register_file_i/rf_reg_292_ ),
    .S(net843),
    .X(\register_file_i/_0216_ ));
 sg13g2_mux2_1 \register_file_i/_6232_  (.A0(net995),
    .A1(\register_file_i/rf_reg_293_ ),
    .S(net842),
    .X(\register_file_i/_0217_ ));
 sg13g2_mux2_1 \register_file_i/_6233_  (.A0(net880),
    .A1(\register_file_i/rf_reg_294_ ),
    .S(net843),
    .X(\register_file_i/_0218_ ));
 sg13g2_mux2_1 \register_file_i/_6234_  (.A0(net991),
    .A1(\register_file_i/rf_reg_295_ ),
    .S(net843),
    .X(\register_file_i/_0219_ ));
 sg13g2_mux2_1 \register_file_i/_6235_  (.A0(net875),
    .A1(\register_file_i/rf_reg_296_ ),
    .S(net843),
    .X(\register_file_i/_0220_ ));
 sg13g2_mux2_1 \register_file_i/_6236_  (.A0(net804),
    .A1(\register_file_i/rf_reg_297_ ),
    .S(net842),
    .X(\register_file_i/_0221_ ));
 sg13g2_buf_1 fanout116 (.A(net120),
    .X(net116));
 sg13g2_mux2_1 \register_file_i/_6238_  (.A0(net795),
    .A1(\register_file_i/rf_reg_298_ ),
    .S(net842),
    .X(\register_file_i/_0222_ ));
 sg13g2_mux2_1 \register_file_i/_6239_  (.A0(net790),
    .A1(\register_file_i/rf_reg_299_ ),
    .S(net842),
    .X(\register_file_i/_0223_ ));
 sg13g2_mux2_1 \register_file_i/_6240_  (.A0(net799),
    .A1(\register_file_i/rf_reg_300_ ),
    .S(net842),
    .X(\register_file_i/_0224_ ));
 sg13g2_mux2_1 \register_file_i/_6241_  (.A0(net785),
    .A1(\register_file_i/rf_reg_301_ ),
    .S(net842),
    .X(\register_file_i/_0225_ ));
 sg13g2_mux2_1 \register_file_i/_6242_  (.A0(net747),
    .A1(\register_file_i/rf_reg_302_ ),
    .S(net845),
    .X(\register_file_i/_0226_ ));
 sg13g2_mux2_1 \register_file_i/_6243_  (.A0(net780),
    .A1(\register_file_i/rf_reg_303_ ),
    .S(net845),
    .X(\register_file_i/_0227_ ));
 sg13g2_mux2_1 \register_file_i/_6244_  (.A0(net708),
    .A1(\register_file_i/rf_reg_304_ ),
    .S(net846),
    .X(\register_file_i/_0228_ ));
 sg13g2_mux2_1 \register_file_i/_6245_  (.A0(net724),
    .A1(\register_file_i/rf_reg_305_ ),
    .S(net845),
    .X(\register_file_i/_0229_ ));
 sg13g2_mux2_1 \register_file_i/_6246_  (.A0(net703),
    .A1(\register_file_i/rf_reg_306_ ),
    .S(net845),
    .X(\register_file_i/_0230_ ));
 sg13g2_mux2_1 \register_file_i/_6247_  (.A0(net699),
    .A1(\register_file_i/rf_reg_307_ ),
    .S(net845),
    .X(\register_file_i/_0231_ ));
 sg13g2_buf_2 fanout115 (.A(net120),
    .X(net115));
 sg13g2_mux2_1 \register_file_i/_6249_  (.A0(net736),
    .A1(\register_file_i/rf_reg_308_ ),
    .S(net846),
    .X(\register_file_i/_0232_ ));
 sg13g2_mux2_1 \register_file_i/_6250_  (.A0(net670),
    .A1(\register_file_i/rf_reg_309_ ),
    .S(net846),
    .X(\register_file_i/_0233_ ));
 sg13g2_mux2_1 \register_file_i/_6251_  (.A0(net694),
    .A1(\register_file_i/rf_reg_310_ ),
    .S(net846),
    .X(\register_file_i/_0234_ ));
 sg13g2_mux2_1 \register_file_i/_6252_  (.A0(net689),
    .A1(\register_file_i/rf_reg_311_ ),
    .S(net846),
    .X(\register_file_i/_0235_ ));
 sg13g2_mux2_1 \register_file_i/_6253_  (.A0(net684),
    .A1(\register_file_i/rf_reg_312_ ),
    .S(net845),
    .X(\register_file_i/_0236_ ));
 sg13g2_mux2_1 \register_file_i/_6254_  (.A0(net599),
    .A1(\register_file_i/rf_reg_313_ ),
    .S(net844),
    .X(\register_file_i/_0237_ ));
 sg13g2_mux2_1 \register_file_i/_6255_  (.A0(net665),
    .A1(\register_file_i/rf_reg_314_ ),
    .S(net844),
    .X(\register_file_i/_0238_ ));
 sg13g2_mux2_1 \register_file_i/_6256_  (.A0(net581),
    .A1(\register_file_i/rf_reg_315_ ),
    .S(net842),
    .X(\register_file_i/_0239_ ));
 sg13g2_mux2_1 \register_file_i/_6257_  (.A0(net577),
    .A1(\register_file_i/rf_reg_316_ ),
    .S(net844),
    .X(\register_file_i/_0240_ ));
 sg13g2_mux2_1 \register_file_i/_6258_  (.A0(net567),
    .A1(\register_file_i/rf_reg_317_ ),
    .S(net842),
    .X(\register_file_i/_0241_ ));
 sg13g2_mux2_1 \register_file_i/_6259_  (.A0(net576),
    .A1(\register_file_i/rf_reg_318_ ),
    .S(net845),
    .X(\register_file_i/_0242_ ));
 sg13g2_mux2_1 \register_file_i/_6260_  (.A0(net562),
    .A1(\register_file_i/rf_reg_319_ ),
    .S(net845),
    .X(\register_file_i/_0243_ ));
 sg13g2_nand2_2 \register_file_i/_6261_  (.Y(\register_file_i/_2911_ ),
    .A(\register_file_i/_2884_ ),
    .B(\register_file_i/_2902_ ));
 sg13g2_buf_8 fanout114 (.A(net120),
    .X(net114));
 sg13g2_mux2_1 \register_file_i/_6263_  (.A0(net755),
    .A1(\register_file_i/rf_reg_320_ ),
    .S(net838),
    .X(\register_file_i/_0244_ ));
 sg13g2_mux2_1 \register_file_i/_6264_  (.A0(net1002),
    .A1(\register_file_i/rf_reg_321_ ),
    .S(net838),
    .X(\register_file_i/_0245_ ));
 sg13g2_mux2_1 \register_file_i/_6265_  (.A0(net886),
    .A1(\register_file_i/rf_reg_322_ ),
    .S(net838),
    .X(\register_file_i/_0246_ ));
 sg13g2_mux2_1 \register_file_i/_6266_  (.A0(net1020),
    .A1(\register_file_i/rf_reg_323_ ),
    .S(net838),
    .X(\register_file_i/_0247_ ));
 sg13g2_mux2_1 \register_file_i/_6267_  (.A0(net1015),
    .A1(\register_file_i/rf_reg_324_ ),
    .S(net838),
    .X(\register_file_i/_0248_ ));
 sg13g2_mux2_1 \register_file_i/_6268_  (.A0(net995),
    .A1(\register_file_i/rf_reg_325_ ),
    .S(net837),
    .X(\register_file_i/_0249_ ));
 sg13g2_mux2_1 \register_file_i/_6269_  (.A0(net880),
    .A1(\register_file_i/rf_reg_326_ ),
    .S(net838),
    .X(\register_file_i/_0250_ ));
 sg13g2_mux2_1 \register_file_i/_6270_  (.A0(net991),
    .A1(\register_file_i/rf_reg_327_ ),
    .S(net838),
    .X(\register_file_i/_0251_ ));
 sg13g2_mux2_1 \register_file_i/_6271_  (.A0(net875),
    .A1(\register_file_i/rf_reg_328_ ),
    .S(net838),
    .X(\register_file_i/_0252_ ));
 sg13g2_mux2_1 \register_file_i/_6272_  (.A0(net804),
    .A1(\register_file_i/rf_reg_329_ ),
    .S(net837),
    .X(\register_file_i/_0253_ ));
 sg13g2_nand2_2 \register_file_i/_6273_  (.Y(\register_file_i/_2913_ ),
    .A(\register_file_i/_2816_ ),
    .B(\register_file_i/_2878_ ));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(net120));
 sg13g2_mux2_1 \register_file_i/_6275_  (.A0(net755),
    .A1(\register_file_i/rf_reg_32_ ),
    .S(net834),
    .X(\register_file_i/_0254_ ));
 sg13g2_buf_16 fanout112 (.X(net112),
    .A(net120));
 sg13g2_mux2_1 \register_file_i/_6277_  (.A0(net795),
    .A1(\register_file_i/rf_reg_330_ ),
    .S(net837),
    .X(\register_file_i/_0255_ ));
 sg13g2_mux2_1 \register_file_i/_6278_  (.A0(net790),
    .A1(\register_file_i/rf_reg_331_ ),
    .S(net837),
    .X(\register_file_i/_0256_ ));
 sg13g2_mux2_1 \register_file_i/_6279_  (.A0(net800),
    .A1(\register_file_i/rf_reg_332_ ),
    .S(net837),
    .X(\register_file_i/_0257_ ));
 sg13g2_mux2_1 \register_file_i/_6280_  (.A0(net785),
    .A1(\register_file_i/rf_reg_333_ ),
    .S(net839),
    .X(\register_file_i/_0258_ ));
 sg13g2_mux2_1 \register_file_i/_6281_  (.A0(net747),
    .A1(\register_file_i/rf_reg_334_ ),
    .S(net837),
    .X(\register_file_i/_0259_ ));
 sg13g2_mux2_1 \register_file_i/_6282_  (.A0(net780),
    .A1(\register_file_i/rf_reg_335_ ),
    .S(net840),
    .X(\register_file_i/_0260_ ));
 sg13g2_mux2_1 \register_file_i/_6283_  (.A0(net708),
    .A1(\register_file_i/rf_reg_336_ ),
    .S(net840),
    .X(\register_file_i/_0261_ ));
 sg13g2_mux2_1 \register_file_i/_6284_  (.A0(net723),
    .A1(\register_file_i/rf_reg_337_ ),
    .S(net840),
    .X(\register_file_i/_0262_ ));
 sg13g2_mux2_1 \register_file_i/_6285_  (.A0(net703),
    .A1(\register_file_i/rf_reg_338_ ),
    .S(net840),
    .X(\register_file_i/_0263_ ));
 sg13g2_mux2_1 \register_file_i/_6286_  (.A0(net699),
    .A1(\register_file_i/rf_reg_339_ ),
    .S(net840),
    .X(\register_file_i/_0264_ ));
 sg13g2_mux2_1 \register_file_i/_6287_  (.A0(net1003),
    .A1(\register_file_i/rf_reg_33_ ),
    .S(net832),
    .X(\register_file_i/_0265_ ));
 sg13g2_buf_16 fanout111 (.X(net111),
    .A(net120));
 sg13g2_mux2_1 \register_file_i/_6289_  (.A0(net736),
    .A1(\register_file_i/rf_reg_340_ ),
    .S(net841),
    .X(\register_file_i/_0266_ ));
 sg13g2_mux2_1 \register_file_i/_6290_  (.A0(net670),
    .A1(\register_file_i/rf_reg_341_ ),
    .S(net841),
    .X(\register_file_i/_0267_ ));
 sg13g2_mux2_1 \register_file_i/_6291_  (.A0(net694),
    .A1(\register_file_i/rf_reg_342_ ),
    .S(net841),
    .X(\register_file_i/_0268_ ));
 sg13g2_mux2_1 \register_file_i/_6292_  (.A0(net689),
    .A1(\register_file_i/rf_reg_343_ ),
    .S(net841),
    .X(\register_file_i/_0269_ ));
 sg13g2_mux2_1 \register_file_i/_6293_  (.A0(net684),
    .A1(\register_file_i/rf_reg_344_ ),
    .S(net840),
    .X(\register_file_i/_0270_ ));
 sg13g2_mux2_1 \register_file_i/_6294_  (.A0(net599),
    .A1(\register_file_i/rf_reg_345_ ),
    .S(net839),
    .X(\register_file_i/_0271_ ));
 sg13g2_mux2_1 \register_file_i/_6295_  (.A0(net665),
    .A1(\register_file_i/rf_reg_346_ ),
    .S(net837),
    .X(\register_file_i/_0272_ ));
 sg13g2_mux2_1 \register_file_i/_6296_  (.A0(net581),
    .A1(\register_file_i/rf_reg_347_ ),
    .S(net839),
    .X(\register_file_i/_0273_ ));
 sg13g2_mux2_1 \register_file_i/_6297_  (.A0(net578),
    .A1(\register_file_i/rf_reg_348_ ),
    .S(net839),
    .X(\register_file_i/_0274_ ));
 sg13g2_mux2_1 \register_file_i/_6298_  (.A0(net567),
    .A1(\register_file_i/rf_reg_349_ ),
    .S(net837),
    .X(\register_file_i/_0275_ ));
 sg13g2_mux2_1 \register_file_i/_6299_  (.A0(net886),
    .A1(\register_file_i/rf_reg_34_ ),
    .S(net832),
    .X(\register_file_i/_0276_ ));
 sg13g2_mux2_1 \register_file_i/_6300_  (.A0(net575),
    .A1(\register_file_i/rf_reg_350_ ),
    .S(net840),
    .X(\register_file_i/_0277_ ));
 sg13g2_mux2_1 \register_file_i/_6301_  (.A0(net562),
    .A1(\register_file_i/rf_reg_351_ ),
    .S(net840),
    .X(\register_file_i/_0278_ ));
 sg13g2_nor3_2 \register_file_i/_6302_  (.A(\register_file_i/_2813_ ),
    .B(\register_file_i/_2867_ ),
    .C(\register_file_i/_2901_ ),
    .Y(\register_file_i/_2917_ ));
 sg13g2_buf_4 fanout110 (.X(net110),
    .A(_01868_));
 sg13g2_mux2_1 \register_file_i/_6304_  (.A0(\register_file_i/rf_reg_352_ ),
    .A1(net756),
    .S(net975),
    .X(\register_file_i/_0279_ ));
 sg13g2_mux2_1 \register_file_i/_6305_  (.A0(\register_file_i/rf_reg_353_ ),
    .A1(net1003),
    .S(net975),
    .X(\register_file_i/_0280_ ));
 sg13g2_mux2_1 \register_file_i/_6306_  (.A0(\register_file_i/rf_reg_354_ ),
    .A1(net886),
    .S(net975),
    .X(\register_file_i/_0281_ ));
 sg13g2_mux2_1 \register_file_i/_6307_  (.A0(\register_file_i/rf_reg_355_ ),
    .A1(net1021),
    .S(net975),
    .X(\register_file_i/_0282_ ));
 sg13g2_mux2_1 \register_file_i/_6308_  (.A0(\register_file_i/rf_reg_356_ ),
    .A1(net1015),
    .S(net975),
    .X(\register_file_i/_0283_ ));
 sg13g2_mux2_1 \register_file_i/_6309_  (.A0(\register_file_i/rf_reg_357_ ),
    .A1(net995),
    .S(net974),
    .X(\register_file_i/_0284_ ));
 sg13g2_mux2_1 \register_file_i/_6310_  (.A0(\register_file_i/rf_reg_358_ ),
    .A1(net880),
    .S(net975),
    .X(\register_file_i/_0285_ ));
 sg13g2_mux2_1 \register_file_i/_6311_  (.A0(\register_file_i/rf_reg_359_ ),
    .A1(net991),
    .S(net975),
    .X(\register_file_i/_0286_ ));
 sg13g2_mux2_1 \register_file_i/_6312_  (.A0(net1023),
    .A1(\register_file_i/rf_reg_35_ ),
    .S(net832),
    .X(\register_file_i/_0287_ ));
 sg13g2_mux2_1 \register_file_i/_6313_  (.A0(\register_file_i/rf_reg_360_ ),
    .A1(net875),
    .S(net975),
    .X(\register_file_i/_0288_ ));
 sg13g2_mux2_1 \register_file_i/_6314_  (.A0(\register_file_i/rf_reg_361_ ),
    .A1(net804),
    .S(net974),
    .X(\register_file_i/_0289_ ));
 sg13g2_buf_2 fanout109 (.A(_03283_),
    .X(net109));
 sg13g2_mux2_1 \register_file_i/_6316_  (.A0(\register_file_i/rf_reg_362_ ),
    .A1(net795),
    .S(net974),
    .X(\register_file_i/_0290_ ));
 sg13g2_mux2_1 \register_file_i/_6317_  (.A0(\register_file_i/rf_reg_363_ ),
    .A1(net790),
    .S(net974),
    .X(\register_file_i/_0291_ ));
 sg13g2_mux2_1 \register_file_i/_6318_  (.A0(\register_file_i/rf_reg_364_ ),
    .A1(net800),
    .S(net974),
    .X(\register_file_i/_0292_ ));
 sg13g2_mux2_1 \register_file_i/_6319_  (.A0(\register_file_i/rf_reg_365_ ),
    .A1(net785),
    .S(net976),
    .X(\register_file_i/_0293_ ));
 sg13g2_mux2_1 \register_file_i/_6320_  (.A0(\register_file_i/rf_reg_366_ ),
    .A1(net747),
    .S(net974),
    .X(\register_file_i/_0294_ ));
 sg13g2_mux2_1 \register_file_i/_6321_  (.A0(\register_file_i/rf_reg_367_ ),
    .A1(net780),
    .S(net977),
    .X(\register_file_i/_0295_ ));
 sg13g2_mux2_1 \register_file_i/_6322_  (.A0(\register_file_i/rf_reg_368_ ),
    .A1(net708),
    .S(net977),
    .X(\register_file_i/_0296_ ));
 sg13g2_mux2_1 \register_file_i/_6323_  (.A0(\register_file_i/rf_reg_369_ ),
    .A1(net723),
    .S(net977),
    .X(\register_file_i/_0297_ ));
 sg13g2_mux2_1 \register_file_i/_6324_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_36_ ),
    .S(net833),
    .X(\register_file_i/_0298_ ));
 sg13g2_mux2_1 \register_file_i/_6325_  (.A0(\register_file_i/rf_reg_370_ ),
    .A1(net703),
    .S(net977),
    .X(\register_file_i/_0299_ ));
 sg13g2_mux2_1 \register_file_i/_6326_  (.A0(\register_file_i/rf_reg_371_ ),
    .A1(net698),
    .S(net977),
    .X(\register_file_i/_0300_ ));
 sg13g2_buf_4 fanout108 (.X(net108),
    .A(net109));
 sg13g2_mux2_1 \register_file_i/_6328_  (.A0(\register_file_i/rf_reg_372_ ),
    .A1(net736),
    .S(net978),
    .X(\register_file_i/_0301_ ));
 sg13g2_mux2_1 \register_file_i/_6329_  (.A0(\register_file_i/rf_reg_373_ ),
    .A1(net670),
    .S(net978),
    .X(\register_file_i/_0302_ ));
 sg13g2_mux2_1 \register_file_i/_6330_  (.A0(\register_file_i/rf_reg_374_ ),
    .A1(net694),
    .S(net978),
    .X(\register_file_i/_0303_ ));
 sg13g2_mux2_1 \register_file_i/_6331_  (.A0(\register_file_i/rf_reg_375_ ),
    .A1(net689),
    .S(net978),
    .X(\register_file_i/_0304_ ));
 sg13g2_mux2_1 \register_file_i/_6332_  (.A0(\register_file_i/rf_reg_376_ ),
    .A1(net684),
    .S(net977),
    .X(\register_file_i/_0305_ ));
 sg13g2_mux2_1 \register_file_i/_6333_  (.A0(\register_file_i/rf_reg_377_ ),
    .A1(net599),
    .S(net976),
    .X(\register_file_i/_0306_ ));
 sg13g2_mux2_1 \register_file_i/_6334_  (.A0(\register_file_i/rf_reg_378_ ),
    .A1(net665),
    .S(net974),
    .X(\register_file_i/_0307_ ));
 sg13g2_mux2_1 \register_file_i/_6335_  (.A0(\register_file_i/rf_reg_379_ ),
    .A1(net581),
    .S(net976),
    .X(\register_file_i/_0308_ ));
 sg13g2_mux2_1 \register_file_i/_6336_  (.A0(net998),
    .A1(\register_file_i/rf_reg_37_ ),
    .S(net833),
    .X(\register_file_i/_0309_ ));
 sg13g2_mux2_1 \register_file_i/_6337_  (.A0(\register_file_i/rf_reg_380_ ),
    .A1(net577),
    .S(net976),
    .X(\register_file_i/_0310_ ));
 sg13g2_mux2_1 \register_file_i/_6338_  (.A0(\register_file_i/rf_reg_381_ ),
    .A1(net567),
    .S(net974),
    .X(\register_file_i/_0311_ ));
 sg13g2_mux2_1 \register_file_i/_6339_  (.A0(\register_file_i/rf_reg_382_ ),
    .A1(net575),
    .S(net977),
    .X(\register_file_i/_0312_ ));
 sg13g2_mux2_1 \register_file_i/_6340_  (.A0(\register_file_i/rf_reg_383_ ),
    .A1(net562),
    .S(net977),
    .X(\register_file_i/_0313_ ));
 sg13g2_nand4_1 \register_file_i/_6341_  (.B(net2099),
    .C(\register_file_i/_2814_ ),
    .A(net1991),
    .Y(\register_file_i/_2921_ ),
    .D(\register_file_i/_2866_ ));
 sg13g2_buf_4 fanout107 (.X(net107),
    .A(net109));
 sg13g2_buf_4 fanout106 (.X(net106),
    .A(net109));
 sg13g2_mux2_1 \register_file_i/_6344_  (.A0(net755),
    .A1(\register_file_i/rf_reg_384_ ),
    .S(net969),
    .X(\register_file_i/_0314_ ));
 sg13g2_mux2_1 \register_file_i/_6345_  (.A0(net1002),
    .A1(\register_file_i/rf_reg_385_ ),
    .S(net969),
    .X(\register_file_i/_0315_ ));
 sg13g2_mux2_1 \register_file_i/_6346_  (.A0(net885),
    .A1(\register_file_i/rf_reg_386_ ),
    .S(net969),
    .X(\register_file_i/_0316_ ));
 sg13g2_mux2_1 \register_file_i/_6347_  (.A0(net1020),
    .A1(\register_file_i/rf_reg_387_ ),
    .S(net969),
    .X(\register_file_i/_0317_ ));
 sg13g2_mux2_1 \register_file_i/_6348_  (.A0(net1015),
    .A1(\register_file_i/rf_reg_388_ ),
    .S(net969),
    .X(\register_file_i/_0318_ ));
 sg13g2_mux2_1 \register_file_i/_6349_  (.A0(net995),
    .A1(\register_file_i/rf_reg_389_ ),
    .S(net968),
    .X(\register_file_i/_0319_ ));
 sg13g2_mux2_1 \register_file_i/_6350_  (.A0(net883),
    .A1(\register_file_i/rf_reg_38_ ),
    .S(net833),
    .X(\register_file_i/_0320_ ));
 sg13g2_mux2_1 \register_file_i/_6351_  (.A0(net880),
    .A1(\register_file_i/rf_reg_390_ ),
    .S(net969),
    .X(\register_file_i/_0321_ ));
 sg13g2_mux2_1 \register_file_i/_6352_  (.A0(net991),
    .A1(\register_file_i/rf_reg_391_ ),
    .S(net969),
    .X(\register_file_i/_0322_ ));
 sg13g2_mux2_1 \register_file_i/_6353_  (.A0(net875),
    .A1(\register_file_i/rf_reg_392_ ),
    .S(net969),
    .X(\register_file_i/_0323_ ));
 sg13g2_mux2_1 \register_file_i/_6354_  (.A0(net804),
    .A1(\register_file_i/rf_reg_393_ ),
    .S(net968),
    .X(\register_file_i/_0324_ ));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(net109));
 sg13g2_mux2_1 \register_file_i/_6356_  (.A0(net795),
    .A1(\register_file_i/rf_reg_394_ ),
    .S(net968),
    .X(\register_file_i/_0325_ ));
 sg13g2_mux2_1 \register_file_i/_6357_  (.A0(net790),
    .A1(\register_file_i/rf_reg_395_ ),
    .S(net968),
    .X(\register_file_i/_0326_ ));
 sg13g2_mux2_1 \register_file_i/_6358_  (.A0(net800),
    .A1(\register_file_i/rf_reg_396_ ),
    .S(net968),
    .X(\register_file_i/_0327_ ));
 sg13g2_mux2_1 \register_file_i/_6359_  (.A0(net786),
    .A1(\register_file_i/rf_reg_397_ ),
    .S(net971),
    .X(\register_file_i/_0328_ ));
 sg13g2_mux2_1 \register_file_i/_6360_  (.A0(net747),
    .A1(\register_file_i/rf_reg_398_ ),
    .S(net971),
    .X(\register_file_i/_0329_ ));
 sg13g2_mux2_1 \register_file_i/_6361_  (.A0(net780),
    .A1(\register_file_i/rf_reg_399_ ),
    .S(net971),
    .X(\register_file_i/_0330_ ));
 sg13g2_mux2_1 \register_file_i/_6362_  (.A0(net994),
    .A1(\register_file_i/rf_reg_39_ ),
    .S(net833),
    .X(\register_file_i/_0331_ ));
 sg13g2_mux2_1 \register_file_i/_6363_  (.A0(net708),
    .A1(\register_file_i/rf_reg_400_ ),
    .S(net971),
    .X(\register_file_i/_0332_ ));
 sg13g2_mux2_1 \register_file_i/_6364_  (.A0(net724),
    .A1(\register_file_i/rf_reg_401_ ),
    .S(net972),
    .X(\register_file_i/_0333_ ));
 sg13g2_mux2_1 \register_file_i/_6365_  (.A0(net703),
    .A1(\register_file_i/rf_reg_402_ ),
    .S(net971),
    .X(\register_file_i/_0334_ ));
 sg13g2_mux2_1 \register_file_i/_6366_  (.A0(net698),
    .A1(\register_file_i/rf_reg_403_ ),
    .S(net972),
    .X(\register_file_i/_0335_ ));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(net109));
 sg13g2_mux2_1 \register_file_i/_6368_  (.A0(net736),
    .A1(\register_file_i/rf_reg_404_ ),
    .S(net972),
    .X(\register_file_i/_0336_ ));
 sg13g2_mux2_1 \register_file_i/_6369_  (.A0(net670),
    .A1(\register_file_i/rf_reg_405_ ),
    .S(net972),
    .X(\register_file_i/_0337_ ));
 sg13g2_mux2_1 \register_file_i/_6370_  (.A0(net694),
    .A1(\register_file_i/rf_reg_406_ ),
    .S(net973),
    .X(\register_file_i/_0338_ ));
 sg13g2_mux2_1 \register_file_i/_6371_  (.A0(net689),
    .A1(\register_file_i/rf_reg_407_ ),
    .S(net971),
    .X(\register_file_i/_0339_ ));
 sg13g2_mux2_1 \register_file_i/_6372_  (.A0(net684),
    .A1(\register_file_i/rf_reg_408_ ),
    .S(net971),
    .X(\register_file_i/_0340_ ));
 sg13g2_mux2_1 \register_file_i/_6373_  (.A0(net599),
    .A1(\register_file_i/rf_reg_409_ ),
    .S(net970),
    .X(\register_file_i/_0341_ ));
 sg13g2_mux2_1 \register_file_i/_6374_  (.A0(net878),
    .A1(\register_file_i/rf_reg_40_ ),
    .S(net833),
    .X(\register_file_i/_0342_ ));
 sg13g2_mux2_1 \register_file_i/_6375_  (.A0(net665),
    .A1(\register_file_i/rf_reg_410_ ),
    .S(net968),
    .X(\register_file_i/_0343_ ));
 sg13g2_mux2_1 \register_file_i/_6376_  (.A0(net581),
    .A1(\register_file_i/rf_reg_411_ ),
    .S(net968),
    .X(\register_file_i/_0344_ ));
 sg13g2_mux2_1 \register_file_i/_6377_  (.A0(net577),
    .A1(\register_file_i/rf_reg_412_ ),
    .S(net970),
    .X(\register_file_i/_0345_ ));
 sg13g2_mux2_1 \register_file_i/_6378_  (.A0(net567),
    .A1(\register_file_i/rf_reg_413_ ),
    .S(net968),
    .X(\register_file_i/_0346_ ));
 sg13g2_mux2_1 \register_file_i/_6379_  (.A0(net575),
    .A1(\register_file_i/rf_reg_414_ ),
    .S(net972),
    .X(\register_file_i/_0347_ ));
 sg13g2_mux2_1 \register_file_i/_6380_  (.A0(net562),
    .A1(\register_file_i/rf_reg_415_ ),
    .S(net971),
    .X(\register_file_i/_0348_ ));
 sg13g2_nand2b_2 \register_file_i/_6381_  (.Y(\register_file_i/_2926_ ),
    .B(\register_file_i/_2814_ ),
    .A_N(\register_file_i/_2799_ ));
 sg13g2_nor3_2 \register_file_i/_6382_  (.A(\id_stage_i.controller_i.instr_i_8_ ),
    .B(\register_file_i/_2877_ ),
    .C(\register_file_i/_2926_ ),
    .Y(\register_file_i/_2927_ ));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net109));
 sg13g2_mux2_1 \register_file_i/_6384_  (.A0(\register_file_i/rf_reg_416_ ),
    .A1(net755),
    .S(net827),
    .X(\register_file_i/_0349_ ));
 sg13g2_mux2_1 \register_file_i/_6385_  (.A0(\register_file_i/rf_reg_417_ ),
    .A1(net1002),
    .S(net827),
    .X(\register_file_i/_0350_ ));
 sg13g2_mux2_1 \register_file_i/_6386_  (.A0(\register_file_i/rf_reg_418_ ),
    .A1(net884),
    .S(net827),
    .X(\register_file_i/_0351_ ));
 sg13g2_mux2_1 \register_file_i/_6387_  (.A0(\register_file_i/rf_reg_419_ ),
    .A1(net1021),
    .S(net827),
    .X(\register_file_i/_0352_ ));
 sg13g2_mux2_1 \register_file_i/_6388_  (.A0(net807),
    .A1(\register_file_i/rf_reg_41_ ),
    .S(net832),
    .X(\register_file_i/_0353_ ));
 sg13g2_mux2_1 \register_file_i/_6389_  (.A0(\register_file_i/rf_reg_420_ ),
    .A1(net1015),
    .S(net827),
    .X(\register_file_i/_0354_ ));
 sg13g2_mux2_1 \register_file_i/_6390_  (.A0(\register_file_i/rf_reg_421_ ),
    .A1(net995),
    .S(net826),
    .X(\register_file_i/_0355_ ));
 sg13g2_mux2_1 \register_file_i/_6391_  (.A0(\register_file_i/rf_reg_422_ ),
    .A1(net880),
    .S(net827),
    .X(\register_file_i/_0356_ ));
 sg13g2_mux2_1 \register_file_i/_6392_  (.A0(\register_file_i/rf_reg_423_ ),
    .A1(net991),
    .S(net827),
    .X(\register_file_i/_0357_ ));
 sg13g2_mux2_1 \register_file_i/_6393_  (.A0(\register_file_i/rf_reg_424_ ),
    .A1(net875),
    .S(net827),
    .X(\register_file_i/_0358_ ));
 sg13g2_mux2_1 \register_file_i/_6394_  (.A0(\register_file_i/rf_reg_425_ ),
    .A1(net804),
    .S(net826),
    .X(\register_file_i/_0359_ ));
 sg13g2_buf_2 fanout102 (.A(csr_addr_2_),
    .X(net102));
 sg13g2_mux2_1 \register_file_i/_6396_  (.A0(\register_file_i/rf_reg_426_ ),
    .A1(net795),
    .S(net826),
    .X(\register_file_i/_0360_ ));
 sg13g2_mux2_1 \register_file_i/_6397_  (.A0(\register_file_i/rf_reg_427_ ),
    .A1(net790),
    .S(net826),
    .X(\register_file_i/_0361_ ));
 sg13g2_mux2_1 \register_file_i/_6398_  (.A0(\register_file_i/rf_reg_428_ ),
    .A1(net800),
    .S(net826),
    .X(\register_file_i/_0362_ ));
 sg13g2_mux2_1 \register_file_i/_6399_  (.A0(\register_file_i/rf_reg_429_ ),
    .A1(net786),
    .S(net829),
    .X(\register_file_i/_0363_ ));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(csr_addr_2_));
 sg13g2_mux2_1 \register_file_i/_6401_  (.A0(net798),
    .A1(\register_file_i/rf_reg_42_ ),
    .S(net832),
    .X(\register_file_i/_0364_ ));
 sg13g2_mux2_1 \register_file_i/_6402_  (.A0(\register_file_i/rf_reg_430_ ),
    .A1(net747),
    .S(net829),
    .X(\register_file_i/_0365_ ));
 sg13g2_mux2_1 \register_file_i/_6403_  (.A0(\register_file_i/rf_reg_431_ ),
    .A1(net780),
    .S(net829),
    .X(\register_file_i/_0366_ ));
 sg13g2_mux2_1 \register_file_i/_6404_  (.A0(\register_file_i/rf_reg_432_ ),
    .A1(net709),
    .S(net829),
    .X(\register_file_i/_0367_ ));
 sg13g2_mux2_1 \register_file_i/_6405_  (.A0(\register_file_i/rf_reg_433_ ),
    .A1(net724),
    .S(net830),
    .X(\register_file_i/_0368_ ));
 sg13g2_mux2_1 \register_file_i/_6406_  (.A0(\register_file_i/rf_reg_434_ ),
    .A1(net703),
    .S(net829),
    .X(\register_file_i/_0369_ ));
 sg13g2_mux2_1 \register_file_i/_6407_  (.A0(\register_file_i/rf_reg_435_ ),
    .A1(net698),
    .S(net830),
    .X(\register_file_i/_0370_ ));
 sg13g2_buf_2 fanout100 (.A(csr_addr_2_),
    .X(net100));
 sg13g2_mux2_1 \register_file_i/_6409_  (.A0(\register_file_i/rf_reg_436_ ),
    .A1(net736),
    .S(net830),
    .X(\register_file_i/_0371_ ));
 sg13g2_mux2_1 \register_file_i/_6410_  (.A0(\register_file_i/rf_reg_437_ ),
    .A1(net670),
    .S(net830),
    .X(\register_file_i/_0372_ ));
 sg13g2_mux2_1 \register_file_i/_6411_  (.A0(\register_file_i/rf_reg_438_ ),
    .A1(net694),
    .S(net831),
    .X(\register_file_i/_0373_ ));
 sg13g2_mux2_1 \register_file_i/_6412_  (.A0(\register_file_i/rf_reg_439_ ),
    .A1(net689),
    .S(net829),
    .X(\register_file_i/_0374_ ));
 sg13g2_mux2_1 \register_file_i/_6413_  (.A0(net793),
    .A1(\register_file_i/rf_reg_43_ ),
    .S(net832),
    .X(\register_file_i/_0375_ ));
 sg13g2_mux2_1 \register_file_i/_6414_  (.A0(\register_file_i/rf_reg_440_ ),
    .A1(net684),
    .S(net829),
    .X(\register_file_i/_0376_ ));
 sg13g2_mux2_1 \register_file_i/_6415_  (.A0(\register_file_i/rf_reg_441_ ),
    .A1(net599),
    .S(net828),
    .X(\register_file_i/_0377_ ));
 sg13g2_mux2_1 \register_file_i/_6416_  (.A0(\register_file_i/rf_reg_442_ ),
    .A1(net665),
    .S(net826),
    .X(\register_file_i/_0378_ ));
 sg13g2_mux2_1 \register_file_i/_6417_  (.A0(\register_file_i/rf_reg_443_ ),
    .A1(net581),
    .S(net826),
    .X(\register_file_i/_0379_ ));
 sg13g2_mux2_1 \register_file_i/_6418_  (.A0(\register_file_i/rf_reg_444_ ),
    .A1(net577),
    .S(net828),
    .X(\register_file_i/_0380_ ));
 sg13g2_mux2_1 \register_file_i/_6419_  (.A0(\register_file_i/rf_reg_445_ ),
    .A1(net567),
    .S(net826),
    .X(\register_file_i/_0381_ ));
 sg13g2_mux2_1 \register_file_i/_6420_  (.A0(\register_file_i/rf_reg_446_ ),
    .A1(net575),
    .S(net829),
    .X(\register_file_i/_0382_ ));
 sg13g2_mux2_1 \register_file_i/_6421_  (.A0(\register_file_i/rf_reg_447_ ),
    .A1(net562),
    .S(net830),
    .X(\register_file_i/_0383_ ));
 sg13g2_nor3_2 \register_file_i/_6422_  (.A(\register_file_i/_2883_ ),
    .B(net1993),
    .C(\register_file_i/_2926_ ),
    .Y(\register_file_i/_2932_ ));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(csr_addr_2_));
 sg13g2_mux2_1 \register_file_i/_6424_  (.A0(\register_file_i/rf_reg_448_ ),
    .A1(net755),
    .S(net821),
    .X(\register_file_i/_0384_ ));
 sg13g2_mux2_1 \register_file_i/_6425_  (.A0(\register_file_i/rf_reg_449_ ),
    .A1(net1002),
    .S(net821),
    .X(\register_file_i/_0385_ ));
 sg13g2_mux2_1 \register_file_i/_6426_  (.A0(net802),
    .A1(\register_file_i/rf_reg_44_ ),
    .S(net832),
    .X(\register_file_i/_0386_ ));
 sg13g2_mux2_1 \register_file_i/_6427_  (.A0(\register_file_i/rf_reg_450_ ),
    .A1(net885),
    .S(net821),
    .X(\register_file_i/_0387_ ));
 sg13g2_mux2_1 \register_file_i/_6428_  (.A0(\register_file_i/rf_reg_451_ ),
    .A1(net1021),
    .S(net821),
    .X(\register_file_i/_0388_ ));
 sg13g2_mux2_1 \register_file_i/_6429_  (.A0(\register_file_i/rf_reg_452_ ),
    .A1(net1015),
    .S(net821),
    .X(\register_file_i/_0389_ ));
 sg13g2_mux2_1 \register_file_i/_6430_  (.A0(\register_file_i/rf_reg_453_ ),
    .A1(net995),
    .S(net820),
    .X(\register_file_i/_0390_ ));
 sg13g2_mux2_1 \register_file_i/_6431_  (.A0(\register_file_i/rf_reg_454_ ),
    .A1(net880),
    .S(net821),
    .X(\register_file_i/_0391_ ));
 sg13g2_mux2_1 \register_file_i/_6432_  (.A0(\register_file_i/rf_reg_455_ ),
    .A1(net991),
    .S(net821),
    .X(\register_file_i/_0392_ ));
 sg13g2_mux2_1 \register_file_i/_6433_  (.A0(\register_file_i/rf_reg_456_ ),
    .A1(net875),
    .S(net821),
    .X(\register_file_i/_0393_ ));
 sg13g2_mux2_1 \register_file_i/_6434_  (.A0(\register_file_i/rf_reg_457_ ),
    .A1(net804),
    .S(net820),
    .X(\register_file_i/_0394_ ));
 sg13g2_buf_1 fanout98 (.A(_04166_),
    .X(net98));
 sg13g2_mux2_1 \register_file_i/_6436_  (.A0(\register_file_i/rf_reg_458_ ),
    .A1(net795),
    .S(net820),
    .X(\register_file_i/_0395_ ));
 sg13g2_mux2_1 \register_file_i/_6437_  (.A0(\register_file_i/rf_reg_459_ ),
    .A1(net790),
    .S(net820),
    .X(\register_file_i/_0396_ ));
 sg13g2_mux2_1 \register_file_i/_6438_  (.A0(net789),
    .A1(\register_file_i/rf_reg_45_ ),
    .S(net835),
    .X(\register_file_i/_0397_ ));
 sg13g2_mux2_1 \register_file_i/_6439_  (.A0(\register_file_i/rf_reg_460_ ),
    .A1(net800),
    .S(net820),
    .X(\register_file_i/_0398_ ));
 sg13g2_mux2_1 \register_file_i/_6440_  (.A0(\register_file_i/rf_reg_461_ ),
    .A1(net786),
    .S(net823),
    .X(\register_file_i/_0399_ ));
 sg13g2_mux2_1 \register_file_i/_6441_  (.A0(\register_file_i/rf_reg_462_ ),
    .A1(net747),
    .S(net823),
    .X(\register_file_i/_0400_ ));
 sg13g2_mux2_1 \register_file_i/_6442_  (.A0(\register_file_i/rf_reg_463_ ),
    .A1(net780),
    .S(net823),
    .X(\register_file_i/_0401_ ));
 sg13g2_mux2_1 \register_file_i/_6443_  (.A0(\register_file_i/rf_reg_464_ ),
    .A1(net708),
    .S(net824),
    .X(\register_file_i/_0402_ ));
 sg13g2_mux2_1 \register_file_i/_6444_  (.A0(\register_file_i/rf_reg_465_ ),
    .A1(net723),
    .S(net824),
    .X(\register_file_i/_0403_ ));
 sg13g2_mux2_1 \register_file_i/_6445_  (.A0(\register_file_i/rf_reg_466_ ),
    .A1(net703),
    .S(net823),
    .X(\register_file_i/_0404_ ));
 sg13g2_mux2_1 \register_file_i/_6446_  (.A0(\register_file_i/rf_reg_467_ ),
    .A1(net698),
    .S(net823),
    .X(\register_file_i/_0405_ ));
 sg13g2_buf_2 fanout97 (.A(net98),
    .X(net97));
 sg13g2_mux2_1 \register_file_i/_6448_  (.A0(\register_file_i/rf_reg_468_ ),
    .A1(net736),
    .S(net824),
    .X(\register_file_i/_0406_ ));
 sg13g2_mux2_1 \register_file_i/_6449_  (.A0(\register_file_i/rf_reg_469_ ),
    .A1(net670),
    .S(net824),
    .X(\register_file_i/_0407_ ));
 sg13g2_mux2_1 \register_file_i/_6450_  (.A0(net751),
    .A1(\register_file_i/rf_reg_46_ ),
    .S(net835),
    .X(\register_file_i/_0408_ ));
 sg13g2_mux2_1 \register_file_i/_6451_  (.A0(\register_file_i/rf_reg_470_ ),
    .A1(net694),
    .S(net825),
    .X(\register_file_i/_0409_ ));
 sg13g2_mux2_1 \register_file_i/_6452_  (.A0(\register_file_i/rf_reg_471_ ),
    .A1(net689),
    .S(net825),
    .X(\register_file_i/_0410_ ));
 sg13g2_mux2_1 \register_file_i/_6453_  (.A0(\register_file_i/rf_reg_472_ ),
    .A1(net684),
    .S(net823),
    .X(\register_file_i/_0411_ ));
 sg13g2_mux2_1 \register_file_i/_6454_  (.A0(\register_file_i/rf_reg_473_ ),
    .A1(net600),
    .S(net822),
    .X(\register_file_i/_0412_ ));
 sg13g2_mux2_1 \register_file_i/_6455_  (.A0(\register_file_i/rf_reg_474_ ),
    .A1(net665),
    .S(net820),
    .X(\register_file_i/_0413_ ));
 sg13g2_mux2_1 \register_file_i/_6456_  (.A0(\register_file_i/rf_reg_475_ ),
    .A1(net581),
    .S(net820),
    .X(\register_file_i/_0414_ ));
 sg13g2_mux2_1 \register_file_i/_6457_  (.A0(\register_file_i/rf_reg_476_ ),
    .A1(net577),
    .S(net822),
    .X(\register_file_i/_0415_ ));
 sg13g2_mux2_1 \register_file_i/_6458_  (.A0(\register_file_i/rf_reg_477_ ),
    .A1(net567),
    .S(net820),
    .X(\register_file_i/_0416_ ));
 sg13g2_mux2_1 \register_file_i/_6459_  (.A0(\register_file_i/rf_reg_478_ ),
    .A1(net575),
    .S(net823),
    .X(\register_file_i/_0417_ ));
 sg13g2_mux2_1 \register_file_i/_6460_  (.A0(\register_file_i/rf_reg_479_ ),
    .A1(net562),
    .S(net823),
    .X(\register_file_i/_0418_ ));
 sg13g2_mux2_1 \register_file_i/_6461_  (.A0(net783),
    .A1(\register_file_i/rf_reg_47_ ),
    .S(net835),
    .X(\register_file_i/_0419_ ));
 sg13g2_nor2_2 \register_file_i/_6462_  (.A(\register_file_i/_2813_ ),
    .B(\register_file_i/_2926_ ),
    .Y(\register_file_i/_2936_ ));
 sg13g2_buf_2 fanout96 (.A(net98),
    .X(net96));
 sg13g2_mux2_1 \register_file_i/_6464_  (.A0(\register_file_i/rf_reg_480_ ),
    .A1(net755),
    .S(net815),
    .X(\register_file_i/_0420_ ));
 sg13g2_mux2_1 \register_file_i/_6465_  (.A0(\register_file_i/rf_reg_481_ ),
    .A1(net1002),
    .S(net815),
    .X(\register_file_i/_0421_ ));
 sg13g2_mux2_1 \register_file_i/_6466_  (.A0(\register_file_i/rf_reg_482_ ),
    .A1(net885),
    .S(net815),
    .X(\register_file_i/_0422_ ));
 sg13g2_mux2_1 \register_file_i/_6467_  (.A0(\register_file_i/rf_reg_483_ ),
    .A1(net1020),
    .S(net815),
    .X(\register_file_i/_0423_ ));
 sg13g2_mux2_1 \register_file_i/_6468_  (.A0(\register_file_i/rf_reg_484_ ),
    .A1(net1015),
    .S(net815),
    .X(\register_file_i/_0424_ ));
 sg13g2_mux2_1 \register_file_i/_6469_  (.A0(\register_file_i/rf_reg_485_ ),
    .A1(net995),
    .S(net814),
    .X(\register_file_i/_0425_ ));
 sg13g2_mux2_1 \register_file_i/_6470_  (.A0(\register_file_i/rf_reg_486_ ),
    .A1(net880),
    .S(net815),
    .X(\register_file_i/_0426_ ));
 sg13g2_mux2_1 \register_file_i/_6471_  (.A0(\register_file_i/rf_reg_487_ ),
    .A1(net991),
    .S(net815),
    .X(\register_file_i/_0427_ ));
 sg13g2_mux2_1 \register_file_i/_6472_  (.A0(\register_file_i/rf_reg_488_ ),
    .A1(net875),
    .S(net815),
    .X(\register_file_i/_0428_ ));
 sg13g2_mux2_1 \register_file_i/_6473_  (.A0(\register_file_i/rf_reg_489_ ),
    .A1(net804),
    .S(net814),
    .X(\register_file_i/_0429_ ));
 sg13g2_mux2_1 \register_file_i/_6474_  (.A0(net710),
    .A1(\register_file_i/rf_reg_48_ ),
    .S(net835),
    .X(\register_file_i/_0430_ ));
 sg13g2_buf_2 fanout95 (.A(net98),
    .X(net95));
 sg13g2_mux2_1 \register_file_i/_6476_  (.A0(\register_file_i/rf_reg_490_ ),
    .A1(net795),
    .S(net814),
    .X(\register_file_i/_0431_ ));
 sg13g2_mux2_1 \register_file_i/_6477_  (.A0(\register_file_i/rf_reg_491_ ),
    .A1(net790),
    .S(net814),
    .X(\register_file_i/_0432_ ));
 sg13g2_mux2_1 \register_file_i/_6478_  (.A0(\register_file_i/rf_reg_492_ ),
    .A1(net800),
    .S(net814),
    .X(\register_file_i/_0433_ ));
 sg13g2_mux2_1 \register_file_i/_6479_  (.A0(\register_file_i/rf_reg_493_ ),
    .A1(net786),
    .S(net817),
    .X(\register_file_i/_0434_ ));
 sg13g2_mux2_1 \register_file_i/_6480_  (.A0(\register_file_i/rf_reg_494_ ),
    .A1(net747),
    .S(net817),
    .X(\register_file_i/_0435_ ));
 sg13g2_mux2_1 \register_file_i/_6481_  (.A0(\register_file_i/rf_reg_495_ ),
    .A1(net780),
    .S(net817),
    .X(\register_file_i/_0436_ ));
 sg13g2_mux2_1 \register_file_i/_6482_  (.A0(\register_file_i/rf_reg_496_ ),
    .A1(net708),
    .S(net818),
    .X(\register_file_i/_0437_ ));
 sg13g2_mux2_1 \register_file_i/_6483_  (.A0(\register_file_i/rf_reg_497_ ),
    .A1(net723),
    .S(net818),
    .X(\register_file_i/_0438_ ));
 sg13g2_mux2_1 \register_file_i/_6484_  (.A0(\register_file_i/rf_reg_498_ ),
    .A1(net703),
    .S(net817),
    .X(\register_file_i/_0439_ ));
 sg13g2_mux2_1 \register_file_i/_6485_  (.A0(\register_file_i/rf_reg_499_ ),
    .A1(net698),
    .S(net817),
    .X(\register_file_i/_0440_ ));
 sg13g2_mux2_1 \register_file_i/_6486_  (.A0(net726),
    .A1(\register_file_i/rf_reg_49_ ),
    .S(net836),
    .X(\register_file_i/_0441_ ));
 sg13g2_buf_2 fanout94 (.A(net98),
    .X(net94));
 sg13g2_mux2_1 \register_file_i/_6488_  (.A0(\register_file_i/rf_reg_500_ ),
    .A1(net736),
    .S(net818),
    .X(\register_file_i/_0442_ ));
 sg13g2_mux2_1 \register_file_i/_6489_  (.A0(\register_file_i/rf_reg_501_ ),
    .A1(net670),
    .S(net818),
    .X(\register_file_i/_0443_ ));
 sg13g2_mux2_1 \register_file_i/_6490_  (.A0(\register_file_i/rf_reg_502_ ),
    .A1(net693),
    .S(net819),
    .X(\register_file_i/_0444_ ));
 sg13g2_mux2_1 \register_file_i/_6491_  (.A0(\register_file_i/rf_reg_503_ ),
    .A1(net689),
    .S(net819),
    .X(\register_file_i/_0445_ ));
 sg13g2_mux2_1 \register_file_i/_6492_  (.A0(\register_file_i/rf_reg_504_ ),
    .A1(net684),
    .S(net817),
    .X(\register_file_i/_0446_ ));
 sg13g2_mux2_1 \register_file_i/_6493_  (.A0(\register_file_i/rf_reg_505_ ),
    .A1(net599),
    .S(net816),
    .X(\register_file_i/_0447_ ));
 sg13g2_mux2_1 \register_file_i/_6494_  (.A0(\register_file_i/rf_reg_506_ ),
    .A1(net665),
    .S(net814),
    .X(\register_file_i/_0448_ ));
 sg13g2_mux2_1 \register_file_i/_6495_  (.A0(\register_file_i/rf_reg_507_ ),
    .A1(net581),
    .S(net814),
    .X(\register_file_i/_0449_ ));
 sg13g2_mux2_1 \register_file_i/_6496_  (.A0(\register_file_i/rf_reg_508_ ),
    .A1(net577),
    .S(net816),
    .X(\register_file_i/_0450_ ));
 sg13g2_mux2_1 \register_file_i/_6497_  (.A0(\register_file_i/rf_reg_509_ ),
    .A1(net567),
    .S(net814),
    .X(\register_file_i/_0451_ ));
 sg13g2_mux2_1 \register_file_i/_6498_  (.A0(net706),
    .A1(\register_file_i/rf_reg_50_ ),
    .S(net836),
    .X(\register_file_i/_0452_ ));
 sg13g2_mux2_1 \register_file_i/_6499_  (.A0(\register_file_i/rf_reg_510_ ),
    .A1(net575),
    .S(net817),
    .X(\register_file_i/_0453_ ));
 sg13g2_mux2_1 \register_file_i/_6500_  (.A0(\register_file_i/rf_reg_511_ ),
    .A1(net562),
    .S(net817),
    .X(\register_file_i/_0454_ ));
 sg13g2_and3_2 \register_file_i/_6501_  (.X(\register_file_i/_2940_ ),
    .A(net553),
    .B(rf_we_wb),
    .C(\register_file_i/_2866_ ));
 sg13g2_nand2_2 \register_file_i/_6502_  (.Y(\register_file_i/_2941_ ),
    .A(\register_file_i/_2815_ ),
    .B(\register_file_i/_2940_ ));
 sg13g2_buf_2 fanout93 (.A(net98),
    .X(net93));
 sg13g2_mux2_1 \register_file_i/_6504_  (.A0(net752),
    .A1(\register_file_i/rf_reg_512_ ),
    .S(net965),
    .X(\register_file_i/_0455_ ));
 sg13g2_mux2_1 \register_file_i/_6505_  (.A0(net1000),
    .A1(\register_file_i/rf_reg_513_ ),
    .S(net964),
    .X(\register_file_i/_0456_ ));
 sg13g2_mux2_1 \register_file_i/_6506_  (.A0(net885),
    .A1(\register_file_i/rf_reg_514_ ),
    .S(net964),
    .X(\register_file_i/_0457_ ));
 sg13g2_mux2_1 \register_file_i/_6507_  (.A0(net1023),
    .A1(\register_file_i/rf_reg_515_ ),
    .S(net964),
    .X(\register_file_i/_0458_ ));
 sg13g2_mux2_1 \register_file_i/_6508_  (.A0(net1016),
    .A1(\register_file_i/rf_reg_516_ ),
    .S(net964),
    .X(\register_file_i/_0459_ ));
 sg13g2_mux2_1 \register_file_i/_6509_  (.A0(net996),
    .A1(\register_file_i/rf_reg_517_ ),
    .S(net963),
    .X(\register_file_i/_0460_ ));
 sg13g2_mux2_1 \register_file_i/_6510_  (.A0(net881),
    .A1(\register_file_i/rf_reg_518_ ),
    .S(net964),
    .X(\register_file_i/_0461_ ));
 sg13g2_mux2_1 \register_file_i/_6511_  (.A0(net992),
    .A1(\register_file_i/rf_reg_519_ ),
    .S(net964),
    .X(\register_file_i/_0462_ ));
 sg13g2_mux2_1 \register_file_i/_6512_  (.A0(net701),
    .A1(\register_file_i/rf_reg_51_ ),
    .S(net836),
    .X(\register_file_i/_0463_ ));
 sg13g2_mux2_1 \register_file_i/_6513_  (.A0(net876),
    .A1(\register_file_i/rf_reg_520_ ),
    .S(net964),
    .X(\register_file_i/_0464_ ));
 sg13g2_mux2_1 \register_file_i/_6514_  (.A0(net805),
    .A1(\register_file_i/rf_reg_521_ ),
    .S(net963),
    .X(\register_file_i/_0465_ ));
 sg13g2_buf_2 fanout92 (.A(_05522_),
    .X(net92));
 sg13g2_mux2_1 \register_file_i/_6516_  (.A0(net796),
    .A1(\register_file_i/rf_reg_522_ ),
    .S(net963),
    .X(\register_file_i/_0466_ ));
 sg13g2_mux2_1 \register_file_i/_6517_  (.A0(net791),
    .A1(\register_file_i/rf_reg_523_ ),
    .S(net963),
    .X(\register_file_i/_0467_ ));
 sg13g2_mux2_1 \register_file_i/_6518_  (.A0(net799),
    .A1(\register_file_i/rf_reg_524_ ),
    .S(net963),
    .X(\register_file_i/_0468_ ));
 sg13g2_mux2_1 \register_file_i/_6519_  (.A0(net785),
    .A1(\register_file_i/rf_reg_525_ ),
    .S(net963),
    .X(\register_file_i/_0469_ ));
 sg13g2_mux2_1 \register_file_i/_6520_  (.A0(net748),
    .A1(\register_file_i/rf_reg_526_ ),
    .S(net966),
    .X(\register_file_i/_0470_ ));
 sg13g2_mux2_1 \register_file_i/_6521_  (.A0(net781),
    .A1(\register_file_i/rf_reg_527_ ),
    .S(net966),
    .X(\register_file_i/_0471_ ));
 sg13g2_mux2_1 \register_file_i/_6522_  (.A0(net709),
    .A1(\register_file_i/rf_reg_528_ ),
    .S(net966),
    .X(\register_file_i/_0472_ ));
 sg13g2_mux2_1 \register_file_i/_6523_  (.A0(net723),
    .A1(\register_file_i/rf_reg_529_ ),
    .S(net966),
    .X(\register_file_i/_0473_ ));
 sg13g2_buf_2 fanout91 (.A(net92),
    .X(net91));
 sg13g2_mux2_1 \register_file_i/_6525_  (.A0(net740),
    .A1(\register_file_i/rf_reg_52_ ),
    .S(net836),
    .X(\register_file_i/_0474_ ));
 sg13g2_mux2_1 \register_file_i/_6526_  (.A0(net704),
    .A1(\register_file_i/rf_reg_530_ ),
    .S(net966),
    .X(\register_file_i/_0475_ ));
 sg13g2_mux2_1 \register_file_i/_6527_  (.A0(net698),
    .A1(\register_file_i/rf_reg_531_ ),
    .S(net966),
    .X(\register_file_i/_0476_ ));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net92));
 sg13g2_mux2_1 \register_file_i/_6529_  (.A0(net736),
    .A1(\register_file_i/rf_reg_532_ ),
    .S(net967),
    .X(\register_file_i/_0477_ ));
 sg13g2_mux2_1 \register_file_i/_6530_  (.A0(net671),
    .A1(\register_file_i/rf_reg_533_ ),
    .S(net967),
    .X(\register_file_i/_0478_ ));
 sg13g2_mux2_1 \register_file_i/_6531_  (.A0(net693),
    .A1(\register_file_i/rf_reg_534_ ),
    .S(net967),
    .X(\register_file_i/_0479_ ));
 sg13g2_mux2_1 \register_file_i/_6532_  (.A0(net690),
    .A1(\register_file_i/rf_reg_535_ ),
    .S(net967),
    .X(\register_file_i/_0480_ ));
 sg13g2_mux2_1 \register_file_i/_6533_  (.A0(net683),
    .A1(\register_file_i/rf_reg_536_ ),
    .S(net965),
    .X(\register_file_i/_0481_ ));
 sg13g2_mux2_1 \register_file_i/_6534_  (.A0(net600),
    .A1(\register_file_i/rf_reg_537_ ),
    .S(net965),
    .X(\register_file_i/_0482_ ));
 sg13g2_mux2_1 \register_file_i/_6535_  (.A0(net666),
    .A1(\register_file_i/rf_reg_538_ ),
    .S(net963),
    .X(\register_file_i/_0483_ ));
 sg13g2_mux2_1 \register_file_i/_6536_  (.A0(net582),
    .A1(\register_file_i/rf_reg_539_ ),
    .S(net965),
    .X(\register_file_i/_0484_ ));
 sg13g2_mux2_1 \register_file_i/_6537_  (.A0(net673),
    .A1(\register_file_i/rf_reg_53_ ),
    .S(net836),
    .X(\register_file_i/_0485_ ));
 sg13g2_mux2_1 \register_file_i/_6538_  (.A0(net578),
    .A1(\register_file_i/rf_reg_540_ ),
    .S(net964),
    .X(\register_file_i/_0486_ ));
 sg13g2_mux2_1 \register_file_i/_6539_  (.A0(net568),
    .A1(\register_file_i/rf_reg_541_ ),
    .S(net963),
    .X(\register_file_i/_0487_ ));
 sg13g2_mux2_1 \register_file_i/_6540_  (.A0(net573),
    .A1(\register_file_i/rf_reg_542_ ),
    .S(net966),
    .X(\register_file_i/_0488_ ));
 sg13g2_mux2_1 \register_file_i/_6541_  (.A0(net563),
    .A1(\register_file_i/rf_reg_543_ ),
    .S(net966),
    .X(\register_file_i/_0489_ ));
 sg13g2_nand3_1 \register_file_i/_6542_  (.B(rf_we_wb),
    .C(\register_file_i/_2878_ ),
    .A(\id_stage_i.controller_i.instr_i_11_ ),
    .Y(\register_file_i/_2946_ ));
 sg13g2_nor3_2 \register_file_i/_6543_  (.A(net1991),
    .B(net2099),
    .C(\register_file_i/_2946_ ),
    .Y(\register_file_i/_2947_ ));
 sg13g2_buf_2 fanout89 (.A(_05924_),
    .X(net89));
 sg13g2_mux2_1 \register_file_i/_6545_  (.A0(\register_file_i/rf_reg_544_ ),
    .A1(net752),
    .S(net960),
    .X(\register_file_i/_0490_ ));
 sg13g2_mux2_1 \register_file_i/_6546_  (.A0(\register_file_i/rf_reg_545_ ),
    .A1(net1000),
    .S(net959),
    .X(\register_file_i/_0491_ ));
 sg13g2_mux2_1 \register_file_i/_6547_  (.A0(\register_file_i/rf_reg_546_ ),
    .A1(net885),
    .S(net959),
    .X(\register_file_i/_0492_ ));
 sg13g2_mux2_1 \register_file_i/_6548_  (.A0(\register_file_i/rf_reg_547_ ),
    .A1(net1023),
    .S(net959),
    .X(\register_file_i/_0493_ ));
 sg13g2_mux2_1 \register_file_i/_6549_  (.A0(\register_file_i/rf_reg_548_ ),
    .A1(net1016),
    .S(net959),
    .X(\register_file_i/_0494_ ));
 sg13g2_mux2_1 \register_file_i/_6550_  (.A0(\register_file_i/rf_reg_549_ ),
    .A1(net996),
    .S(net958),
    .X(\register_file_i/_0495_ ));
 sg13g2_mux2_1 \register_file_i/_6551_  (.A0(net695),
    .A1(\register_file_i/rf_reg_54_ ),
    .S(net835),
    .X(\register_file_i/_0496_ ));
 sg13g2_mux2_1 \register_file_i/_6552_  (.A0(\register_file_i/rf_reg_550_ ),
    .A1(net881),
    .S(net959),
    .X(\register_file_i/_0497_ ));
 sg13g2_mux2_1 \register_file_i/_6553_  (.A0(\register_file_i/rf_reg_551_ ),
    .A1(net992),
    .S(net959),
    .X(\register_file_i/_0498_ ));
 sg13g2_mux2_1 \register_file_i/_6554_  (.A0(\register_file_i/rf_reg_552_ ),
    .A1(net876),
    .S(net959),
    .X(\register_file_i/_0499_ ));
 sg13g2_mux2_1 \register_file_i/_6555_  (.A0(\register_file_i/rf_reg_553_ ),
    .A1(net805),
    .S(net958),
    .X(\register_file_i/_0500_ ));
 sg13g2_buf_2 fanout88 (.A(alu_operand_a_ex_26_),
    .X(net88));
 sg13g2_mux2_1 \register_file_i/_6557_  (.A0(\register_file_i/rf_reg_554_ ),
    .A1(net796),
    .S(net958),
    .X(\register_file_i/_0501_ ));
 sg13g2_mux2_1 \register_file_i/_6558_  (.A0(\register_file_i/rf_reg_555_ ),
    .A1(net791),
    .S(net958),
    .X(\register_file_i/_0502_ ));
 sg13g2_mux2_1 \register_file_i/_6559_  (.A0(\register_file_i/rf_reg_556_ ),
    .A1(net799),
    .S(net958),
    .X(\register_file_i/_0503_ ));
 sg13g2_mux2_1 \register_file_i/_6560_  (.A0(\register_file_i/rf_reg_557_ ),
    .A1(net785),
    .S(net958),
    .X(\register_file_i/_0504_ ));
 sg13g2_mux2_1 \register_file_i/_6561_  (.A0(\register_file_i/rf_reg_558_ ),
    .A1(net748),
    .S(net961),
    .X(\register_file_i/_0505_ ));
 sg13g2_mux2_1 \register_file_i/_6562_  (.A0(\register_file_i/rf_reg_559_ ),
    .A1(net781),
    .S(net961),
    .X(\register_file_i/_0506_ ));
 sg13g2_mux2_1 \register_file_i/_6563_  (.A0(net692),
    .A1(\register_file_i/rf_reg_55_ ),
    .S(net835),
    .X(\register_file_i/_0507_ ));
 sg13g2_mux2_1 \register_file_i/_6564_  (.A0(\register_file_i/rf_reg_560_ ),
    .A1(net708),
    .S(net961),
    .X(\register_file_i/_0508_ ));
 sg13g2_mux2_1 \register_file_i/_6565_  (.A0(\register_file_i/rf_reg_561_ ),
    .A1(net723),
    .S(net961),
    .X(\register_file_i/_0509_ ));
 sg13g2_mux2_1 \register_file_i/_6566_  (.A0(\register_file_i/rf_reg_562_ ),
    .A1(net704),
    .S(net961),
    .X(\register_file_i/_0510_ ));
 sg13g2_mux2_1 \register_file_i/_6567_  (.A0(\register_file_i/rf_reg_563_ ),
    .A1(net698),
    .S(net961),
    .X(\register_file_i/_0511_ ));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(net88));
 sg13g2_mux2_1 \register_file_i/_6569_  (.A0(\register_file_i/rf_reg_564_ ),
    .A1(net737),
    .S(net962),
    .X(\register_file_i/_0512_ ));
 sg13g2_mux2_1 \register_file_i/_6570_  (.A0(\register_file_i/rf_reg_565_ ),
    .A1(net671),
    .S(net962),
    .X(\register_file_i/_0513_ ));
 sg13g2_mux2_1 \register_file_i/_6571_  (.A0(\register_file_i/rf_reg_566_ ),
    .A1(net693),
    .S(net962),
    .X(\register_file_i/_0514_ ));
 sg13g2_mux2_1 \register_file_i/_6572_  (.A0(\register_file_i/rf_reg_567_ ),
    .A1(net690),
    .S(net962),
    .X(\register_file_i/_0515_ ));
 sg13g2_mux2_1 \register_file_i/_6573_  (.A0(\register_file_i/rf_reg_568_ ),
    .A1(net683),
    .S(net960),
    .X(\register_file_i/_0516_ ));
 sg13g2_mux2_1 \register_file_i/_6574_  (.A0(\register_file_i/rf_reg_569_ ),
    .A1(net601),
    .S(net960),
    .X(\register_file_i/_0517_ ));
 sg13g2_mux2_1 \register_file_i/_6575_  (.A0(net686),
    .A1(\register_file_i/rf_reg_56_ ),
    .S(net834),
    .X(\register_file_i/_0518_ ));
 sg13g2_mux2_1 \register_file_i/_6576_  (.A0(\register_file_i/rf_reg_570_ ),
    .A1(net666),
    .S(net958),
    .X(\register_file_i/_0519_ ));
 sg13g2_mux2_1 \register_file_i/_6577_  (.A0(\register_file_i/rf_reg_571_ ),
    .A1(net582),
    .S(net960),
    .X(\register_file_i/_0520_ ));
 sg13g2_mux2_1 \register_file_i/_6578_  (.A0(\register_file_i/rf_reg_572_ ),
    .A1(net577),
    .S(net959),
    .X(\register_file_i/_0521_ ));
 sg13g2_mux2_1 \register_file_i/_6579_  (.A0(\register_file_i/rf_reg_573_ ),
    .A1(net568),
    .S(net958),
    .X(\register_file_i/_0522_ ));
 sg13g2_mux2_1 \register_file_i/_6580_  (.A0(\register_file_i/rf_reg_574_ ),
    .A1(net573),
    .S(net961),
    .X(\register_file_i/_0523_ ));
 sg13g2_mux2_1 \register_file_i/_6581_  (.A0(\register_file_i/rf_reg_575_ ),
    .A1(net563),
    .S(net961),
    .X(\register_file_i/_0524_ ));
 sg13g2_nand3_1 \register_file_i/_6582_  (.B(rf_we_wb),
    .C(\register_file_i/_2884_ ),
    .A(\id_stage_i.controller_i.instr_i_11_ ),
    .Y(\register_file_i/_2951_ ));
 sg13g2_nor3_2 \register_file_i/_6583_  (.A(net1991),
    .B(net2099),
    .C(\register_file_i/_2951_ ),
    .Y(\register_file_i/_2952_ ));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(_03234_));
 sg13g2_mux2_1 \register_file_i/_6585_  (.A0(\register_file_i/rf_reg_576_ ),
    .A1(net753),
    .S(net955),
    .X(\register_file_i/_0525_ ));
 sg13g2_mux2_1 \register_file_i/_6586_  (.A0(\register_file_i/rf_reg_577_ ),
    .A1(net1000),
    .S(net954),
    .X(\register_file_i/_0526_ ));
 sg13g2_mux2_1 \register_file_i/_6587_  (.A0(\register_file_i/rf_reg_578_ ),
    .A1(net885),
    .S(net954),
    .X(\register_file_i/_0527_ ));
 sg13g2_mux2_1 \register_file_i/_6588_  (.A0(\register_file_i/rf_reg_579_ ),
    .A1(net1023),
    .S(net954),
    .X(\register_file_i/_0528_ ));
 sg13g2_mux2_1 \register_file_i/_6589_  (.A0(net602),
    .A1(\register_file_i/rf_reg_57_ ),
    .S(net834),
    .X(\register_file_i/_0529_ ));
 sg13g2_mux2_1 \register_file_i/_6590_  (.A0(\register_file_i/rf_reg_580_ ),
    .A1(net1016),
    .S(net954),
    .X(\register_file_i/_0530_ ));
 sg13g2_mux2_1 \register_file_i/_6591_  (.A0(\register_file_i/rf_reg_581_ ),
    .A1(net996),
    .S(net952),
    .X(\register_file_i/_0531_ ));
 sg13g2_mux2_1 \register_file_i/_6592_  (.A0(\register_file_i/rf_reg_582_ ),
    .A1(net881),
    .S(net954),
    .X(\register_file_i/_0532_ ));
 sg13g2_mux2_1 \register_file_i/_6593_  (.A0(\register_file_i/rf_reg_583_ ),
    .A1(net992),
    .S(net954),
    .X(\register_file_i/_0533_ ));
 sg13g2_buf_4 fanout85 (.X(net85),
    .A(net86));
 sg13g2_mux2_1 \register_file_i/_6595_  (.A0(\register_file_i/rf_reg_584_ ),
    .A1(net876),
    .S(net954),
    .X(\register_file_i/_0534_ ));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net86));
 sg13g2_mux2_1 \register_file_i/_6597_  (.A0(\register_file_i/rf_reg_585_ ),
    .A1(net805),
    .S(net952),
    .X(\register_file_i/_0535_ ));
 sg13g2_buf_2 fanout83 (.A(net86),
    .X(net83));
 sg13g2_buf_4 fanout82 (.X(net82),
    .A(net86));
 sg13g2_mux2_1 \register_file_i/_6600_  (.A0(\register_file_i/rf_reg_586_ ),
    .A1(net796),
    .S(net952),
    .X(\register_file_i/_0536_ ));
 sg13g2_buf_2 fanout81 (.A(alu_operand_a_ex_31_),
    .X(net81));
 sg13g2_mux2_1 \register_file_i/_6602_  (.A0(\register_file_i/rf_reg_587_ ),
    .A1(net791),
    .S(net952),
    .X(\register_file_i/_0537_ ));
 sg13g2_buf_2 fanout80 (.A(csr_addr_1_),
    .X(net80));
 sg13g2_mux2_1 \register_file_i/_6604_  (.A0(\register_file_i/rf_reg_588_ ),
    .A1(net799),
    .S(net952),
    .X(\register_file_i/_0538_ ));
 sg13g2_buf_4 fanout79 (.X(net79),
    .A(net80));
 sg13g2_mux2_1 \register_file_i/_6606_  (.A0(\register_file_i/rf_reg_589_ ),
    .A1(net785),
    .S(net953),
    .X(\register_file_i/_0539_ ));
 sg13g2_mux2_1 \register_file_i/_6607_  (.A0(net667),
    .A1(\register_file_i/rf_reg_58_ ),
    .S(net833),
    .X(\register_file_i/_0540_ ));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(net80));
 sg13g2_mux2_1 \register_file_i/_6609_  (.A0(\register_file_i/rf_reg_590_ ),
    .A1(net748),
    .S(net953),
    .X(\register_file_i/_0541_ ));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(net79));
 sg13g2_mux2_1 \register_file_i/_6611_  (.A0(\register_file_i/rf_reg_591_ ),
    .A1(net781),
    .S(net956),
    .X(\register_file_i/_0542_ ));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(net79));
 sg13g2_mux2_1 \register_file_i/_6613_  (.A0(\register_file_i/rf_reg_592_ ),
    .A1(net708),
    .S(net956),
    .X(\register_file_i/_0543_ ));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(net79));
 sg13g2_mux2_1 \register_file_i/_6615_  (.A0(\register_file_i/rf_reg_593_ ),
    .A1(net724),
    .S(net956),
    .X(\register_file_i/_0544_ ));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(net80));
 sg13g2_mux2_1 \register_file_i/_6617_  (.A0(\register_file_i/rf_reg_594_ ),
    .A1(net704),
    .S(net956),
    .X(\register_file_i/_0545_ ));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(net78));
 sg13g2_mux2_1 \register_file_i/_6619_  (.A0(\register_file_i/rf_reg_595_ ),
    .A1(net702),
    .S(net956),
    .X(\register_file_i/_0546_ ));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(net78));
 sg13g2_buf_8 fanout71 (.A(net78),
    .X(net71));
 sg13g2_mux2_1 \register_file_i/_6622_  (.A0(\register_file_i/rf_reg_596_ ),
    .A1(net737),
    .S(net957),
    .X(\register_file_i/_0547_ ));
 sg13g2_buf_8 fanout70 (.A(net78),
    .X(net70));
 sg13g2_mux2_1 \register_file_i/_6624_  (.A0(\register_file_i/rf_reg_597_ ),
    .A1(net671),
    .S(net956),
    .X(\register_file_i/_0548_ ));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(net78));
 sg13g2_mux2_1 \register_file_i/_6626_  (.A0(\register_file_i/rf_reg_598_ ),
    .A1(net693),
    .S(net957),
    .X(\register_file_i/_0549_ ));
 sg13g2_buf_8 fanout68 (.A(net78),
    .X(net68));
 sg13g2_mux2_1 \register_file_i/_6628_  (.A0(\register_file_i/rf_reg_599_ ),
    .A1(net690),
    .S(net957),
    .X(\register_file_i/_0550_ ));
 sg13g2_mux2_1 \register_file_i/_6629_  (.A0(net585),
    .A1(\register_file_i/rf_reg_59_ ),
    .S(net833),
    .X(\register_file_i/_0551_ ));
 sg13g2_buf_8 fanout67 (.A(net78),
    .X(net67));
 sg13g2_mux2_1 \register_file_i/_6631_  (.A0(\register_file_i/rf_reg_600_ ),
    .A1(net683),
    .S(net953),
    .X(\register_file_i/_0552_ ));
 sg13g2_buf_8 fanout66 (.A(net78),
    .X(net66));
 sg13g2_mux2_1 \register_file_i/_6633_  (.A0(\register_file_i/rf_reg_601_ ),
    .A1(net601),
    .S(net953),
    .X(\register_file_i/_0553_ ));
 sg13g2_buf_8 fanout65 (.A(net79),
    .X(net65));
 sg13g2_mux2_1 \register_file_i/_6635_  (.A0(\register_file_i/rf_reg_602_ ),
    .A1(net666),
    .S(net952),
    .X(\register_file_i/_0554_ ));
 sg13g2_buf_4 fanout64 (.X(net64),
    .A(net79));
 sg13g2_mux2_1 \register_file_i/_6637_  (.A0(\register_file_i/rf_reg_603_ ),
    .A1(net582),
    .S(net952),
    .X(\register_file_i/_0555_ ));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(net79));
 sg13g2_mux2_1 \register_file_i/_6639_  (.A0(\register_file_i/rf_reg_604_ ),
    .A1(net578),
    .S(net954),
    .X(\register_file_i/_0556_ ));
 sg13g2_buf_8 fanout62 (.A(net79),
    .X(net62));
 sg13g2_mux2_1 \register_file_i/_6641_  (.A0(\register_file_i/rf_reg_605_ ),
    .A1(net568),
    .S(net952),
    .X(\register_file_i/_0557_ ));
 sg13g2_buf_2 fanout61 (.A(net79),
    .X(net61));
 sg13g2_mux2_1 \register_file_i/_6643_  (.A0(\register_file_i/rf_reg_606_ ),
    .A1(net573),
    .S(net956),
    .X(\register_file_i/_0558_ ));
 sg13g2_buf_2 fanout60 (.A(\cs_registers_i/_0486_ ),
    .X(net60));
 sg13g2_mux2_1 \register_file_i/_6645_  (.A0(\register_file_i/rf_reg_607_ ),
    .A1(net563),
    .S(net956),
    .X(\register_file_i/_0559_ ));
 sg13g2_buf_2 fanout59 (.A(\cs_registers_i/_0486_ ),
    .X(net59));
 sg13g2_nor2b_2 \register_file_i/_6647_  (.A(\register_file_i/_2800_ ),
    .B_N(\register_file_i/_2815_ ),
    .Y(\register_file_i/_2981_ ));
 sg13g2_buf_2 fanout58 (.A(\cs_registers_i/_0510_ ),
    .X(net58));
 sg13g2_mux2_1 \register_file_i/_6649_  (.A0(\register_file_i/rf_reg_608_ ),
    .A1(net752),
    .S(net949),
    .X(\register_file_i/_0560_ ));
 sg13g2_buf_2 fanout57 (.A(\cs_registers_i/_0510_ ),
    .X(net57));
 sg13g2_mux2_1 \register_file_i/_6651_  (.A0(\register_file_i/rf_reg_609_ ),
    .A1(net1001),
    .S(net948),
    .X(\register_file_i/_0561_ ));
 sg13g2_mux2_1 \register_file_i/_6652_  (.A0(net579),
    .A1(\register_file_i/rf_reg_60_ ),
    .S(net833),
    .X(\register_file_i/_0562_ ));
 sg13g2_buf_2 fanout56 (.A(\cs_registers_i/_0510_ ),
    .X(net56));
 sg13g2_mux2_1 \register_file_i/_6654_  (.A0(\register_file_i/rf_reg_610_ ),
    .A1(net887),
    .S(net948),
    .X(\register_file_i/_0563_ ));
 sg13g2_buf_1 fanout55 (.A(\cs_registers_i/_0562_ ),
    .X(net55));
 sg13g2_mux2_1 \register_file_i/_6656_  (.A0(\register_file_i/rf_reg_611_ ),
    .A1(net1023),
    .S(net948),
    .X(\register_file_i/_0564_ ));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(\cs_registers_i/_0562_ ));
 sg13g2_mux2_1 \register_file_i/_6658_  (.A0(\register_file_i/rf_reg_612_ ),
    .A1(net1016),
    .S(net948),
    .X(\register_file_i/_0565_ ));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(\cs_registers_i/_0562_ ));
 sg13g2_mux2_1 \register_file_i/_6660_  (.A0(\register_file_i/rf_reg_613_ ),
    .A1(net996),
    .S(net947),
    .X(\register_file_i/_0566_ ));
 sg13g2_buf_2 fanout52 (.A(_04541_),
    .X(net52));
 sg13g2_mux2_1 \register_file_i/_6662_  (.A0(\register_file_i/rf_reg_614_ ),
    .A1(net881),
    .S(net948),
    .X(\register_file_i/_0567_ ));
 sg13g2_buf_2 fanout51 (.A(net52),
    .X(net51));
 sg13g2_mux2_1 \register_file_i/_6664_  (.A0(\register_file_i/rf_reg_615_ ),
    .A1(net992),
    .S(net948),
    .X(\register_file_i/_0568_ ));
 sg13g2_mux2_1 \register_file_i/_6665_  (.A0(\register_file_i/rf_reg_616_ ),
    .A1(net876),
    .S(net948),
    .X(\register_file_i/_0569_ ));
 sg13g2_mux2_1 \register_file_i/_6666_  (.A0(\register_file_i/rf_reg_617_ ),
    .A1(net805),
    .S(net947),
    .X(\register_file_i/_0570_ ));
 sg13g2_buf_2 fanout50 (.A(_08068_),
    .X(net50));
 sg13g2_mux2_1 \register_file_i/_6668_  (.A0(\register_file_i/rf_reg_618_ ),
    .A1(net796),
    .S(net947),
    .X(\register_file_i/_0571_ ));
 sg13g2_mux2_1 \register_file_i/_6669_  (.A0(\register_file_i/rf_reg_619_ ),
    .A1(net791),
    .S(net947),
    .X(\register_file_i/_0572_ ));
 sg13g2_mux2_1 \register_file_i/_6670_  (.A0(net572),
    .A1(\register_file_i/rf_reg_61_ ),
    .S(net832),
    .X(\register_file_i/_0573_ ));
 sg13g2_mux2_1 \register_file_i/_6671_  (.A0(\register_file_i/rf_reg_620_ ),
    .A1(net799),
    .S(net947),
    .X(\register_file_i/_0574_ ));
 sg13g2_mux2_1 \register_file_i/_6672_  (.A0(\register_file_i/rf_reg_621_ ),
    .A1(net785),
    .S(net947),
    .X(\register_file_i/_0575_ ));
 sg13g2_mux2_1 \register_file_i/_6673_  (.A0(\register_file_i/rf_reg_622_ ),
    .A1(net748),
    .S(net950),
    .X(\register_file_i/_0576_ ));
 sg13g2_mux2_1 \register_file_i/_6674_  (.A0(\register_file_i/rf_reg_623_ ),
    .A1(net781),
    .S(net950),
    .X(\register_file_i/_0577_ ));
 sg13g2_mux2_1 \register_file_i/_6675_  (.A0(\register_file_i/rf_reg_624_ ),
    .A1(net709),
    .S(net950),
    .X(\register_file_i/_0578_ ));
 sg13g2_mux2_1 \register_file_i/_6676_  (.A0(\register_file_i/rf_reg_625_ ),
    .A1(net727),
    .S(net950),
    .X(\register_file_i/_0579_ ));
 sg13g2_mux2_1 \register_file_i/_6677_  (.A0(\register_file_i/rf_reg_626_ ),
    .A1(net704),
    .S(net950),
    .X(\register_file_i/_0580_ ));
 sg13g2_mux2_1 \register_file_i/_6678_  (.A0(\register_file_i/rf_reg_627_ ),
    .A1(net699),
    .S(net950),
    .X(\register_file_i/_0581_ ));
 sg13g2_buf_2 fanout49 (.A(net50),
    .X(net49));
 sg13g2_mux2_1 \register_file_i/_6680_  (.A0(\register_file_i/rf_reg_628_ ),
    .A1(net737),
    .S(net951),
    .X(\register_file_i/_0582_ ));
 sg13g2_mux2_1 \register_file_i/_6681_  (.A0(\register_file_i/rf_reg_629_ ),
    .A1(net671),
    .S(net951),
    .X(\register_file_i/_0583_ ));
 sg13g2_mux2_1 \register_file_i/_6682_  (.A0(net576),
    .A1(\register_file_i/rf_reg_62_ ),
    .S(net835),
    .X(\register_file_i/_0584_ ));
 sg13g2_mux2_1 \register_file_i/_6683_  (.A0(\register_file_i/rf_reg_630_ ),
    .A1(net693),
    .S(net951),
    .X(\register_file_i/_0585_ ));
 sg13g2_mux2_1 \register_file_i/_6684_  (.A0(\register_file_i/rf_reg_631_ ),
    .A1(net690),
    .S(net951),
    .X(\register_file_i/_0586_ ));
 sg13g2_mux2_1 \register_file_i/_6685_  (.A0(\register_file_i/rf_reg_632_ ),
    .A1(net683),
    .S(net949),
    .X(\register_file_i/_0587_ ));
 sg13g2_mux2_1 \register_file_i/_6686_  (.A0(\register_file_i/rf_reg_633_ ),
    .A1(net601),
    .S(net949),
    .X(\register_file_i/_0588_ ));
 sg13g2_mux2_1 \register_file_i/_6687_  (.A0(\register_file_i/rf_reg_634_ ),
    .A1(net666),
    .S(net947),
    .X(\register_file_i/_0589_ ));
 sg13g2_mux2_1 \register_file_i/_6688_  (.A0(\register_file_i/rf_reg_635_ ),
    .A1(net583),
    .S(net949),
    .X(\register_file_i/_0590_ ));
 sg13g2_mux2_1 \register_file_i/_6689_  (.A0(\register_file_i/rf_reg_636_ ),
    .A1(net578),
    .S(net948),
    .X(\register_file_i/_0591_ ));
 sg13g2_mux2_1 \register_file_i/_6690_  (.A0(\register_file_i/rf_reg_637_ ),
    .A1(net568),
    .S(net947),
    .X(\register_file_i/_0592_ ));
 sg13g2_mux2_1 \register_file_i/_6691_  (.A0(\register_file_i/rf_reg_638_ ),
    .A1(net573),
    .S(net950),
    .X(\register_file_i/_0593_ ));
 sg13g2_mux2_1 \register_file_i/_6692_  (.A0(\register_file_i/rf_reg_639_ ),
    .A1(net563),
    .S(net950),
    .X(\register_file_i/_0594_ ));
 sg13g2_mux2_1 \register_file_i/_6693_  (.A0(net565),
    .A1(\register_file_i/rf_reg_63_ ),
    .S(net835),
    .X(\register_file_i/_0595_ ));
 sg13g2_nand2b_1 \register_file_i/_6694_  (.Y(\register_file_i/_2992_ ),
    .B(\register_file_i/_2940_ ),
    .A_N(\register_file_i/_2868_ ));
 sg13g2_buf_2 fanout48 (.A(net50),
    .X(net48));
 sg13g2_buf_2 fanout47 (.A(_08502_),
    .X(net47));
 sg13g2_mux2_1 \register_file_i/_6697_  (.A0(net752),
    .A1(\register_file_i/rf_reg_640_ ),
    .S(net942),
    .X(\register_file_i/_0596_ ));
 sg13g2_mux2_1 \register_file_i/_6698_  (.A0(net1000),
    .A1(\register_file_i/rf_reg_641_ ),
    .S(net941),
    .X(\register_file_i/_0597_ ));
 sg13g2_mux2_1 \register_file_i/_6699_  (.A0(net885),
    .A1(\register_file_i/rf_reg_642_ ),
    .S(net943),
    .X(\register_file_i/_0598_ ));
 sg13g2_mux2_1 \register_file_i/_6700_  (.A0(net1020),
    .A1(\register_file_i/rf_reg_643_ ),
    .S(net943),
    .X(\register_file_i/_0599_ ));
 sg13g2_mux2_1 \register_file_i/_6701_  (.A0(net1016),
    .A1(\register_file_i/rf_reg_644_ ),
    .S(net943),
    .X(\register_file_i/_0600_ ));
 sg13g2_mux2_1 \register_file_i/_6702_  (.A0(net996),
    .A1(\register_file_i/rf_reg_645_ ),
    .S(net941),
    .X(\register_file_i/_0601_ ));
 sg13g2_mux2_1 \register_file_i/_6703_  (.A0(net881),
    .A1(\register_file_i/rf_reg_646_ ),
    .S(net943),
    .X(\register_file_i/_0602_ ));
 sg13g2_mux2_1 \register_file_i/_6704_  (.A0(net992),
    .A1(\register_file_i/rf_reg_647_ ),
    .S(net943),
    .X(\register_file_i/_0603_ ));
 sg13g2_mux2_1 \register_file_i/_6705_  (.A0(net876),
    .A1(\register_file_i/rf_reg_648_ ),
    .S(net941),
    .X(\register_file_i/_0604_ ));
 sg13g2_mux2_1 \register_file_i/_6706_  (.A0(net805),
    .A1(\register_file_i/rf_reg_649_ ),
    .S(net941),
    .X(\register_file_i/_0605_ ));
 sg13g2_nand2_2 \register_file_i/_6707_  (.Y(\register_file_i/_2995_ ),
    .A(\register_file_i/_2816_ ),
    .B(\register_file_i/_2884_ ));
 sg13g2_buf_1 fanout46 (.A(net47),
    .X(net46));
 sg13g2_mux2_1 \register_file_i/_6709_  (.A0(net756),
    .A1(\register_file_i/rf_reg_64_ ),
    .S(net809),
    .X(\register_file_i/_0606_ ));
 sg13g2_buf_2 fanout45 (.A(net47),
    .X(net45));
 sg13g2_mux2_1 \register_file_i/_6711_  (.A0(net796),
    .A1(\register_file_i/rf_reg_650_ ),
    .S(net941),
    .X(\register_file_i/_0607_ ));
 sg13g2_mux2_1 \register_file_i/_6712_  (.A0(net791),
    .A1(\register_file_i/rf_reg_651_ ),
    .S(net941),
    .X(\register_file_i/_0608_ ));
 sg13g2_mux2_1 \register_file_i/_6713_  (.A0(net799),
    .A1(\register_file_i/rf_reg_652_ ),
    .S(net941),
    .X(\register_file_i/_0609_ ));
 sg13g2_mux2_1 \register_file_i/_6714_  (.A0(net787),
    .A1(\register_file_i/rf_reg_653_ ),
    .S(net944),
    .X(\register_file_i/_0610_ ));
 sg13g2_mux2_1 \register_file_i/_6715_  (.A0(net749),
    .A1(\register_file_i/rf_reg_654_ ),
    .S(net944),
    .X(\register_file_i/_0611_ ));
 sg13g2_mux2_1 \register_file_i/_6716_  (.A0(net781),
    .A1(\register_file_i/rf_reg_655_ ),
    .S(net944),
    .X(\register_file_i/_0612_ ));
 sg13g2_mux2_1 \register_file_i/_6717_  (.A0(net709),
    .A1(\register_file_i/rf_reg_656_ ),
    .S(net945),
    .X(\register_file_i/_0613_ ));
 sg13g2_mux2_1 \register_file_i/_6718_  (.A0(net723),
    .A1(\register_file_i/rf_reg_657_ ),
    .S(net945),
    .X(\register_file_i/_0614_ ));
 sg13g2_mux2_1 \register_file_i/_6719_  (.A0(net704),
    .A1(\register_file_i/rf_reg_658_ ),
    .S(net945),
    .X(\register_file_i/_0615_ ));
 sg13g2_mux2_1 \register_file_i/_6720_  (.A0(net698),
    .A1(\register_file_i/rf_reg_659_ ),
    .S(net944),
    .X(\register_file_i/_0616_ ));
 sg13g2_mux2_1 \register_file_i/_6721_  (.A0(net1003),
    .A1(\register_file_i/rf_reg_65_ ),
    .S(net809),
    .X(\register_file_i/_0617_ ));
 sg13g2_buf_1 fanout44 (.A(_08575_),
    .X(net44));
 sg13g2_mux2_1 \register_file_i/_6723_  (.A0(net738),
    .A1(\register_file_i/rf_reg_660_ ),
    .S(net945),
    .X(\register_file_i/_0618_ ));
 sg13g2_mux2_1 \register_file_i/_6724_  (.A0(net672),
    .A1(\register_file_i/rf_reg_661_ ),
    .S(net945),
    .X(\register_file_i/_0619_ ));
 sg13g2_mux2_1 \register_file_i/_6725_  (.A0(net693),
    .A1(\register_file_i/rf_reg_662_ ),
    .S(net946),
    .X(\register_file_i/_0620_ ));
 sg13g2_mux2_1 \register_file_i/_6726_  (.A0(net687),
    .A1(\register_file_i/rf_reg_663_ ),
    .S(net944),
    .X(\register_file_i/_0621_ ));
 sg13g2_mux2_1 \register_file_i/_6727_  (.A0(net683),
    .A1(\register_file_i/rf_reg_664_ ),
    .S(net944),
    .X(\register_file_i/_0622_ ));
 sg13g2_mux2_1 \register_file_i/_6728_  (.A0(net599),
    .A1(\register_file_i/rf_reg_665_ ),
    .S(net942),
    .X(\register_file_i/_0623_ ));
 sg13g2_mux2_1 \register_file_i/_6729_  (.A0(net666),
    .A1(\register_file_i/rf_reg_666_ ),
    .S(net941),
    .X(\register_file_i/_0624_ ));
 sg13g2_mux2_1 \register_file_i/_6730_  (.A0(net582),
    .A1(\register_file_i/rf_reg_667_ ),
    .S(net942),
    .X(\register_file_i/_0625_ ));
 sg13g2_mux2_1 \register_file_i/_6731_  (.A0(net578),
    .A1(\register_file_i/rf_reg_668_ ),
    .S(net943),
    .X(\register_file_i/_0626_ ));
 sg13g2_mux2_1 \register_file_i/_6732_  (.A0(net568),
    .A1(\register_file_i/rf_reg_669_ ),
    .S(net942),
    .X(\register_file_i/_0627_ ));
 sg13g2_mux2_1 \register_file_i/_6733_  (.A0(net887),
    .A1(\register_file_i/rf_reg_66_ ),
    .S(net809),
    .X(\register_file_i/_0628_ ));
 sg13g2_mux2_1 \register_file_i/_6734_  (.A0(net573),
    .A1(\register_file_i/rf_reg_670_ ),
    .S(net944),
    .X(\register_file_i/_0629_ ));
 sg13g2_mux2_1 \register_file_i/_6735_  (.A0(net563),
    .A1(\register_file_i/rf_reg_671_ ),
    .S(net944),
    .X(\register_file_i/_0630_ ));
 sg13g2_nor2_2 \register_file_i/_6736_  (.A(\register_file_i/_2868_ ),
    .B(\register_file_i/_2946_ ),
    .Y(\register_file_i/_2999_ ));
 sg13g2_buf_2 fanout43 (.A(net44),
    .X(net43));
 sg13g2_mux2_1 \register_file_i/_6738_  (.A0(\register_file_i/rf_reg_672_ ),
    .A1(net752),
    .S(net937),
    .X(\register_file_i/_0631_ ));
 sg13g2_mux2_1 \register_file_i/_6739_  (.A0(\register_file_i/rf_reg_673_ ),
    .A1(net1000),
    .S(net936),
    .X(\register_file_i/_0632_ ));
 sg13g2_mux2_1 \register_file_i/_6740_  (.A0(\register_file_i/rf_reg_674_ ),
    .A1(net887),
    .S(net938),
    .X(\register_file_i/_0633_ ));
 sg13g2_mux2_1 \register_file_i/_6741_  (.A0(\register_file_i/rf_reg_675_ ),
    .A1(net1023),
    .S(net938),
    .X(\register_file_i/_0634_ ));
 sg13g2_mux2_1 \register_file_i/_6742_  (.A0(\register_file_i/rf_reg_676_ ),
    .A1(net1016),
    .S(net938),
    .X(\register_file_i/_0635_ ));
 sg13g2_mux2_1 \register_file_i/_6743_  (.A0(\register_file_i/rf_reg_677_ ),
    .A1(net996),
    .S(net936),
    .X(\register_file_i/_0636_ ));
 sg13g2_mux2_1 \register_file_i/_6744_  (.A0(\register_file_i/rf_reg_678_ ),
    .A1(net881),
    .S(net938),
    .X(\register_file_i/_0637_ ));
 sg13g2_mux2_1 \register_file_i/_6745_  (.A0(\register_file_i/rf_reg_679_ ),
    .A1(net992),
    .S(net938),
    .X(\register_file_i/_0638_ ));
 sg13g2_mux2_1 \register_file_i/_6746_  (.A0(net1024),
    .A1(\register_file_i/rf_reg_67_ ),
    .S(net809),
    .X(\register_file_i/_0639_ ));
 sg13g2_mux2_1 \register_file_i/_6747_  (.A0(\register_file_i/rf_reg_680_ ),
    .A1(net876),
    .S(net936),
    .X(\register_file_i/_0640_ ));
 sg13g2_mux2_1 \register_file_i/_6748_  (.A0(\register_file_i/rf_reg_681_ ),
    .A1(net805),
    .S(net936),
    .X(\register_file_i/_0641_ ));
 sg13g2_buf_2 fanout42 (.A(net43),
    .X(net42));
 sg13g2_mux2_1 \register_file_i/_6750_  (.A0(\register_file_i/rf_reg_682_ ),
    .A1(net796),
    .S(net936),
    .X(\register_file_i/_0642_ ));
 sg13g2_mux2_1 \register_file_i/_6751_  (.A0(\register_file_i/rf_reg_683_ ),
    .A1(net791),
    .S(net936),
    .X(\register_file_i/_0643_ ));
 sg13g2_mux2_1 \register_file_i/_6752_  (.A0(\register_file_i/rf_reg_684_ ),
    .A1(net799),
    .S(net936),
    .X(\register_file_i/_0644_ ));
 sg13g2_mux2_1 \register_file_i/_6753_  (.A0(\register_file_i/rf_reg_685_ ),
    .A1(net787),
    .S(net937),
    .X(\register_file_i/_0645_ ));
 sg13g2_mux2_1 \register_file_i/_6754_  (.A0(\register_file_i/rf_reg_686_ ),
    .A1(net749),
    .S(net939),
    .X(\register_file_i/_0646_ ));
 sg13g2_mux2_1 \register_file_i/_6755_  (.A0(\register_file_i/rf_reg_687_ ),
    .A1(net781),
    .S(net939),
    .X(\register_file_i/_0647_ ));
 sg13g2_mux2_1 \register_file_i/_6756_  (.A0(\register_file_i/rf_reg_688_ ),
    .A1(net709),
    .S(net939),
    .X(\register_file_i/_0648_ ));
 sg13g2_mux2_1 \register_file_i/_6757_  (.A0(\register_file_i/rf_reg_689_ ),
    .A1(net724),
    .S(net940),
    .X(\register_file_i/_0649_ ));
 sg13g2_mux2_1 \register_file_i/_6758_  (.A0(net1018),
    .A1(\register_file_i/rf_reg_68_ ),
    .S(net810),
    .X(\register_file_i/_0650_ ));
 sg13g2_mux2_1 \register_file_i/_6759_  (.A0(\register_file_i/rf_reg_690_ ),
    .A1(net704),
    .S(net940),
    .X(\register_file_i/_0651_ ));
 sg13g2_mux2_1 \register_file_i/_6760_  (.A0(\register_file_i/rf_reg_691_ ),
    .A1(net699),
    .S(net939),
    .X(\register_file_i/_0652_ ));
 sg13g2_buf_4 fanout41 (.X(net41),
    .A(net43));
 sg13g2_mux2_1 \register_file_i/_6762_  (.A0(\register_file_i/rf_reg_692_ ),
    .A1(net738),
    .S(net940),
    .X(\register_file_i/_0653_ ));
 sg13g2_mux2_1 \register_file_i/_6763_  (.A0(\register_file_i/rf_reg_693_ ),
    .A1(net672),
    .S(net940),
    .X(\register_file_i/_0654_ ));
 sg13g2_mux2_1 \register_file_i/_6764_  (.A0(\register_file_i/rf_reg_694_ ),
    .A1(net693),
    .S(net940),
    .X(\register_file_i/_0655_ ));
 sg13g2_mux2_1 \register_file_i/_6765_  (.A0(\register_file_i/rf_reg_695_ ),
    .A1(net687),
    .S(net939),
    .X(\register_file_i/_0656_ ));
 sg13g2_mux2_1 \register_file_i/_6766_  (.A0(\register_file_i/rf_reg_696_ ),
    .A1(net683),
    .S(net939),
    .X(\register_file_i/_0657_ ));
 sg13g2_mux2_1 \register_file_i/_6767_  (.A0(\register_file_i/rf_reg_697_ ),
    .A1(net600),
    .S(net937),
    .X(\register_file_i/_0658_ ));
 sg13g2_mux2_1 \register_file_i/_6768_  (.A0(\register_file_i/rf_reg_698_ ),
    .A1(net666),
    .S(net936),
    .X(\register_file_i/_0659_ ));
 sg13g2_mux2_1 \register_file_i/_6769_  (.A0(\register_file_i/rf_reg_699_ ),
    .A1(net582),
    .S(net937),
    .X(\register_file_i/_0660_ ));
 sg13g2_mux2_1 \register_file_i/_6770_  (.A0(net998),
    .A1(\register_file_i/rf_reg_69_ ),
    .S(net810),
    .X(\register_file_i/_0661_ ));
 sg13g2_mux2_1 \register_file_i/_6771_  (.A0(\register_file_i/rf_reg_700_ ),
    .A1(net578),
    .S(net938),
    .X(\register_file_i/_0662_ ));
 sg13g2_mux2_1 \register_file_i/_6772_  (.A0(\register_file_i/rf_reg_701_ ),
    .A1(net569),
    .S(net937),
    .X(\register_file_i/_0663_ ));
 sg13g2_mux2_1 \register_file_i/_6773_  (.A0(\register_file_i/rf_reg_702_ ),
    .A1(net574),
    .S(net939),
    .X(\register_file_i/_0664_ ));
 sg13g2_mux2_1 \register_file_i/_6774_  (.A0(\register_file_i/rf_reg_703_ ),
    .A1(net563),
    .S(net939),
    .X(\register_file_i/_0665_ ));
 sg13g2_nor2_1 \register_file_i/_6775_  (.A(\register_file_i/_2868_ ),
    .B(\register_file_i/_2951_ ),
    .Y(\register_file_i/_3003_ ));
 sg13g2_buf_2 fanout40 (.A(\cs_registers_i/_0519_ ),
    .X(net40));
 sg13g2_mux2_1 \register_file_i/_6777_  (.A0(\register_file_i/rf_reg_704_ ),
    .A1(net752),
    .S(net931),
    .X(\register_file_i/_0666_ ));
 sg13g2_mux2_1 \register_file_i/_6778_  (.A0(\register_file_i/rf_reg_705_ ),
    .A1(net1001),
    .S(net931),
    .X(\register_file_i/_0667_ ));
 sg13g2_mux2_1 \register_file_i/_6779_  (.A0(\register_file_i/rf_reg_706_ ),
    .A1(net887),
    .S(net932),
    .X(\register_file_i/_0668_ ));
 sg13g2_mux2_1 \register_file_i/_6780_  (.A0(\register_file_i/rf_reg_707_ ),
    .A1(net1020),
    .S(net932),
    .X(\register_file_i/_0669_ ));
 sg13g2_mux2_1 \register_file_i/_6781_  (.A0(\register_file_i/rf_reg_708_ ),
    .A1(net1016),
    .S(net932),
    .X(\register_file_i/_0670_ ));
 sg13g2_mux2_1 \register_file_i/_6782_  (.A0(\register_file_i/rf_reg_709_ ),
    .A1(net996),
    .S(net930),
    .X(\register_file_i/_0671_ ));
 sg13g2_mux2_1 \register_file_i/_6783_  (.A0(net883),
    .A1(\register_file_i/rf_reg_70_ ),
    .S(net810),
    .X(\register_file_i/_0672_ ));
 sg13g2_mux2_1 \register_file_i/_6784_  (.A0(\register_file_i/rf_reg_710_ ),
    .A1(net881),
    .S(net932),
    .X(\register_file_i/_0673_ ));
 sg13g2_mux2_1 \register_file_i/_6785_  (.A0(\register_file_i/rf_reg_711_ ),
    .A1(net992),
    .S(net932),
    .X(\register_file_i/_0674_ ));
 sg13g2_mux2_1 \register_file_i/_6786_  (.A0(\register_file_i/rf_reg_712_ ),
    .A1(net876),
    .S(net930),
    .X(\register_file_i/_0675_ ));
 sg13g2_mux2_1 \register_file_i/_6787_  (.A0(\register_file_i/rf_reg_713_ ),
    .A1(net805),
    .S(net930),
    .X(\register_file_i/_0676_ ));
 sg13g2_buf_4 fanout39 (.X(net39),
    .A(\cs_registers_i/_1824_ ));
 sg13g2_mux2_1 \register_file_i/_6789_  (.A0(\register_file_i/rf_reg_714_ ),
    .A1(net796),
    .S(net930),
    .X(\register_file_i/_0677_ ));
 sg13g2_mux2_1 \register_file_i/_6790_  (.A0(\register_file_i/rf_reg_715_ ),
    .A1(net791),
    .S(net930),
    .X(\register_file_i/_0678_ ));
 sg13g2_mux2_1 \register_file_i/_6791_  (.A0(\register_file_i/rf_reg_716_ ),
    .A1(net800),
    .S(net930),
    .X(\register_file_i/_0679_ ));
 sg13g2_mux2_1 \register_file_i/_6792_  (.A0(\register_file_i/rf_reg_717_ ),
    .A1(net787),
    .S(net933),
    .X(\register_file_i/_0680_ ));
 sg13g2_mux2_1 \register_file_i/_6793_  (.A0(\register_file_i/rf_reg_718_ ),
    .A1(net749),
    .S(net933),
    .X(\register_file_i/_0681_ ));
 sg13g2_mux2_1 \register_file_i/_6794_  (.A0(\register_file_i/rf_reg_719_ ),
    .A1(net781),
    .S(net933),
    .X(\register_file_i/_0682_ ));
 sg13g2_mux2_1 \register_file_i/_6795_  (.A0(net994),
    .A1(\register_file_i/rf_reg_71_ ),
    .S(net810),
    .X(\register_file_i/_0683_ ));
 sg13g2_mux2_1 \register_file_i/_6796_  (.A0(\register_file_i/rf_reg_720_ ),
    .A1(net709),
    .S(net934),
    .X(\register_file_i/_0684_ ));
 sg13g2_mux2_1 \register_file_i/_6797_  (.A0(\register_file_i/rf_reg_721_ ),
    .A1(net723),
    .S(net934),
    .X(\register_file_i/_0685_ ));
 sg13g2_mux2_1 \register_file_i/_6798_  (.A0(\register_file_i/rf_reg_722_ ),
    .A1(net704),
    .S(net934),
    .X(\register_file_i/_0686_ ));
 sg13g2_mux2_1 \register_file_i/_6799_  (.A0(\register_file_i/rf_reg_723_ ),
    .A1(net699),
    .S(net933),
    .X(\register_file_i/_0687_ ));
 sg13g2_buf_4 fanout38 (.X(net38),
    .A(\cs_registers_i/_1824_ ));
 sg13g2_mux2_1 \register_file_i/_6801_  (.A0(\register_file_i/rf_reg_724_ ),
    .A1(net738),
    .S(net934),
    .X(\register_file_i/_0688_ ));
 sg13g2_mux2_1 \register_file_i/_6802_  (.A0(\register_file_i/rf_reg_725_ ),
    .A1(net672),
    .S(net934),
    .X(\register_file_i/_0689_ ));
 sg13g2_mux2_1 \register_file_i/_6803_  (.A0(\register_file_i/rf_reg_726_ ),
    .A1(net693),
    .S(net935),
    .X(\register_file_i/_0690_ ));
 sg13g2_mux2_1 \register_file_i/_6804_  (.A0(\register_file_i/rf_reg_727_ ),
    .A1(net687),
    .S(net933),
    .X(\register_file_i/_0691_ ));
 sg13g2_mux2_1 \register_file_i/_6805_  (.A0(\register_file_i/rf_reg_728_ ),
    .A1(net683),
    .S(net933),
    .X(\register_file_i/_0692_ ));
 sg13g2_mux2_1 \register_file_i/_6806_  (.A0(\register_file_i/rf_reg_729_ ),
    .A1(net601),
    .S(net931),
    .X(\register_file_i/_0693_ ));
 sg13g2_mux2_1 \register_file_i/_6807_  (.A0(net878),
    .A1(\register_file_i/rf_reg_72_ ),
    .S(net810),
    .X(\register_file_i/_0694_ ));
 sg13g2_mux2_1 \register_file_i/_6808_  (.A0(\register_file_i/rf_reg_730_ ),
    .A1(net666),
    .S(net930),
    .X(\register_file_i/_0695_ ));
 sg13g2_mux2_1 \register_file_i/_6809_  (.A0(\register_file_i/rf_reg_731_ ),
    .A1(net582),
    .S(net930),
    .X(\register_file_i/_0696_ ));
 sg13g2_mux2_1 \register_file_i/_6810_  (.A0(\register_file_i/rf_reg_732_ ),
    .A1(net578),
    .S(net932),
    .X(\register_file_i/_0697_ ));
 sg13g2_mux2_1 \register_file_i/_6811_  (.A0(\register_file_i/rf_reg_733_ ),
    .A1(net569),
    .S(net931),
    .X(\register_file_i/_0698_ ));
 sg13g2_mux2_1 \register_file_i/_6812_  (.A0(\register_file_i/rf_reg_734_ ),
    .A1(net574),
    .S(net933),
    .X(\register_file_i/_0699_ ));
 sg13g2_mux2_1 \register_file_i/_6813_  (.A0(\register_file_i/rf_reg_735_ ),
    .A1(net563),
    .S(net933),
    .X(\register_file_i/_0700_ ));
 sg13g2_nor2_2 \register_file_i/_6814_  (.A(\register_file_i/_2800_ ),
    .B(\register_file_i/_2868_ ),
    .Y(\register_file_i/_3007_ ));
 sg13g2_buf_8 fanout37 (.A(data_addr_o_31_),
    .X(net37));
 sg13g2_mux2_1 \register_file_i/_6816_  (.A0(\register_file_i/rf_reg_736_ ),
    .A1(net753),
    .S(net926),
    .X(\register_file_i/_0701_ ));
 sg13g2_mux2_1 \register_file_i/_6817_  (.A0(\register_file_i/rf_reg_737_ ),
    .A1(net1001),
    .S(net925),
    .X(\register_file_i/_0702_ ));
 sg13g2_mux2_1 \register_file_i/_6818_  (.A0(\register_file_i/rf_reg_738_ ),
    .A1(net885),
    .S(net927),
    .X(\register_file_i/_0703_ ));
 sg13g2_mux2_1 \register_file_i/_6819_  (.A0(\register_file_i/rf_reg_739_ ),
    .A1(net1020),
    .S(net927),
    .X(\register_file_i/_0704_ ));
 sg13g2_mux2_1 \register_file_i/_6820_  (.A0(net807),
    .A1(\register_file_i/rf_reg_73_ ),
    .S(net809),
    .X(\register_file_i/_0705_ ));
 sg13g2_mux2_1 \register_file_i/_6821_  (.A0(\register_file_i/rf_reg_740_ ),
    .A1(net1016),
    .S(net927),
    .X(\register_file_i/_0706_ ));
 sg13g2_mux2_1 \register_file_i/_6822_  (.A0(\register_file_i/rf_reg_741_ ),
    .A1(net996),
    .S(net925),
    .X(\register_file_i/_0707_ ));
 sg13g2_mux2_1 \register_file_i/_6823_  (.A0(\register_file_i/rf_reg_742_ ),
    .A1(net881),
    .S(net927),
    .X(\register_file_i/_0708_ ));
 sg13g2_mux2_1 \register_file_i/_6824_  (.A0(\register_file_i/rf_reg_743_ ),
    .A1(net992),
    .S(net927),
    .X(\register_file_i/_0709_ ));
 sg13g2_mux2_1 \register_file_i/_6825_  (.A0(\register_file_i/rf_reg_744_ ),
    .A1(net876),
    .S(net925),
    .X(\register_file_i/_0710_ ));
 sg13g2_mux2_1 \register_file_i/_6826_  (.A0(\register_file_i/rf_reg_745_ ),
    .A1(net805),
    .S(net925),
    .X(\register_file_i/_0711_ ));
 sg13g2_buf_8 fanout36 (.A(net37),
    .X(net36));
 sg13g2_mux2_1 \register_file_i/_6828_  (.A0(\register_file_i/rf_reg_746_ ),
    .A1(net796),
    .S(net925),
    .X(\register_file_i/_0712_ ));
 sg13g2_mux2_1 \register_file_i/_6829_  (.A0(\register_file_i/rf_reg_747_ ),
    .A1(net791),
    .S(net925),
    .X(\register_file_i/_0713_ ));
 sg13g2_mux2_1 \register_file_i/_6830_  (.A0(\register_file_i/rf_reg_748_ ),
    .A1(net803),
    .S(net925),
    .X(\register_file_i/_0714_ ));
 sg13g2_mux2_1 \register_file_i/_6831_  (.A0(\register_file_i/rf_reg_749_ ),
    .A1(net787),
    .S(net929),
    .X(\register_file_i/_0715_ ));
 sg13g2_buf_2 fanout35 (.A(_05613_),
    .X(net35));
 sg13g2_mux2_1 \register_file_i/_6833_  (.A0(net798),
    .A1(\register_file_i/rf_reg_74_ ),
    .S(net809),
    .X(\register_file_i/_0716_ ));
 sg13g2_mux2_1 \register_file_i/_6834_  (.A0(\register_file_i/rf_reg_750_ ),
    .A1(net749),
    .S(net929),
    .X(\register_file_i/_0717_ ));
 sg13g2_mux2_1 \register_file_i/_6835_  (.A0(\register_file_i/rf_reg_751_ ),
    .A1(net784),
    .S(net929),
    .X(\register_file_i/_0718_ ));
 sg13g2_mux2_1 \register_file_i/_6836_  (.A0(\register_file_i/rf_reg_752_ ),
    .A1(net709),
    .S(net928),
    .X(\register_file_i/_0719_ ));
 sg13g2_mux2_1 \register_file_i/_6837_  (.A0(\register_file_i/rf_reg_753_ ),
    .A1(net727),
    .S(net928),
    .X(\register_file_i/_0720_ ));
 sg13g2_mux2_1 \register_file_i/_6838_  (.A0(\register_file_i/rf_reg_754_ ),
    .A1(net704),
    .S(net928),
    .X(\register_file_i/_0721_ ));
 sg13g2_mux2_1 \register_file_i/_6839_  (.A0(\register_file_i/rf_reg_755_ ),
    .A1(net699),
    .S(net928),
    .X(\register_file_i/_0722_ ));
 sg13g2_buf_8 fanout34 (.A(\cs_registers_i/_1761_ ),
    .X(net34));
 sg13g2_mux2_1 \register_file_i/_6841_  (.A0(\register_file_i/rf_reg_756_ ),
    .A1(net738),
    .S(net929),
    .X(\register_file_i/_0723_ ));
 sg13g2_mux2_1 \register_file_i/_6842_  (.A0(\register_file_i/rf_reg_757_ ),
    .A1(rf_wdata_wb_21_),
    .S(net928),
    .X(\register_file_i/_0724_ ));
 sg13g2_mux2_1 \register_file_i/_6843_  (.A0(\register_file_i/rf_reg_758_ ),
    .A1(net697),
    .S(net928),
    .X(\register_file_i/_0725_ ));
 sg13g2_mux2_1 \register_file_i/_6844_  (.A0(\register_file_i/rf_reg_759_ ),
    .A1(net687),
    .S(net929),
    .X(\register_file_i/_0726_ ));
 sg13g2_mux2_1 \register_file_i/_6845_  (.A0(net793),
    .A1(\register_file_i/rf_reg_75_ ),
    .S(net809),
    .X(\register_file_i/_0727_ ));
 sg13g2_mux2_1 \register_file_i/_6846_  (.A0(\register_file_i/rf_reg_760_ ),
    .A1(net683),
    .S(net929),
    .X(\register_file_i/_0728_ ));
 sg13g2_mux2_1 \register_file_i/_6847_  (.A0(\register_file_i/rf_reg_761_ ),
    .A1(net601),
    .S(net926),
    .X(\register_file_i/_0729_ ));
 sg13g2_mux2_1 \register_file_i/_6848_  (.A0(\register_file_i/rf_reg_762_ ),
    .A1(net666),
    .S(net925),
    .X(\register_file_i/_0730_ ));
 sg13g2_mux2_1 \register_file_i/_6849_  (.A0(\register_file_i/rf_reg_763_ ),
    .A1(net583),
    .S(net926),
    .X(\register_file_i/_0731_ ));
 sg13g2_mux2_1 \register_file_i/_6850_  (.A0(\register_file_i/rf_reg_764_ ),
    .A1(net578),
    .S(net927),
    .X(\register_file_i/_0732_ ));
 sg13g2_mux2_1 \register_file_i/_6851_  (.A0(\register_file_i/rf_reg_765_ ),
    .A1(net569),
    .S(net926),
    .X(\register_file_i/_0733_ ));
 sg13g2_mux2_1 \register_file_i/_6852_  (.A0(\register_file_i/rf_reg_766_ ),
    .A1(net573),
    .S(net928),
    .X(\register_file_i/_0734_ ));
 sg13g2_mux2_1 \register_file_i/_6853_  (.A0(\register_file_i/rf_reg_767_ ),
    .A1(net563),
    .S(net928),
    .X(\register_file_i/_0735_ ));
 sg13g2_nand2b_2 \register_file_i/_6854_  (.Y(\register_file_i/_3012_ ),
    .B(\register_file_i/_2940_ ),
    .A_N(\register_file_i/_2901_ ));
 sg13g2_buf_4 fanout33 (.X(net33),
    .A(net34));
 sg13g2_buf_4 fanout32 (.X(net32),
    .A(net34));
 sg13g2_mux2_1 \register_file_i/_6857_  (.A0(net753),
    .A1(\register_file_i/rf_reg_768_ ),
    .S(net922),
    .X(\register_file_i/_0736_ ));
 sg13g2_mux2_1 \register_file_i/_6858_  (.A0(net1000),
    .A1(\register_file_i/rf_reg_769_ ),
    .S(net921),
    .X(\register_file_i/_0737_ ));
 sg13g2_mux2_1 \register_file_i/_6859_  (.A0(net802),
    .A1(\register_file_i/rf_reg_76_ ),
    .S(net809),
    .X(\register_file_i/_0738_ ));
 sg13g2_mux2_1 \register_file_i/_6860_  (.A0(net884),
    .A1(\register_file_i/rf_reg_770_ ),
    .S(net921),
    .X(\register_file_i/_0739_ ));
 sg13g2_mux2_1 \register_file_i/_6861_  (.A0(net1022),
    .A1(\register_file_i/rf_reg_771_ ),
    .S(net921),
    .X(\register_file_i/_0740_ ));
 sg13g2_mux2_1 \register_file_i/_6862_  (.A0(net1017),
    .A1(\register_file_i/rf_reg_772_ ),
    .S(net920),
    .X(\register_file_i/_0741_ ));
 sg13g2_mux2_1 \register_file_i/_6863_  (.A0(net998),
    .A1(\register_file_i/rf_reg_773_ ),
    .S(net920),
    .X(\register_file_i/_0742_ ));
 sg13g2_mux2_1 \register_file_i/_6864_  (.A0(net882),
    .A1(\register_file_i/rf_reg_774_ ),
    .S(net920),
    .X(\register_file_i/_0743_ ));
 sg13g2_mux2_1 \register_file_i/_6865_  (.A0(net994),
    .A1(\register_file_i/rf_reg_775_ ),
    .S(net920),
    .X(\register_file_i/_0744_ ));
 sg13g2_mux2_1 \register_file_i/_6866_  (.A0(net877),
    .A1(\register_file_i/rf_reg_776_ ),
    .S(net920),
    .X(\register_file_i/_0745_ ));
 sg13g2_mux2_1 \register_file_i/_6867_  (.A0(net806),
    .A1(\register_file_i/rf_reg_777_ ),
    .S(net920),
    .X(\register_file_i/_0746_ ));
 sg13g2_buf_16 fanout31 (.X(net31),
    .A(net34));
 sg13g2_mux2_1 \register_file_i/_6869_  (.A0(net797),
    .A1(\register_file_i/rf_reg_778_ ),
    .S(net920),
    .X(\register_file_i/_0747_ ));
 sg13g2_mux2_1 \register_file_i/_6870_  (.A0(net792),
    .A1(\register_file_i/rf_reg_779_ ),
    .S(net920),
    .X(\register_file_i/_0748_ ));
 sg13g2_mux2_1 \register_file_i/_6871_  (.A0(net789),
    .A1(\register_file_i/rf_reg_77_ ),
    .S(net812),
    .X(\register_file_i/_0749_ ));
 sg13g2_mux2_1 \register_file_i/_6872_  (.A0(net801),
    .A1(\register_file_i/rf_reg_780_ ),
    .S(net921),
    .X(\register_file_i/_0750_ ));
 sg13g2_mux2_1 \register_file_i/_6873_  (.A0(net788),
    .A1(\register_file_i/rf_reg_781_ ),
    .S(net922),
    .X(\register_file_i/_0751_ ));
 sg13g2_mux2_1 \register_file_i/_6874_  (.A0(net750),
    .A1(\register_file_i/rf_reg_782_ ),
    .S(net922),
    .X(\register_file_i/_0752_ ));
 sg13g2_mux2_1 \register_file_i/_6875_  (.A0(net782),
    .A1(\register_file_i/rf_reg_783_ ),
    .S(net922),
    .X(\register_file_i/_0753_ ));
 sg13g2_mux2_1 \register_file_i/_6876_  (.A0(net711),
    .A1(\register_file_i/rf_reg_784_ ),
    .S(net922),
    .X(\register_file_i/_0754_ ));
 sg13g2_mux2_1 \register_file_i/_6877_  (.A0(net725),
    .A1(\register_file_i/rf_reg_785_ ),
    .S(net923),
    .X(\register_file_i/_0755_ ));
 sg13g2_mux2_1 \register_file_i/_6878_  (.A0(net705),
    .A1(\register_file_i/rf_reg_786_ ),
    .S(net922),
    .X(\register_file_i/_0756_ ));
 sg13g2_mux2_1 \register_file_i/_6879_  (.A0(net700),
    .A1(\register_file_i/rf_reg_787_ ),
    .S(net923),
    .X(\register_file_i/_0757_ ));
 sg13g2_buf_16 fanout30 (.X(net30),
    .A(net34));
 sg13g2_mux2_1 \register_file_i/_6881_  (.A0(net739),
    .A1(\register_file_i/rf_reg_788_ ),
    .S(net923),
    .X(\register_file_i/_0758_ ));
 sg13g2_mux2_1 \register_file_i/_6882_  (.A0(net674),
    .A1(\register_file_i/rf_reg_789_ ),
    .S(net923),
    .X(\register_file_i/_0759_ ));
 sg13g2_mux2_1 \register_file_i/_6883_  (.A0(net751),
    .A1(\register_file_i/rf_reg_78_ ),
    .S(net812),
    .X(\register_file_i/_0760_ ));
 sg13g2_mux2_1 \register_file_i/_6884_  (.A0(net695),
    .A1(\register_file_i/rf_reg_790_ ),
    .S(net924),
    .X(\register_file_i/_0761_ ));
 sg13g2_mux2_1 \register_file_i/_6885_  (.A0(net687),
    .A1(\register_file_i/rf_reg_791_ ),
    .S(net921),
    .X(\register_file_i/_0762_ ));
 sg13g2_mux2_1 \register_file_i/_6886_  (.A0(net685),
    .A1(\register_file_i/rf_reg_792_ ),
    .S(net924),
    .X(\register_file_i/_0763_ ));
 sg13g2_mux2_1 \register_file_i/_6887_  (.A0(net602),
    .A1(\register_file_i/rf_reg_793_ ),
    .S(net924),
    .X(\register_file_i/_0764_ ));
 sg13g2_mux2_1 \register_file_i/_6888_  (.A0(net669),
    .A1(\register_file_i/rf_reg_794_ ),
    .S(net924),
    .X(\register_file_i/_0765_ ));
 sg13g2_mux2_1 \register_file_i/_6889_  (.A0(net584),
    .A1(\register_file_i/rf_reg_795_ ),
    .S(net921),
    .X(\register_file_i/_0766_ ));
 sg13g2_mux2_1 \register_file_i/_6890_  (.A0(net580),
    .A1(\register_file_i/rf_reg_796_ ),
    .S(net921),
    .X(\register_file_i/_0767_ ));
 sg13g2_mux2_1 \register_file_i/_6891_  (.A0(net570),
    .A1(\register_file_i/rf_reg_797_ ),
    .S(\register_file_i/_3012_ ),
    .X(\register_file_i/_0768_ ));
 sg13g2_mux2_1 \register_file_i/_6892_  (.A0(net574),
    .A1(\register_file_i/rf_reg_798_ ),
    .S(net922),
    .X(\register_file_i/_0769_ ));
 sg13g2_mux2_1 \register_file_i/_6893_  (.A0(net564),
    .A1(\register_file_i/rf_reg_799_ ),
    .S(net922),
    .X(\register_file_i/_0770_ ));
 sg13g2_mux2_1 \register_file_i/_6894_  (.A0(net783),
    .A1(\register_file_i/rf_reg_79_ ),
    .S(net812),
    .X(\register_file_i/_0771_ ));
 sg13g2_nor2_2 \register_file_i/_6895_  (.A(\register_file_i/_2901_ ),
    .B(\register_file_i/_2946_ ),
    .Y(\register_file_i/_3017_ ));
 sg13g2_buf_8 fanout29 (.A(\cs_registers_i/_1771_ ),
    .X(net29));
 sg13g2_mux2_1 \register_file_i/_6897_  (.A0(\register_file_i/rf_reg_800_ ),
    .A1(net753),
    .S(net917),
    .X(\register_file_i/_0772_ ));
 sg13g2_mux2_1 \register_file_i/_6898_  (.A0(\register_file_i/rf_reg_801_ ),
    .A1(net1001),
    .S(net916),
    .X(\register_file_i/_0773_ ));
 sg13g2_mux2_1 \register_file_i/_6899_  (.A0(\register_file_i/rf_reg_802_ ),
    .A1(rf_wdata_wb_2_),
    .S(net916),
    .X(\register_file_i/_0774_ ));
 sg13g2_mux2_1 \register_file_i/_6900_  (.A0(\register_file_i/rf_reg_803_ ),
    .A1(net1022),
    .S(net916),
    .X(\register_file_i/_0775_ ));
 sg13g2_mux2_1 \register_file_i/_6901_  (.A0(\register_file_i/rf_reg_804_ ),
    .A1(net1017),
    .S(net914),
    .X(\register_file_i/_0776_ ));
 sg13g2_mux2_1 \register_file_i/_6902_  (.A0(\register_file_i/rf_reg_805_ ),
    .A1(net997),
    .S(net914),
    .X(\register_file_i/_0777_ ));
 sg13g2_mux2_1 \register_file_i/_6903_  (.A0(\register_file_i/rf_reg_806_ ),
    .A1(net882),
    .S(net914),
    .X(\register_file_i/_0778_ ));
 sg13g2_mux2_1 \register_file_i/_6904_  (.A0(\register_file_i/rf_reg_807_ ),
    .A1(net994),
    .S(net914),
    .X(\register_file_i/_0779_ ));
 sg13g2_mux2_1 \register_file_i/_6905_  (.A0(\register_file_i/rf_reg_808_ ),
    .A1(net877),
    .S(net914),
    .X(\register_file_i/_0780_ ));
 sg13g2_mux2_1 \register_file_i/_6906_  (.A0(\register_file_i/rf_reg_809_ ),
    .A1(net807),
    .S(net914),
    .X(\register_file_i/_0781_ ));
 sg13g2_mux2_1 \register_file_i/_6907_  (.A0(net710),
    .A1(\register_file_i/rf_reg_80_ ),
    .S(net813),
    .X(\register_file_i/_0782_ ));
 sg13g2_buf_8 fanout28 (.A(\cs_registers_i/_1771_ ),
    .X(net28));
 sg13g2_mux2_1 \register_file_i/_6909_  (.A0(\register_file_i/rf_reg_810_ ),
    .A1(net798),
    .S(net914),
    .X(\register_file_i/_0783_ ));
 sg13g2_mux2_1 \register_file_i/_6910_  (.A0(\register_file_i/rf_reg_811_ ),
    .A1(net792),
    .S(net915),
    .X(\register_file_i/_0784_ ));
 sg13g2_mux2_1 \register_file_i/_6911_  (.A0(\register_file_i/rf_reg_812_ ),
    .A1(net801),
    .S(net914),
    .X(\register_file_i/_0785_ ));
 sg13g2_mux2_1 \register_file_i/_6912_  (.A0(\register_file_i/rf_reg_813_ ),
    .A1(net788),
    .S(net917),
    .X(\register_file_i/_0786_ ));
 sg13g2_mux2_1 \register_file_i/_6913_  (.A0(\register_file_i/rf_reg_814_ ),
    .A1(net750),
    .S(net917),
    .X(\register_file_i/_0787_ ));
 sg13g2_mux2_1 \register_file_i/_6914_  (.A0(\register_file_i/rf_reg_815_ ),
    .A1(net782),
    .S(net917),
    .X(\register_file_i/_0788_ ));
 sg13g2_mux2_1 \register_file_i/_6915_  (.A0(\register_file_i/rf_reg_816_ ),
    .A1(net711),
    .S(net917),
    .X(\register_file_i/_0789_ ));
 sg13g2_mux2_1 \register_file_i/_6916_  (.A0(\register_file_i/rf_reg_817_ ),
    .A1(net725),
    .S(net918),
    .X(\register_file_i/_0790_ ));
 sg13g2_mux2_1 \register_file_i/_6917_  (.A0(\register_file_i/rf_reg_818_ ),
    .A1(net705),
    .S(net917),
    .X(\register_file_i/_0791_ ));
 sg13g2_mux2_1 \register_file_i/_6918_  (.A0(\register_file_i/rf_reg_819_ ),
    .A1(net700),
    .S(net918),
    .X(\register_file_i/_0792_ ));
 sg13g2_mux2_1 \register_file_i/_6919_  (.A0(net726),
    .A1(\register_file_i/rf_reg_81_ ),
    .S(net812),
    .X(\register_file_i/_0793_ ));
 sg13g2_buf_8 fanout27 (.A(\cs_registers_i/_1771_ ),
    .X(net27));
 sg13g2_mux2_1 \register_file_i/_6921_  (.A0(\register_file_i/rf_reg_820_ ),
    .A1(net740),
    .S(net918),
    .X(\register_file_i/_0794_ ));
 sg13g2_mux2_1 \register_file_i/_6922_  (.A0(\register_file_i/rf_reg_821_ ),
    .A1(net675),
    .S(net918),
    .X(\register_file_i/_0795_ ));
 sg13g2_mux2_1 \register_file_i/_6923_  (.A0(\register_file_i/rf_reg_822_ ),
    .A1(net695),
    .S(net919),
    .X(\register_file_i/_0796_ ));
 sg13g2_mux2_1 \register_file_i/_6924_  (.A0(\register_file_i/rf_reg_823_ ),
    .A1(net688),
    .S(net916),
    .X(\register_file_i/_0797_ ));
 sg13g2_mux2_1 \register_file_i/_6925_  (.A0(\register_file_i/rf_reg_824_ ),
    .A1(net686),
    .S(net919),
    .X(\register_file_i/_0798_ ));
 sg13g2_mux2_1 \register_file_i/_6926_  (.A0(\register_file_i/rf_reg_825_ ),
    .A1(net603),
    .S(net919),
    .X(\register_file_i/_0799_ ));
 sg13g2_mux2_1 \register_file_i/_6927_  (.A0(\register_file_i/rf_reg_826_ ),
    .A1(net669),
    .S(net915),
    .X(\register_file_i/_0800_ ));
 sg13g2_mux2_1 \register_file_i/_6928_  (.A0(\register_file_i/rf_reg_827_ ),
    .A1(net584),
    .S(net915),
    .X(\register_file_i/_0801_ ));
 sg13g2_mux2_1 \register_file_i/_6929_  (.A0(\register_file_i/rf_reg_828_ ),
    .A1(net580),
    .S(net915),
    .X(\register_file_i/_0802_ ));
 sg13g2_mux2_1 \register_file_i/_6930_  (.A0(\register_file_i/rf_reg_829_ ),
    .A1(net571),
    .S(net915),
    .X(\register_file_i/_0803_ ));
 sg13g2_mux2_1 \register_file_i/_6931_  (.A0(net706),
    .A1(\register_file_i/rf_reg_82_ ),
    .S(net812),
    .X(\register_file_i/_0804_ ));
 sg13g2_mux2_1 \register_file_i/_6932_  (.A0(\register_file_i/rf_reg_830_ ),
    .A1(net575),
    .S(net917),
    .X(\register_file_i/_0805_ ));
 sg13g2_mux2_1 \register_file_i/_6933_  (.A0(\register_file_i/rf_reg_831_ ),
    .A1(net564),
    .S(net917),
    .X(\register_file_i/_0806_ ));
 sg13g2_nor2_2 \register_file_i/_6934_  (.A(\register_file_i/_2901_ ),
    .B(\register_file_i/_2951_ ),
    .Y(\register_file_i/_3021_ ));
 sg13g2_buf_8 fanout26 (.A(\cs_registers_i/_1771_ ),
    .X(net26));
 sg13g2_mux2_1 \register_file_i/_6936_  (.A0(\register_file_i/rf_reg_832_ ),
    .A1(net754),
    .S(net911),
    .X(\register_file_i/_0807_ ));
 sg13g2_mux2_1 \register_file_i/_6937_  (.A0(\register_file_i/rf_reg_833_ ),
    .A1(net1004),
    .S(net910),
    .X(\register_file_i/_0808_ ));
 sg13g2_mux2_1 \register_file_i/_6938_  (.A0(\register_file_i/rf_reg_834_ ),
    .A1(net884),
    .S(net910),
    .X(\register_file_i/_0809_ ));
 sg13g2_mux2_1 \register_file_i/_6939_  (.A0(\register_file_i/rf_reg_835_ ),
    .A1(net1022),
    .S(net910),
    .X(\register_file_i/_0810_ ));
 sg13g2_mux2_1 \register_file_i/_6940_  (.A0(\register_file_i/rf_reg_836_ ),
    .A1(net1017),
    .S(net909),
    .X(\register_file_i/_0811_ ));
 sg13g2_mux2_1 \register_file_i/_6941_  (.A0(\register_file_i/rf_reg_837_ ),
    .A1(net997),
    .S(net909),
    .X(\register_file_i/_0812_ ));
 sg13g2_mux2_1 \register_file_i/_6942_  (.A0(\register_file_i/rf_reg_838_ ),
    .A1(net882),
    .S(net909),
    .X(\register_file_i/_0813_ ));
 sg13g2_mux2_1 \register_file_i/_6943_  (.A0(\register_file_i/rf_reg_839_ ),
    .A1(net993),
    .S(net909),
    .X(\register_file_i/_0814_ ));
 sg13g2_mux2_1 \register_file_i/_6944_  (.A0(net701),
    .A1(\register_file_i/rf_reg_83_ ),
    .S(net812),
    .X(\register_file_i/_0815_ ));
 sg13g2_mux2_1 \register_file_i/_6945_  (.A0(\register_file_i/rf_reg_840_ ),
    .A1(net877),
    .S(net909),
    .X(\register_file_i/_0816_ ));
 sg13g2_mux2_1 \register_file_i/_6946_  (.A0(\register_file_i/rf_reg_841_ ),
    .A1(net807),
    .S(net909),
    .X(\register_file_i/_0817_ ));
 sg13g2_buf_8 fanout25 (.A(\cs_registers_i/_1771_ ),
    .X(net25));
 sg13g2_mux2_1 \register_file_i/_6948_  (.A0(\register_file_i/rf_reg_842_ ),
    .A1(net797),
    .S(net909),
    .X(\register_file_i/_0818_ ));
 sg13g2_mux2_1 \register_file_i/_6949_  (.A0(\register_file_i/rf_reg_843_ ),
    .A1(net792),
    .S(net909),
    .X(\register_file_i/_0819_ ));
 sg13g2_mux2_1 \register_file_i/_6950_  (.A0(\register_file_i/rf_reg_844_ ),
    .A1(net801),
    .S(net910),
    .X(\register_file_i/_0820_ ));
 sg13g2_mux2_1 \register_file_i/_6951_  (.A0(\register_file_i/rf_reg_845_ ),
    .A1(net788),
    .S(net911),
    .X(\register_file_i/_0821_ ));
 sg13g2_mux2_1 \register_file_i/_6952_  (.A0(\register_file_i/rf_reg_846_ ),
    .A1(net750),
    .S(net911),
    .X(\register_file_i/_0822_ ));
 sg13g2_mux2_1 \register_file_i/_6953_  (.A0(\register_file_i/rf_reg_847_ ),
    .A1(net782),
    .S(net911),
    .X(\register_file_i/_0823_ ));
 sg13g2_mux2_1 \register_file_i/_6954_  (.A0(\register_file_i/rf_reg_848_ ),
    .A1(net711),
    .S(net912),
    .X(\register_file_i/_0824_ ));
 sg13g2_mux2_1 \register_file_i/_6955_  (.A0(\register_file_i/rf_reg_849_ ),
    .A1(net725),
    .S(net912),
    .X(\register_file_i/_0825_ ));
 sg13g2_buf_2 fanout24 (.A(\cs_registers_i/_2067_ ),
    .X(net24));
 sg13g2_mux2_1 \register_file_i/_6957_  (.A0(net740),
    .A1(\register_file_i/rf_reg_84_ ),
    .S(net813),
    .X(\register_file_i/_0826_ ));
 sg13g2_mux2_1 \register_file_i/_6958_  (.A0(\register_file_i/rf_reg_850_ ),
    .A1(net705),
    .S(net912),
    .X(\register_file_i/_0827_ ));
 sg13g2_mux2_1 \register_file_i/_6959_  (.A0(\register_file_i/rf_reg_851_ ),
    .A1(net700),
    .S(net911),
    .X(\register_file_i/_0828_ ));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(net24));
 sg13g2_mux2_1 \register_file_i/_6961_  (.A0(\register_file_i/rf_reg_852_ ),
    .A1(net739),
    .S(net912),
    .X(\register_file_i/_0829_ ));
 sg13g2_mux2_1 \register_file_i/_6962_  (.A0(\register_file_i/rf_reg_853_ ),
    .A1(net673),
    .S(net912),
    .X(\register_file_i/_0830_ ));
 sg13g2_mux2_1 \register_file_i/_6963_  (.A0(\register_file_i/rf_reg_854_ ),
    .A1(net696),
    .S(net913),
    .X(\register_file_i/_0831_ ));
 sg13g2_mux2_1 \register_file_i/_6964_  (.A0(\register_file_i/rf_reg_855_ ),
    .A1(net688),
    .S(net911),
    .X(\register_file_i/_0832_ ));
 sg13g2_mux2_1 \register_file_i/_6965_  (.A0(\register_file_i/rf_reg_856_ ),
    .A1(net685),
    .S(net913),
    .X(\register_file_i/_0833_ ));
 sg13g2_mux2_1 \register_file_i/_6966_  (.A0(\register_file_i/rf_reg_857_ ),
    .A1(net603),
    .S(net913),
    .X(\register_file_i/_0834_ ));
 sg13g2_mux2_1 \register_file_i/_6967_  (.A0(\register_file_i/rf_reg_858_ ),
    .A1(net668),
    .S(net913),
    .X(\register_file_i/_0835_ ));
 sg13g2_mux2_1 \register_file_i/_6968_  (.A0(\register_file_i/rf_reg_859_ ),
    .A1(net584),
    .S(net910),
    .X(\register_file_i/_0836_ ));
 sg13g2_mux2_1 \register_file_i/_6969_  (.A0(net673),
    .A1(\register_file_i/rf_reg_85_ ),
    .S(net813),
    .X(\register_file_i/_0837_ ));
 sg13g2_mux2_1 \register_file_i/_6970_  (.A0(\register_file_i/rf_reg_860_ ),
    .A1(net580),
    .S(net910),
    .X(\register_file_i/_0838_ ));
 sg13g2_mux2_1 \register_file_i/_6971_  (.A0(\register_file_i/rf_reg_861_ ),
    .A1(net571),
    .S(net910),
    .X(\register_file_i/_0839_ ));
 sg13g2_mux2_1 \register_file_i/_6972_  (.A0(\register_file_i/rf_reg_862_ ),
    .A1(net573),
    .S(net911),
    .X(\register_file_i/_0840_ ));
 sg13g2_mux2_1 \register_file_i/_6973_  (.A0(\register_file_i/rf_reg_863_ ),
    .A1(net564),
    .S(net911),
    .X(\register_file_i/_0841_ ));
 sg13g2_nor2_2 \register_file_i/_6974_  (.A(\register_file_i/_2800_ ),
    .B(\register_file_i/_2901_ ),
    .Y(\register_file_i/_3026_ ));
 sg13g2_buf_8 fanout22 (.A(net24),
    .X(net22));
 sg13g2_mux2_1 \register_file_i/_6976_  (.A0(\register_file_i/rf_reg_864_ ),
    .A1(net754),
    .S(net907),
    .X(\register_file_i/_0842_ ));
 sg13g2_mux2_1 \register_file_i/_6977_  (.A0(\register_file_i/rf_reg_865_ ),
    .A1(net1004),
    .S(net905),
    .X(\register_file_i/_0843_ ));
 sg13g2_mux2_1 \register_file_i/_6978_  (.A0(\register_file_i/rf_reg_866_ ),
    .A1(net884),
    .S(net905),
    .X(\register_file_i/_0844_ ));
 sg13g2_mux2_1 \register_file_i/_6979_  (.A0(\register_file_i/rf_reg_867_ ),
    .A1(net1022),
    .S(net905),
    .X(\register_file_i/_0845_ ));
 sg13g2_mux2_1 \register_file_i/_6980_  (.A0(\register_file_i/rf_reg_868_ ),
    .A1(net1017),
    .S(net904),
    .X(\register_file_i/_0846_ ));
 sg13g2_mux2_1 \register_file_i/_6981_  (.A0(\register_file_i/rf_reg_869_ ),
    .A1(net997),
    .S(net904),
    .X(\register_file_i/_0847_ ));
 sg13g2_mux2_1 \register_file_i/_6982_  (.A0(net695),
    .A1(\register_file_i/rf_reg_86_ ),
    .S(net812),
    .X(\register_file_i/_0848_ ));
 sg13g2_mux2_1 \register_file_i/_6983_  (.A0(\register_file_i/rf_reg_870_ ),
    .A1(net882),
    .S(net904),
    .X(\register_file_i/_0849_ ));
 sg13g2_mux2_1 \register_file_i/_6984_  (.A0(\register_file_i/rf_reg_871_ ),
    .A1(net993),
    .S(net904),
    .X(\register_file_i/_0850_ ));
 sg13g2_mux2_1 \register_file_i/_6985_  (.A0(\register_file_i/rf_reg_872_ ),
    .A1(net877),
    .S(net904),
    .X(\register_file_i/_0851_ ));
 sg13g2_mux2_1 \register_file_i/_6986_  (.A0(\register_file_i/rf_reg_873_ ),
    .A1(net806),
    .S(net904),
    .X(\register_file_i/_0852_ ));
 sg13g2_buf_8 fanout21 (.A(net24),
    .X(net21));
 sg13g2_mux2_1 \register_file_i/_6988_  (.A0(\register_file_i/rf_reg_874_ ),
    .A1(net797),
    .S(net904),
    .X(\register_file_i/_0853_ ));
 sg13g2_mux2_1 \register_file_i/_6989_  (.A0(\register_file_i/rf_reg_875_ ),
    .A1(net792),
    .S(net904),
    .X(\register_file_i/_0854_ ));
 sg13g2_mux2_1 \register_file_i/_6990_  (.A0(\register_file_i/rf_reg_876_ ),
    .A1(net801),
    .S(net905),
    .X(\register_file_i/_0855_ ));
 sg13g2_mux2_1 \register_file_i/_6991_  (.A0(\register_file_i/rf_reg_877_ ),
    .A1(net788),
    .S(net907),
    .X(\register_file_i/_0856_ ));
 sg13g2_mux2_1 \register_file_i/_6992_  (.A0(\register_file_i/rf_reg_878_ ),
    .A1(net750),
    .S(net906),
    .X(\register_file_i/_0857_ ));
 sg13g2_mux2_1 \register_file_i/_6993_  (.A0(\register_file_i/rf_reg_879_ ),
    .A1(net782),
    .S(net907),
    .X(\register_file_i/_0858_ ));
 sg13g2_mux2_1 \register_file_i/_6994_  (.A0(net692),
    .A1(\register_file_i/rf_reg_87_ ),
    .S(net811),
    .X(\register_file_i/_0859_ ));
 sg13g2_mux2_1 \register_file_i/_6995_  (.A0(\register_file_i/rf_reg_880_ ),
    .A1(net710),
    .S(net906),
    .X(\register_file_i/_0860_ ));
 sg13g2_mux2_1 \register_file_i/_6996_  (.A0(\register_file_i/rf_reg_881_ ),
    .A1(net725),
    .S(net906),
    .X(\register_file_i/_0861_ ));
 sg13g2_mux2_1 \register_file_i/_6997_  (.A0(\register_file_i/rf_reg_882_ ),
    .A1(net705),
    .S(net906),
    .X(\register_file_i/_0862_ ));
 sg13g2_mux2_1 \register_file_i/_6998_  (.A0(\register_file_i/rf_reg_883_ ),
    .A1(net700),
    .S(net906),
    .X(\register_file_i/_0863_ ));
 sg13g2_buf_2 fanout20 (.A(net24),
    .X(net20));
 sg13g2_mux2_1 \register_file_i/_7000_  (.A0(\register_file_i/rf_reg_884_ ),
    .A1(net739),
    .S(net907),
    .X(\register_file_i/_0864_ ));
 sg13g2_mux2_1 \register_file_i/_7001_  (.A0(\register_file_i/rf_reg_885_ ),
    .A1(net675),
    .S(net906),
    .X(\register_file_i/_0865_ ));
 sg13g2_mux2_1 \register_file_i/_7002_  (.A0(\register_file_i/rf_reg_886_ ),
    .A1(net696),
    .S(net908),
    .X(\register_file_i/_0866_ ));
 sg13g2_mux2_1 \register_file_i/_7003_  (.A0(\register_file_i/rf_reg_887_ ),
    .A1(net688),
    .S(net905),
    .X(\register_file_i/_0867_ ));
 sg13g2_mux2_1 \register_file_i/_7004_  (.A0(\register_file_i/rf_reg_888_ ),
    .A1(net685),
    .S(net908),
    .X(\register_file_i/_0868_ ));
 sg13g2_mux2_1 \register_file_i/_7005_  (.A0(\register_file_i/rf_reg_889_ ),
    .A1(net603),
    .S(net908),
    .X(\register_file_i/_0869_ ));
 sg13g2_mux2_1 \register_file_i/_7006_  (.A0(net685),
    .A1(\register_file_i/rf_reg_88_ ),
    .S(net813),
    .X(\register_file_i/_0870_ ));
 sg13g2_mux2_1 \register_file_i/_7007_  (.A0(\register_file_i/rf_reg_890_ ),
    .A1(net668),
    .S(net908),
    .X(\register_file_i/_0871_ ));
 sg13g2_mux2_1 \register_file_i/_7008_  (.A0(\register_file_i/rf_reg_891_ ),
    .A1(net584),
    .S(net905),
    .X(\register_file_i/_0872_ ));
 sg13g2_mux2_1 \register_file_i/_7009_  (.A0(\register_file_i/rf_reg_892_ ),
    .A1(net580),
    .S(net905),
    .X(\register_file_i/_0873_ ));
 sg13g2_mux2_1 \register_file_i/_7010_  (.A0(\register_file_i/rf_reg_893_ ),
    .A1(net571),
    .S(\register_file_i/_3026_ ),
    .X(\register_file_i/_0874_ ));
 sg13g2_mux2_1 \register_file_i/_7011_  (.A0(\register_file_i/rf_reg_894_ ),
    .A1(net573),
    .S(net906),
    .X(\register_file_i/_0875_ ));
 sg13g2_mux2_1 \register_file_i/_7012_  (.A0(\register_file_i/rf_reg_895_ ),
    .A1(net564),
    .S(net906),
    .X(\register_file_i/_0876_ ));
 sg13g2_nor2b_2 \register_file_i/_7013_  (.A(\register_file_i/_2799_ ),
    .B_N(\register_file_i/_2940_ ),
    .Y(\register_file_i/_3030_ ));
 sg13g2_buf_8 fanout19 (.A(net24),
    .X(net19));
 sg13g2_mux2_1 \register_file_i/_7015_  (.A0(\register_file_i/rf_reg_896_ ),
    .A1(net753),
    .S(net901),
    .X(\register_file_i/_0877_ ));
 sg13g2_mux2_1 \register_file_i/_7016_  (.A0(\register_file_i/rf_reg_897_ ),
    .A1(net1000),
    .S(net901),
    .X(\register_file_i/_0878_ ));
 sg13g2_mux2_1 \register_file_i/_7017_  (.A0(\register_file_i/rf_reg_898_ ),
    .A1(net884),
    .S(net901),
    .X(\register_file_i/_0879_ ));
 sg13g2_mux2_1 \register_file_i/_7018_  (.A0(\register_file_i/rf_reg_899_ ),
    .A1(net1020),
    .S(net901),
    .X(\register_file_i/_0880_ ));
 sg13g2_mux2_1 \register_file_i/_7019_  (.A0(net602),
    .A1(\register_file_i/rf_reg_89_ ),
    .S(net811),
    .X(\register_file_i/_0881_ ));
 sg13g2_mux2_1 \register_file_i/_7020_  (.A0(\register_file_i/rf_reg_900_ ),
    .A1(net1017),
    .S(net899),
    .X(\register_file_i/_0882_ ));
 sg13g2_mux2_1 \register_file_i/_7021_  (.A0(\register_file_i/rf_reg_901_ ),
    .A1(net997),
    .S(net899),
    .X(\register_file_i/_0883_ ));
 sg13g2_mux2_1 \register_file_i/_7022_  (.A0(\register_file_i/rf_reg_902_ ),
    .A1(net883),
    .S(net899),
    .X(\register_file_i/_0884_ ));
 sg13g2_mux2_1 \register_file_i/_7023_  (.A0(\register_file_i/rf_reg_903_ ),
    .A1(net993),
    .S(net899),
    .X(\register_file_i/_0885_ ));
 sg13g2_mux2_1 \register_file_i/_7024_  (.A0(\register_file_i/rf_reg_904_ ),
    .A1(net877),
    .S(net899),
    .X(\register_file_i/_0886_ ));
 sg13g2_mux2_1 \register_file_i/_7025_  (.A0(\register_file_i/rf_reg_905_ ),
    .A1(net806),
    .S(net899),
    .X(\register_file_i/_0887_ ));
 sg13g2_buf_8 fanout18 (.A(\cs_registers_i/_1769_ ),
    .X(net18));
 sg13g2_mux2_1 \register_file_i/_7027_  (.A0(\register_file_i/rf_reg_906_ ),
    .A1(net797),
    .S(net899),
    .X(\register_file_i/_0888_ ));
 sg13g2_mux2_1 \register_file_i/_7028_  (.A0(\register_file_i/rf_reg_907_ ),
    .A1(net792),
    .S(net899),
    .X(\register_file_i/_0889_ ));
 sg13g2_mux2_1 \register_file_i/_7029_  (.A0(\register_file_i/rf_reg_908_ ),
    .A1(net801),
    .S(net901),
    .X(\register_file_i/_0890_ ));
 sg13g2_mux2_1 \register_file_i/_7030_  (.A0(\register_file_i/rf_reg_909_ ),
    .A1(net788),
    .S(net902),
    .X(\register_file_i/_0891_ ));
 sg13g2_mux2_1 \register_file_i/_7031_  (.A0(net667),
    .A1(\register_file_i/rf_reg_90_ ),
    .S(net811),
    .X(\register_file_i/_0892_ ));
 sg13g2_mux2_1 \register_file_i/_7032_  (.A0(\register_file_i/rf_reg_910_ ),
    .A1(net750),
    .S(net902),
    .X(\register_file_i/_0893_ ));
 sg13g2_mux2_1 \register_file_i/_7033_  (.A0(\register_file_i/rf_reg_911_ ),
    .A1(net782),
    .S(net902),
    .X(\register_file_i/_0894_ ));
 sg13g2_mux2_1 \register_file_i/_7034_  (.A0(\register_file_i/rf_reg_912_ ),
    .A1(net711),
    .S(net902),
    .X(\register_file_i/_0895_ ));
 sg13g2_mux2_1 \register_file_i/_7035_  (.A0(\register_file_i/rf_reg_913_ ),
    .A1(net725),
    .S(net903),
    .X(\register_file_i/_0896_ ));
 sg13g2_mux2_1 \register_file_i/_7036_  (.A0(\register_file_i/rf_reg_914_ ),
    .A1(net705),
    .S(net902),
    .X(\register_file_i/_0897_ ));
 sg13g2_mux2_1 \register_file_i/_7037_  (.A0(\register_file_i/rf_reg_915_ ),
    .A1(net700),
    .S(net902),
    .X(\register_file_i/_0898_ ));
 sg13g2_buf_16 fanout17 (.X(net17),
    .A(net18));
 sg13g2_mux2_1 \register_file_i/_7039_  (.A0(\register_file_i/rf_reg_916_ ),
    .A1(net739),
    .S(net903),
    .X(\register_file_i/_0899_ ));
 sg13g2_mux2_1 \register_file_i/_7040_  (.A0(\register_file_i/rf_reg_917_ ),
    .A1(net674),
    .S(net903),
    .X(\register_file_i/_0900_ ));
 sg13g2_mux2_1 \register_file_i/_7041_  (.A0(\register_file_i/rf_reg_918_ ),
    .A1(net696),
    .S(net903),
    .X(\register_file_i/_0901_ ));
 sg13g2_mux2_1 \register_file_i/_7042_  (.A0(\register_file_i/rf_reg_919_ ),
    .A1(net688),
    .S(net901),
    .X(\register_file_i/_0902_ ));
 sg13g2_mux2_1 \register_file_i/_7043_  (.A0(net585),
    .A1(\register_file_i/rf_reg_91_ ),
    .S(net810),
    .X(\register_file_i/_0903_ ));
 sg13g2_mux2_1 \register_file_i/_7044_  (.A0(\register_file_i/rf_reg_920_ ),
    .A1(net685),
    .S(net903),
    .X(\register_file_i/_0904_ ));
 sg13g2_mux2_1 \register_file_i/_7045_  (.A0(\register_file_i/rf_reg_921_ ),
    .A1(net603),
    .S(net903),
    .X(\register_file_i/_0905_ ));
 sg13g2_mux2_1 \register_file_i/_7046_  (.A0(\register_file_i/rf_reg_922_ ),
    .A1(net668),
    .S(net900),
    .X(\register_file_i/_0906_ ));
 sg13g2_mux2_1 \register_file_i/_7047_  (.A0(\register_file_i/rf_reg_923_ ),
    .A1(net584),
    .S(net900),
    .X(\register_file_i/_0907_ ));
 sg13g2_mux2_1 \register_file_i/_7048_  (.A0(\register_file_i/rf_reg_924_ ),
    .A1(net580),
    .S(net900),
    .X(\register_file_i/_0908_ ));
 sg13g2_mux2_1 \register_file_i/_7049_  (.A0(\register_file_i/rf_reg_925_ ),
    .A1(net571),
    .S(net900),
    .X(\register_file_i/_0909_ ));
 sg13g2_mux2_1 \register_file_i/_7050_  (.A0(\register_file_i/rf_reg_926_ ),
    .A1(net574),
    .S(net902),
    .X(\register_file_i/_0910_ ));
 sg13g2_mux2_1 \register_file_i/_7051_  (.A0(\register_file_i/rf_reg_927_ ),
    .A1(net564),
    .S(net902),
    .X(\register_file_i/_0911_ ));
 sg13g2_nor2_1 \register_file_i/_7052_  (.A(\register_file_i/_2799_ ),
    .B(\register_file_i/_2946_ ),
    .Y(\register_file_i/_3034_ ));
 sg13g2_buf_2 fanout16 (.A(net18),
    .X(net16));
 sg13g2_mux2_1 \register_file_i/_7054_  (.A0(\register_file_i/rf_reg_928_ ),
    .A1(net753),
    .S(net895),
    .X(\register_file_i/_0912_ ));
 sg13g2_mux2_1 \register_file_i/_7055_  (.A0(\register_file_i/rf_reg_929_ ),
    .A1(net1000),
    .S(net894),
    .X(\register_file_i/_0913_ ));
 sg13g2_mux2_1 \register_file_i/_7056_  (.A0(net579),
    .A1(\register_file_i/rf_reg_92_ ),
    .S(net810),
    .X(\register_file_i/_0914_ ));
 sg13g2_mux2_1 \register_file_i/_7057_  (.A0(\register_file_i/rf_reg_930_ ),
    .A1(net884),
    .S(net894),
    .X(\register_file_i/_0915_ ));
 sg13g2_mux2_1 \register_file_i/_7058_  (.A0(\register_file_i/rf_reg_931_ ),
    .A1(net1020),
    .S(net894),
    .X(\register_file_i/_0916_ ));
 sg13g2_mux2_1 \register_file_i/_7059_  (.A0(\register_file_i/rf_reg_932_ ),
    .A1(net1017),
    .S(net893),
    .X(\register_file_i/_0917_ ));
 sg13g2_mux2_1 \register_file_i/_7060_  (.A0(\register_file_i/rf_reg_933_ ),
    .A1(net997),
    .S(net893),
    .X(\register_file_i/_0918_ ));
 sg13g2_mux2_1 \register_file_i/_7061_  (.A0(\register_file_i/rf_reg_934_ ),
    .A1(net883),
    .S(net893),
    .X(\register_file_i/_0919_ ));
 sg13g2_mux2_1 \register_file_i/_7062_  (.A0(\register_file_i/rf_reg_935_ ),
    .A1(net993),
    .S(net893),
    .X(\register_file_i/_0920_ ));
 sg13g2_mux2_1 \register_file_i/_7063_  (.A0(\register_file_i/rf_reg_936_ ),
    .A1(net877),
    .S(net893),
    .X(\register_file_i/_0921_ ));
 sg13g2_mux2_1 \register_file_i/_7064_  (.A0(\register_file_i/rf_reg_937_ ),
    .A1(net806),
    .S(net893),
    .X(\register_file_i/_0922_ ));
 sg13g2_buf_1 fanout15 (.A(\cs_registers_i/_2184_ ),
    .X(net15));
 sg13g2_mux2_1 \register_file_i/_7066_  (.A0(\register_file_i/rf_reg_938_ ),
    .A1(net797),
    .S(net894),
    .X(\register_file_i/_0923_ ));
 sg13g2_mux2_1 \register_file_i/_7067_  (.A0(\register_file_i/rf_reg_939_ ),
    .A1(net792),
    .S(net893),
    .X(\register_file_i/_0924_ ));
 sg13g2_mux2_1 \register_file_i/_7068_  (.A0(net570),
    .A1(\register_file_i/rf_reg_93_ ),
    .S(net810),
    .X(\register_file_i/_0925_ ));
 sg13g2_mux2_1 \register_file_i/_7069_  (.A0(\register_file_i/rf_reg_940_ ),
    .A1(net801),
    .S(net894),
    .X(\register_file_i/_0926_ ));
 sg13g2_mux2_1 \register_file_i/_7070_  (.A0(\register_file_i/rf_reg_941_ ),
    .A1(net788),
    .S(net895),
    .X(\register_file_i/_0927_ ));
 sg13g2_mux2_1 \register_file_i/_7071_  (.A0(\register_file_i/rf_reg_942_ ),
    .A1(net750),
    .S(net895),
    .X(\register_file_i/_0928_ ));
 sg13g2_mux2_1 \register_file_i/_7072_  (.A0(\register_file_i/rf_reg_943_ ),
    .A1(net782),
    .S(net895),
    .X(\register_file_i/_0929_ ));
 sg13g2_mux2_1 \register_file_i/_7073_  (.A0(\register_file_i/rf_reg_944_ ),
    .A1(net711),
    .S(net895),
    .X(\register_file_i/_0930_ ));
 sg13g2_mux2_1 \register_file_i/_7074_  (.A0(\register_file_i/rf_reg_945_ ),
    .A1(net725),
    .S(net896),
    .X(\register_file_i/_0931_ ));
 sg13g2_mux2_1 \register_file_i/_7075_  (.A0(\register_file_i/rf_reg_946_ ),
    .A1(net705),
    .S(net896),
    .X(\register_file_i/_0932_ ));
 sg13g2_mux2_1 \register_file_i/_7076_  (.A0(\register_file_i/rf_reg_947_ ),
    .A1(net700),
    .S(net895),
    .X(\register_file_i/_0933_ ));
 sg13g2_buf_2 fanout14 (.A(net15),
    .X(net14));
 sg13g2_mux2_1 \register_file_i/_7078_  (.A0(\register_file_i/rf_reg_948_ ),
    .A1(net739),
    .S(net896),
    .X(\register_file_i/_0934_ ));
 sg13g2_mux2_1 \register_file_i/_7079_  (.A0(\register_file_i/rf_reg_949_ ),
    .A1(net674),
    .S(net896),
    .X(\register_file_i/_0935_ ));
 sg13g2_mux2_1 \register_file_i/_7080_  (.A0(net576),
    .A1(\register_file_i/rf_reg_94_ ),
    .S(net813),
    .X(\register_file_i/_0936_ ));
 sg13g2_mux2_1 \register_file_i/_7081_  (.A0(\register_file_i/rf_reg_950_ ),
    .A1(net696),
    .S(net897),
    .X(\register_file_i/_0937_ ));
 sg13g2_mux2_1 \register_file_i/_7082_  (.A0(\register_file_i/rf_reg_951_ ),
    .A1(net687),
    .S(net894),
    .X(\register_file_i/_0938_ ));
 sg13g2_mux2_1 \register_file_i/_7083_  (.A0(\register_file_i/rf_reg_952_ ),
    .A1(net685),
    .S(net897),
    .X(\register_file_i/_0939_ ));
 sg13g2_mux2_1 \register_file_i/_7084_  (.A0(\register_file_i/rf_reg_953_ ),
    .A1(net603),
    .S(net897),
    .X(\register_file_i/_0940_ ));
 sg13g2_mux2_1 \register_file_i/_7085_  (.A0(\register_file_i/rf_reg_954_ ),
    .A1(net668),
    .S(net894),
    .X(\register_file_i/_0941_ ));
 sg13g2_mux2_1 \register_file_i/_7086_  (.A0(\register_file_i/rf_reg_955_ ),
    .A1(net584),
    .S(net898),
    .X(\register_file_i/_0942_ ));
 sg13g2_mux2_1 \register_file_i/_7087_  (.A0(\register_file_i/rf_reg_956_ ),
    .A1(net579),
    .S(net898),
    .X(\register_file_i/_0943_ ));
 sg13g2_mux2_1 \register_file_i/_7088_  (.A0(\register_file_i/rf_reg_957_ ),
    .A1(net570),
    .S(net893),
    .X(\register_file_i/_0944_ ));
 sg13g2_mux2_1 \register_file_i/_7089_  (.A0(\register_file_i/rf_reg_958_ ),
    .A1(net574),
    .S(net895),
    .X(\register_file_i/_0945_ ));
 sg13g2_mux2_1 \register_file_i/_7090_  (.A0(\register_file_i/rf_reg_959_ ),
    .A1(net564),
    .S(net895),
    .X(\register_file_i/_0946_ ));
 sg13g2_mux2_1 \register_file_i/_7091_  (.A0(net565),
    .A1(\register_file_i/rf_reg_95_ ),
    .S(net812),
    .X(\register_file_i/_0947_ ));
 sg13g2_nor2_1 \register_file_i/_7092_  (.A(\register_file_i/_2799_ ),
    .B(\register_file_i/_2951_ ),
    .Y(\register_file_i/_3038_ ));
 sg13g2_buf_4 fanout13 (.X(net13),
    .A(net15));
 sg13g2_mux2_1 \register_file_i/_7094_  (.A0(\register_file_i/rf_reg_960_ ),
    .A1(net752),
    .S(net889),
    .X(\register_file_i/_0948_ ));
 sg13g2_mux2_1 \register_file_i/_7095_  (.A0(\register_file_i/rf_reg_961_ ),
    .A1(net1001),
    .S(net889),
    .X(\register_file_i/_0949_ ));
 sg13g2_mux2_1 \register_file_i/_7096_  (.A0(\register_file_i/rf_reg_962_ ),
    .A1(net884),
    .S(net889),
    .X(\register_file_i/_0950_ ));
 sg13g2_mux2_1 \register_file_i/_7097_  (.A0(\register_file_i/rf_reg_963_ ),
    .A1(net1022),
    .S(net889),
    .X(\register_file_i/_0951_ ));
 sg13g2_mux2_1 \register_file_i/_7098_  (.A0(\register_file_i/rf_reg_964_ ),
    .A1(net1017),
    .S(net888),
    .X(\register_file_i/_0952_ ));
 sg13g2_mux2_1 \register_file_i/_7099_  (.A0(\register_file_i/rf_reg_965_ ),
    .A1(net997),
    .S(net888),
    .X(\register_file_i/_0953_ ));
 sg13g2_mux2_1 \register_file_i/_7100_  (.A0(\register_file_i/rf_reg_966_ ),
    .A1(net882),
    .S(net888),
    .X(\register_file_i/_0954_ ));
 sg13g2_mux2_1 \register_file_i/_7101_  (.A0(\register_file_i/rf_reg_967_ ),
    .A1(net993),
    .S(net888),
    .X(\register_file_i/_0955_ ));
 sg13g2_mux2_1 \register_file_i/_7102_  (.A0(\register_file_i/rf_reg_968_ ),
    .A1(net877),
    .S(net888),
    .X(\register_file_i/_0956_ ));
 sg13g2_mux2_1 \register_file_i/_7103_  (.A0(\register_file_i/rf_reg_969_ ),
    .A1(net806),
    .S(net888),
    .X(\register_file_i/_0957_ ));
 sg13g2_mux2_1 \register_file_i/_7104_  (.A0(net756),
    .A1(\register_file_i/rf_reg_96_ ),
    .S(net870),
    .X(\register_file_i/_0958_ ));
 sg13g2_buf_2 fanout12 (.A(net15),
    .X(net12));
 sg13g2_mux2_1 \register_file_i/_7106_  (.A0(\register_file_i/rf_reg_970_ ),
    .A1(net797),
    .S(net889),
    .X(\register_file_i/_0959_ ));
 sg13g2_mux2_1 \register_file_i/_7107_  (.A0(\register_file_i/rf_reg_971_ ),
    .A1(net792),
    .S(net888),
    .X(\register_file_i/_0960_ ));
 sg13g2_mux2_1 \register_file_i/_7108_  (.A0(\register_file_i/rf_reg_972_ ),
    .A1(net801),
    .S(net889),
    .X(\register_file_i/_0961_ ));
 sg13g2_mux2_1 \register_file_i/_7109_  (.A0(\register_file_i/rf_reg_973_ ),
    .A1(net788),
    .S(net889),
    .X(\register_file_i/_0962_ ));
 sg13g2_mux2_1 \register_file_i/_7110_  (.A0(\register_file_i/rf_reg_974_ ),
    .A1(net750),
    .S(net890),
    .X(\register_file_i/_0963_ ));
 sg13g2_mux2_1 \register_file_i/_7111_  (.A0(\register_file_i/rf_reg_975_ ),
    .A1(net782),
    .S(net890),
    .X(\register_file_i/_0964_ ));
 sg13g2_mux2_1 \register_file_i/_7112_  (.A0(\register_file_i/rf_reg_976_ ),
    .A1(net711),
    .S(net891),
    .X(\register_file_i/_0965_ ));
 sg13g2_mux2_1 \register_file_i/_7113_  (.A0(\register_file_i/rf_reg_977_ ),
    .A1(net725),
    .S(net890),
    .X(\register_file_i/_0966_ ));
 sg13g2_mux2_1 \register_file_i/_7114_  (.A0(\register_file_i/rf_reg_978_ ),
    .A1(net705),
    .S(net890),
    .X(\register_file_i/_0967_ ));
 sg13g2_mux2_1 \register_file_i/_7115_  (.A0(\register_file_i/rf_reg_979_ ),
    .A1(net700),
    .S(net890),
    .X(\register_file_i/_0968_ ));
 sg13g2_mux2_1 \register_file_i/_7116_  (.A0(net1003),
    .A1(\register_file_i/rf_reg_97_ ),
    .S(net870),
    .X(\register_file_i/_0969_ ));
 sg13g2_buf_4 fanout11 (.X(net11),
    .A(net15));
 sg13g2_mux2_1 \register_file_i/_7118_  (.A0(\register_file_i/rf_reg_980_ ),
    .A1(net739),
    .S(net891),
    .X(\register_file_i/_0970_ ));
 sg13g2_mux2_1 \register_file_i/_7119_  (.A0(\register_file_i/rf_reg_981_ ),
    .A1(net674),
    .S(net891),
    .X(\register_file_i/_0971_ ));
 sg13g2_mux2_1 \register_file_i/_7120_  (.A0(\register_file_i/rf_reg_982_ ),
    .A1(net697),
    .S(net891),
    .X(\register_file_i/_0972_ ));
 sg13g2_mux2_1 \register_file_i/_7121_  (.A0(\register_file_i/rf_reg_983_ ),
    .A1(net687),
    .S(net890),
    .X(\register_file_i/_0973_ ));
 sg13g2_mux2_1 \register_file_i/_7122_  (.A0(\register_file_i/rf_reg_984_ ),
    .A1(net685),
    .S(net891),
    .X(\register_file_i/_0974_ ));
 sg13g2_mux2_1 \register_file_i/_7123_  (.A0(\register_file_i/rf_reg_985_ ),
    .A1(net603),
    .S(net891),
    .X(\register_file_i/_0975_ ));
 sg13g2_mux2_1 \register_file_i/_7124_  (.A0(\register_file_i/rf_reg_986_ ),
    .A1(net667),
    .S(net892),
    .X(\register_file_i/_0976_ ));
 sg13g2_mux2_1 \register_file_i/_7125_  (.A0(\register_file_i/rf_reg_987_ ),
    .A1(net584),
    .S(net892),
    .X(\register_file_i/_0977_ ));
 sg13g2_mux2_1 \register_file_i/_7126_  (.A0(\register_file_i/rf_reg_988_ ),
    .A1(net579),
    .S(net892),
    .X(\register_file_i/_0978_ ));
 sg13g2_mux2_1 \register_file_i/_7127_  (.A0(\register_file_i/rf_reg_989_ ),
    .A1(net570),
    .S(net888),
    .X(\register_file_i/_0979_ ));
 sg13g2_mux2_1 \register_file_i/_7128_  (.A0(net887),
    .A1(\register_file_i/rf_reg_98_ ),
    .S(net869),
    .X(\register_file_i/_0980_ ));
 sg13g2_mux2_1 \register_file_i/_7129_  (.A0(\register_file_i/rf_reg_990_ ),
    .A1(net574),
    .S(net890),
    .X(\register_file_i/_0981_ ));
 sg13g2_mux2_1 \register_file_i/_7130_  (.A0(\register_file_i/rf_reg_991_ ),
    .A1(net564),
    .S(net890),
    .X(\register_file_i/_0982_ ));
 sg13g2_mux2_1 \register_file_i/_7131_  (.A0(\register_file_i/rf_reg_992_ ),
    .A1(net752),
    .S(net986),
    .X(\register_file_i/_0983_ ));
 sg13g2_mux2_1 \register_file_i/_7132_  (.A0(\register_file_i/rf_reg_993_ ),
    .A1(net1001),
    .S(net986),
    .X(\register_file_i/_0984_ ));
 sg13g2_mux2_1 \register_file_i/_7133_  (.A0(\register_file_i/rf_reg_994_ ),
    .A1(net884),
    .S(net986),
    .X(\register_file_i/_0985_ ));
 sg13g2_mux2_1 \register_file_i/_7134_  (.A0(\register_file_i/rf_reg_995_ ),
    .A1(net1022),
    .S(net986),
    .X(\register_file_i/_0986_ ));
 sg13g2_mux2_1 \register_file_i/_7135_  (.A0(\register_file_i/rf_reg_996_ ),
    .A1(net1017),
    .S(net985),
    .X(\register_file_i/_0987_ ));
 sg13g2_mux2_1 \register_file_i/_7136_  (.A0(\register_file_i/rf_reg_997_ ),
    .A1(net997),
    .S(net985),
    .X(\register_file_i/_0988_ ));
 sg13g2_mux2_1 \register_file_i/_7137_  (.A0(\register_file_i/rf_reg_998_ ),
    .A1(net882),
    .S(net985),
    .X(\register_file_i/_0989_ ));
 sg13g2_mux2_1 \register_file_i/_7138_  (.A0(\register_file_i/rf_reg_999_ ),
    .A1(net993),
    .S(net985),
    .X(\register_file_i/_0990_ ));
 sg13g2_mux2_1 \register_file_i/_7139_  (.A0(net1024),
    .A1(\register_file_i/rf_reg_99_ ),
    .S(net869),
    .X(\register_file_i/_0991_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1000__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0000_ ),
    .Q_N(\register_file_i/_4033_ ),
    .Q(\register_file_i/rf_reg_1000_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1001__reg  (.CLK(clknet_leaf_341_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0001_ ),
    .Q_N(\register_file_i/_4032_ ),
    .Q(\register_file_i/rf_reg_1001_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1002__reg  (.CLK(clknet_leaf_339_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0002_ ),
    .Q_N(\register_file_i/_4031_ ),
    .Q(\register_file_i/rf_reg_1002_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1003__reg  (.CLK(clknet_leaf_341_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0003_ ),
    .Q_N(\register_file_i/_4030_ ),
    .Q(\register_file_i/rf_reg_1003_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1004__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0004_ ),
    .Q_N(\register_file_i/_4029_ ),
    .Q(\register_file_i/rf_reg_1004_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1005__reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0005_ ),
    .Q_N(\register_file_i/_4028_ ),
    .Q(\register_file_i/rf_reg_1005_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1006__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0006_ ),
    .Q_N(\register_file_i/_4027_ ),
    .Q(\register_file_i/rf_reg_1006_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1007__reg  (.CLK(clknet_leaf_160_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0007_ ),
    .Q_N(\register_file_i/_4026_ ),
    .Q(\register_file_i/rf_reg_1007_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1008__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0008_ ),
    .Q_N(\register_file_i/_4025_ ),
    .Q(\register_file_i/rf_reg_1008_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1009__reg  (.CLK(clknet_leaf_135_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0009_ ),
    .Q_N(\register_file_i/_4024_ ),
    .Q(\register_file_i/rf_reg_1009_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_100__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0010_ ),
    .Q_N(\register_file_i/_4023_ ),
    .Q(\register_file_i/rf_reg_100_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1010__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2216),
    .D(\register_file_i/_0011_ ),
    .Q_N(\register_file_i/_4022_ ),
    .Q(\register_file_i/rf_reg_1010_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1011__reg  (.CLK(clknet_leaf_134_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0012_ ),
    .Q_N(\register_file_i/_4021_ ),
    .Q(\register_file_i/rf_reg_1011_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1012__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0013_ ),
    .Q_N(\register_file_i/_4020_ ),
    .Q(\register_file_i/rf_reg_1012_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1013__reg  (.CLK(clknet_leaf_155_clk_i),
    .RESET_B(net2264),
    .D(\register_file_i/_0014_ ),
    .Q_N(\register_file_i/_4019_ ),
    .Q(\register_file_i/rf_reg_1013_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1014__reg  (.CLK(clknet_leaf_171_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0015_ ),
    .Q_N(\register_file_i/_4018_ ),
    .Q(\register_file_i/rf_reg_1014_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1015__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0016_ ),
    .Q_N(\register_file_i/_4017_ ),
    .Q(\register_file_i/rf_reg_1015_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1016__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0017_ ),
    .Q_N(\register_file_i/_4016_ ),
    .Q(\register_file_i/rf_reg_1016_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1017__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0018_ ),
    .Q_N(\register_file_i/_4015_ ),
    .Q(\register_file_i/rf_reg_1017_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1018__reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0019_ ),
    .Q_N(\register_file_i/_4014_ ),
    .Q(\register_file_i/rf_reg_1018_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1019__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0020_ ),
    .Q_N(\register_file_i/_4013_ ),
    .Q(\register_file_i/rf_reg_1019_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_101__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0021_ ),
    .Q_N(\register_file_i/_4012_ ),
    .Q(\register_file_i/rf_reg_101_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1020__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0022_ ),
    .Q_N(\register_file_i/_4011_ ),
    .Q(\register_file_i/rf_reg_1020_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1021__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0023_ ),
    .Q_N(\register_file_i/_4010_ ),
    .Q(\register_file_i/rf_reg_1021_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1022__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0024_ ),
    .Q_N(\register_file_i/_4009_ ),
    .Q(\register_file_i/rf_reg_1022_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_1023__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0025_ ),
    .Q_N(\register_file_i/_4008_ ),
    .Q(\register_file_i/rf_reg_1023_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_102__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0026_ ),
    .Q_N(\register_file_i/_4007_ ),
    .Q(\register_file_i/rf_reg_102_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_103__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0027_ ),
    .Q_N(\register_file_i/_4006_ ),
    .Q(\register_file_i/rf_reg_103_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_104__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0028_ ),
    .Q_N(\register_file_i/_4005_ ),
    .Q(\register_file_i/rf_reg_104_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_105__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0029_ ),
    .Q_N(\register_file_i/_4004_ ),
    .Q(\register_file_i/rf_reg_105_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_106__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0030_ ),
    .Q_N(\register_file_i/_4003_ ),
    .Q(\register_file_i/rf_reg_106_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_107__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0031_ ),
    .Q_N(\register_file_i/_4002_ ),
    .Q(\register_file_i/rf_reg_107_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_108__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0032_ ),
    .Q_N(\register_file_i/_4001_ ),
    .Q(\register_file_i/rf_reg_108_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_109__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0033_ ),
    .Q_N(\register_file_i/_4000_ ),
    .Q(\register_file_i/rf_reg_109_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_110__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0034_ ),
    .Q_N(\register_file_i/_3999_ ),
    .Q(\register_file_i/rf_reg_110_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_111__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0035_ ),
    .Q_N(\register_file_i/_3998_ ),
    .Q(\register_file_i/rf_reg_111_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_112__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0036_ ),
    .Q_N(\register_file_i/_3997_ ),
    .Q(\register_file_i/rf_reg_112_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_113__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0037_ ),
    .Q_N(\register_file_i/_3996_ ),
    .Q(\register_file_i/rf_reg_113_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_114__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0038_ ),
    .Q_N(\register_file_i/_3995_ ),
    .Q(\register_file_i/rf_reg_114_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_115__reg  (.CLK(clknet_leaf_164_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0039_ ),
    .Q_N(\register_file_i/_3994_ ),
    .Q(\register_file_i/rf_reg_115_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_116__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0040_ ),
    .Q_N(\register_file_i/_3993_ ),
    .Q(\register_file_i/rf_reg_116_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_117__reg  (.CLK(clknet_leaf_166_clk_i),
    .RESET_B(net2266),
    .D(\register_file_i/_0041_ ),
    .Q_N(\register_file_i/_3992_ ),
    .Q(\register_file_i/rf_reg_117_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_118__reg  (.CLK(clknet_leaf_170_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0042_ ),
    .Q_N(\register_file_i/_3991_ ),
    .Q(\register_file_i/rf_reg_118_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_119__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0043_ ),
    .Q_N(\register_file_i/_3990_ ),
    .Q(\register_file_i/rf_reg_119_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_120__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0044_ ),
    .Q_N(\register_file_i/_3989_ ),
    .Q(\register_file_i/rf_reg_120_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_121__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0045_ ),
    .Q_N(\register_file_i/_3988_ ),
    .Q(\register_file_i/rf_reg_121_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_122__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0046_ ),
    .Q_N(\register_file_i/_3987_ ),
    .Q(\register_file_i/rf_reg_122_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_123__reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(net2300),
    .D(\register_file_i/_0047_ ),
    .Q_N(\register_file_i/_3986_ ),
    .Q(\register_file_i/rf_reg_123_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_124__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0048_ ),
    .Q_N(\register_file_i/_3985_ ),
    .Q(\register_file_i/rf_reg_124_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_125__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0049_ ),
    .Q_N(\register_file_i/_3984_ ),
    .Q(\register_file_i/rf_reg_125_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_126__reg  (.CLK(clknet_leaf_167_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0050_ ),
    .Q_N(\register_file_i/_3983_ ),
    .Q(\register_file_i/rf_reg_126_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_127__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0051_ ),
    .Q_N(\register_file_i/_3982_ ),
    .Q(\register_file_i/rf_reg_127_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_128__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0052_ ),
    .Q_N(\register_file_i/_3981_ ),
    .Q(\register_file_i/rf_reg_128_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_129__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0053_ ),
    .Q_N(\register_file_i/_3980_ ),
    .Q(\register_file_i/rf_reg_129_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_130__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0054_ ),
    .Q_N(\register_file_i/_3979_ ),
    .Q(\register_file_i/rf_reg_130_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_131__reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0055_ ),
    .Q_N(\register_file_i/_3978_ ),
    .Q(\register_file_i/rf_reg_131_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_132__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0056_ ),
    .Q_N(\register_file_i/_3977_ ),
    .Q(\register_file_i/rf_reg_132_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_133__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0057_ ),
    .Q_N(\register_file_i/_3976_ ),
    .Q(\register_file_i/rf_reg_133_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_134__reg  (.CLK(clknet_leaf_312_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0058_ ),
    .Q_N(\register_file_i/_3975_ ),
    .Q(\register_file_i/rf_reg_134_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_135__reg  (.CLK(clknet_leaf_312_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0059_ ),
    .Q_N(\register_file_i/_3974_ ),
    .Q(\register_file_i/rf_reg_135_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_136__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0060_ ),
    .Q_N(\register_file_i/_3973_ ),
    .Q(\register_file_i/rf_reg_136_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_137__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0061_ ),
    .Q_N(\register_file_i/_3972_ ),
    .Q(\register_file_i/rf_reg_137_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_138__reg  (.CLK(clknet_leaf_337_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0062_ ),
    .Q_N(\register_file_i/_3971_ ),
    .Q(\register_file_i/rf_reg_138_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_139__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0063_ ),
    .Q_N(\register_file_i/_3970_ ),
    .Q(\register_file_i/rf_reg_139_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_140__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0064_ ),
    .Q_N(\register_file_i/_3969_ ),
    .Q(\register_file_i/rf_reg_140_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_141__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0065_ ),
    .Q_N(\register_file_i/_3968_ ),
    .Q(\register_file_i/rf_reg_141_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_142__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0066_ ),
    .Q_N(\register_file_i/_3967_ ),
    .Q(\register_file_i/rf_reg_142_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_143__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0067_ ),
    .Q_N(\register_file_i/_3966_ ),
    .Q(\register_file_i/rf_reg_143_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_144__reg  (.CLK(clknet_leaf_160_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0068_ ),
    .Q_N(\register_file_i/_3965_ ),
    .Q(\register_file_i/rf_reg_144_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_145__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0069_ ),
    .Q_N(\register_file_i/_3964_ ),
    .Q(\register_file_i/rf_reg_145_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_146__reg  (.CLK(clknet_leaf_157_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0070_ ),
    .Q_N(\register_file_i/_3963_ ),
    .Q(\register_file_i/rf_reg_146_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_147__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0071_ ),
    .Q_N(\register_file_i/_3962_ ),
    .Q(\register_file_i/rf_reg_147_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_148__reg  (.CLK(clknet_leaf_151_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0072_ ),
    .Q_N(\register_file_i/_3961_ ),
    .Q(\register_file_i/rf_reg_148_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_149__reg  (.CLK(clknet_leaf_157_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0073_ ),
    .Q_N(\register_file_i/_3960_ ),
    .Q(\register_file_i/rf_reg_149_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_150__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0074_ ),
    .Q_N(\register_file_i/_3959_ ),
    .Q(\register_file_i/rf_reg_150_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_151__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0075_ ),
    .Q_N(\register_file_i/_3958_ ),
    .Q(\register_file_i/rf_reg_151_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_152__reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0076_ ),
    .Q_N(\register_file_i/_3957_ ),
    .Q(\register_file_i/rf_reg_152_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_153__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0077_ ),
    .Q_N(\register_file_i/_3956_ ),
    .Q(\register_file_i/rf_reg_153_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_154__reg  (.CLK(clknet_leaf_55_clk_i),
    .RESET_B(net2300),
    .D(\register_file_i/_0078_ ),
    .Q_N(\register_file_i/_3955_ ),
    .Q(\register_file_i/rf_reg_154_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_155__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0079_ ),
    .Q_N(\register_file_i/_3954_ ),
    .Q(\register_file_i/rf_reg_155_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_156__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0080_ ),
    .Q_N(\register_file_i/_3953_ ),
    .Q(\register_file_i/rf_reg_156_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_157__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0081_ ),
    .Q_N(\register_file_i/_3952_ ),
    .Q(\register_file_i/rf_reg_157_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_158__reg  (.CLK(clknet_leaf_167_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0082_ ),
    .Q_N(\register_file_i/_3951_ ),
    .Q(\register_file_i/rf_reg_158_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_159__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0083_ ),
    .Q_N(\register_file_i/_3950_ ),
    .Q(\register_file_i/rf_reg_159_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_160__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0084_ ),
    .Q_N(\register_file_i/_3949_ ),
    .Q(\register_file_i/rf_reg_160_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_161__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0085_ ),
    .Q_N(\register_file_i/_3948_ ),
    .Q(\register_file_i/rf_reg_161_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_162__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0086_ ),
    .Q_N(\register_file_i/_3947_ ),
    .Q(\register_file_i/rf_reg_162_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_163__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0087_ ),
    .Q_N(\register_file_i/_3946_ ),
    .Q(\register_file_i/rf_reg_163_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_164__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0088_ ),
    .Q_N(\register_file_i/_3945_ ),
    .Q(\register_file_i/rf_reg_164_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_165__reg  (.CLK(clknet_leaf_312_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0089_ ),
    .Q_N(\register_file_i/_3944_ ),
    .Q(\register_file_i/rf_reg_165_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_166__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0090_ ),
    .Q_N(\register_file_i/_3943_ ),
    .Q(\register_file_i/rf_reg_166_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_167__reg  (.CLK(clknet_leaf_313_clk_i),
    .RESET_B(net2289),
    .D(\register_file_i/_0091_ ),
    .Q_N(\register_file_i/_3942_ ),
    .Q(\register_file_i/rf_reg_167_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_168__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0092_ ),
    .Q_N(\register_file_i/_3941_ ),
    .Q(\register_file_i/rf_reg_168_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_169__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0093_ ),
    .Q_N(\register_file_i/_3940_ ),
    .Q(\register_file_i/rf_reg_169_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_170__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0094_ ),
    .Q_N(\register_file_i/_3939_ ),
    .Q(\register_file_i/rf_reg_170_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_171__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0095_ ),
    .Q_N(\register_file_i/_3938_ ),
    .Q(\register_file_i/rf_reg_171_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_172__reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0096_ ),
    .Q_N(\register_file_i/_3937_ ),
    .Q(\register_file_i/rf_reg_172_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_173__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0097_ ),
    .Q_N(\register_file_i/_3936_ ),
    .Q(\register_file_i/rf_reg_173_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_174__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0098_ ),
    .Q_N(\register_file_i/_3935_ ),
    .Q(\register_file_i/rf_reg_174_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_175__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0099_ ),
    .Q_N(\register_file_i/_3934_ ),
    .Q(\register_file_i/rf_reg_175_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_176__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0100_ ),
    .Q_N(\register_file_i/_3933_ ),
    .Q(\register_file_i/rf_reg_176_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_177__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0101_ ),
    .Q_N(\register_file_i/_3932_ ),
    .Q(\register_file_i/rf_reg_177_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_178__reg  (.CLK(clknet_leaf_157_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0102_ ),
    .Q_N(\register_file_i/_3931_ ),
    .Q(\register_file_i/rf_reg_178_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_179__reg  (.CLK(clknet_leaf_153_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0103_ ),
    .Q_N(\register_file_i/_3930_ ),
    .Q(\register_file_i/rf_reg_179_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_180__reg  (.CLK(clknet_leaf_153_clk_i),
    .RESET_B(net2255),
    .D(\register_file_i/_0104_ ),
    .Q_N(\register_file_i/_3929_ ),
    .Q(\register_file_i/rf_reg_180_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_181__reg  (.CLK(clknet_leaf_157_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0105_ ),
    .Q_N(\register_file_i/_3928_ ),
    .Q(\register_file_i/rf_reg_181_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_182__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0106_ ),
    .Q_N(\register_file_i/_3927_ ),
    .Q(\register_file_i/rf_reg_182_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_183__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0107_ ),
    .Q_N(\register_file_i/_3926_ ),
    .Q(\register_file_i/rf_reg_183_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_184__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0108_ ),
    .Q_N(\register_file_i/_3925_ ),
    .Q(\register_file_i/rf_reg_184_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_185__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0109_ ),
    .Q_N(\register_file_i/_3924_ ),
    .Q(\register_file_i/rf_reg_185_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_186__reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0110_ ),
    .Q_N(\register_file_i/_3923_ ),
    .Q(\register_file_i/rf_reg_186_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_187__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0111_ ),
    .Q_N(\register_file_i/_3922_ ),
    .Q(\register_file_i/rf_reg_187_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_188__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0112_ ),
    .Q_N(\register_file_i/_3921_ ),
    .Q(\register_file_i/rf_reg_188_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_189__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0113_ ),
    .Q_N(\register_file_i/_3920_ ),
    .Q(\register_file_i/rf_reg_189_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_190__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0114_ ),
    .Q_N(\register_file_i/_3919_ ),
    .Q(\register_file_i/rf_reg_190_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_191__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2255),
    .D(\register_file_i/_0115_ ),
    .Q_N(\register_file_i/_3918_ ),
    .Q(\register_file_i/rf_reg_191_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_192__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0116_ ),
    .Q_N(\register_file_i/_3917_ ),
    .Q(\register_file_i/rf_reg_192_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_193__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0117_ ),
    .Q_N(\register_file_i/_3916_ ),
    .Q(\register_file_i/rf_reg_193_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_194__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2188),
    .D(\register_file_i/_0118_ ),
    .Q_N(\register_file_i/_3915_ ),
    .Q(\register_file_i/rf_reg_194_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_195__reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0119_ ),
    .Q_N(\register_file_i/_3914_ ),
    .Q(\register_file_i/rf_reg_195_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_196__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2288),
    .D(\register_file_i/_0120_ ),
    .Q_N(\register_file_i/_3913_ ),
    .Q(\register_file_i/rf_reg_196_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_197__reg  (.CLK(clknet_leaf_309_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0121_ ),
    .Q_N(\register_file_i/_3912_ ),
    .Q(\register_file_i/rf_reg_197_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_198__reg  (.CLK(clknet_leaf_309_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0122_ ),
    .Q_N(\register_file_i/_3911_ ),
    .Q(\register_file_i/rf_reg_198_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_199__reg  (.CLK(clknet_leaf_312_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0123_ ),
    .Q_N(\register_file_i/_3910_ ),
    .Q(\register_file_i/rf_reg_199_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_200__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0124_ ),
    .Q_N(\register_file_i/_3909_ ),
    .Q(\register_file_i/rf_reg_200_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_201__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0125_ ),
    .Q_N(\register_file_i/_3908_ ),
    .Q(\register_file_i/rf_reg_201_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_202__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0126_ ),
    .Q_N(\register_file_i/_3907_ ),
    .Q(\register_file_i/rf_reg_202_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_203__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0127_ ),
    .Q_N(\register_file_i/_3906_ ),
    .Q(\register_file_i/rf_reg_203_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_204__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0128_ ),
    .Q_N(\register_file_i/_3905_ ),
    .Q(\register_file_i/rf_reg_204_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_205__reg  (.CLK(clknet_leaf_171_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0129_ ),
    .Q_N(\register_file_i/_3904_ ),
    .Q(\register_file_i/rf_reg_205_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_206__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0130_ ),
    .Q_N(\register_file_i/_3903_ ),
    .Q(\register_file_i/rf_reg_206_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_207__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2249),
    .D(\register_file_i/_0131_ ),
    .Q_N(\register_file_i/_3902_ ),
    .Q(\register_file_i/rf_reg_207_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_208__reg  (.CLK(clknet_leaf_160_clk_i),
    .RESET_B(net2242),
    .D(\register_file_i/_0132_ ),
    .Q_N(\register_file_i/_3901_ ),
    .Q(\register_file_i/rf_reg_208_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_209__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0133_ ),
    .Q_N(\register_file_i/_3900_ ),
    .Q(\register_file_i/rf_reg_209_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_210__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0134_ ),
    .Q_N(\register_file_i/_3899_ ),
    .Q(\register_file_i/rf_reg_210_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_211__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0135_ ),
    .Q_N(\register_file_i/_3898_ ),
    .Q(\register_file_i/rf_reg_211_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_212__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0136_ ),
    .Q_N(\register_file_i/_3897_ ),
    .Q(\register_file_i/rf_reg_212_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_213__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2246),
    .D(\register_file_i/_0137_ ),
    .Q_N(\register_file_i/_3896_ ),
    .Q(\register_file_i/rf_reg_213_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_214__reg  (.CLK(clknet_leaf_169_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0138_ ),
    .Q_N(\register_file_i/_3895_ ),
    .Q(\register_file_i/rf_reg_214_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_215__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0139_ ),
    .Q_N(\register_file_i/_3894_ ),
    .Q(\register_file_i/rf_reg_215_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_216__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0140_ ),
    .Q_N(\register_file_i/_3893_ ),
    .Q(\register_file_i/rf_reg_216_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_217__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0141_ ),
    .Q_N(\register_file_i/_3892_ ),
    .Q(\register_file_i/rf_reg_217_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_218__reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(net2300),
    .D(\register_file_i/_0142_ ),
    .Q_N(\register_file_i/_3891_ ),
    .Q(\register_file_i/rf_reg_218_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_219__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0143_ ),
    .Q_N(\register_file_i/_3890_ ),
    .Q(\register_file_i/rf_reg_219_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_220__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0144_ ),
    .Q_N(\register_file_i/_3889_ ),
    .Q(\register_file_i/rf_reg_220_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_221__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0145_ ),
    .Q_N(\register_file_i/_3888_ ),
    .Q(\register_file_i/rf_reg_221_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_222__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0146_ ),
    .Q_N(\register_file_i/_3887_ ),
    .Q(\register_file_i/rf_reg_222_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_223__reg  (.CLK(clknet_leaf_170_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0147_ ),
    .Q_N(\register_file_i/_3886_ ),
    .Q(\register_file_i/rf_reg_223_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_224__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0148_ ),
    .Q_N(\register_file_i/_3885_ ),
    .Q(\register_file_i/rf_reg_224_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_225__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0149_ ),
    .Q_N(\register_file_i/_3884_ ),
    .Q(\register_file_i/rf_reg_225_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_226__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2188),
    .D(\register_file_i/_0150_ ),
    .Q_N(\register_file_i/_3883_ ),
    .Q(\register_file_i/rf_reg_226_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_227__reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0151_ ),
    .Q_N(\register_file_i/_3882_ ),
    .Q(\register_file_i/rf_reg_227_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_228__reg  (.CLK(clknet_leaf_307_clk_i),
    .RESET_B(net2288),
    .D(\register_file_i/_0152_ ),
    .Q_N(\register_file_i/_3881_ ),
    .Q(\register_file_i/rf_reg_228_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_229__reg  (.CLK(clknet_leaf_309_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0153_ ),
    .Q_N(\register_file_i/_3880_ ),
    .Q(\register_file_i/rf_reg_229_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_230__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0154_ ),
    .Q_N(\register_file_i/_3879_ ),
    .Q(\register_file_i/rf_reg_230_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_231__reg  (.CLK(clknet_leaf_312_clk_i),
    .RESET_B(net2287),
    .D(\register_file_i/_0155_ ),
    .Q_N(\register_file_i/_3878_ ),
    .Q(\register_file_i/rf_reg_231_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_232__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0156_ ),
    .Q_N(\register_file_i/_3877_ ),
    .Q(\register_file_i/rf_reg_232_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_233__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0157_ ),
    .Q_N(\register_file_i/_3876_ ),
    .Q(\register_file_i/rf_reg_233_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_234__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0158_ ),
    .Q_N(\register_file_i/_3875_ ),
    .Q(\register_file_i/rf_reg_234_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_235__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0159_ ),
    .Q_N(\register_file_i/_3874_ ),
    .Q(\register_file_i/rf_reg_235_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_236__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0160_ ),
    .Q_N(\register_file_i/_3873_ ),
    .Q(\register_file_i/rf_reg_236_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_237__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0161_ ),
    .Q_N(\register_file_i/_3872_ ),
    .Q(\register_file_i/rf_reg_237_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_238__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0162_ ),
    .Q_N(\register_file_i/_3871_ ),
    .Q(\register_file_i/rf_reg_238_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_239__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2249),
    .D(\register_file_i/_0163_ ),
    .Q_N(\register_file_i/_3870_ ),
    .Q(\register_file_i/rf_reg_239_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_240__reg  (.CLK(clknet_leaf_160_clk_i),
    .RESET_B(net2242),
    .D(\register_file_i/_0164_ ),
    .Q_N(\register_file_i/_3869_ ),
    .Q(\register_file_i/rf_reg_240_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_241__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2268),
    .D(\register_file_i/_0165_ ),
    .Q_N(\register_file_i/_3868_ ),
    .Q(\register_file_i/rf_reg_241_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_242__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0166_ ),
    .Q_N(\register_file_i/_3867_ ),
    .Q(\register_file_i/rf_reg_242_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_243__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2260),
    .D(\register_file_i/_0167_ ),
    .Q_N(\register_file_i/_3866_ ),
    .Q(\register_file_i/rf_reg_243_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_244__reg  (.CLK(clknet_leaf_152_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0168_ ),
    .Q_N(\register_file_i/_3865_ ),
    .Q(\register_file_i/rf_reg_244_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_245__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2246),
    .D(\register_file_i/_0169_ ),
    .Q_N(\register_file_i/_3864_ ),
    .Q(\register_file_i/rf_reg_245_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_246__reg  (.CLK(clknet_leaf_169_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0170_ ),
    .Q_N(\register_file_i/_3863_ ),
    .Q(\register_file_i/rf_reg_246_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_247__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0171_ ),
    .Q_N(\register_file_i/_3862_ ),
    .Q(\register_file_i/rf_reg_247_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_248__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0172_ ),
    .Q_N(\register_file_i/_3861_ ),
    .Q(\register_file_i/rf_reg_248_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_249__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0173_ ),
    .Q_N(\register_file_i/_3860_ ),
    .Q(\register_file_i/rf_reg_249_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_250__reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(net2300),
    .D(\register_file_i/_0174_ ),
    .Q_N(\register_file_i/_3859_ ),
    .Q(\register_file_i/rf_reg_250_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_251__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0175_ ),
    .Q_N(\register_file_i/_3858_ ),
    .Q(\register_file_i/rf_reg_251_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_252__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2288),
    .D(\register_file_i/_0176_ ),
    .Q_N(\register_file_i/_3857_ ),
    .Q(\register_file_i/rf_reg_252_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_253__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0177_ ),
    .Q_N(\register_file_i/_3856_ ),
    .Q(\register_file_i/rf_reg_253_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_254__reg  (.CLK(clknet_leaf_167_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0178_ ),
    .Q_N(\register_file_i/_3855_ ),
    .Q(\register_file_i/rf_reg_254_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_255__reg  (.CLK(clknet_leaf_170_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0179_ ),
    .Q_N(\register_file_i/_3854_ ),
    .Q(\register_file_i/rf_reg_255_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_256__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2193),
    .D(\register_file_i/_0180_ ),
    .Q_N(\register_file_i/_3853_ ),
    .Q(\register_file_i/rf_reg_256_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_257__reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0181_ ),
    .Q_N(\register_file_i/_3852_ ),
    .Q(\register_file_i/rf_reg_257_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_258__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0182_ ),
    .Q_N(\register_file_i/_3851_ ),
    .Q(\register_file_i/rf_reg_258_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_259__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0183_ ),
    .Q_N(\register_file_i/_3850_ ),
    .Q(\register_file_i/rf_reg_259_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_260__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0184_ ),
    .Q_N(\register_file_i/_3849_ ),
    .Q(\register_file_i/rf_reg_260_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_261__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0185_ ),
    .Q_N(\register_file_i/_3848_ ),
    .Q(\register_file_i/rf_reg_261_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_262__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0186_ ),
    .Q_N(\register_file_i/_3847_ ),
    .Q(\register_file_i/rf_reg_262_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_263__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0187_ ),
    .Q_N(\register_file_i/_3846_ ),
    .Q(\register_file_i/rf_reg_263_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_264__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0188_ ),
    .Q_N(\register_file_i/_3845_ ),
    .Q(\register_file_i/rf_reg_264_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_265__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0189_ ),
    .Q_N(\register_file_i/_3844_ ),
    .Q(\register_file_i/rf_reg_265_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_266__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0190_ ),
    .Q_N(\register_file_i/_3843_ ),
    .Q(\register_file_i/rf_reg_266_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_267__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2118),
    .D(\register_file_i/_0191_ ),
    .Q_N(\register_file_i/_3842_ ),
    .Q(\register_file_i/rf_reg_267_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_268__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0192_ ),
    .Q_N(\register_file_i/_3841_ ),
    .Q(\register_file_i/rf_reg_268_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_269__reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0193_ ),
    .Q_N(\register_file_i/_3840_ ),
    .Q(\register_file_i/rf_reg_269_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_270__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0194_ ),
    .Q_N(\register_file_i/_3839_ ),
    .Q(\register_file_i/rf_reg_270_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_271__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0195_ ),
    .Q_N(\register_file_i/_3838_ ),
    .Q(\register_file_i/rf_reg_271_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_272__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0196_ ),
    .Q_N(\register_file_i/_3837_ ),
    .Q(\register_file_i/rf_reg_272_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_273__reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0197_ ),
    .Q_N(\register_file_i/_3836_ ),
    .Q(\register_file_i/rf_reg_273_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_274__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0198_ ),
    .Q_N(\register_file_i/_3835_ ),
    .Q(\register_file_i/rf_reg_274_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_275__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0199_ ),
    .Q_N(\register_file_i/_3834_ ),
    .Q(\register_file_i/rf_reg_275_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_276__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0200_ ),
    .Q_N(\register_file_i/_3833_ ),
    .Q(\register_file_i/rf_reg_276_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_277__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0201_ ),
    .Q_N(\register_file_i/_3832_ ),
    .Q(\register_file_i/rf_reg_277_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_278__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0202_ ),
    .Q_N(\register_file_i/_3831_ ),
    .Q(\register_file_i/rf_reg_278_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_279__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0203_ ),
    .Q_N(\register_file_i/_3830_ ),
    .Q(\register_file_i/rf_reg_279_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_280__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0204_ ),
    .Q_N(\register_file_i/_3829_ ),
    .Q(\register_file_i/rf_reg_280_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_281__reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0205_ ),
    .Q_N(\register_file_i/_3828_ ),
    .Q(\register_file_i/rf_reg_281_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_282__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0206_ ),
    .Q_N(\register_file_i/_3827_ ),
    .Q(\register_file_i/rf_reg_282_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_283__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0207_ ),
    .Q_N(\register_file_i/_3826_ ),
    .Q(\register_file_i/rf_reg_283_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_284__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0208_ ),
    .Q_N(\register_file_i/_3825_ ),
    .Q(\register_file_i/rf_reg_284_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_285__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0209_ ),
    .Q_N(\register_file_i/_3824_ ),
    .Q(\register_file_i/rf_reg_285_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_286__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0210_ ),
    .Q_N(\register_file_i/_3823_ ),
    .Q(\register_file_i/rf_reg_286_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_287__reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0211_ ),
    .Q_N(\register_file_i/_3822_ ),
    .Q(\register_file_i/rf_reg_287_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_288__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0212_ ),
    .Q_N(\register_file_i/_3821_ ),
    .Q(\register_file_i/rf_reg_288_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_289__reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0213_ ),
    .Q_N(\register_file_i/_3820_ ),
    .Q(\register_file_i/rf_reg_289_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_290__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0214_ ),
    .Q_N(\register_file_i/_3819_ ),
    .Q(\register_file_i/rf_reg_290_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_291__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0215_ ),
    .Q_N(\register_file_i/_3818_ ),
    .Q(\register_file_i/rf_reg_291_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_292__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0216_ ),
    .Q_N(\register_file_i/_3817_ ),
    .Q(\register_file_i/rf_reg_292_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_293__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0217_ ),
    .Q_N(\register_file_i/_3816_ ),
    .Q(\register_file_i/rf_reg_293_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_294__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0218_ ),
    .Q_N(\register_file_i/_3815_ ),
    .Q(\register_file_i/rf_reg_294_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_295__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0219_ ),
    .Q_N(\register_file_i/_3814_ ),
    .Q(\register_file_i/rf_reg_295_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_296__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0220_ ),
    .Q_N(\register_file_i/_3813_ ),
    .Q(\register_file_i/rf_reg_296_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_297__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0221_ ),
    .Q_N(\register_file_i/_3812_ ),
    .Q(\register_file_i/rf_reg_297_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_298__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2118),
    .D(\register_file_i/_0222_ ),
    .Q_N(\register_file_i/_3811_ ),
    .Q(\register_file_i/rf_reg_298_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_299__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2118),
    .D(\register_file_i/_0223_ ),
    .Q_N(\register_file_i/_3810_ ),
    .Q(\register_file_i/rf_reg_299_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_300__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0224_ ),
    .Q_N(\register_file_i/_3809_ ),
    .Q(\register_file_i/rf_reg_300_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_301__reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0225_ ),
    .Q_N(\register_file_i/_3808_ ),
    .Q(\register_file_i/rf_reg_301_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_302__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0226_ ),
    .Q_N(\register_file_i/_3807_ ),
    .Q(\register_file_i/rf_reg_302_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_303__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0227_ ),
    .Q_N(\register_file_i/_3806_ ),
    .Q(\register_file_i/rf_reg_303_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_304__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0228_ ),
    .Q_N(\register_file_i/_3805_ ),
    .Q(\register_file_i/rf_reg_304_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_305__reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0229_ ),
    .Q_N(\register_file_i/_3804_ ),
    .Q(\register_file_i/rf_reg_305_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_306__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0230_ ),
    .Q_N(\register_file_i/_3803_ ),
    .Q(\register_file_i/rf_reg_306_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_307__reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0231_ ),
    .Q_N(\register_file_i/_3802_ ),
    .Q(\register_file_i/rf_reg_307_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_308__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0232_ ),
    .Q_N(\register_file_i/_3801_ ),
    .Q(\register_file_i/rf_reg_308_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_309__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0233_ ),
    .Q_N(\register_file_i/_3800_ ),
    .Q(\register_file_i/rf_reg_309_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_310__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0234_ ),
    .Q_N(\register_file_i/_3799_ ),
    .Q(\register_file_i/rf_reg_310_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_311__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0235_ ),
    .Q_N(\register_file_i/_3798_ ),
    .Q(\register_file_i/rf_reg_311_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_312__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0236_ ),
    .Q_N(\register_file_i/_3797_ ),
    .Q(\register_file_i/rf_reg_312_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_313__reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0237_ ),
    .Q_N(\register_file_i/_3796_ ),
    .Q(\register_file_i/rf_reg_313_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_314__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0238_ ),
    .Q_N(\register_file_i/_3795_ ),
    .Q(\register_file_i/rf_reg_314_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_315__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0239_ ),
    .Q_N(\register_file_i/_3794_ ),
    .Q(\register_file_i/rf_reg_315_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_316__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0240_ ),
    .Q_N(\register_file_i/_3793_ ),
    .Q(\register_file_i/rf_reg_316_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_317__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0241_ ),
    .Q_N(\register_file_i/_3792_ ),
    .Q(\register_file_i/rf_reg_317_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_318__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0242_ ),
    .Q_N(\register_file_i/_3791_ ),
    .Q(\register_file_i/rf_reg_318_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_319__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0243_ ),
    .Q_N(\register_file_i/_3790_ ),
    .Q(\register_file_i/rf_reg_319_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_320__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2193),
    .D(\register_file_i/_0244_ ),
    .Q_N(\register_file_i/_3789_ ),
    .Q(\register_file_i/rf_reg_320_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_321__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0245_ ),
    .Q_N(\register_file_i/_3788_ ),
    .Q(\register_file_i/rf_reg_321_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_322__reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0246_ ),
    .Q_N(\register_file_i/_3787_ ),
    .Q(\register_file_i/rf_reg_322_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_323__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0247_ ),
    .Q_N(\register_file_i/_3786_ ),
    .Q(\register_file_i/rf_reg_323_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_324__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0248_ ),
    .Q_N(\register_file_i/_3785_ ),
    .Q(\register_file_i/rf_reg_324_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_325__reg  (.CLK(clknet_leaf_342_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0249_ ),
    .Q_N(\register_file_i/_3784_ ),
    .Q(\register_file_i/rf_reg_325_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_326__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0250_ ),
    .Q_N(\register_file_i/_3783_ ),
    .Q(\register_file_i/rf_reg_326_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_327__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0251_ ),
    .Q_N(\register_file_i/_3782_ ),
    .Q(\register_file_i/rf_reg_327_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_328__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0252_ ),
    .Q_N(\register_file_i/_3781_ ),
    .Q(\register_file_i/rf_reg_328_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_329__reg  (.CLK(clknet_leaf_342_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0253_ ),
    .Q_N(\register_file_i/_3780_ ),
    .Q(\register_file_i/rf_reg_329_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_32__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0254_ ),
    .Q_N(\register_file_i/_3779_ ),
    .Q(\register_file_i/rf_reg_32_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_330__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0255_ ),
    .Q_N(\register_file_i/_3778_ ),
    .Q(\register_file_i/rf_reg_330_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_331__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0256_ ),
    .Q_N(\register_file_i/_3777_ ),
    .Q(\register_file_i/rf_reg_331_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_332__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0257_ ),
    .Q_N(\register_file_i/_3776_ ),
    .Q(\register_file_i/rf_reg_332_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_333__reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0258_ ),
    .Q_N(\register_file_i/_3775_ ),
    .Q(\register_file_i/rf_reg_333_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_334__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0259_ ),
    .Q_N(\register_file_i/_3774_ ),
    .Q(\register_file_i/rf_reg_334_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_335__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0260_ ),
    .Q_N(\register_file_i/_3773_ ),
    .Q(\register_file_i/rf_reg_335_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_336__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0261_ ),
    .Q_N(\register_file_i/_3772_ ),
    .Q(\register_file_i/rf_reg_336_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_337__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0262_ ),
    .Q_N(\register_file_i/_3771_ ),
    .Q(\register_file_i/rf_reg_337_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_338__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0263_ ),
    .Q_N(\register_file_i/_3770_ ),
    .Q(\register_file_i/rf_reg_338_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_339__reg  (.CLK(clknet_leaf_113_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0264_ ),
    .Q_N(\register_file_i/_3769_ ),
    .Q(\register_file_i/rf_reg_339_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_33__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0265_ ),
    .Q_N(\register_file_i/_3768_ ),
    .Q(\register_file_i/rf_reg_33_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_340__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0266_ ),
    .Q_N(\register_file_i/_3767_ ),
    .Q(\register_file_i/rf_reg_340_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_341__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0267_ ),
    .Q_N(\register_file_i/_3766_ ),
    .Q(\register_file_i/rf_reg_341_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_342__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0268_ ),
    .Q_N(\register_file_i/_3765_ ),
    .Q(\register_file_i/rf_reg_342_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_343__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net2211),
    .D(\register_file_i/_0269_ ),
    .Q_N(\register_file_i/_3764_ ),
    .Q(\register_file_i/rf_reg_343_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_344__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0270_ ),
    .Q_N(\register_file_i/_3763_ ),
    .Q(\register_file_i/rf_reg_344_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_345__reg  (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0271_ ),
    .Q_N(\register_file_i/_3762_ ),
    .Q(\register_file_i/rf_reg_345_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_346__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0272_ ),
    .Q_N(\register_file_i/_3761_ ),
    .Q(\register_file_i/rf_reg_346_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_347__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0273_ ),
    .Q_N(\register_file_i/_3760_ ),
    .Q(\register_file_i/rf_reg_347_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_348__reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0274_ ),
    .Q_N(\register_file_i/_3759_ ),
    .Q(\register_file_i/rf_reg_348_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_349__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0275_ ),
    .Q_N(\register_file_i/_3758_ ),
    .Q(\register_file_i/rf_reg_349_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_34__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2188),
    .D(\register_file_i/_0276_ ),
    .Q_N(\register_file_i/_3757_ ),
    .Q(\register_file_i/rf_reg_34_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_350__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0277_ ),
    .Q_N(\register_file_i/_3756_ ),
    .Q(\register_file_i/rf_reg_350_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_351__reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0278_ ),
    .Q_N(\register_file_i/_3755_ ),
    .Q(\register_file_i/rf_reg_351_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_352__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2193),
    .D(\register_file_i/_0279_ ),
    .Q_N(\register_file_i/_3754_ ),
    .Q(\register_file_i/rf_reg_352_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_353__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2187),
    .D(\register_file_i/_0280_ ),
    .Q_N(\register_file_i/_3753_ ),
    .Q(\register_file_i/rf_reg_353_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_354__reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0281_ ),
    .Q_N(\register_file_i/_3752_ ),
    .Q(\register_file_i/rf_reg_354_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_355__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0282_ ),
    .Q_N(\register_file_i/_3751_ ),
    .Q(\register_file_i/rf_reg_355_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_356__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0283_ ),
    .Q_N(\register_file_i/_3750_ ),
    .Q(\register_file_i/rf_reg_356_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_357__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0284_ ),
    .Q_N(\register_file_i/_3749_ ),
    .Q(\register_file_i/rf_reg_357_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_358__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2157),
    .D(\register_file_i/_0285_ ),
    .Q_N(\register_file_i/_3748_ ),
    .Q(\register_file_i/rf_reg_358_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_359__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net2128),
    .D(\register_file_i/_0286_ ),
    .Q_N(\register_file_i/_3747_ ),
    .Q(\register_file_i/rf_reg_359_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_35__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0287_ ),
    .Q_N(\register_file_i/_3746_ ),
    .Q(\register_file_i/rf_reg_35_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_360__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0288_ ),
    .Q_N(\register_file_i/_3745_ ),
    .Q(\register_file_i/rf_reg_360_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_361__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2125),
    .D(\register_file_i/_0289_ ),
    .Q_N(\register_file_i/_3744_ ),
    .Q(\register_file_i/rf_reg_361_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_362__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0290_ ),
    .Q_N(\register_file_i/_3743_ ),
    .Q(\register_file_i/rf_reg_362_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_363__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2118),
    .D(\register_file_i/_0291_ ),
    .Q_N(\register_file_i/_3742_ ),
    .Q(\register_file_i/rf_reg_363_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_364__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0292_ ),
    .Q_N(\register_file_i/_3741_ ),
    .Q(\register_file_i/rf_reg_364_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_365__reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0293_ ),
    .Q_N(\register_file_i/_3740_ ),
    .Q(\register_file_i/rf_reg_365_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_366__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0294_ ),
    .Q_N(\register_file_i/_3739_ ),
    .Q(\register_file_i/rf_reg_366_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_367__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0295_ ),
    .Q_N(\register_file_i/_3738_ ),
    .Q(\register_file_i/rf_reg_367_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_368__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0296_ ),
    .Q_N(\register_file_i/_3737_ ),
    .Q(\register_file_i/rf_reg_368_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_369__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0297_ ),
    .Q_N(\register_file_i/_3736_ ),
    .Q(\register_file_i/rf_reg_369_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_36__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0298_ ),
    .Q_N(\register_file_i/_3735_ ),
    .Q(\register_file_i/rf_reg_36_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_370__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0299_ ),
    .Q_N(\register_file_i/_3734_ ),
    .Q(\register_file_i/rf_reg_370_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_371__reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0300_ ),
    .Q_N(\register_file_i/_3733_ ),
    .Q(\register_file_i/rf_reg_371_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_372__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0301_ ),
    .Q_N(\register_file_i/_3732_ ),
    .Q(\register_file_i/rf_reg_372_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_373__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0302_ ),
    .Q_N(\register_file_i/_3731_ ),
    .Q(\register_file_i/rf_reg_373_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_374__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0303_ ),
    .Q_N(\register_file_i/_3730_ ),
    .Q(\register_file_i/rf_reg_374_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_375__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0304_ ),
    .Q_N(\register_file_i/_3729_ ),
    .Q(\register_file_i/rf_reg_375_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_376__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0305_ ),
    .Q_N(\register_file_i/_3728_ ),
    .Q(\register_file_i/rf_reg_376_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_377__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0306_ ),
    .Q_N(\register_file_i/_3727_ ),
    .Q(\register_file_i/rf_reg_377_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_378__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0307_ ),
    .Q_N(\register_file_i/_3726_ ),
    .Q(\register_file_i/rf_reg_378_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_379__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0308_ ),
    .Q_N(\register_file_i/_3725_ ),
    .Q(\register_file_i/rf_reg_379_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_37__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2286),
    .D(\register_file_i/_0309_ ),
    .Q_N(\register_file_i/_3724_ ),
    .Q(\register_file_i/rf_reg_37_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_380__reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0310_ ),
    .Q_N(\register_file_i/_3723_ ),
    .Q(\register_file_i/rf_reg_380_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_381__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0311_ ),
    .Q_N(\register_file_i/_3722_ ),
    .Q(\register_file_i/rf_reg_381_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_382__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0312_ ),
    .Q_N(\register_file_i/_3721_ ),
    .Q(\register_file_i/rf_reg_382_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_383__reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0313_ ),
    .Q_N(\register_file_i/_3720_ ),
    .Q(\register_file_i/rf_reg_383_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_384__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0314_ ),
    .Q_N(\register_file_i/_3719_ ),
    .Q(\register_file_i/rf_reg_384_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_385__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0315_ ),
    .Q_N(\register_file_i/_3718_ ),
    .Q(\register_file_i/rf_reg_385_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_386__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0316_ ),
    .Q_N(\register_file_i/_3717_ ),
    .Q(\register_file_i/rf_reg_386_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_387__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0317_ ),
    .Q_N(\register_file_i/_3716_ ),
    .Q(\register_file_i/rf_reg_387_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_388__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0318_ ),
    .Q_N(\register_file_i/_3715_ ),
    .Q(\register_file_i/rf_reg_388_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_389__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0319_ ),
    .Q_N(\register_file_i/_3714_ ),
    .Q(\register_file_i/rf_reg_389_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_38__reg  (.CLK(clknet_leaf_309_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0320_ ),
    .Q_N(\register_file_i/_3713_ ),
    .Q(\register_file_i/rf_reg_38_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_390__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0321_ ),
    .Q_N(\register_file_i/_3712_ ),
    .Q(\register_file_i/rf_reg_390_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_391__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0322_ ),
    .Q_N(\register_file_i/_3711_ ),
    .Q(\register_file_i/rf_reg_391_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_392__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0323_ ),
    .Q_N(\register_file_i/_3710_ ),
    .Q(\register_file_i/rf_reg_392_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_393__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0324_ ),
    .Q_N(\register_file_i/_3709_ ),
    .Q(\register_file_i/rf_reg_393_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_394__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0325_ ),
    .Q_N(\register_file_i/_3708_ ),
    .Q(\register_file_i/rf_reg_394_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_395__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0326_ ),
    .Q_N(\register_file_i/_3707_ ),
    .Q(\register_file_i/rf_reg_395_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_396__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2119),
    .D(\register_file_i/_0327_ ),
    .Q_N(\register_file_i/_3706_ ),
    .Q(\register_file_i/rf_reg_396_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_397__reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(net2199),
    .D(\register_file_i/_0328_ ),
    .Q_N(\register_file_i/_3705_ ),
    .Q(\register_file_i/rf_reg_397_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_398__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2199),
    .D(\register_file_i/_0329_ ),
    .Q_N(\register_file_i/_3704_ ),
    .Q(\register_file_i/rf_reg_398_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_399__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0330_ ),
    .Q_N(\register_file_i/_3703_ ),
    .Q(\register_file_i/rf_reg_399_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_39__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0331_ ),
    .Q_N(\register_file_i/_3702_ ),
    .Q(\register_file_i/rf_reg_39_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_400__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0332_ ),
    .Q_N(\register_file_i/_3701_ ),
    .Q(\register_file_i/rf_reg_400_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_401__reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0333_ ),
    .Q_N(\register_file_i/_3700_ ),
    .Q(\register_file_i/rf_reg_401_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_402__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0334_ ),
    .Q_N(\register_file_i/_3699_ ),
    .Q(\register_file_i/rf_reg_402_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_403__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0335_ ),
    .Q_N(\register_file_i/_3698_ ),
    .Q(\register_file_i/rf_reg_403_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_404__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0336_ ),
    .Q_N(\register_file_i/_3697_ ),
    .Q(\register_file_i/rf_reg_404_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_405__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0337_ ),
    .Q_N(\register_file_i/_3696_ ),
    .Q(\register_file_i/rf_reg_405_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_406__reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0338_ ),
    .Q_N(\register_file_i/_3695_ ),
    .Q(\register_file_i/rf_reg_406_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_407__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0339_ ),
    .Q_N(\register_file_i/_3694_ ),
    .Q(\register_file_i/rf_reg_407_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_408__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0340_ ),
    .Q_N(\register_file_i/_3693_ ),
    .Q(\register_file_i/rf_reg_408_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_409__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0341_ ),
    .Q_N(\register_file_i/_3692_ ),
    .Q(\register_file_i/rf_reg_409_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_40__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0342_ ),
    .Q_N(\register_file_i/_3691_ ),
    .Q(\register_file_i/rf_reg_40_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_410__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2135),
    .D(\register_file_i/_0343_ ),
    .Q_N(\register_file_i/_3690_ ),
    .Q(\register_file_i/rf_reg_410_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_411__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0344_ ),
    .Q_N(\register_file_i/_3689_ ),
    .Q(\register_file_i/rf_reg_411_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_412__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0345_ ),
    .Q_N(\register_file_i/_3688_ ),
    .Q(\register_file_i/rf_reg_412_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_413__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0346_ ),
    .Q_N(\register_file_i/_3687_ ),
    .Q(\register_file_i/rf_reg_413_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_414__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0347_ ),
    .Q_N(\register_file_i/_3686_ ),
    .Q(\register_file_i/rf_reg_414_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_415__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2226),
    .D(\register_file_i/_0348_ ),
    .Q_N(\register_file_i/_3685_ ),
    .Q(\register_file_i/rf_reg_415_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_416__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0349_ ),
    .Q_N(\register_file_i/_3684_ ),
    .Q(\register_file_i/rf_reg_416_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_417__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0350_ ),
    .Q_N(\register_file_i/_3683_ ),
    .Q(\register_file_i/rf_reg_417_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_418__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0351_ ),
    .Q_N(\register_file_i/_3682_ ),
    .Q(\register_file_i/rf_reg_418_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_419__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0352_ ),
    .Q_N(\register_file_i/_3681_ ),
    .Q(\register_file_i/rf_reg_419_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_41__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net2174),
    .D(\register_file_i/_0353_ ),
    .Q_N(\register_file_i/_3680_ ),
    .Q(\register_file_i/rf_reg_41_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_420__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0354_ ),
    .Q_N(\register_file_i/_3679_ ),
    .Q(\register_file_i/rf_reg_420_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_421__reg  (.CLK(clknet_leaf_342_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0355_ ),
    .Q_N(\register_file_i/_3678_ ),
    .Q(\register_file_i/rf_reg_421_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_422__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0356_ ),
    .Q_N(\register_file_i/_3677_ ),
    .Q(\register_file_i/rf_reg_422_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_423__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0357_ ),
    .Q_N(\register_file_i/_3676_ ),
    .Q(\register_file_i/rf_reg_423_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_424__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0358_ ),
    .Q_N(\register_file_i/_3675_ ),
    .Q(\register_file_i/rf_reg_424_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_425__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0359_ ),
    .Q_N(\register_file_i/_3674_ ),
    .Q(\register_file_i/rf_reg_425_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_426__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0360_ ),
    .Q_N(\register_file_i/_3673_ ),
    .Q(\register_file_i/rf_reg_426_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_427__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0361_ ),
    .Q_N(\register_file_i/_3672_ ),
    .Q(\register_file_i/rf_reg_427_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_428__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2119),
    .D(\register_file_i/_0362_ ),
    .Q_N(\register_file_i/_3671_ ),
    .Q(\register_file_i/rf_reg_428_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_429__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0363_ ),
    .Q_N(\register_file_i/_3670_ ),
    .Q(\register_file_i/rf_reg_429_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_42__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net2174),
    .D(\register_file_i/_0364_ ),
    .Q_N(\register_file_i/_3669_ ),
    .Q(\register_file_i/rf_reg_42_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_430__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0365_ ),
    .Q_N(\register_file_i/_3668_ ),
    .Q(\register_file_i/rf_reg_430_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_431__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2199),
    .D(\register_file_i/_0366_ ),
    .Q_N(\register_file_i/_3667_ ),
    .Q(\register_file_i/rf_reg_431_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_432__reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0367_ ),
    .Q_N(\register_file_i/_3666_ ),
    .Q(\register_file_i/rf_reg_432_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_433__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0368_ ),
    .Q_N(\register_file_i/_3665_ ),
    .Q(\register_file_i/rf_reg_433_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_434__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2203),
    .D(\register_file_i/_0369_ ),
    .Q_N(\register_file_i/_3664_ ),
    .Q(\register_file_i/rf_reg_434_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_435__reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0370_ ),
    .Q_N(\register_file_i/_3663_ ),
    .Q(\register_file_i/rf_reg_435_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_436__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2349),
    .D(\register_file_i/_0371_ ),
    .Q_N(\register_file_i/_3662_ ),
    .Q(\register_file_i/rf_reg_436_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_437__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2224),
    .D(\register_file_i/_0372_ ),
    .Q_N(\register_file_i/_3661_ ),
    .Q(\register_file_i/rf_reg_437_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_438__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0373_ ),
    .Q_N(\register_file_i/_3660_ ),
    .Q(\register_file_i/rf_reg_438_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_439__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0374_ ),
    .Q_N(\register_file_i/_3659_ ),
    .Q(\register_file_i/rf_reg_439_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_43__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0375_ ),
    .Q_N(\register_file_i/_3658_ ),
    .Q(\register_file_i/rf_reg_43_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_440__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0376_ ),
    .Q_N(\register_file_i/_3657_ ),
    .Q(\register_file_i/rf_reg_440_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_441__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0377_ ),
    .Q_N(\register_file_i/_3656_ ),
    .Q(\register_file_i/rf_reg_441_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_442__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2135),
    .D(\register_file_i/_0378_ ),
    .Q_N(\register_file_i/_3655_ ),
    .Q(\register_file_i/rf_reg_442_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_443__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2139),
    .D(\register_file_i/_0379_ ),
    .Q_N(\register_file_i/_3654_ ),
    .Q(\register_file_i/rf_reg_443_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_444__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0380_ ),
    .Q_N(\register_file_i/_3653_ ),
    .Q(\register_file_i/rf_reg_444_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_445__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0381_ ),
    .Q_N(\register_file_i/_3652_ ),
    .Q(\register_file_i/rf_reg_445_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_446__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2349),
    .D(\register_file_i/_0382_ ),
    .Q_N(\register_file_i/_3651_ ),
    .Q(\register_file_i/rf_reg_446_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_447__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2226),
    .D(\register_file_i/_0383_ ),
    .Q_N(\register_file_i/_3650_ ),
    .Q(\register_file_i/rf_reg_447_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_448__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0384_ ),
    .Q_N(\register_file_i/_3649_ ),
    .Q(\register_file_i/rf_reg_448_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_449__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0385_ ),
    .Q_N(\register_file_i/_3648_ ),
    .Q(\register_file_i/rf_reg_449_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_44__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0386_ ),
    .Q_N(\register_file_i/_3647_ ),
    .Q(\register_file_i/rf_reg_44_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_450__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0387_ ),
    .Q_N(\register_file_i/_3646_ ),
    .Q(\register_file_i/rf_reg_450_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_451__reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0388_ ),
    .Q_N(\register_file_i/_3645_ ),
    .Q(\register_file_i/rf_reg_451_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_452__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0389_ ),
    .Q_N(\register_file_i/_3644_ ),
    .Q(\register_file_i/rf_reg_452_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_453__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0390_ ),
    .Q_N(\register_file_i/_3643_ ),
    .Q(\register_file_i/rf_reg_453_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_454__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0391_ ),
    .Q_N(\register_file_i/_3642_ ),
    .Q(\register_file_i/rf_reg_454_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_455__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0392_ ),
    .Q_N(\register_file_i/_3641_ ),
    .Q(\register_file_i/rf_reg_455_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_456__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0393_ ),
    .Q_N(\register_file_i/_3640_ ),
    .Q(\register_file_i/rf_reg_456_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_457__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0394_ ),
    .Q_N(\register_file_i/_3639_ ),
    .Q(\register_file_i/rf_reg_457_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_458__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0395_ ),
    .Q_N(\register_file_i/_3638_ ),
    .Q(\register_file_i/rf_reg_458_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_459__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0396_ ),
    .Q_N(\register_file_i/_3637_ ),
    .Q(\register_file_i/rf_reg_459_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_45__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0397_ ),
    .Q_N(\register_file_i/_3636_ ),
    .Q(\register_file_i/rf_reg_45_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_460__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2119),
    .D(\register_file_i/_0398_ ),
    .Q_N(\register_file_i/_3635_ ),
    .Q(\register_file_i/rf_reg_460_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_461__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0399_ ),
    .Q_N(\register_file_i/_3634_ ),
    .Q(\register_file_i/rf_reg_461_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_462__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0400_ ),
    .Q_N(\register_file_i/_3633_ ),
    .Q(\register_file_i/rf_reg_462_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_463__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2199),
    .D(\register_file_i/_0401_ ),
    .Q_N(\register_file_i/_3632_ ),
    .Q(\register_file_i/rf_reg_463_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_464__reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0402_ ),
    .Q_N(\register_file_i/_3631_ ),
    .Q(\register_file_i/rf_reg_464_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_465__reg  (.CLK(clknet_leaf_110_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0403_ ),
    .Q_N(\register_file_i/_3630_ ),
    .Q(\register_file_i/rf_reg_465_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_466__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0404_ ),
    .Q_N(\register_file_i/_3629_ ),
    .Q(\register_file_i/rf_reg_466_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_467__reg  (.CLK(clknet_leaf_116_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0405_ ),
    .Q_N(\register_file_i/_3628_ ),
    .Q(\register_file_i/rf_reg_467_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_468__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0406_ ),
    .Q_N(\register_file_i/_3627_ ),
    .Q(\register_file_i/rf_reg_468_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_469__reg  (.CLK(clknet_leaf_114_clk_i),
    .RESET_B(net2227),
    .D(\register_file_i/_0407_ ),
    .Q_N(\register_file_i/_3626_ ),
    .Q(\register_file_i/rf_reg_469_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_46__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0408_ ),
    .Q_N(\register_file_i/_3625_ ),
    .Q(\register_file_i/rf_reg_46_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_470__reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0409_ ),
    .Q_N(\register_file_i/_3624_ ),
    .Q(\register_file_i/rf_reg_470_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_471__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2211),
    .D(\register_file_i/_0410_ ),
    .Q_N(\register_file_i/_3623_ ),
    .Q(\register_file_i/rf_reg_471_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_472__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0411_ ),
    .Q_N(\register_file_i/_3622_ ),
    .Q(\register_file_i/rf_reg_472_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_473__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0412_ ),
    .Q_N(\register_file_i/_3621_ ),
    .Q(\register_file_i/rf_reg_473_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_474__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2135),
    .D(\register_file_i/_0413_ ),
    .Q_N(\register_file_i/_3620_ ),
    .Q(\register_file_i/rf_reg_474_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_475__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0414_ ),
    .Q_N(\register_file_i/_3619_ ),
    .Q(\register_file_i/rf_reg_475_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_476__reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0415_ ),
    .Q_N(\register_file_i/_3618_ ),
    .Q(\register_file_i/rf_reg_476_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_477__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0416_ ),
    .Q_N(\register_file_i/_3617_ ),
    .Q(\register_file_i/rf_reg_477_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_478__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0417_ ),
    .Q_N(\register_file_i/_3616_ ),
    .Q(\register_file_i/rf_reg_478_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_479__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2226),
    .D(\register_file_i/_0418_ ),
    .Q_N(\register_file_i/_3615_ ),
    .Q(\register_file_i/rf_reg_479_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_47__reg  (.CLK(clknet_leaf_163_clk_i),
    .RESET_B(net2249),
    .D(\register_file_i/_0419_ ),
    .Q_N(\register_file_i/_3614_ ),
    .Q(\register_file_i/rf_reg_47_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_480__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0420_ ),
    .Q_N(\register_file_i/_3613_ ),
    .Q(\register_file_i/rf_reg_480_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_481__reg  (.CLK(clknet_leaf_33_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0421_ ),
    .Q_N(\register_file_i/_3612_ ),
    .Q(\register_file_i/rf_reg_481_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_482__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0422_ ),
    .Q_N(\register_file_i/_3611_ ),
    .Q(\register_file_i/rf_reg_482_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_483__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0423_ ),
    .Q_N(\register_file_i/_3610_ ),
    .Q(\register_file_i/rf_reg_483_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_484__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0424_ ),
    .Q_N(\register_file_i/_3609_ ),
    .Q(\register_file_i/rf_reg_484_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_485__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0425_ ),
    .Q_N(\register_file_i/_3608_ ),
    .Q(\register_file_i/rf_reg_485_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_486__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2156),
    .D(\register_file_i/_0426_ ),
    .Q_N(\register_file_i/_3607_ ),
    .Q(\register_file_i/rf_reg_486_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_487__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net2127),
    .D(\register_file_i/_0427_ ),
    .Q_N(\register_file_i/_3606_ ),
    .Q(\register_file_i/rf_reg_487_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_488__reg  (.CLK(clknet_leaf_342_clk_i),
    .RESET_B(net2126),
    .D(\register_file_i/_0428_ ),
    .Q_N(\register_file_i/_3605_ ),
    .Q(\register_file_i/rf_reg_488_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_489__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net2124),
    .D(\register_file_i/_0429_ ),
    .Q_N(\register_file_i/_3604_ ),
    .Q(\register_file_i/rf_reg_489_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_48__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2249),
    .D(\register_file_i/_0430_ ),
    .Q_N(\register_file_i/_3603_ ),
    .Q(\register_file_i/rf_reg_48_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_490__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0431_ ),
    .Q_N(\register_file_i/_3602_ ),
    .Q(\register_file_i/rf_reg_490_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_491__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0432_ ),
    .Q_N(\register_file_i/_3601_ ),
    .Q(\register_file_i/rf_reg_491_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_492__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2117),
    .D(\register_file_i/_0433_ ),
    .Q_N(\register_file_i/_3600_ ),
    .Q(\register_file_i/rf_reg_492_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_493__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0434_ ),
    .Q_N(\register_file_i/_3599_ ),
    .Q(\register_file_i/rf_reg_493_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_494__reg  (.CLK(clknet_leaf_107_clk_i),
    .RESET_B(net2198),
    .D(\register_file_i/_0435_ ),
    .Q_N(\register_file_i/_3598_ ),
    .Q(\register_file_i/rf_reg_494_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_495__reg  (.CLK(clknet_leaf_106_clk_i),
    .RESET_B(net2199),
    .D(\register_file_i/_0436_ ),
    .Q_N(\register_file_i/_3597_ ),
    .Q(\register_file_i/rf_reg_495_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_496__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0437_ ),
    .Q_N(\register_file_i/_3596_ ),
    .Q(\register_file_i/rf_reg_496_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_497__reg  (.CLK(clknet_leaf_109_clk_i),
    .RESET_B(net2219),
    .D(\register_file_i/_0438_ ),
    .Q_N(\register_file_i/_3595_ ),
    .Q(\register_file_i/rf_reg_497_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_498__reg  (.CLK(clknet_leaf_108_clk_i),
    .RESET_B(net2204),
    .D(\register_file_i/_0439_ ),
    .Q_N(\register_file_i/_3594_ ),
    .Q(\register_file_i/rf_reg_498_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_499__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2220),
    .D(\register_file_i/_0440_ ),
    .Q_N(\register_file_i/_3593_ ),
    .Q(\register_file_i/rf_reg_499_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_49__reg  (.CLK(clknet_leaf_164_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0441_ ),
    .Q_N(\register_file_i/_3592_ ),
    .Q(\register_file_i/rf_reg_49_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_500__reg  (.CLK(clknet_leaf_118_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0442_ ),
    .Q_N(\register_file_i/_3591_ ),
    .Q(\register_file_i/rf_reg_500_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_501__reg  (.CLK(clknet_leaf_115_clk_i),
    .RESET_B(net2227),
    .D(\register_file_i/_0443_ ),
    .Q_N(\register_file_i/_3590_ ),
    .Q(\register_file_i/rf_reg_501_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_502__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0444_ ),
    .Q_N(\register_file_i/_3589_ ),
    .Q(\register_file_i/rf_reg_502_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_503__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net2211),
    .D(\register_file_i/_0445_ ),
    .Q_N(\register_file_i/_3588_ ),
    .Q(\register_file_i/rf_reg_503_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_504__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0446_ ),
    .Q_N(\register_file_i/_3587_ ),
    .Q(\register_file_i/rf_reg_504_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_505__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0447_ ),
    .Q_N(\register_file_i/_3586_ ),
    .Q(\register_file_i/rf_reg_505_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_506__reg  (.CLK(clknet_6_4_0_clk_i),
    .RESET_B(net2135),
    .D(\register_file_i/_0448_ ),
    .Q_N(\register_file_i/_3585_ ),
    .Q(\register_file_i/rf_reg_506_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_507__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net2140),
    .D(\register_file_i/_0449_ ),
    .Q_N(\register_file_i/_3584_ ),
    .Q(\register_file_i/rf_reg_507_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_508__reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0450_ ),
    .Q_N(\register_file_i/_3583_ ),
    .Q(\register_file_i/rf_reg_508_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_509__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net2122),
    .D(\register_file_i/_0451_ ),
    .Q_N(\register_file_i/_3582_ ),
    .Q(\register_file_i/rf_reg_509_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_50__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0452_ ),
    .Q_N(\register_file_i/_3581_ ),
    .Q(\register_file_i/rf_reg_50_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_510__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2234),
    .D(\register_file_i/_0453_ ),
    .Q_N(\register_file_i/_3580_ ),
    .Q(\register_file_i/rf_reg_510_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_511__reg  (.CLK(clknet_leaf_112_clk_i),
    .RESET_B(net2226),
    .D(\register_file_i/_0454_ ),
    .Q_N(\register_file_i/_3579_ ),
    .Q(\register_file_i/rf_reg_511_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_512__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0455_ ),
    .Q_N(\register_file_i/_3578_ ),
    .Q(\register_file_i/rf_reg_512_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_513__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0456_ ),
    .Q_N(\register_file_i/_3577_ ),
    .Q(\register_file_i/rf_reg_513_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_514__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0457_ ),
    .Q_N(\register_file_i/_3576_ ),
    .Q(\register_file_i/rf_reg_514_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_515__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0458_ ),
    .Q_N(\register_file_i/_3575_ ),
    .Q(\register_file_i/rf_reg_515_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_516__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0459_ ),
    .Q_N(\register_file_i/_3574_ ),
    .Q(\register_file_i/rf_reg_516_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_517__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0460_ ),
    .Q_N(\register_file_i/_3573_ ),
    .Q(\register_file_i/rf_reg_517_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_518__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2162),
    .D(\register_file_i/_0461_ ),
    .Q_N(\register_file_i/_3572_ ),
    .Q(\register_file_i/rf_reg_518_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_519__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2132),
    .D(\register_file_i/_0462_ ),
    .Q_N(\register_file_i/_3571_ ),
    .Q(\register_file_i/rf_reg_519_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_51__reg  (.CLK(clknet_leaf_164_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0463_ ),
    .Q_N(\register_file_i/_3570_ ),
    .Q(\register_file_i/rf_reg_51_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_520__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0464_ ),
    .Q_N(\register_file_i/_3569_ ),
    .Q(\register_file_i/rf_reg_520_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_521__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0465_ ),
    .Q_N(\register_file_i/_3568_ ),
    .Q(\register_file_i/rf_reg_521_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_522__reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0466_ ),
    .Q_N(\register_file_i/_3567_ ),
    .Q(\register_file_i/rf_reg_522_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_523__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0467_ ),
    .Q_N(\register_file_i/_3566_ ),
    .Q(\register_file_i/rf_reg_523_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_524__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2134),
    .D(\register_file_i/_0468_ ),
    .Q_N(\register_file_i/_3565_ ),
    .Q(\register_file_i/rf_reg_524_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_525__reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0469_ ),
    .Q_N(\register_file_i/_3564_ ),
    .Q(\register_file_i/rf_reg_525_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_526__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0470_ ),
    .Q_N(\register_file_i/_3563_ ),
    .Q(\register_file_i/rf_reg_526_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_527__reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0471_ ),
    .Q_N(\register_file_i/_3562_ ),
    .Q(\register_file_i/rf_reg_527_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_528__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0472_ ),
    .Q_N(\register_file_i/_3561_ ),
    .Q(\register_file_i/rf_reg_528_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_529__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0473_ ),
    .Q_N(\register_file_i/_3560_ ),
    .Q(\register_file_i/rf_reg_529_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_52__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0474_ ),
    .Q_N(\register_file_i/_3559_ ),
    .Q(\register_file_i/rf_reg_52_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_530__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0475_ ),
    .Q_N(\register_file_i/_3558_ ),
    .Q(\register_file_i/rf_reg_530_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_531__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0476_ ),
    .Q_N(\register_file_i/_3557_ ),
    .Q(\register_file_i/rf_reg_531_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_532__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0477_ ),
    .Q_N(\register_file_i/_3556_ ),
    .Q(\register_file_i/rf_reg_532_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_533__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0478_ ),
    .Q_N(\register_file_i/_3555_ ),
    .Q(\register_file_i/rf_reg_533_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_534__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0479_ ),
    .Q_N(\register_file_i/_3554_ ),
    .Q(\register_file_i/rf_reg_534_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_535__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0480_ ),
    .Q_N(\register_file_i/_3553_ ),
    .Q(\register_file_i/rf_reg_535_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_536__reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0481_ ),
    .Q_N(\register_file_i/_3552_ ),
    .Q(\register_file_i/rf_reg_536_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_537__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0482_ ),
    .Q_N(\register_file_i/_3551_ ),
    .Q(\register_file_i/rf_reg_537_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_538__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0483_ ),
    .Q_N(\register_file_i/_3550_ ),
    .Q(\register_file_i/rf_reg_538_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_539__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0484_ ),
    .Q_N(\register_file_i/_3549_ ),
    .Q(\register_file_i/rf_reg_539_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_53__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0485_ ),
    .Q_N(\register_file_i/_3548_ ),
    .Q(\register_file_i/rf_reg_53_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_540__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0486_ ),
    .Q_N(\register_file_i/_3547_ ),
    .Q(\register_file_i/rf_reg_540_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_541__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0487_ ),
    .Q_N(\register_file_i/_3546_ ),
    .Q(\register_file_i/rf_reg_541_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_542__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0488_ ),
    .Q_N(\register_file_i/_3545_ ),
    .Q(\register_file_i/rf_reg_542_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_543__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0489_ ),
    .Q_N(\register_file_i/_3544_ ),
    .Q(\register_file_i/rf_reg_543_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_544__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0490_ ),
    .Q_N(\register_file_i/_3543_ ),
    .Q(\register_file_i/rf_reg_544_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_545__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0491_ ),
    .Q_N(\register_file_i/_3542_ ),
    .Q(\register_file_i/rf_reg_545_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_546__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0492_ ),
    .Q_N(\register_file_i/_3541_ ),
    .Q(\register_file_i/rf_reg_546_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_547__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0493_ ),
    .Q_N(\register_file_i/_3540_ ),
    .Q(\register_file_i/rf_reg_547_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_548__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2162),
    .D(\register_file_i/_0494_ ),
    .Q_N(\register_file_i/_3539_ ),
    .Q(\register_file_i/rf_reg_548_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_549__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0495_ ),
    .Q_N(\register_file_i/_3538_ ),
    .Q(\register_file_i/rf_reg_549_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_54__reg  (.CLK(clknet_leaf_169_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0496_ ),
    .Q_N(\register_file_i/_3537_ ),
    .Q(\register_file_i/rf_reg_54_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_550__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2162),
    .D(\register_file_i/_0497_ ),
    .Q_N(\register_file_i/_3536_ ),
    .Q(\register_file_i/rf_reg_550_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_551__reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net2132),
    .D(\register_file_i/_0498_ ),
    .Q_N(\register_file_i/_3535_ ),
    .Q(\register_file_i/rf_reg_551_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_552__reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net2132),
    .D(\register_file_i/_0499_ ),
    .Q_N(\register_file_i/_3534_ ),
    .Q(\register_file_i/rf_reg_552_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_553__reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0500_ ),
    .Q_N(\register_file_i/_3533_ ),
    .Q(\register_file_i/rf_reg_553_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_554__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0501_ ),
    .Q_N(\register_file_i/_3532_ ),
    .Q(\register_file_i/rf_reg_554_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_555__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0502_ ),
    .Q_N(\register_file_i/_3531_ ),
    .Q(\register_file_i/rf_reg_555_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_556__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0503_ ),
    .Q_N(\register_file_i/_3530_ ),
    .Q(\register_file_i/rf_reg_556_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_557__reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0504_ ),
    .Q_N(\register_file_i/_3529_ ),
    .Q(\register_file_i/rf_reg_557_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_558__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0505_ ),
    .Q_N(\register_file_i/_3528_ ),
    .Q(\register_file_i/rf_reg_558_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_559__reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0506_ ),
    .Q_N(\register_file_i/_3527_ ),
    .Q(\register_file_i/rf_reg_559_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_55__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0507_ ),
    .Q_N(\register_file_i/_3526_ ),
    .Q(\register_file_i/rf_reg_55_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_560__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0508_ ),
    .Q_N(\register_file_i/_3525_ ),
    .Q(\register_file_i/rf_reg_560_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_561__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0509_ ),
    .Q_N(\register_file_i/_3524_ ),
    .Q(\register_file_i/rf_reg_561_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_562__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0510_ ),
    .Q_N(\register_file_i/_3523_ ),
    .Q(\register_file_i/rf_reg_562_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_563__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0511_ ),
    .Q_N(\register_file_i/_3522_ ),
    .Q(\register_file_i/rf_reg_563_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_564__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0512_ ),
    .Q_N(\register_file_i/_3521_ ),
    .Q(\register_file_i/rf_reg_564_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_565__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0513_ ),
    .Q_N(\register_file_i/_3520_ ),
    .Q(\register_file_i/rf_reg_565_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_566__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0514_ ),
    .Q_N(\register_file_i/_3519_ ),
    .Q(\register_file_i/rf_reg_566_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_567__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0515_ ),
    .Q_N(\register_file_i/_3518_ ),
    .Q(\register_file_i/rf_reg_567_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_568__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0516_ ),
    .Q_N(\register_file_i/_3517_ ),
    .Q(\register_file_i/rf_reg_568_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_569__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0517_ ),
    .Q_N(\register_file_i/_3516_ ),
    .Q(\register_file_i/rf_reg_569_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_56__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0518_ ),
    .Q_N(\register_file_i/_3515_ ),
    .Q(\register_file_i/rf_reg_56_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_570__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0519_ ),
    .Q_N(\register_file_i/_3514_ ),
    .Q(\register_file_i/rf_reg_570_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_571__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0520_ ),
    .Q_N(\register_file_i/_3513_ ),
    .Q(\register_file_i/rf_reg_571_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_572__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0521_ ),
    .Q_N(\register_file_i/_3512_ ),
    .Q(\register_file_i/rf_reg_572_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_573__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0522_ ),
    .Q_N(\register_file_i/_3511_ ),
    .Q(\register_file_i/rf_reg_573_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_574__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0523_ ),
    .Q_N(\register_file_i/_3510_ ),
    .Q(\register_file_i/rf_reg_574_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_575__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0524_ ),
    .Q_N(\register_file_i/_3509_ ),
    .Q(\register_file_i/rf_reg_575_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_576__reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0525_ ),
    .Q_N(\register_file_i/_3508_ ),
    .Q(\register_file_i/rf_reg_576_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_577__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0526_ ),
    .Q_N(\register_file_i/_3507_ ),
    .Q(\register_file_i/rf_reg_577_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_578__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0527_ ),
    .Q_N(\register_file_i/_3506_ ),
    .Q(\register_file_i/rf_reg_578_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_579__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0528_ ),
    .Q_N(\register_file_i/_3505_ ),
    .Q(\register_file_i/rf_reg_579_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_57__reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0529_ ),
    .Q_N(\register_file_i/_3504_ ),
    .Q(\register_file_i/rf_reg_57_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_580__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0530_ ),
    .Q_N(\register_file_i/_3503_ ),
    .Q(\register_file_i/rf_reg_580_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_581__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0531_ ),
    .Q_N(\register_file_i/_3502_ ),
    .Q(\register_file_i/rf_reg_581_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_582__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0532_ ),
    .Q_N(\register_file_i/_3501_ ),
    .Q(\register_file_i/rf_reg_582_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_583__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0533_ ),
    .Q_N(\register_file_i/_3500_ ),
    .Q(\register_file_i/rf_reg_583_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_584__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0534_ ),
    .Q_N(\register_file_i/_3499_ ),
    .Q(\register_file_i/rf_reg_584_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_585__reg  (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0535_ ),
    .Q_N(\register_file_i/_3498_ ),
    .Q(\register_file_i/rf_reg_585_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_586__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0536_ ),
    .Q_N(\register_file_i/_3497_ ),
    .Q(\register_file_i/rf_reg_586_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_587__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0537_ ),
    .Q_N(\register_file_i/_3496_ ),
    .Q(\register_file_i/rf_reg_587_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_588__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0538_ ),
    .Q_N(\register_file_i/_3495_ ),
    .Q(\register_file_i/rf_reg_588_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_589__reg  (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0539_ ),
    .Q_N(\register_file_i/_3494_ ),
    .Q(\register_file_i/rf_reg_589_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_58__reg  (.CLK(clknet_leaf_54_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0540_ ),
    .Q_N(\register_file_i/_3493_ ),
    .Q(\register_file_i/rf_reg_58_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_590__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0541_ ),
    .Q_N(\register_file_i/_3492_ ),
    .Q(\register_file_i/rf_reg_590_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_591__reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0542_ ),
    .Q_N(\register_file_i/_3491_ ),
    .Q(\register_file_i/rf_reg_591_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_592__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0543_ ),
    .Q_N(\register_file_i/_3490_ ),
    .Q(\register_file_i/rf_reg_592_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_593__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0544_ ),
    .Q_N(\register_file_i/_3489_ ),
    .Q(\register_file_i/rf_reg_593_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_594__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0545_ ),
    .Q_N(\register_file_i/_3488_ ),
    .Q(\register_file_i/rf_reg_594_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_595__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0546_ ),
    .Q_N(\register_file_i/_3487_ ),
    .Q(\register_file_i/rf_reg_595_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_596__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0547_ ),
    .Q_N(\register_file_i/_3486_ ),
    .Q(\register_file_i/rf_reg_596_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_597__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0548_ ),
    .Q_N(\register_file_i/_3485_ ),
    .Q(\register_file_i/rf_reg_597_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_598__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0549_ ),
    .Q_N(\register_file_i/_3484_ ),
    .Q(\register_file_i/rf_reg_598_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_599__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2216),
    .D(\register_file_i/_0550_ ),
    .Q_N(\register_file_i/_3483_ ),
    .Q(\register_file_i/rf_reg_599_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_59__reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0551_ ),
    .Q_N(\register_file_i/_3482_ ),
    .Q(\register_file_i/rf_reg_59_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_600__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0552_ ),
    .Q_N(\register_file_i/_3481_ ),
    .Q(\register_file_i/rf_reg_600_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_601__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0553_ ),
    .Q_N(\register_file_i/_3480_ ),
    .Q(\register_file_i/rf_reg_601_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_602__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0554_ ),
    .Q_N(\register_file_i/_3479_ ),
    .Q(\register_file_i/rf_reg_602_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_603__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0555_ ),
    .Q_N(\register_file_i/_3478_ ),
    .Q(\register_file_i/rf_reg_603_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_604__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0556_ ),
    .Q_N(\register_file_i/_3477_ ),
    .Q(\register_file_i/rf_reg_604_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_605__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0557_ ),
    .Q_N(\register_file_i/_3476_ ),
    .Q(\register_file_i/rf_reg_605_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_606__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0558_ ),
    .Q_N(\register_file_i/_3475_ ),
    .Q(\register_file_i/rf_reg_606_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_607__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0559_ ),
    .Q_N(\register_file_i/_3474_ ),
    .Q(\register_file_i/rf_reg_607_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_608__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0560_ ),
    .Q_N(\register_file_i/_3473_ ),
    .Q(\register_file_i/rf_reg_608_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_609__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0561_ ),
    .Q_N(\register_file_i/_3472_ ),
    .Q(\register_file_i/rf_reg_609_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_60__reg  (.CLK(clknet_leaf_300_clk_i),
    .RESET_B(net2299),
    .D(\register_file_i/_0562_ ),
    .Q_N(\register_file_i/_3471_ ),
    .Q(\register_file_i/rf_reg_60_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_610__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0563_ ),
    .Q_N(\register_file_i/_3470_ ),
    .Q(\register_file_i/rf_reg_610_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_611__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0564_ ),
    .Q_N(\register_file_i/_3469_ ),
    .Q(\register_file_i/rf_reg_611_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_612__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0565_ ),
    .Q_N(\register_file_i/_3468_ ),
    .Q(\register_file_i/rf_reg_612_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_613__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0566_ ),
    .Q_N(\register_file_i/_3467_ ),
    .Q(\register_file_i/rf_reg_613_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_614__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2177),
    .D(\register_file_i/_0567_ ),
    .Q_N(\register_file_i/_3466_ ),
    .Q(\register_file_i/rf_reg_614_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_615__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0568_ ),
    .Q_N(\register_file_i/_3465_ ),
    .Q(\register_file_i/rf_reg_615_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_616__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0569_ ),
    .Q_N(\register_file_i/_3464_ ),
    .Q(\register_file_i/rf_reg_616_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_617__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0570_ ),
    .Q_N(\register_file_i/_3463_ ),
    .Q(\register_file_i/rf_reg_617_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_618__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0571_ ),
    .Q_N(\register_file_i/_3462_ ),
    .Q(\register_file_i/rf_reg_618_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_619__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0572_ ),
    .Q_N(\register_file_i/_3461_ ),
    .Q(\register_file_i/rf_reg_619_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_61__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0573_ ),
    .Q_N(\register_file_i/_3460_ ),
    .Q(\register_file_i/rf_reg_61_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_620__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0574_ ),
    .Q_N(\register_file_i/_3459_ ),
    .Q(\register_file_i/rf_reg_620_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_621__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0575_ ),
    .Q_N(\register_file_i/_3458_ ),
    .Q(\register_file_i/rf_reg_621_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_622__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0576_ ),
    .Q_N(\register_file_i/_3457_ ),
    .Q(\register_file_i/rf_reg_622_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_623__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0577_ ),
    .Q_N(\register_file_i/_3456_ ),
    .Q(\register_file_i/rf_reg_623_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_624__reg  (.CLK(clknet_leaf_105_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0578_ ),
    .Q_N(\register_file_i/_3455_ ),
    .Q(\register_file_i/rf_reg_624_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_625__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0579_ ),
    .Q_N(\register_file_i/_3454_ ),
    .Q(\register_file_i/rf_reg_625_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_626__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0580_ ),
    .Q_N(\register_file_i/_3453_ ),
    .Q(\register_file_i/rf_reg_626_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_627__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0581_ ),
    .Q_N(\register_file_i/_3452_ ),
    .Q(\register_file_i/rf_reg_627_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_628__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0582_ ),
    .Q_N(\register_file_i/_3451_ ),
    .Q(\register_file_i/rf_reg_628_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_629__reg  (.CLK(clknet_leaf_119_clk_i),
    .RESET_B(net2225),
    .D(\register_file_i/_0583_ ),
    .Q_N(\register_file_i/_3450_ ),
    .Q(\register_file_i/rf_reg_629_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_62__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2255),
    .D(\register_file_i/_0584_ ),
    .Q_N(\register_file_i/_3449_ ),
    .Q(\register_file_i/rf_reg_62_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_630__reg  (.CLK(clknet_leaf_120_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0585_ ),
    .Q_N(\register_file_i/_3448_ ),
    .Q(\register_file_i/rf_reg_630_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_631__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0586_ ),
    .Q_N(\register_file_i/_3447_ ),
    .Q(\register_file_i/rf_reg_631_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_632__reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0587_ ),
    .Q_N(\register_file_i/_3446_ ),
    .Q(\register_file_i/rf_reg_632_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_633__reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0588_ ),
    .Q_N(\register_file_i/_3445_ ),
    .Q(\register_file_i/rf_reg_633_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_634__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0589_ ),
    .Q_N(\register_file_i/_3444_ ),
    .Q(\register_file_i/rf_reg_634_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_635__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0590_ ),
    .Q_N(\register_file_i/_3443_ ),
    .Q(\register_file_i/rf_reg_635_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_636__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0591_ ),
    .Q_N(\register_file_i/_3442_ ),
    .Q(\register_file_i/rf_reg_636_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_637__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0592_ ),
    .Q_N(\register_file_i/_3441_ ),
    .Q(\register_file_i/rf_reg_637_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_638__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2216),
    .D(\register_file_i/_0593_ ),
    .Q_N(\register_file_i/_3440_ ),
    .Q(\register_file_i/rf_reg_638_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_639__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2233),
    .D(\register_file_i/_0594_ ),
    .Q_N(\register_file_i/_3439_ ),
    .Q(\register_file_i/rf_reg_639_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_63__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2254),
    .D(\register_file_i/_0595_ ),
    .Q_N(\register_file_i/_3438_ ),
    .Q(\register_file_i/rf_reg_63_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_640__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0596_ ),
    .Q_N(\register_file_i/_3437_ ),
    .Q(\register_file_i/rf_reg_640_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_641__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0597_ ),
    .Q_N(\register_file_i/_3436_ ),
    .Q(\register_file_i/rf_reg_641_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_642__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0598_ ),
    .Q_N(\register_file_i/_3435_ ),
    .Q(\register_file_i/rf_reg_642_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_643__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0599_ ),
    .Q_N(\register_file_i/_3434_ ),
    .Q(\register_file_i/rf_reg_643_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_644__reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0600_ ),
    .Q_N(\register_file_i/_3433_ ),
    .Q(\register_file_i/rf_reg_644_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_645__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0601_ ),
    .Q_N(\register_file_i/_3432_ ),
    .Q(\register_file_i/rf_reg_645_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_646__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0602_ ),
    .Q_N(\register_file_i/_3431_ ),
    .Q(\register_file_i/rf_reg_646_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_647__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0603_ ),
    .Q_N(\register_file_i/_3430_ ),
    .Q(\register_file_i/rf_reg_647_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_648__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0604_ ),
    .Q_N(\register_file_i/_3429_ ),
    .Q(\register_file_i/rf_reg_648_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_649__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0605_ ),
    .Q_N(\register_file_i/_3428_ ),
    .Q(\register_file_i/rf_reg_649_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_64__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0606_ ),
    .Q_N(\register_file_i/_3427_ ),
    .Q(\register_file_i/rf_reg_64_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_650__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0607_ ),
    .Q_N(\register_file_i/_3426_ ),
    .Q(\register_file_i/rf_reg_650_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_651__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0608_ ),
    .Q_N(\register_file_i/_3425_ ),
    .Q(\register_file_i/rf_reg_651_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_652__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0609_ ),
    .Q_N(\register_file_i/_3424_ ),
    .Q(\register_file_i/rf_reg_652_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_653__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0610_ ),
    .Q_N(\register_file_i/_3423_ ),
    .Q(\register_file_i/rf_reg_653_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_654__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0611_ ),
    .Q_N(\register_file_i/_3422_ ),
    .Q(\register_file_i/rf_reg_654_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_655__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0612_ ),
    .Q_N(\register_file_i/_3421_ ),
    .Q(\register_file_i/rf_reg_655_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_656__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0613_ ),
    .Q_N(\register_file_i/_3420_ ),
    .Q(\register_file_i/rf_reg_656_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_657__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0614_ ),
    .Q_N(\register_file_i/_3419_ ),
    .Q(\register_file_i/rf_reg_657_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_658__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0615_ ),
    .Q_N(\register_file_i/_3418_ ),
    .Q(\register_file_i/rf_reg_658_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_659__reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0616_ ),
    .Q_N(\register_file_i/_3417_ ),
    .Q(\register_file_i/rf_reg_659_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_65__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0617_ ),
    .Q_N(\register_file_i/_3416_ ),
    .Q(\register_file_i/rf_reg_65_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_660__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0618_ ),
    .Q_N(\register_file_i/_3415_ ),
    .Q(\register_file_i/rf_reg_660_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_661__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0619_ ),
    .Q_N(\register_file_i/_3414_ ),
    .Q(\register_file_i/rf_reg_661_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_662__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0620_ ),
    .Q_N(\register_file_i/_3413_ ),
    .Q(\register_file_i/rf_reg_662_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_663__reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0621_ ),
    .Q_N(\register_file_i/_3412_ ),
    .Q(\register_file_i/rf_reg_663_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_664__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0622_ ),
    .Q_N(\register_file_i/_3411_ ),
    .Q(\register_file_i/rf_reg_664_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_665__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0623_ ),
    .Q_N(\register_file_i/_3410_ ),
    .Q(\register_file_i/rf_reg_665_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_666__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0624_ ),
    .Q_N(\register_file_i/_3409_ ),
    .Q(\register_file_i/rf_reg_666_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_667__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0625_ ),
    .Q_N(\register_file_i/_3408_ ),
    .Q(\register_file_i/rf_reg_667_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_668__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0626_ ),
    .Q_N(\register_file_i/_3407_ ),
    .Q(\register_file_i/rf_reg_668_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_669__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0627_ ),
    .Q_N(\register_file_i/_3406_ ),
    .Q(\register_file_i/rf_reg_669_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_66__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0628_ ),
    .Q_N(\register_file_i/_3405_ ),
    .Q(\register_file_i/rf_reg_66_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_670__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0629_ ),
    .Q_N(\register_file_i/_3404_ ),
    .Q(\register_file_i/rf_reg_670_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_671__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0630_ ),
    .Q_N(\register_file_i/_3403_ ),
    .Q(\register_file_i/rf_reg_671_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_672__reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0631_ ),
    .Q_N(\register_file_i/_3402_ ),
    .Q(\register_file_i/rf_reg_672_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_673__reg  (.CLK(clknet_leaf_30_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0632_ ),
    .Q_N(\register_file_i/_3401_ ),
    .Q(\register_file_i/rf_reg_673_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_674__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0633_ ),
    .Q_N(\register_file_i/_3400_ ),
    .Q(\register_file_i/rf_reg_674_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_675__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net2164),
    .D(\register_file_i/_0634_ ),
    .Q_N(\register_file_i/_3399_ ),
    .Q(\register_file_i/rf_reg_675_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_676__reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0635_ ),
    .Q_N(\register_file_i/_3398_ ),
    .Q(\register_file_i/rf_reg_676_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_677__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0636_ ),
    .Q_N(\register_file_i/_3397_ ),
    .Q(\register_file_i/rf_reg_677_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_678__reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net2162),
    .D(\register_file_i/_0637_ ),
    .Q_N(\register_file_i/_3396_ ),
    .Q(\register_file_i/rf_reg_678_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_679__reg  (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net2132),
    .D(\register_file_i/_0638_ ),
    .Q_N(\register_file_i/_3395_ ),
    .Q(\register_file_i/rf_reg_679_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_67__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0639_ ),
    .Q_N(\register_file_i/_3394_ ),
    .Q(\register_file_i/rf_reg_67_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_680__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2132),
    .D(\register_file_i/_0640_ ),
    .Q_N(\register_file_i/_3393_ ),
    .Q(\register_file_i/rf_reg_680_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_681__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2130),
    .D(\register_file_i/_0641_ ),
    .Q_N(\register_file_i/_3392_ ),
    .Q(\register_file_i/rf_reg_681_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_682__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0642_ ),
    .Q_N(\register_file_i/_3391_ ),
    .Q(\register_file_i/rf_reg_682_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_683__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0643_ ),
    .Q_N(\register_file_i/_3390_ ),
    .Q(\register_file_i/rf_reg_683_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_684__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0644_ ),
    .Q_N(\register_file_i/_3389_ ),
    .Q(\register_file_i/rf_reg_684_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_685__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2142),
    .D(\register_file_i/_0645_ ),
    .Q_N(\register_file_i/_3388_ ),
    .Q(\register_file_i/rf_reg_685_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_686__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0646_ ),
    .Q_N(\register_file_i/_3387_ ),
    .Q(\register_file_i/rf_reg_686_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_687__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0647_ ),
    .Q_N(\register_file_i/_3386_ ),
    .Q(\register_file_i/rf_reg_687_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_688__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0648_ ),
    .Q_N(\register_file_i/_3385_ ),
    .Q(\register_file_i/rf_reg_688_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_689__reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0649_ ),
    .Q_N(\register_file_i/_3384_ ),
    .Q(\register_file_i/rf_reg_689_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_68__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2283),
    .D(\register_file_i/_0650_ ),
    .Q_N(\register_file_i/_3383_ ),
    .Q(\register_file_i/rf_reg_68_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_690__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0651_ ),
    .Q_N(\register_file_i/_3382_ ),
    .Q(\register_file_i/rf_reg_690_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_691__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0652_ ),
    .Q_N(\register_file_i/_3381_ ),
    .Q(\register_file_i/rf_reg_691_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_692__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0653_ ),
    .Q_N(\register_file_i/_3380_ ),
    .Q(\register_file_i/rf_reg_692_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_693__reg  (.CLK(clknet_leaf_117_clk_i),
    .RESET_B(net2222),
    .D(\register_file_i/_0654_ ),
    .Q_N(\register_file_i/_3379_ ),
    .Q(\register_file_i/rf_reg_693_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_694__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0655_ ),
    .Q_N(\register_file_i/_3378_ ),
    .Q(\register_file_i/rf_reg_694_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_695__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0656_ ),
    .Q_N(\register_file_i/_3377_ ),
    .Q(\register_file_i/rf_reg_695_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_696__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0657_ ),
    .Q_N(\register_file_i/_3376_ ),
    .Q(\register_file_i/rf_reg_696_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_697__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2141),
    .D(\register_file_i/_0658_ ),
    .Q_N(\register_file_i/_3375_ ),
    .Q(\register_file_i/rf_reg_697_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_698__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0659_ ),
    .Q_N(\register_file_i/_3374_ ),
    .Q(\register_file_i/rf_reg_698_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_699__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0660_ ),
    .Q_N(\register_file_i/_3373_ ),
    .Q(\register_file_i/rf_reg_699_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_69__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0661_ ),
    .Q_N(\register_file_i/_3372_ ),
    .Q(\register_file_i/rf_reg_69_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_700__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0662_ ),
    .Q_N(\register_file_i/_3371_ ),
    .Q(\register_file_i/rf_reg_700_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_701__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0663_ ),
    .Q_N(\register_file_i/_3370_ ),
    .Q(\register_file_i/rf_reg_701_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_702__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2217),
    .D(\register_file_i/_0664_ ),
    .Q_N(\register_file_i/_3369_ ),
    .Q(\register_file_i/rf_reg_702_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_703__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0665_ ),
    .Q_N(\register_file_i/_3368_ ),
    .Q(\register_file_i/rf_reg_703_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_704__reg  (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0666_ ),
    .Q_N(\register_file_i/_3367_ ),
    .Q(\register_file_i/rf_reg_704_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_705__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0667_ ),
    .Q_N(\register_file_i/_3366_ ),
    .Q(\register_file_i/rf_reg_705_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_706__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net2180),
    .D(\register_file_i/_0668_ ),
    .Q_N(\register_file_i/_3365_ ),
    .Q(\register_file_i/rf_reg_706_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_707__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0669_ ),
    .Q_N(\register_file_i/_3364_ ),
    .Q(\register_file_i/rf_reg_707_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_708__reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0670_ ),
    .Q_N(\register_file_i/_3363_ ),
    .Q(\register_file_i/rf_reg_708_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_709__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0671_ ),
    .Q_N(\register_file_i/_3362_ ),
    .Q(\register_file_i/rf_reg_709_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_70__reg  (.CLK(clknet_leaf_308_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0672_ ),
    .Q_N(\register_file_i/_3361_ ),
    .Q(\register_file_i/rf_reg_70_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_710__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0673_ ),
    .Q_N(\register_file_i/_3360_ ),
    .Q(\register_file_i/rf_reg_710_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_711__reg  (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0674_ ),
    .Q_N(\register_file_i/_3359_ ),
    .Q(\register_file_i/rf_reg_711_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_712__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0675_ ),
    .Q_N(\register_file_i/_3358_ ),
    .Q(\register_file_i/rf_reg_712_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_713__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0676_ ),
    .Q_N(\register_file_i/_3357_ ),
    .Q(\register_file_i/rf_reg_713_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_714__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0677_ ),
    .Q_N(\register_file_i/_3356_ ),
    .Q(\register_file_i/rf_reg_714_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_715__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0678_ ),
    .Q_N(\register_file_i/_3355_ ),
    .Q(\register_file_i/rf_reg_715_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_716__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net2121),
    .D(\register_file_i/_0679_ ),
    .Q_N(\register_file_i/_3354_ ),
    .Q(\register_file_i/rf_reg_716_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_717__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2200),
    .D(\register_file_i/_0680_ ),
    .Q_N(\register_file_i/_3353_ ),
    .Q(\register_file_i/rf_reg_717_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_718__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0681_ ),
    .Q_N(\register_file_i/_3352_ ),
    .Q(\register_file_i/rf_reg_718_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_719__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net2201),
    .D(\register_file_i/_0682_ ),
    .Q_N(\register_file_i/_3351_ ),
    .Q(\register_file_i/rf_reg_719_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_71__reg  (.CLK(clknet_leaf_310_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0683_ ),
    .Q_N(\register_file_i/_3350_ ),
    .Q(\register_file_i/rf_reg_71_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_720__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net2206),
    .D(\register_file_i/_0684_ ),
    .Q_N(\register_file_i/_3349_ ),
    .Q(\register_file_i/rf_reg_720_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_721__reg  (.CLK(clknet_leaf_111_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0685_ ),
    .Q_N(\register_file_i/_3348_ ),
    .Q(\register_file_i/rf_reg_721_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_722__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2214),
    .D(\register_file_i/_0686_ ),
    .Q_N(\register_file_i/_3347_ ),
    .Q(\register_file_i/rf_reg_722_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_723__reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0687_ ),
    .Q_N(\register_file_i/_3346_ ),
    .Q(\register_file_i/rf_reg_723_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_724__reg  (.CLK(clknet_leaf_121_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0688_ ),
    .Q_N(\register_file_i/_3345_ ),
    .Q(\register_file_i/rf_reg_724_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_725__reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0689_ ),
    .Q_N(\register_file_i/_3344_ ),
    .Q(\register_file_i/rf_reg_725_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_726__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0690_ ),
    .Q_N(\register_file_i/_3343_ ),
    .Q(\register_file_i/rf_reg_726_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_727__reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0691_ ),
    .Q_N(\register_file_i/_3342_ ),
    .Q(\register_file_i/rf_reg_727_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_728__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0692_ ),
    .Q_N(\register_file_i/_3341_ ),
    .Q(\register_file_i/rf_reg_728_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_729__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0693_ ),
    .Q_N(\register_file_i/_3340_ ),
    .Q(\register_file_i/rf_reg_729_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_72__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0694_ ),
    .Q_N(\register_file_i/_3339_ ),
    .Q(\register_file_i/rf_reg_72_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_730__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0695_ ),
    .Q_N(\register_file_i/_3338_ ),
    .Q(\register_file_i/rf_reg_730_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_731__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0696_ ),
    .Q_N(\register_file_i/_3337_ ),
    .Q(\register_file_i/rf_reg_731_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_732__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0697_ ),
    .Q_N(\register_file_i/_3336_ ),
    .Q(\register_file_i/rf_reg_732_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_733__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0698_ ),
    .Q_N(\register_file_i/_3335_ ),
    .Q(\register_file_i/rf_reg_733_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_734__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0699_ ),
    .Q_N(\register_file_i/_3334_ ),
    .Q(\register_file_i/rf_reg_734_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_735__reg  (.CLK(clknet_leaf_125_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0700_ ),
    .Q_N(\register_file_i/_3333_ ),
    .Q(\register_file_i/rf_reg_735_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_736__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0701_ ),
    .Q_N(\register_file_i/_3332_ ),
    .Q(\register_file_i/rf_reg_736_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_737__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2148),
    .D(\register_file_i/_0702_ ),
    .Q_N(\register_file_i/_3331_ ),
    .Q(\register_file_i/rf_reg_737_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_738__reg  (.CLK(clknet_leaf_34_clk_i),
    .RESET_B(net2179),
    .D(\register_file_i/_0703_ ),
    .Q_N(\register_file_i/_3330_ ),
    .Q(\register_file_i/rf_reg_738_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_739__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0704_ ),
    .Q_N(\register_file_i/_3329_ ),
    .Q(\register_file_i/rf_reg_739_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_73__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net2174),
    .D(\register_file_i/_0705_ ),
    .Q_N(\register_file_i/_3328_ ),
    .Q(\register_file_i/rf_reg_73_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_740__reg  (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0706_ ),
    .Q_N(\register_file_i/_3327_ ),
    .Q(\register_file_i/rf_reg_740_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_741__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0707_ ),
    .Q_N(\register_file_i/_3326_ ),
    .Q(\register_file_i/rf_reg_741_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_742__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2161),
    .D(\register_file_i/_0708_ ),
    .Q_N(\register_file_i/_3325_ ),
    .Q(\register_file_i/rf_reg_742_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_743__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0709_ ),
    .Q_N(\register_file_i/_3324_ ),
    .Q(\register_file_i/rf_reg_743_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_744__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2131),
    .D(\register_file_i/_0710_ ),
    .Q_N(\register_file_i/_3323_ ),
    .Q(\register_file_i/rf_reg_744_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_745__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0711_ ),
    .Q_N(\register_file_i/_3322_ ),
    .Q(\register_file_i/rf_reg_745_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_746__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net2129),
    .D(\register_file_i/_0712_ ),
    .Q_N(\register_file_i/_3321_ ),
    .Q(\register_file_i/rf_reg_746_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_747__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net2120),
    .D(\register_file_i/_0713_ ),
    .Q_N(\register_file_i/_3320_ ),
    .Q(\register_file_i/rf_reg_747_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_748__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2136),
    .D(\register_file_i/_0714_ ),
    .Q_N(\register_file_i/_3319_ ),
    .Q(\register_file_i/rf_reg_748_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_749__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net2150),
    .D(\register_file_i/_0715_ ),
    .Q_N(\register_file_i/_3318_ ),
    .Q(\register_file_i/rf_reg_749_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_74__reg  (.CLK(clknet_leaf_38_clk_i),
    .RESET_B(net2172),
    .D(\register_file_i/_0716_ ),
    .Q_N(\register_file_i/_3317_ ),
    .Q(\register_file_i/rf_reg_74_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_750__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0717_ ),
    .Q_N(\register_file_i/_3316_ ),
    .Q(\register_file_i/rf_reg_750_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_751__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2209),
    .D(\register_file_i/_0718_ ),
    .Q_N(\register_file_i/_3315_ ),
    .Q(\register_file_i/rf_reg_751_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_752__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net2205),
    .D(\register_file_i/_0719_ ),
    .Q_N(\register_file_i/_3314_ ),
    .Q(\register_file_i/rf_reg_752_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_753__reg  (.CLK(clknet_leaf_124_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0720_ ),
    .Q_N(\register_file_i/_3313_ ),
    .Q(\register_file_i/rf_reg_753_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_754__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net2213),
    .D(\register_file_i/_0721_ ),
    .Q_N(\register_file_i/_3312_ ),
    .Q(\register_file_i/rf_reg_754_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_755__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2228),
    .D(\register_file_i/_0722_ ),
    .Q_N(\register_file_i/_3311_ ),
    .Q(\register_file_i/rf_reg_755_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_756__reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0723_ ),
    .Q_N(\register_file_i/_3310_ ),
    .Q(\register_file_i/rf_reg_756_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_757__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2221),
    .D(\register_file_i/_0724_ ),
    .Q_N(\register_file_i/_3309_ ),
    .Q(\register_file_i/rf_reg_757_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_758__reg  (.CLK(clknet_leaf_126_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0725_ ),
    .Q_N(\register_file_i/_3308_ ),
    .Q(\register_file_i/rf_reg_758_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_759__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0726_ ),
    .Q_N(\register_file_i/_3307_ ),
    .Q(\register_file_i/rf_reg_759_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_75__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net2174),
    .D(\register_file_i/_0727_ ),
    .Q_N(\register_file_i/_3306_ ),
    .Q(\register_file_i/rf_reg_75_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_760__reg  (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net2208),
    .D(\register_file_i/_0728_ ),
    .Q_N(\register_file_i/_3305_ ),
    .Q(\register_file_i/rf_reg_760_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_761__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2149),
    .D(\register_file_i/_0729_ ),
    .Q_N(\register_file_i/_3304_ ),
    .Q(\register_file_i/rf_reg_761_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_762__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net2144),
    .D(\register_file_i/_0730_ ),
    .Q_N(\register_file_i/_3303_ ),
    .Q(\register_file_i/rf_reg_762_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_763__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net2145),
    .D(\register_file_i/_0731_ ),
    .Q_N(\register_file_i/_3302_ ),
    .Q(\register_file_i/rf_reg_763_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_764__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0732_ ),
    .Q_N(\register_file_i/_3301_ ),
    .Q(\register_file_i/rf_reg_764_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_765__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net2137),
    .D(\register_file_i/_0733_ ),
    .Q_N(\register_file_i/_3300_ ),
    .Q(\register_file_i/rf_reg_765_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_766__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2216),
    .D(\register_file_i/_0734_ ),
    .Q_N(\register_file_i/_3299_ ),
    .Q(\register_file_i/rf_reg_766_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_767__reg  (.CLK(clknet_leaf_123_clk_i),
    .RESET_B(net2229),
    .D(\register_file_i/_0735_ ),
    .Q_N(\register_file_i/_3298_ ),
    .Q(\register_file_i/rf_reg_767_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_768__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0736_ ),
    .Q_N(\register_file_i/_3297_ ),
    .Q(\register_file_i/rf_reg_768_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_769__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2148),
    .D(\register_file_i/_0737_ ),
    .Q_N(\register_file_i/_3296_ ),
    .Q(\register_file_i/rf_reg_769_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_76__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net2189),
    .D(\register_file_i/_0738_ ),
    .Q_N(\register_file_i/_3295_ ),
    .Q(\register_file_i/rf_reg_76_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_770__reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0739_ ),
    .Q_N(\register_file_i/_3294_ ),
    .Q(\register_file_i/rf_reg_770_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_771__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0740_ ),
    .Q_N(\register_file_i/_3293_ ),
    .Q(\register_file_i/rf_reg_771_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_772__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0741_ ),
    .Q_N(\register_file_i/_3292_ ),
    .Q(\register_file_i/rf_reg_772_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_773__reg  (.CLK(clknet_leaf_311_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0742_ ),
    .Q_N(\register_file_i/_3291_ ),
    .Q(\register_file_i/rf_reg_773_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_774__reg  (.CLK(clknet_leaf_331_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0743_ ),
    .Q_N(\register_file_i/_3290_ ),
    .Q(\register_file_i/rf_reg_774_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_775__reg  (.CLK(clknet_leaf_334_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0744_ ),
    .Q_N(\register_file_i/_3289_ ),
    .Q(\register_file_i/rf_reg_775_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_776__reg  (.CLK(clknet_leaf_331_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0745_ ),
    .Q_N(\register_file_i/_3288_ ),
    .Q(\register_file_i/rf_reg_776_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_777__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0746_ ),
    .Q_N(\register_file_i/_3287_ ),
    .Q(\register_file_i/rf_reg_777_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_778__reg  (.CLK(clknet_leaf_337_clk_i),
    .RESET_B(net2170),
    .D(\register_file_i/_0747_ ),
    .Q_N(\register_file_i/_3286_ ),
    .Q(\register_file_i/rf_reg_778_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_779__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0748_ ),
    .Q_N(\register_file_i/_3285_ ),
    .Q(\register_file_i/rf_reg_779_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_77__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net2193),
    .D(\register_file_i/_0749_ ),
    .Q_N(\register_file_i/_3284_ ),
    .Q(\register_file_i/rf_reg_77_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_780__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0750_ ),
    .Q_N(\register_file_i/_3283_ ),
    .Q(\register_file_i/rf_reg_780_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_781__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0751_ ),
    .Q_N(\register_file_i/_3282_ ),
    .Q(\register_file_i/rf_reg_781_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_782__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0752_ ),
    .Q_N(\register_file_i/_3281_ ),
    .Q(\register_file_i/rf_reg_782_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_783__reg  (.CLK(clknet_leaf_157_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0753_ ),
    .Q_N(\register_file_i/_3280_ ),
    .Q(\register_file_i/rf_reg_783_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_784__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0754_ ),
    .Q_N(\register_file_i/_3279_ ),
    .Q(\register_file_i/rf_reg_784_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_785__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0755_ ),
    .Q_N(\register_file_i/_3278_ ),
    .Q(\register_file_i/rf_reg_785_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_786__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net2211),
    .D(\register_file_i/_0756_ ),
    .Q_N(\register_file_i/_3277_ ),
    .Q(\register_file_i/rf_reg_786_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_787__reg  (.CLK(clknet_leaf_134_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0757_ ),
    .Q_N(\register_file_i/_3276_ ),
    .Q(\register_file_i/rf_reg_787_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_788__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0758_ ),
    .Q_N(\register_file_i/_3275_ ),
    .Q(\register_file_i/rf_reg_788_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_789__reg  (.CLK(clknet_leaf_131_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0759_ ),
    .Q_N(\register_file_i/_3274_ ),
    .Q(\register_file_i/rf_reg_789_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_78__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2248),
    .D(\register_file_i/_0760_ ),
    .Q_N(\register_file_i/_3273_ ),
    .Q(\register_file_i/rf_reg_78_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_790__reg  (.CLK(clknet_leaf_169_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0761_ ),
    .Q_N(\register_file_i/_3272_ ),
    .Q(\register_file_i/rf_reg_790_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_791__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0762_ ),
    .Q_N(\register_file_i/_3271_ ),
    .Q(\register_file_i/rf_reg_791_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_792__reg  (.CLK(clknet_leaf_174_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0763_ ),
    .Q_N(\register_file_i/_3270_ ),
    .Q(\register_file_i/rf_reg_792_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_793__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0764_ ),
    .Q_N(\register_file_i/_3269_ ),
    .Q(\register_file_i/rf_reg_793_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_794__reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0765_ ),
    .Q_N(\register_file_i/_3268_ ),
    .Q(\register_file_i/rf_reg_794_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_795__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0766_ ),
    .Q_N(\register_file_i/_3267_ ),
    .Q(\register_file_i/rf_reg_795_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_796__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0767_ ),
    .Q_N(\register_file_i/_3266_ ),
    .Q(\register_file_i/rf_reg_796_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_797__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0768_ ),
    .Q_N(\register_file_i/_3265_ ),
    .Q(\register_file_i/rf_reg_797_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_798__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0769_ ),
    .Q_N(\register_file_i/_3264_ ),
    .Q(\register_file_i/rf_reg_798_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_799__reg  (.CLK(clknet_leaf_155_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0770_ ),
    .Q_N(\register_file_i/_3263_ ),
    .Q(\register_file_i/rf_reg_799_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_79__reg  (.CLK(clknet_leaf_162_clk_i),
    .RESET_B(net2249),
    .D(\register_file_i/_0771_ ),
    .Q_N(\register_file_i/_3262_ ),
    .Q(\register_file_i/rf_reg_79_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_800__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net2210),
    .D(\register_file_i/_0772_ ),
    .Q_N(\register_file_i/_3261_ ),
    .Q(\register_file_i/rf_reg_800_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_801__reg  (.CLK(clknet_leaf_80_clk_i),
    .RESET_B(net2146),
    .D(\register_file_i/_0773_ ),
    .Q_N(\register_file_i/_3260_ ),
    .Q(\register_file_i/rf_reg_801_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_802__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0774_ ),
    .Q_N(\register_file_i/_3259_ ),
    .Q(\register_file_i/rf_reg_802_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_803__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0775_ ),
    .Q_N(\register_file_i/_3258_ ),
    .Q(\register_file_i/rf_reg_803_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_804__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0776_ ),
    .Q_N(\register_file_i/_3257_ ),
    .Q(\register_file_i/rf_reg_804_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_805__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0777_ ),
    .Q_N(\register_file_i/_3256_ ),
    .Q(\register_file_i/rf_reg_805_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_806__reg  (.CLK(clknet_leaf_331_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0778_ ),
    .Q_N(\register_file_i/_3255_ ),
    .Q(\register_file_i/rf_reg_806_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_807__reg  (.CLK(clknet_leaf_334_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0779_ ),
    .Q_N(\register_file_i/_3254_ ),
    .Q(\register_file_i/rf_reg_807_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_808__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0780_ ),
    .Q_N(\register_file_i/_3253_ ),
    .Q(\register_file_i/rf_reg_808_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_809__reg  (.CLK(clknet_leaf_337_clk_i),
    .RESET_B(net2173),
    .D(\register_file_i/_0781_ ),
    .Q_N(\register_file_i/_3252_ ),
    .Q(\register_file_i/rf_reg_809_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_80__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0782_ ),
    .Q_N(\register_file_i/_3251_ ),
    .Q(\register_file_i/rf_reg_80_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_810__reg  (.CLK(clknet_leaf_337_clk_i),
    .RESET_B(net2170),
    .D(\register_file_i/_0783_ ),
    .Q_N(\register_file_i/_3250_ ),
    .Q(\register_file_i/rf_reg_810_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_811__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0784_ ),
    .Q_N(\register_file_i/_3249_ ),
    .Q(\register_file_i/rf_reg_811_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_812__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0785_ ),
    .Q_N(\register_file_i/_3248_ ),
    .Q(\register_file_i/rf_reg_812_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_813__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0786_ ),
    .Q_N(\register_file_i/_3247_ ),
    .Q(\register_file_i/rf_reg_813_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_814__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0787_ ),
    .Q_N(\register_file_i/_3246_ ),
    .Q(\register_file_i/rf_reg_814_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_815__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0788_ ),
    .Q_N(\register_file_i/_3245_ ),
    .Q(\register_file_i/rf_reg_815_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_816__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0789_ ),
    .Q_N(\register_file_i/_3244_ ),
    .Q(\register_file_i/rf_reg_816_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_817__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0790_ ),
    .Q_N(\register_file_i/_3243_ ),
    .Q(\register_file_i/rf_reg_817_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_818__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2211),
    .D(\register_file_i/_0791_ ),
    .Q_N(\register_file_i/_3242_ ),
    .Q(\register_file_i/rf_reg_818_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_819__reg  (.CLK(clknet_leaf_134_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0792_ ),
    .Q_N(\register_file_i/_3241_ ),
    .Q(\register_file_i/rf_reg_819_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_81__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0793_ ),
    .Q_N(\register_file_i/_3240_ ),
    .Q(\register_file_i/rf_reg_81_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_820__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0794_ ),
    .Q_N(\register_file_i/_3239_ ),
    .Q(\register_file_i/rf_reg_820_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_821__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0795_ ),
    .Q_N(\register_file_i/_3238_ ),
    .Q(\register_file_i/rf_reg_821_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_822__reg  (.CLK(clknet_leaf_169_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0796_ ),
    .Q_N(\register_file_i/_3237_ ),
    .Q(\register_file_i/rf_reg_822_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_823__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0797_ ),
    .Q_N(\register_file_i/_3236_ ),
    .Q(\register_file_i/rf_reg_823_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_824__reg  (.CLK(clknet_leaf_174_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0798_ ),
    .Q_N(\register_file_i/_3235_ ),
    .Q(\register_file_i/rf_reg_824_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_825__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0799_ ),
    .Q_N(\register_file_i/_3234_ ),
    .Q(\register_file_i/rf_reg_825_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_826__reg  (.CLK(clknet_leaf_62_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0800_ ),
    .Q_N(\register_file_i/_3233_ ),
    .Q(\register_file_i/rf_reg_826_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_827__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0801_ ),
    .Q_N(\register_file_i/_3232_ ),
    .Q(\register_file_i/rf_reg_827_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_828__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2283),
    .D(\register_file_i/_0802_ ),
    .Q_N(\register_file_i/_3231_ ),
    .Q(\register_file_i/rf_reg_828_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_829__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0803_ ),
    .Q_N(\register_file_i/_3230_ ),
    .Q(\register_file_i/rf_reg_829_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_82__reg  (.CLK(clknet_leaf_161_clk_i),
    .RESET_B(net2252),
    .D(\register_file_i/_0804_ ),
    .Q_N(\register_file_i/_3229_ ),
    .Q(\register_file_i/rf_reg_82_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_830__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2244),
    .D(\register_file_i/_0805_ ),
    .Q_N(\register_file_i/_3228_ ),
    .Q(\register_file_i/rf_reg_830_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_831__reg  (.CLK(clknet_leaf_155_clk_i),
    .RESET_B(net2260),
    .D(\register_file_i/_0806_ ),
    .Q_N(\register_file_i/_3227_ ),
    .Q(\register_file_i/rf_reg_831_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_832__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0807_ ),
    .Q_N(\register_file_i/_3226_ ),
    .Q(\register_file_i/rf_reg_832_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_833__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2178),
    .D(\register_file_i/_0808_ ),
    .Q_N(\register_file_i/_3225_ ),
    .Q(\register_file_i/rf_reg_833_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_834__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0809_ ),
    .Q_N(\register_file_i/_3224_ ),
    .Q(\register_file_i/rf_reg_834_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_835__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0810_ ),
    .Q_N(\register_file_i/_3223_ ),
    .Q(\register_file_i/rf_reg_835_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_836__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0811_ ),
    .Q_N(\register_file_i/_3222_ ),
    .Q(\register_file_i/rf_reg_836_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_837__reg  (.CLK(clknet_leaf_331_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0812_ ),
    .Q_N(\register_file_i/_3221_ ),
    .Q(\register_file_i/rf_reg_837_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_838__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0813_ ),
    .Q_N(\register_file_i/_3220_ ),
    .Q(\register_file_i/rf_reg_838_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_839__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0814_ ),
    .Q_N(\register_file_i/_3219_ ),
    .Q(\register_file_i/rf_reg_839_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_83__reg  (.CLK(clknet_leaf_153_clk_i),
    .RESET_B(net2267),
    .D(\register_file_i/_0815_ ),
    .Q_N(\register_file_i/_3218_ ),
    .Q(\register_file_i/rf_reg_83_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_840__reg  (.CLK(clknet_leaf_331_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0816_ ),
    .Q_N(\register_file_i/_3217_ ),
    .Q(\register_file_i/rf_reg_840_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_841__reg  (.CLK(clknet_leaf_336_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0817_ ),
    .Q_N(\register_file_i/_3216_ ),
    .Q(\register_file_i/rf_reg_841_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_842__reg  (.CLK(clknet_leaf_339_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0818_ ),
    .Q_N(\register_file_i/_3215_ ),
    .Q(\register_file_i/rf_reg_842_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_843__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0819_ ),
    .Q_N(\register_file_i/_3214_ ),
    .Q(\register_file_i/rf_reg_843_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_844__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0820_ ),
    .Q_N(\register_file_i/_3213_ ),
    .Q(\register_file_i/rf_reg_844_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_845__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0821_ ),
    .Q_N(\register_file_i/_3212_ ),
    .Q(\register_file_i/rf_reg_845_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_846__reg  (.CLK(clknet_leaf_159_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0822_ ),
    .Q_N(\register_file_i/_3211_ ),
    .Q(\register_file_i/rf_reg_846_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_847__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0823_ ),
    .Q_N(\register_file_i/_3210_ ),
    .Q(\register_file_i/rf_reg_847_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_848__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2244),
    .D(\register_file_i/_0824_ ),
    .Q_N(\register_file_i/_3209_ ),
    .Q(\register_file_i/rf_reg_848_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_849__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0825_ ),
    .Q_N(\register_file_i/_3208_ ),
    .Q(\register_file_i/rf_reg_849_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_84__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2255),
    .D(\register_file_i/_0826_ ),
    .Q_N(\register_file_i/_3207_ ),
    .Q(\register_file_i/rf_reg_84_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_850__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0827_ ),
    .Q_N(\register_file_i/_3206_ ),
    .Q(\register_file_i/rf_reg_850_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_851__reg  (.CLK(clknet_leaf_134_clk_i),
    .RESET_B(net2231),
    .D(\register_file_i/_0828_ ),
    .Q_N(\register_file_i/_3205_ ),
    .Q(\register_file_i/rf_reg_851_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_852__reg  (.CLK(clknet_leaf_131_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0829_ ),
    .Q_N(\register_file_i/_3204_ ),
    .Q(\register_file_i/rf_reg_852_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_853__reg  (.CLK(clknet_leaf_131_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0830_ ),
    .Q_N(\register_file_i/_3203_ ),
    .Q(\register_file_i/rf_reg_853_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_854__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2250),
    .D(\register_file_i/_0831_ ),
    .Q_N(\register_file_i/_3202_ ),
    .Q(\register_file_i/rf_reg_854_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_855__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2183),
    .D(\register_file_i/_0832_ ),
    .Q_N(\register_file_i/_3201_ ),
    .Q(\register_file_i/rf_reg_855_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_856__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0833_ ),
    .Q_N(\register_file_i/_3200_ ),
    .Q(\register_file_i/rf_reg_856_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_857__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2297),
    .D(\register_file_i/_0834_ ),
    .Q_N(\register_file_i/_3199_ ),
    .Q(\register_file_i/rf_reg_857_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_858__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2297),
    .D(\register_file_i/_0835_ ),
    .Q_N(\register_file_i/_3198_ ),
    .Q(\register_file_i/rf_reg_858_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_859__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0836_ ),
    .Q_N(\register_file_i/_3197_ ),
    .Q(\register_file_i/rf_reg_859_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_85__reg  (.CLK(clknet_leaf_165_clk_i),
    .RESET_B(net2256),
    .D(\register_file_i/_0837_ ),
    .Q_N(\register_file_i/_3196_ ),
    .Q(\register_file_i/rf_reg_85_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_860__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0838_ ),
    .Q_N(\register_file_i/_3195_ ),
    .Q(\register_file_i/rf_reg_860_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_861__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net2281),
    .D(\register_file_i/_0839_ ),
    .Q_N(\register_file_i/_3194_ ),
    .Q(\register_file_i/rf_reg_861_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_862__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0840_ ),
    .Q_N(\register_file_i/_3193_ ),
    .Q(\register_file_i/rf_reg_862_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_863__reg  (.CLK(clknet_leaf_155_clk_i),
    .RESET_B(net2260),
    .D(\register_file_i/_0841_ ),
    .Q_N(\register_file_i/_3192_ ),
    .Q(\register_file_i/rf_reg_863_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_864__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0842_ ),
    .Q_N(\register_file_i/_3191_ ),
    .Q(\register_file_i/rf_reg_864_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_865__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2181),
    .D(\register_file_i/_0843_ ),
    .Q_N(\register_file_i/_3190_ ),
    .Q(\register_file_i/rf_reg_865_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_866__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0844_ ),
    .Q_N(\register_file_i/_3189_ ),
    .Q(\register_file_i/rf_reg_866_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_867__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0845_ ),
    .Q_N(\register_file_i/_3188_ ),
    .Q(\register_file_i/rf_reg_867_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_868__reg  (.CLK(clknet_leaf_335_clk_i),
    .RESET_B(net2280),
    .D(\register_file_i/_0846_ ),
    .Q_N(\register_file_i/_3187_ ),
    .Q(\register_file_i/rf_reg_868_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_869__reg  (.CLK(clknet_leaf_334_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0847_ ),
    .Q_N(\register_file_i/_3186_ ),
    .Q(\register_file_i/rf_reg_869_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_86__reg  (.CLK(clknet_leaf_170_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0848_ ),
    .Q_N(\register_file_i/_3185_ ),
    .Q(\register_file_i/rf_reg_86_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_870__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0849_ ),
    .Q_N(\register_file_i/_3184_ ),
    .Q(\register_file_i/rf_reg_870_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_871__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0850_ ),
    .Q_N(\register_file_i/_3183_ ),
    .Q(\register_file_i/rf_reg_871_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_872__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2277),
    .D(\register_file_i/_0851_ ),
    .Q_N(\register_file_i/_3182_ ),
    .Q(\register_file_i/rf_reg_872_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_873__reg  (.CLK(clknet_leaf_335_clk_i),
    .RESET_B(net2169),
    .D(\register_file_i/_0852_ ),
    .Q_N(\register_file_i/_3181_ ),
    .Q(\register_file_i/rf_reg_873_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_874__reg  (.CLK(clknet_leaf_339_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0853_ ),
    .Q_N(\register_file_i/_3180_ ),
    .Q(\register_file_i/rf_reg_874_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_875__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0854_ ),
    .Q_N(\register_file_i/_3179_ ),
    .Q(\register_file_i/rf_reg_875_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_876__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0855_ ),
    .Q_N(\register_file_i/_3178_ ),
    .Q(\register_file_i/rf_reg_876_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_877__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0856_ ),
    .Q_N(\register_file_i/_3177_ ),
    .Q(\register_file_i/rf_reg_877_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_878__reg  (.CLK(clknet_leaf_159_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0857_ ),
    .Q_N(\register_file_i/_3176_ ),
    .Q(\register_file_i/rf_reg_878_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_879__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0858_ ),
    .Q_N(\register_file_i/_3175_ ),
    .Q(\register_file_i/rf_reg_879_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_87__reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(net2195),
    .D(\register_file_i/_0859_ ),
    .Q_N(\register_file_i/_3174_ ),
    .Q(\register_file_i/rf_reg_87_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_880__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2245),
    .D(\register_file_i/_0860_ ),
    .Q_N(\register_file_i/_3173_ ),
    .Q(\register_file_i/rf_reg_880_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_881__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2244),
    .D(\register_file_i/_0861_ ),
    .Q_N(\register_file_i/_3172_ ),
    .Q(\register_file_i/rf_reg_881_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_882__reg  (.CLK(clknet_leaf_159_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0862_ ),
    .Q_N(\register_file_i/_3171_ ),
    .Q(\register_file_i/rf_reg_882_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_883__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0863_ ),
    .Q_N(\register_file_i/_3170_ ),
    .Q(\register_file_i/rf_reg_883_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_884__reg  (.CLK(clknet_leaf_130_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0864_ ),
    .Q_N(\register_file_i/_3169_ ),
    .Q(\register_file_i/rf_reg_884_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_885__reg  (.CLK(clknet_leaf_131_clk_i),
    .RESET_B(net2259),
    .D(\register_file_i/_0865_ ),
    .Q_N(\register_file_i/_3168_ ),
    .Q(\register_file_i/rf_reg_885_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_886__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2251),
    .D(\register_file_i/_0866_ ),
    .Q_N(\register_file_i/_3167_ ),
    .Q(\register_file_i/rf_reg_886_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_887__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net2184),
    .D(\register_file_i/_0867_ ),
    .Q_N(\register_file_i/_3166_ ),
    .Q(\register_file_i/rf_reg_887_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_888__reg  (.CLK(clknet_leaf_174_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0868_ ),
    .Q_N(\register_file_i/_3165_ ),
    .Q(\register_file_i/rf_reg_888_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_889__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net2322),
    .D(\register_file_i/_0869_ ),
    .Q_N(\register_file_i/_3164_ ),
    .Q(\register_file_i/rf_reg_889_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_88__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2295),
    .D(\register_file_i/_0870_ ),
    .Q_N(\register_file_i/_3163_ ),
    .Q(\register_file_i/rf_reg_88_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_890__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2297),
    .D(\register_file_i/_0871_ ),
    .Q_N(\register_file_i/_3162_ ),
    .Q(\register_file_i/rf_reg_890_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_891__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0872_ ),
    .Q_N(\register_file_i/_3161_ ),
    .Q(\register_file_i/rf_reg_891_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_892__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0873_ ),
    .Q_N(\register_file_i/_3160_ ),
    .Q(\register_file_i/rf_reg_892_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_893__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2290),
    .D(\register_file_i/_0874_ ),
    .Q_N(\register_file_i/_3159_ ),
    .Q(\register_file_i/rf_reg_893_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_894__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2258),
    .D(\register_file_i/_0875_ ),
    .Q_N(\register_file_i/_3158_ ),
    .Q(\register_file_i/rf_reg_894_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_895__reg  (.CLK(clknet_leaf_155_clk_i),
    .RESET_B(net2260),
    .D(\register_file_i/_0876_ ),
    .Q_N(\register_file_i/_3157_ ),
    .Q(\register_file_i/rf_reg_895_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_896__reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0877_ ),
    .Q_N(\register_file_i/_3156_ ),
    .Q(\register_file_i/rf_reg_896_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_897__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0878_ ),
    .Q_N(\register_file_i/_3155_ ),
    .Q(\register_file_i/rf_reg_897_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_898__reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0879_ ),
    .Q_N(\register_file_i/_3154_ ),
    .Q(\register_file_i/rf_reg_898_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_899__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2163),
    .D(\register_file_i/_0880_ ),
    .Q_N(\register_file_i/_3153_ ),
    .Q(\register_file_i/rf_reg_899_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_89__reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(net2294),
    .D(\register_file_i/_0881_ ),
    .Q_N(\register_file_i/_3152_ ),
    .Q(\register_file_i/rf_reg_89_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_900__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0882_ ),
    .Q_N(\register_file_i/_3151_ ),
    .Q(\register_file_i/rf_reg_900_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_901__reg  (.CLK(clknet_leaf_314_clk_i),
    .RESET_B(net2282),
    .D(\register_file_i/_0883_ ),
    .Q_N(\register_file_i/_3150_ ),
    .Q(\register_file_i/rf_reg_901_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_902__reg  (.CLK(clknet_leaf_314_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0884_ ),
    .Q_N(\register_file_i/_3149_ ),
    .Q(\register_file_i/rf_reg_902_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_903__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0885_ ),
    .Q_N(\register_file_i/_3148_ ),
    .Q(\register_file_i/rf_reg_903_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_904__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0886_ ),
    .Q_N(\register_file_i/_3147_ ),
    .Q(\register_file_i/rf_reg_904_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_905__reg  (.CLK(clknet_leaf_339_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0887_ ),
    .Q_N(\register_file_i/_3146_ ),
    .Q(\register_file_i/rf_reg_905_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_906__reg  (.CLK(clknet_leaf_341_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0888_ ),
    .Q_N(\register_file_i/_3145_ ),
    .Q(\register_file_i/rf_reg_906_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_907__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0889_ ),
    .Q_N(\register_file_i/_3144_ ),
    .Q(\register_file_i/rf_reg_907_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_908__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0890_ ),
    .Q_N(\register_file_i/_3143_ ),
    .Q(\register_file_i/rf_reg_908_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_909__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0891_ ),
    .Q_N(\register_file_i/_3142_ ),
    .Q(\register_file_i/rf_reg_909_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_90__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0892_ ),
    .Q_N(\register_file_i/_3141_ ),
    .Q(\register_file_i/rf_reg_90_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_910__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0893_ ),
    .Q_N(\register_file_i/_3140_ ),
    .Q(\register_file_i/rf_reg_910_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_911__reg  (.CLK(clknet_leaf_160_clk_i),
    .RESET_B(net2242),
    .D(\register_file_i/_0894_ ),
    .Q_N(\register_file_i/_3139_ ),
    .Q(\register_file_i/rf_reg_911_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_912__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0895_ ),
    .Q_N(\register_file_i/_3138_ ),
    .Q(\register_file_i/rf_reg_912_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_913__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2262),
    .D(\register_file_i/_0896_ ),
    .Q_N(\register_file_i/_3137_ ),
    .Q(\register_file_i/rf_reg_913_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_914__reg  (.CLK(clknet_leaf_129_clk_i),
    .RESET_B(net2230),
    .D(\register_file_i/_0897_ ),
    .Q_N(\register_file_i/_3136_ ),
    .Q(\register_file_i/rf_reg_914_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_915__reg  (.CLK(clknet_leaf_134_clk_i),
    .RESET_B(net2262),
    .D(\register_file_i/_0898_ ),
    .Q_N(\register_file_i/_3135_ ),
    .Q(\register_file_i/rf_reg_915_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_916__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2262),
    .D(\register_file_i/_0899_ ),
    .Q_N(\register_file_i/_3134_ ),
    .Q(\register_file_i/rf_reg_916_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_917__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2264),
    .D(\register_file_i/_0900_ ),
    .Q_N(\register_file_i/_3133_ ),
    .Q(\register_file_i/rf_reg_917_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_918__reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0901_ ),
    .Q_N(\register_file_i/_3132_ ),
    .Q(\register_file_i/rf_reg_918_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_919__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2185),
    .D(\register_file_i/_0902_ ),
    .Q_N(\register_file_i/_3131_ ),
    .Q(\register_file_i/rf_reg_919_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_91__reg  (.CLK(clknet_leaf_53_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0903_ ),
    .Q_N(\register_file_i/_3130_ ),
    .Q(\register_file_i/rf_reg_91_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_920__reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0904_ ),
    .Q_N(\register_file_i/_3129_ ),
    .Q(\register_file_i/rf_reg_920_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_921__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2322),
    .D(\register_file_i/_0905_ ),
    .Q_N(\register_file_i/_3128_ ),
    .Q(\register_file_i/rf_reg_921_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_922__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2297),
    .D(\register_file_i/_0906_ ),
    .Q_N(\register_file_i/_3127_ ),
    .Q(\register_file_i/rf_reg_922_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_923__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0907_ ),
    .Q_N(\register_file_i/_3126_ ),
    .Q(\register_file_i/rf_reg_923_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_924__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0908_ ),
    .Q_N(\register_file_i/_3125_ ),
    .Q(\register_file_i/rf_reg_924_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_925__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0909_ ),
    .Q_N(\register_file_i/_3124_ ),
    .Q(\register_file_i/rf_reg_925_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_926__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2246),
    .D(\register_file_i/_0910_ ),
    .Q_N(\register_file_i/_3123_ ),
    .Q(\register_file_i/rf_reg_926_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_927__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2263),
    .D(\register_file_i/_0911_ ),
    .Q_N(\register_file_i/_3122_ ),
    .Q(\register_file_i/rf_reg_927_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_928__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net2152),
    .D(\register_file_i/_0912_ ),
    .Q_N(\register_file_i/_3121_ ),
    .Q(\register_file_i/rf_reg_928_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_929__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net2147),
    .D(\register_file_i/_0913_ ),
    .Q_N(\register_file_i/_3120_ ),
    .Q(\register_file_i/rf_reg_929_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_92__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0914_ ),
    .Q_N(\register_file_i/_3119_ ),
    .Q(\register_file_i/rf_reg_92_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_930__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0915_ ),
    .Q_N(\register_file_i/_3118_ ),
    .Q(\register_file_i/rf_reg_930_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_931__reg  (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net2159),
    .D(\register_file_i/_0916_ ),
    .Q_N(\register_file_i/_3117_ ),
    .Q(\register_file_i/rf_reg_931_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_932__reg  (.CLK(clknet_leaf_330_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0917_ ),
    .Q_N(\register_file_i/_3116_ ),
    .Q(\register_file_i/rf_reg_932_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_933__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0918_ ),
    .Q_N(\register_file_i/_3115_ ),
    .Q(\register_file_i/rf_reg_933_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_934__reg  (.CLK(clknet_leaf_314_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0919_ ),
    .Q_N(\register_file_i/_3114_ ),
    .Q(\register_file_i/rf_reg_934_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_935__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0920_ ),
    .Q_N(\register_file_i/_3113_ ),
    .Q(\register_file_i/rf_reg_935_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_936__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0921_ ),
    .Q_N(\register_file_i/_3112_ ),
    .Q(\register_file_i/rf_reg_936_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_937__reg  (.CLK(clknet_leaf_339_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0922_ ),
    .Q_N(\register_file_i/_3111_ ),
    .Q(\register_file_i/rf_reg_937_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_938__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0923_ ),
    .Q_N(\register_file_i/_3110_ ),
    .Q(\register_file_i/rf_reg_938_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_939__reg  (.CLK(clknet_leaf_335_clk_i),
    .RESET_B(net2275),
    .D(\register_file_i/_0924_ ),
    .Q_N(\register_file_i/_3109_ ),
    .Q(\register_file_i/rf_reg_939_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_93__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0925_ ),
    .Q_N(\register_file_i/_3108_ ),
    .Q(\register_file_i/rf_reg_93_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_940__reg  (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net2171),
    .D(\register_file_i/_0926_ ),
    .Q_N(\register_file_i/_3107_ ),
    .Q(\register_file_i/rf_reg_940_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_941__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0927_ ),
    .Q_N(\register_file_i/_3106_ ),
    .Q(\register_file_i/rf_reg_941_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_942__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0928_ ),
    .Q_N(\register_file_i/_3105_ ),
    .Q(\register_file_i/rf_reg_942_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_943__reg  (.CLK(clknet_leaf_159_clk_i),
    .RESET_B(net2240),
    .D(\register_file_i/_0929_ ),
    .Q_N(\register_file_i/_3104_ ),
    .Q(\register_file_i/rf_reg_943_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_944__reg  (.CLK(clknet_leaf_158_clk_i),
    .RESET_B(net2243),
    .D(\register_file_i/_0930_ ),
    .Q_N(\register_file_i/_3103_ ),
    .Q(\register_file_i/rf_reg_944_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_945__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2262),
    .D(\register_file_i/_0931_ ),
    .Q_N(\register_file_i/_3102_ ),
    .Q(\register_file_i/rf_reg_945_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_946__reg  (.CLK(clknet_leaf_127_clk_i),
    .RESET_B(net2216),
    .D(\register_file_i/_0932_ ),
    .Q_N(\register_file_i/_3101_ ),
    .Q(\register_file_i/rf_reg_946_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_947__reg  (.CLK(clknet_leaf_122_clk_i),
    .RESET_B(net2236),
    .D(\register_file_i/_0933_ ),
    .Q_N(\register_file_i/_3100_ ),
    .Q(\register_file_i/rf_reg_947_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_948__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2262),
    .D(\register_file_i/_0934_ ),
    .Q_N(\register_file_i/_3099_ ),
    .Q(\register_file_i/rf_reg_948_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_949__reg  (.CLK(clknet_leaf_154_clk_i),
    .RESET_B(net2264),
    .D(\register_file_i/_0935_ ),
    .Q_N(\register_file_i/_3098_ ),
    .Q(\register_file_i/rf_reg_949_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_94__reg  (.CLK(clknet_leaf_168_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0936_ ),
    .Q_N(\register_file_i/_3097_ ),
    .Q(\register_file_i/rf_reg_94_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_950__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0937_ ),
    .Q_N(\register_file_i/_3096_ ),
    .Q(\register_file_i/rf_reg_950_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_951__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2185),
    .D(\register_file_i/_0938_ ),
    .Q_N(\register_file_i/_3095_ ),
    .Q(\register_file_i/rf_reg_951_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_952__reg  (.CLK(clknet_leaf_173_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0939_ ),
    .Q_N(\register_file_i/_3094_ ),
    .Q(\register_file_i/rf_reg_952_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_953__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2322),
    .D(\register_file_i/_0940_ ),
    .Q_N(\register_file_i/_3093_ ),
    .Q(\register_file_i/rf_reg_953_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_954__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2297),
    .D(\register_file_i/_0941_ ),
    .Q_N(\register_file_i/_3092_ ),
    .Q(\register_file_i/rf_reg_954_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_955__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0942_ ),
    .Q_N(\register_file_i/_3091_ ),
    .Q(\register_file_i/rf_reg_955_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_956__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net2293),
    .D(\register_file_i/_0943_ ),
    .Q_N(\register_file_i/_3090_ ),
    .Q(\register_file_i/rf_reg_956_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_957__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0944_ ),
    .Q_N(\register_file_i/_3089_ ),
    .Q(\register_file_i/rf_reg_957_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_958__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2246),
    .D(\register_file_i/_0945_ ),
    .Q_N(\register_file_i/_3088_ ),
    .Q(\register_file_i/rf_reg_958_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_959__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2263),
    .D(\register_file_i/_0946_ ),
    .Q_N(\register_file_i/_3087_ ),
    .Q(\register_file_i/rf_reg_959_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_95__reg  (.CLK(clknet_leaf_170_clk_i),
    .RESET_B(net2253),
    .D(\register_file_i/_0947_ ),
    .Q_N(\register_file_i/_3086_ ),
    .Q(\register_file_i/rf_reg_95_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_960__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0948_ ),
    .Q_N(\register_file_i/_3085_ ),
    .Q(\register_file_i/rf_reg_960_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_961__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0949_ ),
    .Q_N(\register_file_i/_3084_ ),
    .Q(\register_file_i/rf_reg_961_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_962__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0950_ ),
    .Q_N(\register_file_i/_3083_ ),
    .Q(\register_file_i/rf_reg_962_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_963__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0951_ ),
    .Q_N(\register_file_i/_3082_ ),
    .Q(\register_file_i/rf_reg_963_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_964__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2276),
    .D(\register_file_i/_0952_ ),
    .Q_N(\register_file_i/_3081_ ),
    .Q(\register_file_i/rf_reg_964_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_965__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0953_ ),
    .Q_N(\register_file_i/_3080_ ),
    .Q(\register_file_i/rf_reg_965_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_966__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0954_ ),
    .Q_N(\register_file_i/_3079_ ),
    .Q(\register_file_i/rf_reg_966_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_967__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0955_ ),
    .Q_N(\register_file_i/_3078_ ),
    .Q(\register_file_i/rf_reg_967_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_968__reg  (.CLK(clknet_leaf_332_clk_i),
    .RESET_B(net2278),
    .D(\register_file_i/_0956_ ),
    .Q_N(\register_file_i/_3077_ ),
    .Q(\register_file_i/rf_reg_968_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_969__reg  (.CLK(clknet_leaf_335_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0957_ ),
    .Q_N(\register_file_i/_3076_ ),
    .Q(\register_file_i/rf_reg_969_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_96__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2194),
    .D(\register_file_i/_0958_ ),
    .Q_N(\register_file_i/_3075_ ),
    .Q(\register_file_i/rf_reg_96_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_970__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2167),
    .D(\register_file_i/_0959_ ),
    .Q_N(\register_file_i/_3074_ ),
    .Q(\register_file_i/rf_reg_970_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_971__reg  (.CLK(clknet_leaf_341_clk_i),
    .RESET_B(net2168),
    .D(\register_file_i/_0960_ ),
    .Q_N(\register_file_i/_3073_ ),
    .Q(\register_file_i/rf_reg_971_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_972__reg  (.CLK(clknet_leaf_338_clk_i),
    .RESET_B(net2170),
    .D(\register_file_i/_0961_ ),
    .Q_N(\register_file_i/_3072_ ),
    .Q(\register_file_i/rf_reg_972_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_973__reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net2182),
    .D(\register_file_i/_0962_ ),
    .Q_N(\register_file_i/_3071_ ),
    .Q(\register_file_i/rf_reg_973_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_974__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0963_ ),
    .Q_N(\register_file_i/_3070_ ),
    .Q(\register_file_i/rf_reg_974_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_975__reg  (.CLK(clknet_leaf_159_clk_i),
    .RESET_B(net2239),
    .D(\register_file_i/_0964_ ),
    .Q_N(\register_file_i/_3069_ ),
    .Q(\register_file_i/rf_reg_975_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_976__reg  (.CLK(clknet_leaf_156_clk_i),
    .RESET_B(net2244),
    .D(\register_file_i/_0965_ ),
    .Q_N(\register_file_i/_3068_ ),
    .Q(\register_file_i/rf_reg_976_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_977__reg  (.CLK(clknet_leaf_135_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0966_ ),
    .Q_N(\register_file_i/_3067_ ),
    .Q(\register_file_i/rf_reg_977_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_978__reg  (.CLK(clknet_leaf_128_clk_i),
    .RESET_B(net2215),
    .D(\register_file_i/_0967_ ),
    .Q_N(\register_file_i/_3066_ ),
    .Q(\register_file_i/rf_reg_978_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_979__reg  (.CLK(clknet_leaf_135_clk_i),
    .RESET_B(net2235),
    .D(\register_file_i/_0968_ ),
    .Q_N(\register_file_i/_3065_ ),
    .Q(\register_file_i/rf_reg_979_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_97__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net2192),
    .D(\register_file_i/_0969_ ),
    .Q_N(\register_file_i/_3064_ ),
    .Q(\register_file_i/rf_reg_97_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_980__reg  (.CLK(clknet_leaf_133_clk_i),
    .RESET_B(net2261),
    .D(\register_file_i/_0970_ ),
    .Q_N(\register_file_i/_3063_ ),
    .Q(\register_file_i/rf_reg_980_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_981__reg  (.CLK(clknet_leaf_147_clk_i),
    .RESET_B(net2264),
    .D(\register_file_i/_0971_ ),
    .Q_N(\register_file_i/_3062_ ),
    .Q(\register_file_i/rf_reg_981_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_982__reg  (.CLK(clknet_leaf_171_clk_i),
    .RESET_B(net2321),
    .D(\register_file_i/_0972_ ),
    .Q_N(\register_file_i/_3061_ ),
    .Q(\register_file_i/rf_reg_982_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_983__reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net2241),
    .D(\register_file_i/_0973_ ),
    .Q_N(\register_file_i/_3060_ ),
    .Q(\register_file_i/rf_reg_983_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_984__reg  (.CLK(clknet_leaf_172_clk_i),
    .RESET_B(net2320),
    .D(\register_file_i/_0974_ ),
    .Q_N(\register_file_i/_3059_ ),
    .Q(\register_file_i/rf_reg_984_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_985__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net2319),
    .D(\register_file_i/_0975_ ),
    .Q_N(\register_file_i/_3058_ ),
    .Q(\register_file_i/rf_reg_985_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_986__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0976_ ),
    .Q_N(\register_file_i/_3057_ ),
    .Q(\register_file_i/rf_reg_986_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_987__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2296),
    .D(\register_file_i/_0977_ ),
    .Q_N(\register_file_i/_3056_ ),
    .Q(\register_file_i/rf_reg_987_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_988__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net2292),
    .D(\register_file_i/_0978_ ),
    .Q_N(\register_file_i/_3055_ ),
    .Q(\register_file_i/rf_reg_988_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_989__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net2291),
    .D(\register_file_i/_0979_ ),
    .Q_N(\register_file_i/_3054_ ),
    .Q(\register_file_i/rf_reg_989_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_98__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net2188),
    .D(\register_file_i/_0980_ ),
    .Q_N(\register_file_i/_3053_ ),
    .Q(\register_file_i/rf_reg_98_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_990__reg  (.CLK(clknet_leaf_131_clk_i),
    .RESET_B(net2244),
    .D(\register_file_i/_0981_ ),
    .Q_N(\register_file_i/_3052_ ),
    .Q(\register_file_i/rf_reg_990_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_991__reg  (.CLK(clknet_leaf_132_clk_i),
    .RESET_B(net2264),
    .D(\register_file_i/_0982_ ),
    .Q_N(\register_file_i/_3051_ ),
    .Q(\register_file_i/rf_reg_991_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_992__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0983_ ),
    .Q_N(\register_file_i/_3050_ ),
    .Q(\register_file_i/rf_reg_992_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_993__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net2151),
    .D(\register_file_i/_0984_ ),
    .Q_N(\register_file_i/_3049_ ),
    .Q(\register_file_i/rf_reg_993_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_994__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2166),
    .D(\register_file_i/_0985_ ),
    .Q_N(\register_file_i/_3048_ ),
    .Q(\register_file_i/rf_reg_994_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_995__reg  (.CLK(clknet_leaf_340_clk_i),
    .RESET_B(net2158),
    .D(\register_file_i/_0986_ ),
    .Q_N(\register_file_i/_3047_ ),
    .Q(\register_file_i/rf_reg_995_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_996__reg  (.CLK(clknet_leaf_329_clk_i),
    .RESET_B(net2277),
    .D(\register_file_i/_0987_ ),
    .Q_N(\register_file_i/_3046_ ),
    .Q(\register_file_i/rf_reg_996_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_997__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2279),
    .D(\register_file_i/_0988_ ),
    .Q_N(\register_file_i/_3045_ ),
    .Q(\register_file_i/rf_reg_997_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_998__reg  (.CLK(clknet_leaf_313_clk_i),
    .RESET_B(net2289),
    .D(\register_file_i/_0989_ ),
    .Q_N(\register_file_i/_3044_ ),
    .Q(\register_file_i/rf_reg_998_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_999__reg  (.CLK(clknet_leaf_333_clk_i),
    .RESET_B(net2285),
    .D(\register_file_i/_0990_ ),
    .Q_N(\register_file_i/_3043_ ),
    .Q(\register_file_i/rf_reg_999_ ));
 sg13g2_dfrbp_1 \register_file_i/rf_reg_99__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net2190),
    .D(\register_file_i/_0991_ ),
    .Q_N(\register_file_i/_3042_ ),
    .Q(\register_file_i/rf_reg_99_ ));
 sg13g2_tielo cve2_core_1 (.L_LO(net1));
 sg13g2_tielo cve2_core_2 (.L_LO(net2));
 sg13g2_tielo cve2_core_3 (.L_LO(net3));
 sg13g2_tielo cve2_core_4 (.L_LO(net4));
 sg13g2_tielo cve2_core_5 (.L_LO(net5));
 sg13g2_tielo \cs_registers_i/_3039__6  (.L_LO(net6));
 sg13g2_tielo _12186__8 (.L_LO(net8));
 sg13g2_tielo _12187__9 (.L_LO(net9));
 sg13g2_tielo _12189__10 (.L_LO(net10));
 sg13g2_buf_2 fanout1335 (.A(_05047_),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1337));
 sg13g2_buf_4 fanout1337 (.X(net1337),
    .A(net1338));
 sg13g2_buf_4 fanout1338 (.X(net1338),
    .A(_04807_));
 sg13g2_buf_4 fanout1339 (.X(net1339),
    .A(_04725_));
 sg13g2_buf_2 fanout1340 (.A(_04725_),
    .X(net1340));
 sg13g2_buf_4 fanout1341 (.X(net1341),
    .A(_04431_));
 sg13g2_buf_2 fanout1342 (.A(_04431_),
    .X(net1342));
 sg13g2_buf_2 fanout1343 (.A(_02526_),
    .X(net1343));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(_02039_));
 sg13g2_buf_2 fanout1345 (.A(_01964_),
    .X(net1345));
 sg13g2_buf_2 fanout1346 (.A(_01936_),
    .X(net1346));
 sg13g2_buf_2 fanout1347 (.A(net1348),
    .X(net1347));
 sg13g2_buf_1 fanout1348 (.A(_01814_),
    .X(net1348));
 sg13g2_buf_4 fanout1349 (.X(net1349),
    .A(_01314_));
 sg13g2_buf_2 fanout1350 (.A(_01314_),
    .X(net1350));
 sg13g2_buf_4 fanout1351 (.X(net1351),
    .A(alu_operand_a_ex_15_));
 sg13g2_buf_2 fanout1352 (.A(alu_operand_a_ex_13_),
    .X(net1352));
 sg13g2_buf_2 fanout1353 (.A(net1354),
    .X(net1353));
 sg13g2_buf_2 fanout1354 (.A(net1357),
    .X(net1354));
 sg13g2_buf_2 fanout1355 (.A(net1356),
    .X(net1355));
 sg13g2_buf_2 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_2 fanout1357 (.A(net1363),
    .X(net1357));
 sg13g2_buf_2 fanout1358 (.A(net1363),
    .X(net1358));
 sg13g2_buf_1 fanout1359 (.A(net1363),
    .X(net1359));
 sg13g2_buf_2 fanout1360 (.A(net1362),
    .X(net1360));
 sg13g2_buf_2 fanout1361 (.A(net1362),
    .X(net1361));
 sg13g2_buf_1 fanout1362 (.A(net1363),
    .X(net1362));
 sg13g2_buf_1 fanout1363 (.A(_08519_),
    .X(net1363));
 sg13g2_buf_2 fanout1364 (.A(net1365),
    .X(net1364));
 sg13g2_buf_2 fanout1365 (.A(net1368),
    .X(net1365));
 sg13g2_buf_2 fanout1366 (.A(net1367),
    .X(net1366));
 sg13g2_buf_2 fanout1367 (.A(net1368),
    .X(net1367));
 sg13g2_buf_2 fanout1368 (.A(_08515_),
    .X(net1368));
 sg13g2_buf_2 fanout1369 (.A(net1370),
    .X(net1369));
 sg13g2_buf_1 fanout1370 (.A(_06761_),
    .X(net1370));
 sg13g2_buf_2 fanout1371 (.A(_05658_),
    .X(net1371));
 sg13g2_buf_4 fanout1372 (.X(net1372),
    .A(_05649_));
 sg13g2_buf_2 fanout1373 (.A(_05649_),
    .X(net1373));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(net1375));
 sg13g2_buf_4 fanout1375 (.X(net1375),
    .A(_05041_));
 sg13g2_buf_2 fanout1376 (.A(_04253_),
    .X(net1376));
 sg13g2_buf_2 fanout1377 (.A(net1378),
    .X(net1377));
 sg13g2_buf_2 fanout1378 (.A(_04237_),
    .X(net1378));
 sg13g2_buf_2 fanout1379 (.A(_04051_),
    .X(net1379));
 sg13g2_buf_2 fanout1380 (.A(net1381),
    .X(net1380));
 sg13g2_buf_4 fanout1381 (.X(net1381),
    .A(_03932_));
 sg13g2_buf_2 fanout1382 (.A(net1391),
    .X(net1382));
 sg13g2_buf_1 fanout1383 (.A(net1391),
    .X(net1383));
 sg13g2_buf_2 fanout1384 (.A(net1387),
    .X(net1384));
 sg13g2_buf_2 fanout1385 (.A(net1387),
    .X(net1385));
 sg13g2_buf_1 fanout1386 (.A(net1387),
    .X(net1386));
 sg13g2_buf_2 fanout1387 (.A(net1391),
    .X(net1387));
 sg13g2_buf_2 fanout1388 (.A(net1390),
    .X(net1388));
 sg13g2_buf_1 fanout1389 (.A(net1390),
    .X(net1389));
 sg13g2_buf_1 fanout1390 (.A(net1391),
    .X(net1390));
 sg13g2_buf_2 fanout1391 (.A(csr_mtvec_init),
    .X(net1391));
 sg13g2_buf_2 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_2 fanout1393 (.A(net1394),
    .X(net1393));
 sg13g2_buf_2 fanout1394 (.A(_03457_),
    .X(net1394));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(_03428_));
 sg13g2_buf_2 fanout1396 (.A(_03428_),
    .X(net1396));
 sg13g2_buf_2 fanout1397 (.A(_02642_),
    .X(net1397));
 sg13g2_buf_2 fanout1398 (.A(_02328_),
    .X(net1398));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(_02259_));
 sg13g2_buf_2 fanout1400 (.A(_02164_),
    .X(net1400));
 sg13g2_buf_2 fanout1401 (.A(_02159_),
    .X(net1401));
 sg13g2_buf_4 fanout1402 (.X(net1402),
    .A(net1403));
 sg13g2_buf_4 fanout1403 (.X(net1403),
    .A(_01630_));
 sg13g2_buf_4 fanout1404 (.X(net1404),
    .A(alu_operand_a_ex_5_));
 sg13g2_buf_2 fanout1405 (.A(alu_operand_a_ex_5_),
    .X(net1405));
 sg13g2_buf_8 fanout1406 (.A(_01307_),
    .X(net1406));
 sg13g2_buf_2 fanout1407 (.A(_01307_),
    .X(net1407));
 sg13g2_buf_4 fanout1408 (.X(net1408),
    .A(alu_operand_a_ex_3_));
 sg13g2_buf_4 fanout1409 (.X(net1409),
    .A(alu_operand_a_ex_2_));
 sg13g2_buf_2 fanout1410 (.A(alu_operand_a_ex_2_),
    .X(net1410));
 sg13g2_buf_8 fanout1411 (.A(alu_operand_a_ex_1_),
    .X(net1411));
 sg13g2_buf_4 fanout1412 (.X(net1412),
    .A(_01217_));
 sg13g2_buf_1 fanout1413 (.A(_01217_),
    .X(net1413));
 sg13g2_buf_4 fanout1414 (.X(net1414),
    .A(_01214_));
 sg13g2_buf_2 fanout1415 (.A(_01214_),
    .X(net1415));
 sg13g2_buf_2 fanout1416 (.A(net1420),
    .X(net1416));
 sg13g2_buf_1 fanout1417 (.A(net1420),
    .X(net1417));
 sg13g2_buf_2 fanout1418 (.A(net1420),
    .X(net1418));
 sg13g2_buf_2 fanout1419 (.A(net1420),
    .X(net1419));
 sg13g2_buf_1 fanout1420 (.A(_08535_),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(net1425),
    .X(net1421));
 sg13g2_buf_2 fanout1422 (.A(net1425),
    .X(net1422));
 sg13g2_buf_2 fanout1423 (.A(net1424),
    .X(net1423));
 sg13g2_buf_2 fanout1424 (.A(net1425),
    .X(net1424));
 sg13g2_buf_2 fanout1425 (.A(_08522_),
    .X(net1425));
 sg13g2_buf_2 fanout1426 (.A(_07664_),
    .X(net1426));
 sg13g2_buf_2 fanout1427 (.A(_07664_),
    .X(net1427));
 sg13g2_buf_2 fanout1428 (.A(net1429),
    .X(net1428));
 sg13g2_buf_2 fanout1429 (.A(net1430),
    .X(net1429));
 sg13g2_buf_2 fanout1430 (.A(net1432),
    .X(net1430));
 sg13g2_buf_2 fanout1431 (.A(net1432),
    .X(net1431));
 sg13g2_buf_2 fanout1432 (.A(_07258_),
    .X(net1432));
 sg13g2_buf_2 fanout1433 (.A(net1434),
    .X(net1433));
 sg13g2_buf_4 fanout1434 (.X(net1434),
    .A(_05302_));
 sg13g2_buf_2 fanout1435 (.A(net1436),
    .X(net1435));
 sg13g2_buf_4 fanout1436 (.X(net1436),
    .A(_05192_));
 sg13g2_buf_2 fanout1437 (.A(_04786_),
    .X(net1437));
 sg13g2_buf_4 fanout1438 (.X(net1438),
    .A(_04786_));
 sg13g2_buf_2 fanout1439 (.A(net1440),
    .X(net1439));
 sg13g2_buf_2 fanout1440 (.A(_04174_),
    .X(net1440));
 sg13g2_buf_2 fanout1441 (.A(net1444),
    .X(net1441));
 sg13g2_buf_2 fanout1442 (.A(net1444),
    .X(net1442));
 sg13g2_buf_1 fanout1443 (.A(net1444),
    .X(net1443));
 sg13g2_buf_2 fanout1444 (.A(net1446),
    .X(net1444));
 sg13g2_buf_2 fanout1445 (.A(net1446),
    .X(net1445));
 sg13g2_buf_1 fanout1446 (.A(_04119_),
    .X(net1446));
 sg13g2_buf_2 fanout1447 (.A(net1448),
    .X(net1447));
 sg13g2_buf_2 fanout1448 (.A(_03967_),
    .X(net1448));
 sg13g2_buf_2 fanout1449 (.A(_03967_),
    .X(net1449));
 sg13g2_buf_2 fanout1450 (.A(_03967_),
    .X(net1450));
 sg13g2_buf_4 fanout1451 (.X(net1451),
    .A(net1453));
 sg13g2_buf_1 fanout1452 (.A(net1453),
    .X(net1452));
 sg13g2_buf_2 fanout1453 (.A(_03951_),
    .X(net1453));
 sg13g2_buf_4 fanout1454 (.X(net1454),
    .A(net1455));
 sg13g2_buf_4 fanout1455 (.X(net1455),
    .A(_03951_));
 sg13g2_buf_2 fanout1456 (.A(_03322_),
    .X(net1456));
 sg13g2_buf_4 fanout1457 (.X(net1457),
    .A(_02345_));
 sg13g2_buf_2 fanout1458 (.A(_02345_),
    .X(net1458));
 sg13g2_buf_4 fanout1459 (.X(net1459),
    .A(net1462));
 sg13g2_buf_4 fanout1460 (.X(net1460),
    .A(net1461));
 sg13g2_buf_4 fanout1461 (.X(net1461),
    .A(net1462));
 sg13g2_buf_2 fanout1462 (.A(_02345_),
    .X(net1462));
 sg13g2_buf_4 fanout1463 (.X(net1463),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ));
 sg13g2_buf_2 fanout1464 (.A(net1465),
    .X(net1464));
 sg13g2_buf_1 fanout1465 (.A(net1466),
    .X(net1465));
 sg13g2_buf_4 fanout1466 (.X(net1466),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_9_ ));
 sg13g2_buf_4 fanout1467 (.X(net1467),
    .A(net1468));
 sg13g2_buf_2 fanout1468 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ),
    .X(net1468));
 sg13g2_buf_4 fanout1469 (.X(net1469),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_15_ ));
 sg13g2_buf_2 fanout1470 (.A(net1471),
    .X(net1470));
 sg13g2_buf_4 fanout1471 (.X(net1471),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_16_ ));
 sg13g2_buf_2 fanout1472 (.A(_07195_),
    .X(net1472));
 sg13g2_buf_2 fanout1473 (.A(net1475),
    .X(net1473));
 sg13g2_buf_2 fanout1474 (.A(net1475),
    .X(net1474));
 sg13g2_buf_4 fanout1475 (.X(net1475),
    .A(_04527_));
 sg13g2_buf_2 fanout1476 (.A(net1477),
    .X(net1476));
 sg13g2_buf_2 fanout1477 (.A(_04236_),
    .X(net1477));
 sg13g2_buf_4 fanout1478 (.X(net1478),
    .A(_04134_));
 sg13g2_buf_4 fanout1479 (.X(net1479),
    .A(net1480));
 sg13g2_buf_4 fanout1480 (.X(net1480),
    .A(net1481));
 sg13g2_buf_4 fanout1481 (.X(net1481),
    .A(net1482));
 sg13g2_buf_4 fanout1482 (.X(net1482),
    .A(net1483));
 sg13g2_buf_4 fanout1483 (.X(net1483),
    .A(csr_save_if));
 sg13g2_buf_4 fanout1484 (.X(net1484),
    .A(net1488));
 sg13g2_buf_4 fanout1485 (.X(net1485),
    .A(net1487));
 sg13g2_buf_1 fanout1486 (.A(net1487),
    .X(net1486));
 sg13g2_buf_2 fanout1487 (.A(net1488),
    .X(net1487));
 sg13g2_buf_2 fanout1488 (.A(net1489),
    .X(net1488));
 sg13g2_buf_2 fanout1489 (.A(_03314_),
    .X(net1489));
 sg13g2_buf_2 fanout1490 (.A(_01427_),
    .X(net1490));
 sg13g2_buf_4 fanout1491 (.X(net1491),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_22_ ));
 sg13g2_buf_2 fanout1492 (.A(net1493),
    .X(net1492));
 sg13g2_buf_2 fanout1493 (.A(net1494),
    .X(net1493));
 sg13g2_buf_4 fanout1494 (.X(net1494),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_23_ ));
 sg13g2_buf_2 fanout1495 (.A(net1496),
    .X(net1495));
 sg13g2_buf_2 fanout1496 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_25_ ),
    .X(net1496));
 sg13g2_buf_4 fanout1497 (.X(net1497),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_26_ ));
 sg13g2_buf_4 fanout1498 (.X(net1498),
    .A(net1499));
 sg13g2_buf_4 fanout1499 (.X(net1499),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_27_ ));
 sg13g2_buf_4 fanout1500 (.X(net1500),
    .A(net1501));
 sg13g2_buf_2 fanout1501 (.A(net1502),
    .X(net1501));
 sg13g2_buf_2 fanout1502 (.A(net1503),
    .X(net1502));
 sg13g2_buf_4 fanout1503 (.X(net1503),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_1_ ));
 sg13g2_buf_4 fanout1504 (.X(net1504),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_buf_2 fanout1505 (.A(net1506),
    .X(net1505));
 sg13g2_buf_1 fanout1506 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_3_ ),
    .X(net1506));
 sg13g2_buf_4 fanout1507 (.X(net1507),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_4_ ));
 sg13g2_buf_2 fanout1508 (.A(net1510),
    .X(net1508));
 sg13g2_buf_1 fanout1509 (.A(net1510),
    .X(net1509));
 sg13g2_buf_1 fanout1510 (.A(net1511),
    .X(net1510));
 sg13g2_buf_4 fanout1511 (.X(net1511),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_5_ ));
 sg13g2_buf_2 fanout1512 (.A(net1513),
    .X(net1512));
 sg13g2_buf_4 fanout1513 (.X(net1513),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_6_ ));
 sg13g2_buf_2 fanout1514 (.A(net1515),
    .X(net1514));
 sg13g2_buf_1 fanout1515 (.A(net1516),
    .X(net1515));
 sg13g2_buf_4 fanout1516 (.X(net1516),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_18_ ));
 sg13g2_buf_2 fanout1517 (.A(net1519),
    .X(net1517));
 sg13g2_buf_1 fanout1518 (.A(net1519),
    .X(net1518));
 sg13g2_buf_1 fanout1519 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ),
    .X(net1519));
 sg13g2_buf_4 fanout1520 (.X(net1520),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_21_ ));
 sg13g2_buf_1 fanout1521 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_21_ ),
    .X(net1521));
 sg13g2_buf_2 fanout1522 (.A(net1525),
    .X(net1522));
 sg13g2_buf_2 fanout1523 (.A(net1525),
    .X(net1523));
 sg13g2_buf_4 fanout1524 (.X(net1524),
    .A(net1525));
 sg13g2_buf_2 fanout1525 (.A(_07566_),
    .X(net1525));
 sg13g2_buf_2 fanout1526 (.A(net1528),
    .X(net1526));
 sg13g2_buf_2 fanout1527 (.A(net1528),
    .X(net1527));
 sg13g2_buf_4 fanout1528 (.X(net1528),
    .A(_07563_));
 sg13g2_buf_2 fanout1529 (.A(net1532),
    .X(net1529));
 sg13g2_buf_4 fanout1530 (.X(net1530),
    .A(net1531));
 sg13g2_buf_2 fanout1531 (.A(net1532),
    .X(net1531));
 sg13g2_buf_1 fanout1532 (.A(_07514_),
    .X(net1532));
 sg13g2_buf_2 fanout1533 (.A(net1535),
    .X(net1533));
 sg13g2_buf_1 fanout1534 (.A(net1535),
    .X(net1534));
 sg13g2_buf_2 fanout1535 (.A(net1537),
    .X(net1535));
 sg13g2_buf_2 fanout1536 (.A(net1537),
    .X(net1536));
 sg13g2_buf_2 fanout1537 (.A(_07470_),
    .X(net1537));
 sg13g2_buf_2 fanout1538 (.A(net1540),
    .X(net1538));
 sg13g2_buf_1 fanout1539 (.A(net1540),
    .X(net1539));
 sg13g2_buf_2 fanout1540 (.A(net1543),
    .X(net1540));
 sg13g2_buf_2 fanout1541 (.A(net1543),
    .X(net1541));
 sg13g2_buf_2 fanout1542 (.A(net1543),
    .X(net1542));
 sg13g2_buf_2 fanout1543 (.A(_04041_),
    .X(net1543));
 sg13g2_buf_2 fanout1544 (.A(_03693_),
    .X(net1544));
 sg13g2_buf_2 fanout1545 (.A(net1549),
    .X(net1545));
 sg13g2_buf_2 fanout1546 (.A(net1548),
    .X(net1546));
 sg13g2_buf_1 fanout1547 (.A(net1548),
    .X(net1547));
 sg13g2_buf_2 fanout1548 (.A(net1549),
    .X(net1548));
 sg13g2_buf_2 fanout1549 (.A(net1550),
    .X(net1549));
 sg13g2_buf_2 fanout1550 (.A(_03306_),
    .X(net1550));
 sg13g2_buf_4 fanout1551 (.X(net1551),
    .A(net1556));
 sg13g2_buf_2 fanout1552 (.A(net1553),
    .X(net1552));
 sg13g2_buf_2 fanout1553 (.A(net1554),
    .X(net1553));
 sg13g2_buf_1 fanout1554 (.A(net1555),
    .X(net1554));
 sg13g2_buf_1 fanout1555 (.A(net1556),
    .X(net1555));
 sg13g2_buf_2 fanout1556 (.A(_03299_),
    .X(net1556));
 sg13g2_buf_2 fanout1557 (.A(net1561),
    .X(net1557));
 sg13g2_buf_2 fanout1558 (.A(net1561),
    .X(net1558));
 sg13g2_buf_2 fanout1559 (.A(net1561),
    .X(net1559));
 sg13g2_buf_1 fanout1560 (.A(net1561),
    .X(net1560));
 sg13g2_buf_2 fanout1561 (.A(_01918_),
    .X(net1561));
 sg13g2_buf_2 fanout1562 (.A(_01721_),
    .X(net1562));
 sg13g2_buf_2 fanout1563 (.A(_07693_),
    .X(net1563));
 sg13g2_buf_2 fanout1564 (.A(_07693_),
    .X(net1564));
 sg13g2_buf_2 fanout1565 (.A(net1566),
    .X(net1565));
 sg13g2_buf_2 fanout1566 (.A(_05912_),
    .X(net1566));
 sg13g2_buf_2 fanout1567 (.A(net1568),
    .X(net1567));
 sg13g2_buf_2 fanout1568 (.A(_05910_),
    .X(net1568));
 sg13g2_buf_2 fanout1569 (.A(_04132_),
    .X(net1569));
 sg13g2_buf_1 fanout1570 (.A(net1571),
    .X(net1570));
 sg13g2_buf_2 fanout1571 (.A(_04132_),
    .X(net1571));
 sg13g2_buf_2 fanout1572 (.A(net1574),
    .X(net1572));
 sg13g2_buf_1 fanout1573 (.A(net1574),
    .X(net1573));
 sg13g2_buf_2 fanout1574 (.A(net1575),
    .X(net1574));
 sg13g2_buf_2 fanout1575 (.A(_04132_),
    .X(net1575));
 sg13g2_buf_2 fanout1576 (.A(net1577),
    .X(net1576));
 sg13g2_buf_2 fanout1577 (.A(net1578),
    .X(net1577));
 sg13g2_buf_2 fanout1578 (.A(net1579),
    .X(net1578));
 sg13g2_buf_2 fanout1579 (.A(_04030_),
    .X(net1579));
 sg13g2_buf_2 fanout1580 (.A(_01682_),
    .X(net1580));
 sg13g2_buf_2 fanout1581 (.A(_01669_),
    .X(net1581));
 sg13g2_buf_2 fanout1582 (.A(net1584),
    .X(net1582));
 sg13g2_buf_1 fanout1583 (.A(net1584),
    .X(net1583));
 sg13g2_buf_2 fanout1584 (.A(net1585),
    .X(net1584));
 sg13g2_buf_2 fanout1585 (.A(net1588),
    .X(net1585));
 sg13g2_buf_2 fanout1586 (.A(net1587),
    .X(net1586));
 sg13g2_buf_2 fanout1587 (.A(net1588),
    .X(net1587));
 sg13g2_buf_2 fanout1588 (.A(net1589),
    .X(net1588));
 sg13g2_buf_2 fanout1589 (.A(net1592),
    .X(net1589));
 sg13g2_buf_2 fanout1590 (.A(net1592),
    .X(net1590));
 sg13g2_buf_2 fanout1591 (.A(net1592),
    .X(net1591));
 sg13g2_buf_2 fanout1592 (.A(_01194_),
    .X(net1592));
 sg13g2_buf_2 fanout1593 (.A(net1594),
    .X(net1593));
 sg13g2_buf_2 fanout1594 (.A(net1597),
    .X(net1594));
 sg13g2_buf_2 fanout1595 (.A(net1596),
    .X(net1595));
 sg13g2_buf_2 fanout1596 (.A(net1597),
    .X(net1596));
 sg13g2_buf_1 fanout1597 (.A(net1599),
    .X(net1597));
 sg13g2_buf_4 fanout1598 (.X(net1598),
    .A(net1599));
 sg13g2_buf_2 fanout1599 (.A(_01173_),
    .X(net1599));
 sg13g2_buf_2 fanout1600 (.A(net1601),
    .X(net1600));
 sg13g2_buf_2 fanout1601 (.A(_00583_),
    .X(net1601));
 sg13g2_buf_2 fanout1602 (.A(_08620_),
    .X(net1602));
 sg13g2_buf_2 fanout1603 (.A(net1605),
    .X(net1603));
 sg13g2_buf_2 fanout1604 (.A(net1605),
    .X(net1604));
 sg13g2_buf_2 fanout1605 (.A(_07637_),
    .X(net1605));
 sg13g2_buf_2 fanout1606 (.A(_07592_),
    .X(net1606));
 sg13g2_buf_2 fanout1607 (.A(_07527_),
    .X(net1607));
 sg13g2_buf_1 fanout1608 (.A(_07527_),
    .X(net1608));
 sg13g2_buf_2 fanout1609 (.A(_07523_),
    .X(net1609));
 sg13g2_buf_4 fanout1610 (.X(net1610),
    .A(_07519_));
 sg13g2_buf_1 fanout1611 (.A(_07519_),
    .X(net1611));
 sg13g2_buf_2 fanout1612 (.A(_01880_),
    .X(net1612));
 sg13g2_buf_2 fanout1613 (.A(net1614),
    .X(net1613));
 sg13g2_buf_2 fanout1614 (.A(_01778_),
    .X(net1614));
 sg13g2_buf_2 fanout1615 (.A(net1616),
    .X(net1615));
 sg13g2_buf_4 fanout1616 (.X(net1616),
    .A(_01553_));
 sg13g2_buf_2 fanout1617 (.A(net1619),
    .X(net1617));
 sg13g2_buf_1 fanout1618 (.A(net1619),
    .X(net1618));
 sg13g2_buf_1 fanout1619 (.A(net1621),
    .X(net1619));
 sg13g2_buf_2 fanout1620 (.A(net1621),
    .X(net1620));
 sg13g2_buf_2 fanout1621 (.A(_01176_),
    .X(net1621));
 sg13g2_buf_2 fanout1622 (.A(_07672_),
    .X(net1622));
 sg13g2_buf_4 fanout1623 (.X(net1623),
    .A(net1624));
 sg13g2_buf_2 fanout1624 (.A(_07575_),
    .X(net1624));
 sg13g2_buf_2 fanout1625 (.A(_07535_),
    .X(net1625));
 sg13g2_buf_2 fanout1626 (.A(_07535_),
    .X(net1626));
 sg13g2_buf_2 fanout1627 (.A(net1628),
    .X(net1627));
 sg13g2_buf_2 fanout1628 (.A(_07531_),
    .X(net1628));
 sg13g2_buf_2 fanout1629 (.A(net1631),
    .X(net1629));
 sg13g2_buf_2 fanout1630 (.A(net1631),
    .X(net1630));
 sg13g2_buf_2 fanout1631 (.A(_07508_),
    .X(net1631));
 sg13g2_buf_2 fanout1632 (.A(net1633),
    .X(net1632));
 sg13g2_buf_2 fanout1633 (.A(_07508_),
    .X(net1633));
 sg13g2_buf_2 fanout1634 (.A(net1635),
    .X(net1634));
 sg13g2_buf_2 fanout1635 (.A(_04137_),
    .X(net1635));
 sg13g2_buf_2 fanout1636 (.A(net1639),
    .X(net1636));
 sg13g2_buf_1 fanout1637 (.A(net1639),
    .X(net1637));
 sg13g2_buf_2 fanout1638 (.A(net1639),
    .X(net1638));
 sg13g2_buf_1 fanout1639 (.A(_04137_),
    .X(net1639));
 sg13g2_buf_2 fanout1640 (.A(net1641),
    .X(net1640));
 sg13g2_buf_2 fanout1641 (.A(_03730_),
    .X(net1641));
 sg13g2_buf_2 fanout1642 (.A(net1643),
    .X(net1642));
 sg13g2_buf_2 fanout1643 (.A(net1644),
    .X(net1643));
 sg13g2_buf_2 fanout1644 (.A(net1645),
    .X(net1644));
 sg13g2_buf_2 fanout1645 (.A(_03327_),
    .X(net1645));
 sg13g2_buf_2 fanout1646 (.A(net1647),
    .X(net1646));
 sg13g2_buf_2 fanout1647 (.A(_08634_),
    .X(net1647));
 sg13g2_buf_4 fanout1648 (.X(net1648),
    .A(net1651));
 sg13g2_buf_4 fanout1649 (.X(net1649),
    .A(net1650));
 sg13g2_buf_2 fanout1650 (.A(net1651),
    .X(net1650));
 sg13g2_buf_4 fanout1651 (.X(net1651),
    .A(_08384_));
 sg13g2_buf_4 fanout1652 (.X(net1652),
    .A(net1655));
 sg13g2_buf_2 fanout1653 (.A(net1655),
    .X(net1653));
 sg13g2_buf_4 fanout1654 (.X(net1654),
    .A(net1655));
 sg13g2_buf_2 fanout1655 (.A(_08375_),
    .X(net1655));
 sg13g2_buf_2 fanout1656 (.A(net1658),
    .X(net1656));
 sg13g2_buf_1 fanout1657 (.A(net1658),
    .X(net1657));
 sg13g2_buf_2 fanout1658 (.A(net1660),
    .X(net1658));
 sg13g2_buf_4 fanout1659 (.X(net1659),
    .A(net1660));
 sg13g2_buf_2 fanout1660 (.A(_07568_),
    .X(net1660));
 sg13g2_buf_2 fanout1661 (.A(_07546_),
    .X(net1661));
 sg13g2_buf_2 fanout1662 (.A(_07537_),
    .X(net1662));
 sg13g2_buf_2 fanout1663 (.A(_07537_),
    .X(net1663));
 sg13g2_buf_2 fanout1664 (.A(net1669),
    .X(net1664));
 sg13g2_buf_1 fanout1665 (.A(net1669),
    .X(net1665));
 sg13g2_buf_2 fanout1666 (.A(net1669),
    .X(net1666));
 sg13g2_buf_2 fanout1667 (.A(net1668),
    .X(net1667));
 sg13g2_buf_2 fanout1668 (.A(net1669),
    .X(net1668));
 sg13g2_buf_2 fanout1669 (.A(_07501_),
    .X(net1669));
 sg13g2_buf_2 fanout1670 (.A(net1671),
    .X(net1670));
 sg13g2_buf_2 fanout1671 (.A(net1673),
    .X(net1671));
 sg13g2_buf_4 fanout1672 (.X(net1672),
    .A(net1673));
 sg13g2_buf_2 fanout1673 (.A(_07494_),
    .X(net1673));
 sg13g2_buf_2 fanout1674 (.A(_01848_),
    .X(net1674));
 sg13g2_buf_1 fanout1675 (.A(_01848_),
    .X(net1675));
 sg13g2_buf_4 fanout1676 (.X(net1676),
    .A(net1678));
 sg13g2_buf_4 fanout1677 (.X(net1677),
    .A(net1678));
 sg13g2_buf_2 fanout1678 (.A(net1681),
    .X(net1678));
 sg13g2_buf_2 fanout1679 (.A(net1681),
    .X(net1679));
 sg13g2_buf_2 fanout1680 (.A(net1681),
    .X(net1680));
 sg13g2_buf_2 fanout1681 (.A(_01304_),
    .X(net1681));
 sg13g2_buf_4 fanout1682 (.X(net1682),
    .A(net1683));
 sg13g2_buf_4 fanout1683 (.X(net1683),
    .A(net1687));
 sg13g2_buf_2 fanout1684 (.A(net1687),
    .X(net1684));
 sg13g2_buf_4 fanout1685 (.X(net1685),
    .A(net1687));
 sg13g2_buf_2 fanout1686 (.A(net1687),
    .X(net1686));
 sg13g2_buf_4 fanout1687 (.X(net1687),
    .A(\register_file_i/_1951_ ));
 sg13g2_buf_2 fanout1688 (.A(net1689),
    .X(net1688));
 sg13g2_buf_4 fanout1689 (.X(net1689),
    .A(net1692));
 sg13g2_buf_4 fanout1690 (.X(net1690),
    .A(net1692));
 sg13g2_buf_2 fanout1691 (.A(net1692),
    .X(net1691));
 sg13g2_buf_2 fanout1692 (.A(\register_file_i/_1931_ ),
    .X(net1692));
 sg13g2_buf_4 fanout1693 (.X(net1693),
    .A(net1694));
 sg13g2_buf_4 fanout1694 (.X(net1694),
    .A(net1698));
 sg13g2_buf_2 fanout1695 (.A(net1698),
    .X(net1695));
 sg13g2_buf_4 fanout1696 (.X(net1696),
    .A(net1698));
 sg13g2_buf_1 fanout1697 (.A(net1698),
    .X(net1697));
 sg13g2_buf_4 fanout1698 (.X(net1698),
    .A(\register_file_i/_1049_ ));
 sg13g2_buf_2 fanout1699 (.A(net1700),
    .X(net1699));
 sg13g2_buf_4 fanout1700 (.X(net1700),
    .A(net1703));
 sg13g2_buf_4 fanout1701 (.X(net1701),
    .A(net1703));
 sg13g2_buf_2 fanout1702 (.A(net1703),
    .X(net1702));
 sg13g2_buf_2 fanout1703 (.A(\register_file_i/_1029_ ),
    .X(net1703));
 sg13g2_buf_2 fanout1704 (.A(_08404_),
    .X(net1704));
 sg13g2_buf_2 fanout1705 (.A(net1706),
    .X(net1705));
 sg13g2_buf_2 fanout1706 (.A(_08390_),
    .X(net1706));
 sg13g2_buf_2 fanout1707 (.A(_08390_),
    .X(net1707));
 sg13g2_buf_2 fanout1708 (.A(_04066_),
    .X(net1708));
 sg13g2_buf_2 fanout1709 (.A(net1710),
    .X(net1709));
 sg13g2_buf_1 fanout1710 (.A(net1711),
    .X(net1710));
 sg13g2_buf_2 fanout1711 (.A(_01840_),
    .X(net1711));
 sg13g2_buf_2 fanout1712 (.A(net1714),
    .X(net1712));
 sg13g2_buf_1 fanout1713 (.A(net1714),
    .X(net1713));
 sg13g2_buf_1 fanout1714 (.A(_01840_),
    .X(net1714));
 sg13g2_buf_2 fanout1715 (.A(_01477_),
    .X(net1715));
 sg13g2_buf_4 fanout1716 (.X(net1716),
    .A(_01198_));
 sg13g2_buf_2 fanout1717 (.A(net1718),
    .X(net1717));
 sg13g2_buf_4 fanout1718 (.X(net1718),
    .A(_01146_));
 sg13g2_buf_4 fanout1719 (.X(net1719),
    .A(net1721));
 sg13g2_buf_4 fanout1720 (.X(net1720),
    .A(net1721));
 sg13g2_buf_4 fanout1721 (.X(net1721),
    .A(\register_file_i/_1968_ ));
 sg13g2_buf_4 fanout1722 (.X(net1722),
    .A(net1723));
 sg13g2_buf_4 fanout1723 (.X(net1723),
    .A(\register_file_i/_1968_ ));
 sg13g2_buf_4 fanout1724 (.X(net1724),
    .A(net1725));
 sg13g2_buf_4 fanout1725 (.X(net1725),
    .A(net1729));
 sg13g2_buf_1 fanout1726 (.A(net1729),
    .X(net1726));
 sg13g2_buf_4 fanout1727 (.X(net1727),
    .A(net1729));
 sg13g2_buf_2 fanout1728 (.A(net1729),
    .X(net1728));
 sg13g2_buf_4 fanout1729 (.X(net1729),
    .A(\register_file_i/_1944_ ));
 sg13g2_buf_4 fanout1730 (.X(net1730),
    .A(net1740));
 sg13g2_buf_4 fanout1731 (.X(net1731),
    .A(net1740));
 sg13g2_buf_4 fanout1732 (.X(net1732),
    .A(net1735));
 sg13g2_buf_4 fanout1733 (.X(net1733),
    .A(net1735));
 sg13g2_buf_2 fanout1734 (.A(net1735),
    .X(net1734));
 sg13g2_buf_4 fanout1735 (.X(net1735),
    .A(net1740));
 sg13g2_buf_4 fanout1736 (.X(net1736),
    .A(net1738));
 sg13g2_buf_4 fanout1737 (.X(net1737),
    .A(net1738));
 sg13g2_buf_4 fanout1738 (.X(net1738),
    .A(net1739));
 sg13g2_buf_4 fanout1739 (.X(net1739),
    .A(net1740));
 sg13g2_buf_4 fanout1740 (.X(net1740),
    .A(\register_file_i/_1916_ ));
 sg13g2_buf_4 fanout1741 (.X(net1741),
    .A(net1751));
 sg13g2_buf_4 fanout1742 (.X(net1742),
    .A(net1751));
 sg13g2_buf_4 fanout1743 (.X(net1743),
    .A(net1746));
 sg13g2_buf_4 fanout1744 (.X(net1744),
    .A(net1746));
 sg13g2_buf_2 fanout1745 (.A(net1746),
    .X(net1745));
 sg13g2_buf_4 fanout1746 (.X(net1746),
    .A(net1751));
 sg13g2_buf_4 fanout1747 (.X(net1747),
    .A(net1749));
 sg13g2_buf_4 fanout1748 (.X(net1748),
    .A(net1749));
 sg13g2_buf_4 fanout1749 (.X(net1749),
    .A(net1750));
 sg13g2_buf_4 fanout1750 (.X(net1750),
    .A(net1751));
 sg13g2_buf_4 fanout1751 (.X(net1751),
    .A(\register_file_i/_1910_ ));
 sg13g2_buf_4 fanout1752 (.X(net1752),
    .A(net1754));
 sg13g2_buf_4 fanout1753 (.X(net1753),
    .A(net1754));
 sg13g2_buf_4 fanout1754 (.X(net1754),
    .A(net1769));
 sg13g2_buf_4 fanout1755 (.X(net1755),
    .A(net1759));
 sg13g2_buf_2 fanout1756 (.A(net1759),
    .X(net1756));
 sg13g2_buf_4 fanout1757 (.X(net1757),
    .A(net1759));
 sg13g2_buf_2 fanout1758 (.A(net1759),
    .X(net1758));
 sg13g2_buf_4 fanout1759 (.X(net1759),
    .A(net1769));
 sg13g2_buf_4 fanout1760 (.X(net1760),
    .A(net1761));
 sg13g2_buf_4 fanout1761 (.X(net1761),
    .A(net1765));
 sg13g2_buf_4 fanout1762 (.X(net1762),
    .A(net1763));
 sg13g2_buf_2 fanout1763 (.A(net1764),
    .X(net1763));
 sg13g2_buf_4 fanout1764 (.X(net1764),
    .A(net1765));
 sg13g2_buf_4 fanout1765 (.X(net1765),
    .A(net1769));
 sg13g2_buf_4 fanout1766 (.X(net1766),
    .A(net1767));
 sg13g2_buf_4 fanout1767 (.X(net1767),
    .A(net1768));
 sg13g2_buf_2 fanout1768 (.A(net1769),
    .X(net1768));
 sg13g2_buf_2 fanout1769 (.A(\register_file_i/_1905_ ),
    .X(net1769));
 sg13g2_buf_4 fanout1770 (.X(net1770),
    .A(net1771));
 sg13g2_buf_4 fanout1771 (.X(net1771),
    .A(net1777));
 sg13g2_buf_4 fanout1772 (.X(net1772),
    .A(net1776));
 sg13g2_buf_2 fanout1773 (.A(net1776),
    .X(net1773));
 sg13g2_buf_4 fanout1774 (.X(net1774),
    .A(net1776));
 sg13g2_buf_2 fanout1775 (.A(net1776),
    .X(net1775));
 sg13g2_buf_4 fanout1776 (.X(net1776),
    .A(net1777));
 sg13g2_buf_4 fanout1777 (.X(net1777),
    .A(\register_file_i/_1896_ ));
 sg13g2_buf_4 fanout1778 (.X(net1778),
    .A(net1779));
 sg13g2_buf_4 fanout1779 (.X(net1779),
    .A(net1783));
 sg13g2_buf_4 fanout1780 (.X(net1780),
    .A(net1782));
 sg13g2_buf_2 fanout1781 (.A(net1782),
    .X(net1781));
 sg13g2_buf_4 fanout1782 (.X(net1782),
    .A(net1783));
 sg13g2_buf_4 fanout1783 (.X(net1783),
    .A(\register_file_i/_1896_ ));
 sg13g2_buf_4 fanout1784 (.X(net1784),
    .A(net1786));
 sg13g2_buf_2 fanout1785 (.A(net1786),
    .X(net1785));
 sg13g2_buf_4 fanout1786 (.X(net1786),
    .A(\register_file_i/_1896_ ));
 sg13g2_buf_4 fanout1787 (.X(net1787),
    .A(net1789));
 sg13g2_buf_4 fanout1788 (.X(net1788),
    .A(net1789));
 sg13g2_buf_4 fanout1789 (.X(net1789),
    .A(\register_file_i/_1066_ ));
 sg13g2_buf_4 fanout1790 (.X(net1790),
    .A(net1791));
 sg13g2_buf_4 fanout1791 (.X(net1791),
    .A(\register_file_i/_1066_ ));
 sg13g2_buf_4 fanout1792 (.X(net1792),
    .A(net1793));
 sg13g2_buf_4 fanout1793 (.X(net1793),
    .A(net1797));
 sg13g2_buf_1 fanout1794 (.A(net1797),
    .X(net1794));
 sg13g2_buf_4 fanout1795 (.X(net1795),
    .A(net1797));
 sg13g2_buf_2 fanout1796 (.A(net1797),
    .X(net1796));
 sg13g2_buf_4 fanout1797 (.X(net1797),
    .A(\register_file_i/_1042_ ));
 sg13g2_buf_4 fanout1798 (.X(net1798),
    .A(net1808));
 sg13g2_buf_4 fanout1799 (.X(net1799),
    .A(net1808));
 sg13g2_buf_4 fanout1800 (.X(net1800),
    .A(net1803));
 sg13g2_buf_4 fanout1801 (.X(net1801),
    .A(net1803));
 sg13g2_buf_2 fanout1802 (.A(net1803),
    .X(net1802));
 sg13g2_buf_4 fanout1803 (.X(net1803),
    .A(net1808));
 sg13g2_buf_4 fanout1804 (.X(net1804),
    .A(net1806));
 sg13g2_buf_4 fanout1805 (.X(net1805),
    .A(net1806));
 sg13g2_buf_4 fanout1806 (.X(net1806),
    .A(net1807));
 sg13g2_buf_4 fanout1807 (.X(net1807),
    .A(net1808));
 sg13g2_buf_4 fanout1808 (.X(net1808),
    .A(\register_file_i/_1014_ ));
 sg13g2_buf_4 fanout1809 (.X(net1809),
    .A(net1819));
 sg13g2_buf_4 fanout1810 (.X(net1810),
    .A(net1819));
 sg13g2_buf_4 fanout1811 (.X(net1811),
    .A(net1814));
 sg13g2_buf_4 fanout1812 (.X(net1812),
    .A(net1814));
 sg13g2_buf_2 fanout1813 (.A(net1814),
    .X(net1813));
 sg13g2_buf_4 fanout1814 (.X(net1814),
    .A(net1819));
 sg13g2_buf_4 fanout1815 (.X(net1815),
    .A(net1817));
 sg13g2_buf_4 fanout1816 (.X(net1816),
    .A(net1817));
 sg13g2_buf_4 fanout1817 (.X(net1817),
    .A(net1818));
 sg13g2_buf_4 fanout1818 (.X(net1818),
    .A(net1819));
 sg13g2_buf_4 fanout1819 (.X(net1819),
    .A(\register_file_i/_1008_ ));
 sg13g2_buf_4 fanout1820 (.X(net1820),
    .A(net1822));
 sg13g2_buf_4 fanout1821 (.X(net1821),
    .A(net1822));
 sg13g2_buf_4 fanout1822 (.X(net1822),
    .A(\register_file_i/_1003_ ));
 sg13g2_buf_4 fanout1823 (.X(net1823),
    .A(net1827));
 sg13g2_buf_2 fanout1824 (.A(net1827),
    .X(net1824));
 sg13g2_buf_4 fanout1825 (.X(net1825),
    .A(net1827));
 sg13g2_buf_2 fanout1826 (.A(net1827),
    .X(net1826));
 sg13g2_buf_2 fanout1827 (.A(\register_file_i/_1003_ ),
    .X(net1827));
 sg13g2_buf_4 fanout1828 (.X(net1828),
    .A(net1829));
 sg13g2_buf_4 fanout1829 (.X(net1829),
    .A(net1836));
 sg13g2_buf_2 fanout1830 (.A(net1836),
    .X(net1830));
 sg13g2_buf_4 fanout1831 (.X(net1831),
    .A(net1832));
 sg13g2_buf_2 fanout1832 (.A(net1833),
    .X(net1832));
 sg13g2_buf_4 fanout1833 (.X(net1833),
    .A(net1836));
 sg13g2_buf_4 fanout1834 (.X(net1834),
    .A(net1835));
 sg13g2_buf_4 fanout1835 (.X(net1835),
    .A(net1836));
 sg13g2_buf_2 fanout1836 (.A(\register_file_i/_1003_ ),
    .X(net1836));
 sg13g2_buf_4 fanout1837 (.X(net1837),
    .A(net1839));
 sg13g2_buf_4 fanout1838 (.X(net1838),
    .A(net1839));
 sg13g2_buf_4 fanout1839 (.X(net1839),
    .A(net1854));
 sg13g2_buf_4 fanout1840 (.X(net1840),
    .A(net1844));
 sg13g2_buf_2 fanout1841 (.A(net1844),
    .X(net1841));
 sg13g2_buf_4 fanout1842 (.X(net1842),
    .A(net1844));
 sg13g2_buf_2 fanout1843 (.A(net1844),
    .X(net1843));
 sg13g2_buf_4 fanout1844 (.X(net1844),
    .A(net1854));
 sg13g2_buf_4 fanout1845 (.X(net1845),
    .A(net1846));
 sg13g2_buf_4 fanout1846 (.X(net1846),
    .A(net1850));
 sg13g2_buf_2 fanout1847 (.A(net1850),
    .X(net1847));
 sg13g2_buf_4 fanout1848 (.X(net1848),
    .A(net1849));
 sg13g2_buf_4 fanout1849 (.X(net1849),
    .A(net1850));
 sg13g2_buf_2 fanout1850 (.A(net1854),
    .X(net1850));
 sg13g2_buf_4 fanout1851 (.X(net1851),
    .A(net1853));
 sg13g2_buf_2 fanout1852 (.A(net1853),
    .X(net1852));
 sg13g2_buf_4 fanout1853 (.X(net1853),
    .A(net1854));
 sg13g2_buf_2 fanout1854 (.A(\register_file_i/_0994_ ),
    .X(net1854));
 sg13g2_buf_4 fanout1855 (.X(net1855),
    .A(net1859));
 sg13g2_buf_2 fanout1856 (.A(net1859),
    .X(net1856));
 sg13g2_buf_4 fanout1857 (.X(net1857),
    .A(net1859));
 sg13g2_buf_2 fanout1858 (.A(net1859),
    .X(net1858));
 sg13g2_buf_2 fanout1859 (.A(net1860),
    .X(net1859));
 sg13g2_buf_4 fanout1860 (.X(net1860),
    .A(_08242_));
 sg13g2_buf_4 fanout1861 (.X(net1861),
    .A(_07475_));
 sg13g2_buf_2 fanout1862 (.A(_07475_),
    .X(net1862));
 sg13g2_buf_2 fanout1863 (.A(net1864),
    .X(net1863));
 sg13g2_buf_1 fanout1864 (.A(_07475_),
    .X(net1864));
 sg13g2_buf_2 fanout1865 (.A(net1868),
    .X(net1865));
 sg13g2_buf_2 fanout1866 (.A(net1868),
    .X(net1866));
 sg13g2_buf_1 fanout1867 (.A(net1868),
    .X(net1867));
 sg13g2_buf_1 fanout1868 (.A(net1871),
    .X(net1868));
 sg13g2_buf_4 fanout1869 (.X(net1869),
    .A(net1871));
 sg13g2_buf_2 fanout1870 (.A(net1871),
    .X(net1870));
 sg13g2_buf_2 fanout1871 (.A(_04056_),
    .X(net1871));
 sg13g2_buf_4 fanout1872 (.X(net1872),
    .A(net1873));
 sg13g2_buf_2 fanout1873 (.A(_04050_),
    .X(net1873));
 sg13g2_buf_2 fanout1874 (.A(net1878),
    .X(net1874));
 sg13g2_buf_1 fanout1875 (.A(net1878),
    .X(net1875));
 sg13g2_buf_2 fanout1876 (.A(net1878),
    .X(net1876));
 sg13g2_buf_2 fanout1877 (.A(net1878),
    .X(net1877));
 sg13g2_buf_1 fanout1878 (.A(_04050_),
    .X(net1878));
 sg13g2_buf_2 fanout1879 (.A(net1880),
    .X(net1879));
 sg13g2_buf_1 fanout1880 (.A(_03330_),
    .X(net1880));
 sg13g2_buf_4 fanout1881 (.X(net1881),
    .A(_01906_));
 sg13g2_buf_2 fanout1882 (.A(net1883),
    .X(net1882));
 sg13g2_buf_2 fanout1883 (.A(_01831_),
    .X(net1883));
 sg13g2_buf_2 fanout1884 (.A(net1887),
    .X(net1884));
 sg13g2_buf_1 fanout1885 (.A(net1887),
    .X(net1885));
 sg13g2_buf_2 fanout1886 (.A(net1887),
    .X(net1886));
 sg13g2_buf_2 fanout1887 (.A(_01831_),
    .X(net1887));
 sg13g2_buf_2 fanout1888 (.A(net1891),
    .X(net1888));
 sg13g2_buf_2 fanout1889 (.A(net1890),
    .X(net1889));
 sg13g2_buf_2 fanout1890 (.A(net1891),
    .X(net1890));
 sg13g2_buf_2 fanout1891 (.A(_01830_),
    .X(net1891));
 sg13g2_buf_2 fanout1892 (.A(net1893),
    .X(net1892));
 sg13g2_buf_2 fanout1893 (.A(net1896),
    .X(net1893));
 sg13g2_buf_2 fanout1894 (.A(net1895),
    .X(net1894));
 sg13g2_buf_1 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_2 fanout1896 (.A(_01826_),
    .X(net1896));
 sg13g2_buf_2 fanout1897 (.A(_01590_),
    .X(net1897));
 sg13g2_buf_2 fanout1898 (.A(_01590_),
    .X(net1898));
 sg13g2_buf_2 fanout1899 (.A(net1901),
    .X(net1899));
 sg13g2_buf_2 fanout1900 (.A(net1901),
    .X(net1900));
 sg13g2_buf_2 fanout1901 (.A(net1902),
    .X(net1901));
 sg13g2_buf_2 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_1 fanout1903 (.A(_01590_),
    .X(net1903));
 sg13g2_buf_2 fanout1904 (.A(_01329_),
    .X(net1904));
 sg13g2_buf_2 fanout1905 (.A(net1906),
    .X(net1905));
 sg13g2_buf_1 fanout1906 (.A(_01155_),
    .X(net1906));
 sg13g2_buf_2 fanout1907 (.A(net1909),
    .X(net1907));
 sg13g2_buf_4 fanout1908 (.X(net1908),
    .A(net1912));
 sg13g2_buf_2 fanout1909 (.A(net1912),
    .X(net1909));
 sg13g2_buf_2 fanout1910 (.A(net1911),
    .X(net1910));
 sg13g2_buf_2 fanout1911 (.A(net1912),
    .X(net1911));
 sg13g2_buf_2 fanout1912 (.A(\register_file_i/_1923_ ),
    .X(net1912));
 sg13g2_buf_2 fanout1913 (.A(net1915),
    .X(net1913));
 sg13g2_buf_2 fanout1914 (.A(net1915),
    .X(net1914));
 sg13g2_buf_4 fanout1915 (.X(net1915),
    .A(\register_file_i/_1920_ ));
 sg13g2_buf_4 fanout1916 (.X(net1916),
    .A(net1918));
 sg13g2_buf_1 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_4 fanout1918 (.X(net1918),
    .A(\register_file_i/_1920_ ));
 sg13g2_buf_2 fanout1919 (.A(net1921),
    .X(net1919));
 sg13g2_buf_4 fanout1920 (.X(net1920),
    .A(net1924));
 sg13g2_buf_2 fanout1921 (.A(net1924),
    .X(net1921));
 sg13g2_buf_2 fanout1922 (.A(net1923),
    .X(net1922));
 sg13g2_buf_2 fanout1923 (.A(net1924),
    .X(net1923));
 sg13g2_buf_2 fanout1924 (.A(\register_file_i/_1021_ ),
    .X(net1924));
 sg13g2_buf_2 fanout1925 (.A(net1927),
    .X(net1925));
 sg13g2_buf_1 fanout1926 (.A(net1927),
    .X(net1926));
 sg13g2_buf_4 fanout1927 (.X(net1927),
    .A(\register_file_i/_1018_ ));
 sg13g2_buf_4 fanout1928 (.X(net1928),
    .A(net1930));
 sg13g2_buf_1 fanout1929 (.A(net1930),
    .X(net1929));
 sg13g2_buf_4 fanout1930 (.X(net1930),
    .A(\register_file_i/_1018_ ));
 sg13g2_buf_2 fanout1931 (.A(net1932),
    .X(net1931));
 sg13g2_buf_2 fanout1932 (.A(_08403_),
    .X(net1932));
 sg13g2_buf_2 fanout1933 (.A(_08403_),
    .X(net1933));
 sg13g2_buf_1 fanout1934 (.A(_08403_),
    .X(net1934));
 sg13g2_buf_2 fanout1935 (.A(net1943),
    .X(net1935));
 sg13g2_buf_1 fanout1936 (.A(net1943),
    .X(net1936));
 sg13g2_buf_2 fanout1937 (.A(net1938),
    .X(net1937));
 sg13g2_buf_2 fanout1938 (.A(net1943),
    .X(net1938));
 sg13g2_buf_2 fanout1939 (.A(net1942),
    .X(net1939));
 sg13g2_buf_2 fanout1940 (.A(net1942),
    .X(net1940));
 sg13g2_buf_1 fanout1941 (.A(net1942),
    .X(net1941));
 sg13g2_buf_1 fanout1942 (.A(net1943),
    .X(net1942));
 sg13g2_buf_1 fanout1943 (.A(_08398_),
    .X(net1943));
 sg13g2_buf_2 fanout1944 (.A(net1947),
    .X(net1944));
 sg13g2_buf_2 fanout1945 (.A(net1947),
    .X(net1945));
 sg13g2_buf_1 fanout1946 (.A(net1947),
    .X(net1946));
 sg13g2_buf_1 fanout1947 (.A(_08395_),
    .X(net1947));
 sg13g2_buf_2 fanout1948 (.A(net1950),
    .X(net1948));
 sg13g2_buf_2 fanout1949 (.A(net1950),
    .X(net1949));
 sg13g2_buf_1 fanout1950 (.A(_08395_),
    .X(net1950));
 sg13g2_buf_2 fanout1951 (.A(net1952),
    .X(net1951));
 sg13g2_buf_1 fanout1952 (.A(net1958),
    .X(net1952));
 sg13g2_buf_2 fanout1953 (.A(net1954),
    .X(net1953));
 sg13g2_buf_2 fanout1954 (.A(net1958),
    .X(net1954));
 sg13g2_buf_2 fanout1955 (.A(net1957),
    .X(net1955));
 sg13g2_buf_2 fanout1956 (.A(net1957),
    .X(net1956));
 sg13g2_buf_2 fanout1957 (.A(net1958),
    .X(net1957));
 sg13g2_buf_1 fanout1958 (.A(_08392_),
    .X(net1958));
 sg13g2_buf_2 fanout1959 (.A(_08388_),
    .X(net1959));
 sg13g2_buf_2 fanout1960 (.A(net1963),
    .X(net1960));
 sg13g2_buf_1 fanout1961 (.A(net1963),
    .X(net1961));
 sg13g2_buf_2 fanout1962 (.A(net1963),
    .X(net1962));
 sg13g2_buf_1 fanout1963 (.A(_08386_),
    .X(net1963));
 sg13g2_buf_4 fanout1964 (.X(net1964),
    .A(net1970));
 sg13g2_buf_4 fanout1965 (.X(net1965),
    .A(net1970));
 sg13g2_buf_4 fanout1966 (.X(net1966),
    .A(net1969));
 sg13g2_buf_2 fanout1967 (.A(net1969),
    .X(net1967));
 sg13g2_buf_4 fanout1968 (.X(net1968),
    .A(net1969));
 sg13g2_buf_1 fanout1969 (.A(net1970),
    .X(net1969));
 sg13g2_buf_2 fanout1970 (.A(_08032_),
    .X(net1970));
 sg13g2_buf_2 fanout1971 (.A(net1975),
    .X(net1971));
 sg13g2_buf_2 fanout1972 (.A(net1975),
    .X(net1972));
 sg13g2_buf_2 fanout1973 (.A(net1975),
    .X(net1973));
 sg13g2_buf_2 fanout1974 (.A(net1975),
    .X(net1974));
 sg13g2_buf_2 fanout1975 (.A(_01536_),
    .X(net1975));
 sg13g2_buf_2 fanout1976 (.A(\load_store_unit_i.pmp_err_q ),
    .X(net1976));
 sg13g2_buf_2 fanout1977 (.A(\load_store_unit_i.ls_fsm_cs_0_ ),
    .X(net1977));
 sg13g2_buf_4 fanout1978 (.X(net1978),
    .A(net1982));
 sg13g2_buf_2 fanout1979 (.A(net1982),
    .X(net1979));
 sg13g2_buf_4 fanout1980 (.X(net1980),
    .A(net1981));
 sg13g2_buf_4 fanout1981 (.X(net1981),
    .A(net1982));
 sg13g2_buf_2 fanout1982 (.A(\if_stage_i.prefetch_buffer_i.fifo_i.valid_q_0_ ),
    .X(net1982));
 sg13g2_buf_2 fanout1983 (.A(net1984),
    .X(net1983));
 sg13g2_buf_1 fanout1984 (.A(net1985),
    .X(net1984));
 sg13g2_buf_2 fanout1985 (.A(\if_stage_i.prefetch_buffer_i.fifo_i.valid_q_0_ ),
    .X(net1985));
 sg13g2_buf_4 fanout1986 (.X(net1986),
    .A(net1987));
 sg13g2_buf_4 fanout1987 (.X(net1987),
    .A(net1990));
 sg13g2_buf_4 fanout1988 (.X(net1988),
    .A(net1989));
 sg13g2_buf_4 fanout1989 (.X(net1989),
    .A(net1990));
 sg13g2_buf_4 fanout1990 (.X(net1990),
    .A(\if_stage_i.prefetch_buffer_i.fifo_busy_1_ ));
 sg13g2_buf_4 fanout1991 (.X(net1991),
    .A(net1992));
 sg13g2_buf_2 fanout1992 (.A(\id_stage_i.controller_i.instr_i_9_ ),
    .X(net1992));
 sg13g2_buf_4 fanout1993 (.X(net1993),
    .A(net1994));
 sg13g2_buf_2 fanout1994 (.A(\id_stage_i.controller_i.instr_i_7_ ),
    .X(net1994));
 sg13g2_buf_2 fanout1995 (.A(\id_stage_i.controller_i.instr_i_6_ ),
    .X(net1995));
 sg13g2_buf_4 fanout1996 (.X(net1996),
    .A(\id_stage_i.controller_i.instr_i_5_ ));
 sg13g2_buf_2 fanout1997 (.A(\id_stage_i.controller_i.instr_i_4_ ),
    .X(net1997));
 sg13g2_buf_2 fanout1998 (.A(\id_stage_i.controller_i.instr_i_3_ ),
    .X(net1998));
 sg13g2_buf_2 fanout1999 (.A(net2001),
    .X(net1999));
 sg13g2_buf_1 fanout2000 (.A(net2001),
    .X(net2000));
 sg13g2_buf_2 fanout2001 (.A(net2002),
    .X(net2001));
 sg13g2_buf_4 fanout2002 (.X(net2002),
    .A(\id_stage_i.controller_i.instr_i_31_ ));
 sg13g2_buf_2 fanout2003 (.A(\id_stage_i.controller_i.instr_i_26_ ),
    .X(net2003));
 sg13g2_buf_2 fanout2004 (.A(net2005),
    .X(net2004));
 sg13g2_buf_1 fanout2005 (.A(net2006),
    .X(net2005));
 sg13g2_buf_2 fanout2006 (.A(\id_stage_i.controller_i.instr_i_25_ ),
    .X(net2006));
 sg13g2_buf_4 fanout2007 (.X(net2007),
    .A(\id_stage_i.controller_i.instr_i_23_ ));
 sg13g2_buf_2 fanout2008 (.A(\id_stage_i.controller_i.instr_i_23_ ),
    .X(net2008));
 sg13g2_buf_4 fanout2009 (.X(net2009),
    .A(\id_stage_i.controller_i.instr_i_18_ ));
 sg13g2_buf_4 fanout2010 (.X(net2010),
    .A(net2019));
 sg13g2_buf_2 fanout2011 (.A(net2019),
    .X(net2011));
 sg13g2_buf_4 fanout2012 (.X(net2012),
    .A(net2013));
 sg13g2_buf_4 fanout2013 (.X(net2013),
    .A(net2019));
 sg13g2_buf_4 fanout2014 (.X(net2014),
    .A(net2016));
 sg13g2_buf_4 fanout2015 (.X(net2015),
    .A(net2018));
 sg13g2_buf_2 fanout2016 (.A(net2018),
    .X(net2016));
 sg13g2_buf_8 fanout2017 (.A(net2018),
    .X(net2017));
 sg13g2_buf_4 fanout2018 (.X(net2018),
    .A(net2019));
 sg13g2_buf_2 fanout2019 (.A(net2030),
    .X(net2019));
 sg13g2_buf_4 fanout2020 (.X(net2020),
    .A(net2021));
 sg13g2_buf_4 fanout2021 (.X(net2021),
    .A(net2030));
 sg13g2_buf_4 fanout2022 (.X(net2022),
    .A(net2024));
 sg13g2_buf_2 fanout2023 (.A(net2024),
    .X(net2023));
 sg13g2_buf_4 fanout2024 (.X(net2024),
    .A(net2030));
 sg13g2_buf_4 fanout2025 (.X(net2025),
    .A(net2029));
 sg13g2_buf_2 fanout2026 (.A(net2029),
    .X(net2026));
 sg13g2_buf_4 fanout2027 (.X(net2027),
    .A(net2029));
 sg13g2_buf_4 fanout2028 (.X(net2028),
    .A(net2029));
 sg13g2_buf_2 fanout2029 (.A(net2030),
    .X(net2029));
 sg13g2_buf_4 fanout2030 (.X(net2030),
    .A(net2085));
 sg13g2_buf_4 fanout2031 (.X(net2031),
    .A(net2033));
 sg13g2_buf_4 fanout2032 (.X(net2032),
    .A(net2033));
 sg13g2_buf_4 fanout2033 (.X(net2033),
    .A(net2041));
 sg13g2_buf_4 fanout2034 (.X(net2034),
    .A(net2041));
 sg13g2_buf_4 fanout2035 (.X(net2035),
    .A(net2041));
 sg13g2_buf_4 fanout2036 (.X(net2036),
    .A(net2040));
 sg13g2_buf_4 fanout2037 (.X(net2037),
    .A(net2040));
 sg13g2_buf_4 fanout2038 (.X(net2038),
    .A(net2039));
 sg13g2_buf_4 fanout2039 (.X(net2039),
    .A(net2040));
 sg13g2_buf_2 fanout2040 (.A(net2041),
    .X(net2040));
 sg13g2_buf_2 fanout2041 (.A(net2085),
    .X(net2041));
 sg13g2_buf_4 fanout2042 (.X(net2042),
    .A(net2052));
 sg13g2_buf_4 fanout2043 (.X(net2043),
    .A(net2052));
 sg13g2_buf_4 fanout2044 (.X(net2044),
    .A(net2046));
 sg13g2_buf_4 fanout2045 (.X(net2045),
    .A(net2046));
 sg13g2_buf_2 fanout2046 (.A(net2052),
    .X(net2046));
 sg13g2_buf_4 fanout2047 (.X(net2047),
    .A(net2048));
 sg13g2_buf_4 fanout2048 (.X(net2048),
    .A(net2052));
 sg13g2_buf_4 fanout2049 (.X(net2049),
    .A(net2051));
 sg13g2_buf_4 fanout2050 (.X(net2050),
    .A(net2051));
 sg13g2_buf_2 fanout2051 (.A(net2052),
    .X(net2051));
 sg13g2_buf_2 fanout2052 (.A(net2085),
    .X(net2052));
 sg13g2_buf_4 fanout2053 (.X(net2053),
    .A(net2055));
 sg13g2_buf_4 fanout2054 (.X(net2054),
    .A(net2055));
 sg13g2_buf_2 fanout2055 (.A(net2059),
    .X(net2055));
 sg13g2_buf_4 fanout2056 (.X(net2056),
    .A(net2058));
 sg13g2_buf_2 fanout2057 (.A(net2058),
    .X(net2057));
 sg13g2_buf_4 fanout2058 (.X(net2058),
    .A(net2059));
 sg13g2_buf_2 fanout2059 (.A(net2065),
    .X(net2059));
 sg13g2_buf_4 fanout2060 (.X(net2060),
    .A(net2065));
 sg13g2_buf_2 fanout2061 (.A(net2065),
    .X(net2061));
 sg13g2_buf_4 fanout2062 (.X(net2062),
    .A(net2064));
 sg13g2_buf_2 fanout2063 (.A(net2064),
    .X(net2063));
 sg13g2_buf_2 fanout2064 (.A(net2065),
    .X(net2064));
 sg13g2_buf_2 fanout2065 (.A(net2084),
    .X(net2065));
 sg13g2_buf_4 fanout2066 (.X(net2066),
    .A(net2067));
 sg13g2_buf_4 fanout2067 (.X(net2067),
    .A(net2071));
 sg13g2_buf_4 fanout2068 (.X(net2068),
    .A(net2070));
 sg13g2_buf_4 fanout2069 (.X(net2069),
    .A(net2070));
 sg13g2_buf_4 fanout2070 (.X(net2070),
    .A(net2071));
 sg13g2_buf_2 fanout2071 (.A(net2084),
    .X(net2071));
 sg13g2_buf_4 fanout2072 (.X(net2072),
    .A(net2073));
 sg13g2_buf_4 fanout2073 (.X(net2073),
    .A(net2075));
 sg13g2_buf_4 fanout2074 (.X(net2074),
    .A(net2075));
 sg13g2_buf_4 fanout2075 (.X(net2075),
    .A(net2084));
 sg13g2_buf_4 fanout2076 (.X(net2076),
    .A(net2080));
 sg13g2_buf_4 fanout2077 (.X(net2077),
    .A(net2080));
 sg13g2_buf_4 fanout2078 (.X(net2078),
    .A(net2080));
 sg13g2_buf_2 fanout2079 (.A(net2080),
    .X(net2079));
 sg13g2_buf_2 fanout2080 (.A(net2081),
    .X(net2080));
 sg13g2_buf_4 fanout2081 (.X(net2081),
    .A(net2084));
 sg13g2_buf_4 fanout2082 (.X(net2082),
    .A(net2083));
 sg13g2_buf_4 fanout2083 (.X(net2083),
    .A(net2084));
 sg13g2_buf_4 fanout2084 (.X(net2084),
    .A(net2085));
 sg13g2_buf_4 fanout2085 (.X(net2085),
    .A(\id_stage_i.controller_i.instr_i_15_ ));
 sg13g2_buf_2 fanout2086 (.A(net2087),
    .X(net2086));
 sg13g2_buf_2 fanout2087 (.A(net2088),
    .X(net2087));
 sg13g2_buf_2 fanout2088 (.A(\id_stage_i.alu_op_b_mux_sel_dec_$_MUX__Y_B_$_OR__Y_A_$_AND__Y_A ),
    .X(net2088));
 sg13g2_buf_2 fanout2089 (.A(net2090),
    .X(net2089));
 sg13g2_buf_1 fanout2090 (.A(net2093),
    .X(net2090));
 sg13g2_buf_2 fanout2091 (.A(net2093),
    .X(net2091));
 sg13g2_buf_1 fanout2092 (.A(net2093),
    .X(net2092));
 sg13g2_buf_4 fanout2093 (.X(net2093),
    .A(\id_stage_i.controller_i.instr_i_14_ ));
 sg13g2_buf_2 fanout2094 (.A(net2095),
    .X(net2094));
 sg13g2_buf_2 fanout2095 (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .X(net2095));
 sg13g2_buf_1 fanout2096 (.A(\div_sel_ex_$_AND__Y_B_$_MUX__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .X(net2096));
 sg13g2_buf_2 fanout2097 (.A(net2098),
    .X(net2097));
 sg13g2_buf_2 fanout2098 (.A(\id_stage_i.controller_i.instr_i_12_ ),
    .X(net2098));
 sg13g2_buf_4 fanout2099 (.X(net2099),
    .A(\id_stage_i.controller_i.instr_i_10_ ));
 sg13g2_buf_2 fanout2100 (.A(net2101),
    .X(net2100));
 sg13g2_buf_1 fanout2101 (.A(\id_stage_i.controller_i.illegal_insn_q ),
    .X(net2101));
 sg13g2_buf_2 fanout2102 (.A(net2103),
    .X(net2102));
 sg13g2_buf_2 fanout2103 (.A(\csr_save_id_$_AND__Y_B_$_NOT__Y_A_$_OR__Y_A_$_OR__Y_A ),
    .X(net2103));
 sg13g2_buf_2 fanout2104 (.A(\id_stage_i.controller_i.ctrl_fsm_cs_0_ ),
    .X(net2104));
 sg13g2_buf_2 fanout2105 (.A(net2106),
    .X(net2105));
 sg13g2_buf_2 fanout2106 (.A(net2107),
    .X(net2106));
 sg13g2_buf_4 fanout2107 (.X(net2107),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2_ ));
 sg13g2_buf_2 fanout2108 (.A(net2109),
    .X(net2108));
 sg13g2_buf_2 fanout2109 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_2_ ),
    .X(net2109));
 sg13g2_buf_2 fanout2110 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_1_ ),
    .X(net2110));
 sg13g2_buf_2 fanout2111 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.md_state_q_0_ ),
    .X(net2111));
 sg13g2_buf_4 fanout2112 (.X(net2112),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_q_3_ ));
 sg13g2_buf_4 fanout2113 (.X(net2113),
    .A(\ex_block_i.gen_multdiv_fast.multdiv_i.div_counter_d_4__$_MUX__Y_A_$_XOR__Y_B_$_OR__Y_B_$_AND__Y_B_$_OR__Y_B_$_AND__Y_A ));
 sg13g2_buf_4 fanout2114 (.X(net2114),
    .A(\ex_block_i.alu_i.imd_val_q_i_44_ ));
 sg13g2_buf_4 fanout2115 (.X(net2115),
    .A(\ex_block_i.alu_i.imd_val_q_i_41_ ));
 sg13g2_buf_2 fanout2116 (.A(\id_stage_i.controller_i.priv_mode_i_1_ ),
    .X(net2116));
 sg13g2_buf_4 fanout2117 (.X(net2117),
    .A(net2119));
 sg13g2_buf_2 fanout2118 (.A(net2119),
    .X(net2118));
 sg13g2_buf_2 fanout2119 (.A(net2123),
    .X(net2119));
 sg13g2_buf_4 fanout2120 (.X(net2120),
    .A(net2123));
 sg13g2_buf_4 fanout2121 (.X(net2121),
    .A(net2123));
 sg13g2_buf_4 fanout2122 (.X(net2122),
    .A(net2123));
 sg13g2_buf_2 fanout2123 (.A(net2155),
    .X(net2123));
 sg13g2_buf_4 fanout2124 (.X(net2124),
    .A(net2128));
 sg13g2_buf_4 fanout2125 (.X(net2125),
    .A(net2128));
 sg13g2_buf_4 fanout2126 (.X(net2126),
    .A(net2127));
 sg13g2_buf_4 fanout2127 (.X(net2127),
    .A(net2128));
 sg13g2_buf_2 fanout2128 (.A(net2155),
    .X(net2128));
 sg13g2_buf_4 fanout2129 (.X(net2129),
    .A(net2133));
 sg13g2_buf_4 fanout2130 (.X(net2130),
    .A(net2133));
 sg13g2_buf_4 fanout2131 (.X(net2131),
    .A(net2133));
 sg13g2_buf_2 fanout2132 (.A(net2133),
    .X(net2132));
 sg13g2_buf_2 fanout2133 (.A(net2155),
    .X(net2133));
 sg13g2_buf_4 fanout2134 (.X(net2134),
    .A(net2138));
 sg13g2_buf_2 fanout2135 (.A(net2138),
    .X(net2135));
 sg13g2_buf_4 fanout2136 (.X(net2136),
    .A(net2138));
 sg13g2_buf_4 fanout2137 (.X(net2137),
    .A(net2138));
 sg13g2_buf_1 fanout2138 (.A(net2154),
    .X(net2138));
 sg13g2_buf_4 fanout2139 (.X(net2139),
    .A(net2143));
 sg13g2_buf_4 fanout2140 (.X(net2140),
    .A(net2143));
 sg13g2_buf_4 fanout2141 (.X(net2141),
    .A(net2143));
 sg13g2_buf_4 fanout2142 (.X(net2142),
    .A(net2143));
 sg13g2_buf_2 fanout2143 (.A(net2154),
    .X(net2143));
 sg13g2_buf_4 fanout2144 (.X(net2144),
    .A(net2145));
 sg13g2_buf_4 fanout2145 (.X(net2145),
    .A(net2148));
 sg13g2_buf_4 fanout2146 (.X(net2146),
    .A(net2147));
 sg13g2_buf_4 fanout2147 (.X(net2147),
    .A(net2148));
 sg13g2_buf_2 fanout2148 (.A(net2154),
    .X(net2148));
 sg13g2_buf_4 fanout2149 (.X(net2149),
    .A(net2153));
 sg13g2_buf_4 fanout2150 (.X(net2150),
    .A(net2153));
 sg13g2_buf_4 fanout2151 (.X(net2151),
    .A(net2153));
 sg13g2_buf_4 fanout2152 (.X(net2152),
    .A(net2153));
 sg13g2_buf_2 fanout2153 (.A(net2154),
    .X(net2153));
 sg13g2_buf_2 fanout2154 (.A(net2155),
    .X(net2154));
 sg13g2_buf_2 fanout2155 (.A(net2274),
    .X(net2155));
 sg13g2_buf_4 fanout2156 (.X(net2156),
    .A(net2160));
 sg13g2_buf_4 fanout2157 (.X(net2157),
    .A(net2160));
 sg13g2_buf_4 fanout2158 (.X(net2158),
    .A(net2160));
 sg13g2_buf_4 fanout2159 (.X(net2159),
    .A(net2160));
 sg13g2_buf_2 fanout2160 (.A(net2176),
    .X(net2160));
 sg13g2_buf_4 fanout2161 (.X(net2161),
    .A(net2165));
 sg13g2_buf_2 fanout2162 (.A(net2165),
    .X(net2162));
 sg13g2_buf_4 fanout2163 (.X(net2163),
    .A(net2165));
 sg13g2_buf_4 fanout2164 (.X(net2164),
    .A(net2165));
 sg13g2_buf_1 fanout2165 (.A(net2176),
    .X(net2165));
 sg13g2_buf_4 fanout2166 (.X(net2166),
    .A(net2167));
 sg13g2_buf_4 fanout2167 (.X(net2167),
    .A(net2170));
 sg13g2_buf_4 fanout2168 (.X(net2168),
    .A(net2170));
 sg13g2_buf_4 fanout2169 (.X(net2169),
    .A(net2170));
 sg13g2_buf_4 fanout2170 (.X(net2170),
    .A(net2176));
 sg13g2_buf_4 fanout2171 (.X(net2171),
    .A(net2175));
 sg13g2_buf_4 fanout2172 (.X(net2172),
    .A(net2175));
 sg13g2_buf_4 fanout2173 (.X(net2173),
    .A(net2175));
 sg13g2_buf_2 fanout2174 (.A(net2175),
    .X(net2174));
 sg13g2_buf_2 fanout2175 (.A(net2176),
    .X(net2175));
 sg13g2_buf_2 fanout2176 (.A(net2197),
    .X(net2176));
 sg13g2_buf_4 fanout2177 (.X(net2177),
    .A(net2186));
 sg13g2_buf_4 fanout2178 (.X(net2178),
    .A(net2186));
 sg13g2_buf_4 fanout2179 (.X(net2179),
    .A(net2180));
 sg13g2_buf_4 fanout2180 (.X(net2180),
    .A(net2186));
 sg13g2_buf_4 fanout2181 (.X(net2181),
    .A(net2185));
 sg13g2_buf_4 fanout2182 (.X(net2182),
    .A(net2185));
 sg13g2_buf_4 fanout2183 (.X(net2183),
    .A(net2184));
 sg13g2_buf_4 fanout2184 (.X(net2184),
    .A(net2185));
 sg13g2_buf_2 fanout2185 (.A(net2186),
    .X(net2185));
 sg13g2_buf_2 fanout2186 (.A(net2197),
    .X(net2186));
 sg13g2_buf_4 fanout2187 (.X(net2187),
    .A(net2191));
 sg13g2_buf_2 fanout2188 (.A(net2191),
    .X(net2188));
 sg13g2_buf_4 fanout2189 (.X(net2189),
    .A(net2191));
 sg13g2_buf_4 fanout2190 (.X(net2190),
    .A(net2191));
 sg13g2_buf_1 fanout2191 (.A(net2197),
    .X(net2191));
 sg13g2_buf_4 fanout2192 (.X(net2192),
    .A(net2196));
 sg13g2_buf_2 fanout2193 (.A(net2196),
    .X(net2193));
 sg13g2_buf_4 fanout2194 (.X(net2194),
    .A(net2196));
 sg13g2_buf_4 fanout2195 (.X(net2195),
    .A(net2196));
 sg13g2_buf_2 fanout2196 (.A(net2197),
    .X(net2196));
 sg13g2_buf_2 fanout2197 (.A(net2274),
    .X(net2197));
 sg13g2_buf_4 fanout2198 (.X(net2198),
    .A(net2202));
 sg13g2_buf_2 fanout2199 (.A(net2202),
    .X(net2199));
 sg13g2_buf_4 fanout2200 (.X(net2200),
    .A(net2202));
 sg13g2_buf_4 fanout2201 (.X(net2201),
    .A(net2202));
 sg13g2_buf_2 fanout2202 (.A(net2218),
    .X(net2202));
 sg13g2_buf_4 fanout2203 (.X(net2203),
    .A(net2207));
 sg13g2_buf_4 fanout2204 (.X(net2204),
    .A(net2207));
 sg13g2_buf_4 fanout2205 (.X(net2205),
    .A(net2207));
 sg13g2_buf_4 fanout2206 (.X(net2206),
    .A(net2207));
 sg13g2_buf_2 fanout2207 (.A(net2218),
    .X(net2207));
 sg13g2_buf_4 fanout2208 (.X(net2208),
    .A(net2212));
 sg13g2_buf_4 fanout2209 (.X(net2209),
    .A(net2212));
 sg13g2_buf_4 fanout2210 (.X(net2210),
    .A(net2212));
 sg13g2_buf_2 fanout2211 (.A(net2212),
    .X(net2211));
 sg13g2_buf_2 fanout2212 (.A(net2218),
    .X(net2212));
 sg13g2_buf_4 fanout2213 (.X(net2213),
    .A(net2214));
 sg13g2_buf_4 fanout2214 (.X(net2214),
    .A(net2217));
 sg13g2_buf_4 fanout2215 (.X(net2215),
    .A(net2217));
 sg13g2_buf_2 fanout2216 (.A(net2217),
    .X(net2216));
 sg13g2_buf_2 fanout2217 (.A(net2218),
    .X(net2217));
 sg13g2_buf_2 fanout2218 (.A(net2274),
    .X(net2218));
 sg13g2_buf_4 fanout2219 (.X(net2219),
    .A(net2223));
 sg13g2_buf_4 fanout2220 (.X(net2220),
    .A(net2223));
 sg13g2_buf_4 fanout2221 (.X(net2221),
    .A(net2223));
 sg13g2_buf_4 fanout2222 (.X(net2222),
    .A(net2223));
 sg13g2_buf_2 fanout2223 (.A(net2238),
    .X(net2223));
 sg13g2_buf_4 fanout2224 (.X(net2224),
    .A(net2227));
 sg13g2_buf_4 fanout2225 (.X(net2225),
    .A(net2227));
 sg13g2_buf_2 fanout2226 (.A(net2227),
    .X(net2226));
 sg13g2_buf_2 fanout2227 (.A(net2238),
    .X(net2227));
 sg13g2_buf_4 fanout2228 (.X(net2228),
    .A(net2232));
 sg13g2_buf_4 fanout2229 (.X(net2229),
    .A(net2232));
 sg13g2_buf_4 fanout2230 (.X(net2230),
    .A(net2232));
 sg13g2_buf_4 fanout2231 (.X(net2231),
    .A(net2232));
 sg13g2_buf_2 fanout2232 (.A(net2238),
    .X(net2232));
 sg13g2_buf_4 fanout2233 (.X(net2233),
    .A(net2237));
 sg13g2_buf_4 fanout2234 (.X(net2234),
    .A(net2237));
 sg13g2_buf_4 fanout2235 (.X(net2235),
    .A(net2237));
 sg13g2_buf_4 fanout2236 (.X(net2236),
    .A(net2237));
 sg13g2_buf_2 fanout2237 (.A(net2238),
    .X(net2237));
 sg13g2_buf_2 fanout2238 (.A(net2274),
    .X(net2238));
 sg13g2_buf_4 fanout2239 (.X(net2239),
    .A(net2242));
 sg13g2_buf_4 fanout2240 (.X(net2240),
    .A(net2242));
 sg13g2_buf_4 fanout2241 (.X(net2241),
    .A(net2242));
 sg13g2_buf_4 fanout2242 (.X(net2242),
    .A(net2273));
 sg13g2_buf_4 fanout2243 (.X(net2243),
    .A(net2247));
 sg13g2_buf_2 fanout2244 (.A(net2247),
    .X(net2244));
 sg13g2_buf_4 fanout2245 (.X(net2245),
    .A(net2247));
 sg13g2_buf_2 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_1 fanout2247 (.A(net2273),
    .X(net2247));
 sg13g2_buf_4 fanout2248 (.X(net2248),
    .A(net2257));
 sg13g2_buf_2 fanout2249 (.A(net2257),
    .X(net2249));
 sg13g2_buf_4 fanout2250 (.X(net2250),
    .A(net2251));
 sg13g2_buf_4 fanout2251 (.X(net2251),
    .A(net2257));
 sg13g2_buf_4 fanout2252 (.X(net2252),
    .A(net2253));
 sg13g2_buf_4 fanout2253 (.X(net2253),
    .A(net2256));
 sg13g2_buf_4 fanout2254 (.X(net2254),
    .A(net2256));
 sg13g2_buf_2 fanout2255 (.A(net2256),
    .X(net2255));
 sg13g2_buf_2 fanout2256 (.A(net2257),
    .X(net2256));
 sg13g2_buf_2 fanout2257 (.A(net2273),
    .X(net2257));
 sg13g2_buf_4 fanout2258 (.X(net2258),
    .A(net2259));
 sg13g2_buf_4 fanout2259 (.X(net2259),
    .A(net2272));
 sg13g2_buf_2 fanout2260 (.A(net2272),
    .X(net2260));
 sg13g2_buf_4 fanout2261 (.X(net2261),
    .A(net2265));
 sg13g2_buf_4 fanout2262 (.X(net2262),
    .A(net2265));
 sg13g2_buf_4 fanout2263 (.X(net2263),
    .A(net2264));
 sg13g2_buf_4 fanout2264 (.X(net2264),
    .A(net2265));
 sg13g2_buf_2 fanout2265 (.A(net2272),
    .X(net2265));
 sg13g2_buf_4 fanout2266 (.X(net2266),
    .A(net2267));
 sg13g2_buf_4 fanout2267 (.X(net2267),
    .A(net2268));
 sg13g2_buf_4 fanout2268 (.X(net2268),
    .A(net2272));
 sg13g2_buf_4 fanout2269 (.X(net2269),
    .A(net2270));
 sg13g2_buf_4 fanout2270 (.X(net2270),
    .A(net2271));
 sg13g2_buf_4 fanout2271 (.X(net2271),
    .A(net2272));
 sg13g2_buf_2 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_2 fanout2273 (.A(net2274),
    .X(net2273));
 sg13g2_buf_4 fanout2274 (.X(net2274),
    .A(net2465));
 sg13g2_buf_4 fanout2275 (.X(net2275),
    .A(net2277));
 sg13g2_buf_4 fanout2276 (.X(net2276),
    .A(net2277));
 sg13g2_buf_2 fanout2277 (.A(net2284),
    .X(net2277));
 sg13g2_buf_4 fanout2278 (.X(net2278),
    .A(net2284));
 sg13g2_buf_4 fanout2279 (.X(net2279),
    .A(net2284));
 sg13g2_buf_4 fanout2280 (.X(net2280),
    .A(net2283));
 sg13g2_buf_4 fanout2281 (.X(net2281),
    .A(net2283));
 sg13g2_buf_4 fanout2282 (.X(net2282),
    .A(net2283));
 sg13g2_buf_2 fanout2283 (.A(net2284),
    .X(net2283));
 sg13g2_buf_2 fanout2284 (.A(net2318),
    .X(net2284));
 sg13g2_buf_4 fanout2285 (.X(net2285),
    .A(net2289));
 sg13g2_buf_4 fanout2286 (.X(net2286),
    .A(net2287));
 sg13g2_buf_4 fanout2287 (.X(net2287),
    .A(net2288));
 sg13g2_buf_2 fanout2288 (.A(net2289),
    .X(net2288));
 sg13g2_buf_2 fanout2289 (.A(net2318),
    .X(net2289));
 sg13g2_buf_4 fanout2290 (.X(net2290),
    .A(net2293));
 sg13g2_buf_4 fanout2291 (.X(net2291),
    .A(net2293));
 sg13g2_buf_4 fanout2292 (.X(net2292),
    .A(net2293));
 sg13g2_buf_2 fanout2293 (.A(net2301),
    .X(net2293));
 sg13g2_buf_4 fanout2294 (.X(net2294),
    .A(net2298));
 sg13g2_buf_4 fanout2295 (.X(net2295),
    .A(net2298));
 sg13g2_buf_4 fanout2296 (.X(net2296),
    .A(net2298));
 sg13g2_buf_2 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_2 fanout2298 (.A(net2301),
    .X(net2298));
 sg13g2_buf_4 fanout2299 (.X(net2299),
    .A(net2301));
 sg13g2_buf_2 fanout2300 (.A(net2301),
    .X(net2300));
 sg13g2_buf_2 fanout2301 (.A(net2318),
    .X(net2301));
 sg13g2_buf_4 fanout2302 (.X(net2302),
    .A(net2317));
 sg13g2_buf_4 fanout2303 (.X(net2303),
    .A(net2317));
 sg13g2_buf_4 fanout2304 (.X(net2304),
    .A(net2307));
 sg13g2_buf_4 fanout2305 (.X(net2305),
    .A(net2307));
 sg13g2_buf_4 fanout2306 (.X(net2306),
    .A(net2307));
 sg13g2_buf_2 fanout2307 (.A(net2308),
    .X(net2307));
 sg13g2_buf_4 fanout2308 (.X(net2308),
    .A(net2317));
 sg13g2_buf_4 fanout2309 (.X(net2309),
    .A(net2311));
 sg13g2_buf_2 fanout2310 (.A(net2311),
    .X(net2310));
 sg13g2_buf_4 fanout2311 (.X(net2311),
    .A(net2316));
 sg13g2_buf_4 fanout2312 (.X(net2312),
    .A(net2316));
 sg13g2_buf_4 fanout2313 (.X(net2313),
    .A(net2315));
 sg13g2_buf_4 fanout2314 (.X(net2314),
    .A(net2315));
 sg13g2_buf_2 fanout2315 (.A(net2316),
    .X(net2315));
 sg13g2_buf_2 fanout2316 (.A(net2317),
    .X(net2316));
 sg13g2_buf_2 fanout2317 (.A(net2318),
    .X(net2317));
 sg13g2_buf_4 fanout2318 (.X(net2318),
    .A(net2465));
 sg13g2_buf_4 fanout2319 (.X(net2319),
    .A(net2320));
 sg13g2_buf_4 fanout2320 (.X(net2320),
    .A(net2322));
 sg13g2_buf_4 fanout2321 (.X(net2321),
    .A(net2322));
 sg13g2_buf_4 fanout2322 (.X(net2322),
    .A(net2348));
 sg13g2_buf_4 fanout2323 (.X(net2323),
    .A(net2348));
 sg13g2_buf_4 fanout2324 (.X(net2324),
    .A(net2325));
 sg13g2_buf_4 fanout2325 (.X(net2325),
    .A(net2326));
 sg13g2_buf_4 fanout2326 (.X(net2326),
    .A(net2337));
 sg13g2_buf_4 fanout2327 (.X(net2327),
    .A(net2329));
 sg13g2_buf_4 fanout2328 (.X(net2328),
    .A(net2329));
 sg13g2_buf_4 fanout2329 (.X(net2329),
    .A(net2330));
 sg13g2_buf_4 fanout2330 (.X(net2330),
    .A(net2337));
 sg13g2_buf_4 fanout2331 (.X(net2331),
    .A(net2335));
 sg13g2_buf_2 fanout2332 (.A(net2335),
    .X(net2332));
 sg13g2_buf_4 fanout2333 (.X(net2333),
    .A(net2335));
 sg13g2_buf_2 fanout2334 (.A(net2335),
    .X(net2334));
 sg13g2_buf_1 fanout2335 (.A(net2337),
    .X(net2335));
 sg13g2_buf_4 fanout2336 (.X(net2336),
    .A(net2337));
 sg13g2_buf_4 fanout2337 (.X(net2337),
    .A(net2348));
 sg13g2_buf_4 fanout2338 (.X(net2338),
    .A(net2339));
 sg13g2_buf_4 fanout2339 (.X(net2339),
    .A(net2347));
 sg13g2_buf_4 fanout2340 (.X(net2340),
    .A(net2343));
 sg13g2_buf_4 fanout2341 (.X(net2341),
    .A(net2343));
 sg13g2_buf_4 fanout2342 (.X(net2342),
    .A(net2347));
 sg13g2_buf_2 fanout2343 (.A(net2347),
    .X(net2343));
 sg13g2_buf_4 fanout2344 (.X(net2344),
    .A(net2346));
 sg13g2_buf_4 fanout2345 (.X(net2345),
    .A(net2346));
 sg13g2_buf_4 fanout2346 (.X(net2346),
    .A(net2347));
 sg13g2_buf_2 fanout2347 (.A(net2348),
    .X(net2347));
 sg13g2_buf_4 fanout2348 (.X(net2348),
    .A(net2465));
 sg13g2_buf_4 fanout2349 (.X(net2349),
    .A(net2351));
 sg13g2_buf_4 fanout2350 (.X(net2350),
    .A(net2351));
 sg13g2_buf_2 fanout2351 (.A(net2357),
    .X(net2351));
 sg13g2_buf_4 fanout2352 (.X(net2352),
    .A(net2353));
 sg13g2_buf_4 fanout2353 (.X(net2353),
    .A(net2357));
 sg13g2_buf_4 fanout2354 (.X(net2354),
    .A(net2356));
 sg13g2_buf_4 fanout2355 (.X(net2355),
    .A(net2356));
 sg13g2_buf_4 fanout2356 (.X(net2356),
    .A(net2357));
 sg13g2_buf_2 fanout2357 (.A(net2394),
    .X(net2357));
 sg13g2_buf_4 fanout2358 (.X(net2358),
    .A(net2382));
 sg13g2_buf_4 fanout2359 (.X(net2359),
    .A(net2382));
 sg13g2_buf_4 fanout2360 (.X(net2360),
    .A(net2365));
 sg13g2_buf_4 fanout2361 (.X(net2361),
    .A(net2365));
 sg13g2_buf_4 fanout2362 (.X(net2362),
    .A(net2364));
 sg13g2_buf_2 fanout2363 (.A(net2364),
    .X(net2363));
 sg13g2_buf_4 fanout2364 (.X(net2364),
    .A(net2365));
 sg13g2_buf_2 fanout2365 (.A(net2382),
    .X(net2365));
 sg13g2_buf_4 fanout2366 (.X(net2366),
    .A(net2369));
 sg13g2_buf_2 fanout2367 (.A(net2369),
    .X(net2367));
 sg13g2_buf_4 fanout2368 (.X(net2368),
    .A(net2369));
 sg13g2_buf_2 fanout2369 (.A(net2381),
    .X(net2369));
 sg13g2_buf_4 fanout2370 (.X(net2370),
    .A(net2372));
 sg13g2_buf_2 fanout2371 (.A(net2372),
    .X(net2371));
 sg13g2_buf_2 fanout2372 (.A(net2381),
    .X(net2372));
 sg13g2_buf_4 fanout2373 (.X(net2373),
    .A(net2377));
 sg13g2_buf_2 fanout2374 (.A(net2377),
    .X(net2374));
 sg13g2_buf_4 fanout2375 (.X(net2375),
    .A(net2377));
 sg13g2_buf_2 fanout2376 (.A(net2377),
    .X(net2376));
 sg13g2_buf_1 fanout2377 (.A(net2381),
    .X(net2377));
 sg13g2_buf_4 fanout2378 (.X(net2378),
    .A(net2379));
 sg13g2_buf_4 fanout2379 (.X(net2379),
    .A(net2380));
 sg13g2_buf_4 fanout2380 (.X(net2380),
    .A(net2381));
 sg13g2_buf_2 fanout2381 (.A(net2382),
    .X(net2381));
 sg13g2_buf_2 fanout2382 (.A(net2394),
    .X(net2382));
 sg13g2_buf_4 fanout2383 (.X(net2383),
    .A(net2394));
 sg13g2_buf_4 fanout2384 (.X(net2384),
    .A(net2385));
 sg13g2_buf_4 fanout2385 (.X(net2385),
    .A(net2386));
 sg13g2_buf_4 fanout2386 (.X(net2386),
    .A(net2393));
 sg13g2_buf_4 fanout2387 (.X(net2387),
    .A(net2389));
 sg13g2_buf_4 fanout2388 (.X(net2388),
    .A(net2393));
 sg13g2_buf_4 fanout2389 (.X(net2389),
    .A(net2393));
 sg13g2_buf_4 fanout2390 (.X(net2390),
    .A(net2391));
 sg13g2_buf_4 fanout2391 (.X(net2391),
    .A(net2393));
 sg13g2_buf_4 fanout2392 (.X(net2392),
    .A(net2393));
 sg13g2_buf_4 fanout2393 (.X(net2393),
    .A(net2394));
 sg13g2_buf_2 fanout2394 (.A(net2465),
    .X(net2394));
 sg13g2_buf_4 fanout2395 (.X(net2395),
    .A(net2398));
 sg13g2_buf_2 fanout2396 (.A(net2398),
    .X(net2396));
 sg13g2_buf_4 fanout2397 (.X(net2397),
    .A(net2398));
 sg13g2_buf_2 fanout2398 (.A(net2425),
    .X(net2398));
 sg13g2_buf_4 fanout2399 (.X(net2399),
    .A(net2402));
 sg13g2_buf_4 fanout2400 (.X(net2400),
    .A(net2402));
 sg13g2_buf_4 fanout2401 (.X(net2401),
    .A(net2402));
 sg13g2_buf_2 fanout2402 (.A(net2425),
    .X(net2402));
 sg13g2_buf_4 fanout2403 (.X(net2403),
    .A(net2409));
 sg13g2_buf_4 fanout2404 (.X(net2404),
    .A(net2405));
 sg13g2_buf_4 fanout2405 (.X(net2405),
    .A(net2409));
 sg13g2_buf_4 fanout2406 (.X(net2406),
    .A(net2408));
 sg13g2_buf_2 fanout2407 (.A(net2408),
    .X(net2407));
 sg13g2_buf_4 fanout2408 (.X(net2408),
    .A(net2409));
 sg13g2_buf_2 fanout2409 (.A(net2425),
    .X(net2409));
 sg13g2_buf_4 fanout2410 (.X(net2410),
    .A(net2413));
 sg13g2_buf_2 fanout2411 (.A(net2413),
    .X(net2411));
 sg13g2_buf_4 fanout2412 (.X(net2412),
    .A(net2413));
 sg13g2_buf_2 fanout2413 (.A(net2414),
    .X(net2413));
 sg13g2_buf_4 fanout2414 (.X(net2414),
    .A(net2424));
 sg13g2_buf_4 fanout2415 (.X(net2415),
    .A(net2416));
 sg13g2_buf_4 fanout2416 (.X(net2416),
    .A(net2419));
 sg13g2_buf_4 fanout2417 (.X(net2417),
    .A(net2419));
 sg13g2_buf_4 fanout2418 (.X(net2418),
    .A(net2419));
 sg13g2_buf_2 fanout2419 (.A(net2424),
    .X(net2419));
 sg13g2_buf_4 fanout2420 (.X(net2420),
    .A(net2422));
 sg13g2_buf_4 fanout2421 (.X(net2421),
    .A(net2422));
 sg13g2_buf_2 fanout2422 (.A(net2424),
    .X(net2422));
 sg13g2_buf_4 fanout2423 (.X(net2423),
    .A(net2424));
 sg13g2_buf_2 fanout2424 (.A(net2425),
    .X(net2424));
 sg13g2_buf_2 fanout2425 (.A(net2436),
    .X(net2425));
 sg13g2_buf_4 fanout2426 (.X(net2426),
    .A(net2436));
 sg13g2_buf_4 fanout2427 (.X(net2427),
    .A(net2428));
 sg13g2_buf_4 fanout2428 (.X(net2428),
    .A(net2429));
 sg13g2_buf_4 fanout2429 (.X(net2429),
    .A(net2436));
 sg13g2_buf_4 fanout2430 (.X(net2430),
    .A(net2431));
 sg13g2_buf_4 fanout2431 (.X(net2431),
    .A(net2434));
 sg13g2_buf_4 fanout2432 (.X(net2432),
    .A(net2433));
 sg13g2_buf_4 fanout2433 (.X(net2433),
    .A(net2434));
 sg13g2_buf_2 fanout2434 (.A(net2435),
    .X(net2434));
 sg13g2_buf_4 fanout2435 (.X(net2435),
    .A(net2436));
 sg13g2_buf_4 fanout2436 (.X(net2436),
    .A(net2465));
 sg13g2_buf_4 fanout2437 (.X(net2437),
    .A(net2441));
 sg13g2_buf_4 fanout2438 (.X(net2438),
    .A(net2441));
 sg13g2_buf_4 fanout2439 (.X(net2439),
    .A(net2441));
 sg13g2_buf_4 fanout2440 (.X(net2440),
    .A(net2441));
 sg13g2_buf_4 fanout2441 (.X(net2441),
    .A(net2464));
 sg13g2_buf_4 fanout2442 (.X(net2442),
    .A(net2443));
 sg13g2_buf_2 fanout2443 (.A(net2451),
    .X(net2443));
 sg13g2_buf_4 fanout2444 (.X(net2444),
    .A(net2451));
 sg13g2_buf_4 fanout2445 (.X(net2445),
    .A(net2451));
 sg13g2_buf_4 fanout2446 (.X(net2446),
    .A(net2451));
 sg13g2_buf_4 fanout2447 (.X(net2447),
    .A(net2451));
 sg13g2_buf_4 fanout2448 (.X(net2448),
    .A(net2450));
 sg13g2_buf_4 fanout2449 (.X(net2449),
    .A(net2450));
 sg13g2_buf_2 fanout2450 (.A(net2451),
    .X(net2450));
 sg13g2_buf_2 fanout2451 (.A(net2464),
    .X(net2451));
 sg13g2_buf_4 fanout2452 (.X(net2452),
    .A(net2454));
 sg13g2_buf_4 fanout2453 (.X(net2453),
    .A(net2454));
 sg13g2_buf_2 fanout2454 (.A(net2459),
    .X(net2454));
 sg13g2_buf_4 fanout2455 (.X(net2455),
    .A(net2459));
 sg13g2_buf_4 fanout2456 (.X(net2456),
    .A(net2459));
 sg13g2_buf_4 fanout2457 (.X(net2457),
    .A(net2458));
 sg13g2_buf_4 fanout2458 (.X(net2458),
    .A(net2459));
 sg13g2_buf_2 fanout2459 (.A(net2463),
    .X(net2459));
 sg13g2_buf_4 fanout2460 (.X(net2460),
    .A(net2462));
 sg13g2_buf_2 fanout2461 (.A(net2462),
    .X(net2461));
 sg13g2_buf_4 fanout2462 (.X(net2462),
    .A(net2463));
 sg13g2_buf_2 fanout2463 (.A(net2464),
    .X(net2463));
 sg13g2_buf_4 fanout2464 (.X(net2464),
    .A(net2465));
 sg13g2_buf_8 fanout2465 (.A(rst_ni),
    .X(net2465));
 sg13g2_buf_2 fanout2466 (.A(data_rvalid_i),
    .X(net2466));
 sg13g2_dlygate4sd1_1 rebuffer2470 (.A(_03646_),
    .X(net2470));
 sg13g2_xnor2_1 clone2487 (.Y(net2487),
    .A(_01926_),
    .B(_02868_));
 sg13g2_buf_8 rebuffer2488 (.A(_03375_),
    .X(net2488));
 sg13g2_buf_1 rebuffer2489 (.A(net2488),
    .X(net2489));
 sg13g2_buf_16 clkbuf_leaf_0_clk_i (.X(clknet_leaf_0_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_1_clk_i (.X(clknet_leaf_1_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_2_clk_i (.X(clknet_leaf_2_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_3_clk_i (.X(clknet_leaf_3_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_4_clk_i (.X(clknet_leaf_4_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_5_clk_i (.X(clknet_leaf_5_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_6_clk_i (.X(clknet_leaf_6_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_7_clk_i (.X(clknet_leaf_7_clk_i),
    .A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_8_clk_i (.X(clknet_leaf_8_clk_i),
    .A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_9_clk_i (.X(clknet_leaf_9_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_10_clk_i (.X(clknet_leaf_10_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_11_clk_i (.X(clknet_leaf_11_clk_i),
    .A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_12_clk_i (.X(clknet_leaf_12_clk_i),
    .A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_13_clk_i (.X(clknet_leaf_13_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_14_clk_i (.X(clknet_leaf_14_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_15_clk_i (.X(clknet_leaf_15_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_16_clk_i (.X(clknet_leaf_16_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_17_clk_i (.X(clknet_leaf_17_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_18_clk_i (.X(clknet_leaf_18_clk_i),
    .A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_19_clk_i (.X(clknet_leaf_19_clk_i),
    .A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_20_clk_i (.X(clknet_leaf_20_clk_i),
    .A(clknet_6_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_21_clk_i (.X(clknet_leaf_21_clk_i),
    .A(clknet_6_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_22_clk_i (.X(clknet_leaf_22_clk_i),
    .A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_23_clk_i (.X(clknet_leaf_23_clk_i),
    .A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_24_clk_i (.X(clknet_leaf_24_clk_i),
    .A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_25_clk_i (.X(clknet_leaf_25_clk_i),
    .A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_26_clk_i (.X(clknet_leaf_26_clk_i),
    .A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_27_clk_i (.X(clknet_leaf_27_clk_i),
    .A(clknet_6_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_28_clk_i (.X(clknet_leaf_28_clk_i),
    .A(clknet_6_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_29_clk_i (.X(clknet_leaf_29_clk_i),
    .A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_30_clk_i (.X(clknet_leaf_30_clk_i),
    .A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_31_clk_i (.X(clknet_leaf_31_clk_i),
    .A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_32_clk_i (.X(clknet_leaf_32_clk_i),
    .A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_33_clk_i (.X(clknet_leaf_33_clk_i),
    .A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_34_clk_i (.X(clknet_leaf_34_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_35_clk_i (.X(clknet_leaf_35_clk_i),
    .A(clknet_6_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_36_clk_i (.X(clknet_leaf_36_clk_i),
    .A(clknet_6_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_37_clk_i (.X(clknet_leaf_37_clk_i),
    .A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_38_clk_i (.X(clknet_leaf_38_clk_i),
    .A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_39_clk_i (.X(clknet_leaf_39_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_40_clk_i (.X(clknet_leaf_40_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_41_clk_i (.X(clknet_leaf_41_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_42_clk_i (.X(clknet_leaf_42_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_43_clk_i (.X(clknet_leaf_43_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_44_clk_i (.X(clknet_leaf_44_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_45_clk_i (.X(clknet_leaf_45_clk_i),
    .A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_46_clk_i (.X(clknet_leaf_46_clk_i),
    .A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_47_clk_i (.X(clknet_leaf_47_clk_i),
    .A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_48_clk_i (.X(clknet_leaf_48_clk_i),
    .A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_49_clk_i (.X(clknet_leaf_49_clk_i),
    .A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_50_clk_i (.X(clknet_leaf_50_clk_i),
    .A(clknet_6_36_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_51_clk_i (.X(clknet_leaf_51_clk_i),
    .A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_52_clk_i (.X(clknet_leaf_52_clk_i),
    .A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_53_clk_i (.X(clknet_leaf_53_clk_i),
    .A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_54_clk_i (.X(clknet_leaf_54_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_55_clk_i (.X(clknet_leaf_55_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_56_clk_i (.X(clknet_leaf_56_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_57_clk_i (.X(clknet_leaf_57_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_58_clk_i (.X(clknet_leaf_58_clk_i),
    .A(clknet_6_49_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_59_clk_i (.X(clknet_leaf_59_clk_i),
    .A(clknet_6_49_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_60_clk_i (.X(clknet_leaf_60_clk_i),
    .A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_61_clk_i (.X(clknet_leaf_61_clk_i),
    .A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_62_clk_i (.X(clknet_leaf_62_clk_i),
    .A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_63_clk_i (.X(clknet_leaf_63_clk_i),
    .A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_64_clk_i (.X(clknet_leaf_64_clk_i),
    .A(clknet_6_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_65_clk_i (.X(clknet_leaf_65_clk_i),
    .A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_66_clk_i (.X(clknet_leaf_66_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_67_clk_i (.X(clknet_leaf_67_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_68_clk_i (.X(clknet_leaf_68_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_69_clk_i (.X(clknet_leaf_69_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_70_clk_i (.X(clknet_leaf_70_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_71_clk_i (.X(clknet_leaf_71_clk_i),
    .A(clknet_6_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_72_clk_i (.X(clknet_leaf_72_clk_i),
    .A(clknet_6_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_73_clk_i (.X(clknet_leaf_73_clk_i),
    .A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_74_clk_i (.X(clknet_leaf_74_clk_i),
    .A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_75_clk_i (.X(clknet_leaf_75_clk_i),
    .A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_76_clk_i (.X(clknet_leaf_76_clk_i),
    .A(clknet_6_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_77_clk_i (.X(clknet_leaf_77_clk_i),
    .A(clknet_6_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_78_clk_i (.X(clknet_leaf_78_clk_i),
    .A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_79_clk_i (.X(clknet_leaf_79_clk_i),
    .A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_80_clk_i (.X(clknet_leaf_80_clk_i),
    .A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_81_clk_i (.X(clknet_leaf_81_clk_i),
    .A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_82_clk_i (.X(clknet_leaf_82_clk_i),
    .A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_83_clk_i (.X(clknet_leaf_83_clk_i),
    .A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_84_clk_i (.X(clknet_leaf_84_clk_i),
    .A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_86_clk_i (.X(clknet_leaf_86_clk_i),
    .A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_87_clk_i (.X(clknet_leaf_87_clk_i),
    .A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_88_clk_i (.X(clknet_leaf_88_clk_i),
    .A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_89_clk_i (.X(clknet_leaf_89_clk_i),
    .A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_91_clk_i (.X(clknet_leaf_91_clk_i),
    .A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_92_clk_i (.X(clknet_leaf_92_clk_i),
    .A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_93_clk_i (.X(clknet_leaf_93_clk_i),
    .A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_94_clk_i (.X(clknet_leaf_94_clk_i),
    .A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_95_clk_i (.X(clknet_leaf_95_clk_i),
    .A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_96_clk_i (.X(clknet_leaf_96_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_97_clk_i (.X(clknet_leaf_97_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_98_clk_i (.X(clknet_leaf_98_clk_i),
    .A(clknet_6_18_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_99_clk_i (.X(clknet_leaf_99_clk_i),
    .A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_100_clk_i (.X(clknet_leaf_100_clk_i),
    .A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_101_clk_i (.X(clknet_leaf_101_clk_i),
    .A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_102_clk_i (.X(clknet_leaf_102_clk_i),
    .A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_103_clk_i (.X(clknet_leaf_103_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_104_clk_i (.X(clknet_leaf_104_clk_i),
    .A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_105_clk_i (.X(clknet_leaf_105_clk_i),
    .A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_106_clk_i (.X(clknet_leaf_106_clk_i),
    .A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_107_clk_i (.X(clknet_leaf_107_clk_i),
    .A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_108_clk_i (.X(clknet_leaf_108_clk_i),
    .A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_109_clk_i (.X(clknet_leaf_109_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_110_clk_i (.X(clknet_leaf_110_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_111_clk_i (.X(clknet_leaf_111_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_112_clk_i (.X(clknet_leaf_112_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_113_clk_i (.X(clknet_leaf_113_clk_i),
    .A(clknet_6_20_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_114_clk_i (.X(clknet_leaf_114_clk_i),
    .A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_115_clk_i (.X(clknet_leaf_115_clk_i),
    .A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_116_clk_i (.X(clknet_leaf_116_clk_i),
    .A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_117_clk_i (.X(clknet_leaf_117_clk_i),
    .A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_118_clk_i (.X(clknet_leaf_118_clk_i),
    .A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_119_clk_i (.X(clknet_leaf_119_clk_i),
    .A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_120_clk_i (.X(clknet_leaf_120_clk_i),
    .A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_121_clk_i (.X(clknet_leaf_121_clk_i),
    .A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_122_clk_i (.X(clknet_leaf_122_clk_i),
    .A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_123_clk_i (.X(clknet_leaf_123_clk_i),
    .A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_124_clk_i (.X(clknet_leaf_124_clk_i),
    .A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_125_clk_i (.X(clknet_leaf_125_clk_i),
    .A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_126_clk_i (.X(clknet_leaf_126_clk_i),
    .A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_127_clk_i (.X(clknet_leaf_127_clk_i),
    .A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_128_clk_i (.X(clknet_leaf_128_clk_i),
    .A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_129_clk_i (.X(clknet_leaf_129_clk_i),
    .A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_130_clk_i (.X(clknet_leaf_130_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_131_clk_i (.X(clknet_leaf_131_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_132_clk_i (.X(clknet_leaf_132_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_133_clk_i (.X(clknet_leaf_133_clk_i),
    .A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_134_clk_i (.X(clknet_leaf_134_clk_i),
    .A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_135_clk_i (.X(clknet_leaf_135_clk_i),
    .A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_136_clk_i (.X(clknet_leaf_136_clk_i),
    .A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_137_clk_i (.X(clknet_leaf_137_clk_i),
    .A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_138_clk_i (.X(clknet_leaf_138_clk_i),
    .A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_139_clk_i (.X(clknet_leaf_139_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_140_clk_i (.X(clknet_leaf_140_clk_i),
    .A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_141_clk_i (.X(clknet_leaf_141_clk_i),
    .A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_142_clk_i (.X(clknet_leaf_142_clk_i),
    .A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_143_clk_i (.X(clknet_leaf_143_clk_i),
    .A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_144_clk_i (.X(clknet_leaf_144_clk_i),
    .A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_145_clk_i (.X(clknet_leaf_145_clk_i),
    .A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_146_clk_i (.X(clknet_leaf_146_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_147_clk_i (.X(clknet_leaf_147_clk_i),
    .A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_148_clk_i (.X(clknet_leaf_148_clk_i),
    .A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_149_clk_i (.X(clknet_leaf_149_clk_i),
    .A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_151_clk_i (.X(clknet_leaf_151_clk_i),
    .A(clknet_6_27_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_152_clk_i (.X(clknet_leaf_152_clk_i),
    .A(clknet_6_27_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_153_clk_i (.X(clknet_leaf_153_clk_i),
    .A(clknet_6_27_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_154_clk_i (.X(clknet_leaf_154_clk_i),
    .A(clknet_6_27_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_155_clk_i (.X(clknet_leaf_155_clk_i),
    .A(clknet_6_28_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_156_clk_i (.X(clknet_leaf_156_clk_i),
    .A(clknet_6_25_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_157_clk_i (.X(clknet_leaf_157_clk_i),
    .A(clknet_6_25_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_158_clk_i (.X(clknet_leaf_158_clk_i),
    .A(clknet_6_25_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_159_clk_i (.X(clknet_leaf_159_clk_i),
    .A(clknet_6_25_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_160_clk_i (.X(clknet_leaf_160_clk_i),
    .A(clknet_6_25_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_161_clk_i (.X(clknet_leaf_161_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_162_clk_i (.X(clknet_leaf_162_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_163_clk_i (.X(clknet_leaf_163_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_164_clk_i (.X(clknet_leaf_164_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_165_clk_i (.X(clknet_leaf_165_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_166_clk_i (.X(clknet_leaf_166_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_167_clk_i (.X(clknet_leaf_167_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_168_clk_i (.X(clknet_leaf_168_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_169_clk_i (.X(clknet_leaf_169_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_170_clk_i (.X(clknet_leaf_170_clk_i),
    .A(clknet_6_26_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_171_clk_i (.X(clknet_leaf_171_clk_i),
    .A(clknet_6_24_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_172_clk_i (.X(clknet_leaf_172_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_173_clk_i (.X(clknet_leaf_173_clk_i),
    .A(clknet_6_49_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_174_clk_i (.X(clknet_leaf_174_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_175_clk_i (.X(clknet_leaf_175_clk_i),
    .A(clknet_6_49_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_176_clk_i (.X(clknet_leaf_176_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_177_clk_i (.X(clknet_leaf_177_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_178_clk_i (.X(clknet_leaf_178_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_179_clk_i (.X(clknet_leaf_179_clk_i),
    .A(clknet_6_52_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_180_clk_i (.X(clknet_leaf_180_clk_i),
    .A(clknet_6_53_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_181_clk_i (.X(clknet_leaf_181_clk_i),
    .A(clknet_6_53_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_183_clk_i (.X(clknet_leaf_183_clk_i),
    .A(clknet_6_55_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_184_clk_i (.X(clknet_leaf_184_clk_i),
    .A(clknet_6_55_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_185_clk_i (.X(clknet_leaf_185_clk_i),
    .A(clknet_6_55_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_186_clk_i (.X(clknet_leaf_186_clk_i),
    .A(clknet_6_53_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_187_clk_i (.X(clknet_leaf_187_clk_i),
    .A(clknet_6_53_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_188_clk_i (.X(clknet_leaf_188_clk_i),
    .A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_189_clk_i (.X(clknet_leaf_189_clk_i),
    .A(clknet_6_55_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_190_clk_i (.X(clknet_leaf_190_clk_i),
    .A(clknet_6_63_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_191_clk_i (.X(clknet_leaf_191_clk_i),
    .A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_192_clk_i (.X(clknet_leaf_192_clk_i),
    .A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_193_clk_i (.X(clknet_leaf_193_clk_i),
    .A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_194_clk_i (.X(clknet_leaf_194_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_195_clk_i (.X(clknet_leaf_195_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_196_clk_i (.X(clknet_leaf_196_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_197_clk_i (.X(clknet_leaf_197_clk_i),
    .A(clknet_6_63_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_198_clk_i (.X(clknet_leaf_198_clk_i),
    .A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_199_clk_i (.X(clknet_leaf_199_clk_i),
    .A(clknet_6_63_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_200_clk_i (.X(clknet_leaf_200_clk_i),
    .A(clknet_6_63_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_201_clk_i (.X(clknet_leaf_201_clk_i),
    .A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_202_clk_i (.X(clknet_leaf_202_clk_i),
    .A(clknet_6_63_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_203_clk_i (.X(clknet_leaf_203_clk_i),
    .A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_204_clk_i (.X(clknet_leaf_204_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_205_clk_i (.X(clknet_leaf_205_clk_i),
    .A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_206_clk_i (.X(clknet_leaf_206_clk_i),
    .A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_207_clk_i (.X(clknet_leaf_207_clk_i),
    .A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_208_clk_i (.X(clknet_leaf_208_clk_i),
    .A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_209_clk_i (.X(clknet_leaf_209_clk_i),
    .A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_210_clk_i (.X(clknet_leaf_210_clk_i),
    .A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_211_clk_i (.X(clknet_leaf_211_clk_i),
    .A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_212_clk_i (.X(clknet_leaf_212_clk_i),
    .A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_213_clk_i (.X(clknet_leaf_213_clk_i),
    .A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_214_clk_i (.X(clknet_leaf_214_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_215_clk_i (.X(clknet_leaf_215_clk_i),
    .A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_216_clk_i (.X(clknet_leaf_216_clk_i),
    .A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_217_clk_i (.X(clknet_leaf_217_clk_i),
    .A(clknet_6_60_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_218_clk_i (.X(clknet_leaf_218_clk_i),
    .A(clknet_6_55_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_219_clk_i (.X(clknet_leaf_219_clk_i),
    .A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_220_clk_i (.X(clknet_leaf_220_clk_i),
    .A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_221_clk_i (.X(clknet_leaf_221_clk_i),
    .A(clknet_6_49_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_222_clk_i (.X(clknet_leaf_222_clk_i),
    .A(clknet_6_51_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_223_clk_i (.X(clknet_leaf_223_clk_i),
    .A(clknet_6_51_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_224_clk_i (.X(clknet_leaf_224_clk_i),
    .A(clknet_6_51_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_225_clk_i (.X(clknet_leaf_225_clk_i),
    .A(clknet_6_51_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_226_clk_i (.X(clknet_leaf_226_clk_i),
    .A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_228_clk_i (.X(clknet_leaf_228_clk_i),
    .A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_230_clk_i (.X(clknet_leaf_230_clk_i),
    .A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_231_clk_i (.X(clknet_leaf_231_clk_i),
    .A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_232_clk_i (.X(clknet_leaf_232_clk_i),
    .A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_233_clk_i (.X(clknet_leaf_233_clk_i),
    .A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_234_clk_i (.X(clknet_leaf_234_clk_i),
    .A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_235_clk_i (.X(clknet_leaf_235_clk_i),
    .A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_236_clk_i (.X(clknet_leaf_236_clk_i),
    .A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_237_clk_i (.X(clknet_leaf_237_clk_i),
    .A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_238_clk_i (.X(clknet_leaf_238_clk_i),
    .A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_239_clk_i (.X(clknet_leaf_239_clk_i),
    .A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_240_clk_i (.X(clknet_leaf_240_clk_i),
    .A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_241_clk_i (.X(clknet_leaf_241_clk_i),
    .A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_242_clk_i (.X(clknet_leaf_242_clk_i),
    .A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_243_clk_i (.X(clknet_leaf_243_clk_i),
    .A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_244_clk_i (.X(clknet_leaf_244_clk_i),
    .A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_245_clk_i (.X(clknet_leaf_245_clk_i),
    .A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_246_clk_i (.X(clknet_leaf_246_clk_i),
    .A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_247_clk_i (.X(clknet_leaf_247_clk_i),
    .A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_248_clk_i (.X(clknet_leaf_248_clk_i),
    .A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_249_clk_i (.X(clknet_leaf_249_clk_i),
    .A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_250_clk_i (.X(clknet_leaf_250_clk_i),
    .A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_251_clk_i (.X(clknet_leaf_251_clk_i),
    .A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_252_clk_i (.X(clknet_leaf_252_clk_i),
    .A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_253_clk_i (.X(clknet_leaf_253_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_254_clk_i (.X(clknet_leaf_254_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_255_clk_i (.X(clknet_leaf_255_clk_i),
    .A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_256_clk_i (.X(clknet_leaf_256_clk_i),
    .A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_257_clk_i (.X(clknet_leaf_257_clk_i),
    .A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_258_clk_i (.X(clknet_leaf_258_clk_i),
    .A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_259_clk_i (.X(clknet_leaf_259_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_260_clk_i (.X(clknet_leaf_260_clk_i),
    .A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_261_clk_i (.X(clknet_leaf_261_clk_i),
    .A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_262_clk_i (.X(clknet_leaf_262_clk_i),
    .A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_263_clk_i (.X(clknet_leaf_263_clk_i),
    .A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_264_clk_i (.X(clknet_leaf_264_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_265_clk_i (.X(clknet_leaf_265_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_266_clk_i (.X(clknet_leaf_266_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_267_clk_i (.X(clknet_leaf_267_clk_i),
    .A(clknet_6_42_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_268_clk_i (.X(clknet_leaf_268_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_269_clk_i (.X(clknet_leaf_269_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_270_clk_i (.X(clknet_leaf_270_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_271_clk_i (.X(clknet_leaf_271_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_272_clk_i (.X(clknet_leaf_272_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_273_clk_i (.X(clknet_leaf_273_clk_i),
    .A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_274_clk_i (.X(clknet_leaf_274_clk_i),
    .A(clknet_6_40_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_275_clk_i (.X(clknet_leaf_275_clk_i),
    .A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_276_clk_i (.X(clknet_leaf_276_clk_i),
    .A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_277_clk_i (.X(clknet_leaf_277_clk_i),
    .A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_278_clk_i (.X(clknet_leaf_278_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_279_clk_i (.X(clknet_leaf_279_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_280_clk_i (.X(clknet_leaf_280_clk_i),
    .A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_281_clk_i (.X(clknet_leaf_281_clk_i),
    .A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_282_clk_i (.X(clknet_leaf_282_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_283_clk_i (.X(clknet_leaf_283_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_284_clk_i (.X(clknet_leaf_284_clk_i),
    .A(clknet_6_44_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_285_clk_i (.X(clknet_leaf_285_clk_i),
    .A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_286_clk_i (.X(clknet_leaf_286_clk_i),
    .A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_287_clk_i (.X(clknet_leaf_287_clk_i),
    .A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_288_clk_i (.X(clknet_leaf_288_clk_i),
    .A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_289_clk_i (.X(clknet_leaf_289_clk_i),
    .A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_290_clk_i (.X(clknet_leaf_290_clk_i),
    .A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_291_clk_i (.X(clknet_leaf_291_clk_i),
    .A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_292_clk_i (.X(clknet_leaf_292_clk_i),
    .A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_293_clk_i (.X(clknet_leaf_293_clk_i),
    .A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_294_clk_i (.X(clknet_leaf_294_clk_i),
    .A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_295_clk_i (.X(clknet_leaf_295_clk_i),
    .A(clknet_6_51_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_296_clk_i (.X(clknet_leaf_296_clk_i),
    .A(clknet_6_48_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_297_clk_i (.X(clknet_leaf_297_clk_i),
    .A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_298_clk_i (.X(clknet_leaf_298_clk_i),
    .A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_299_clk_i (.X(clknet_leaf_299_clk_i),
    .A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_300_clk_i (.X(clknet_leaf_300_clk_i),
    .A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_301_clk_i (.X(clknet_leaf_301_clk_i),
    .A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_302_clk_i (.X(clknet_leaf_302_clk_i),
    .A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_303_clk_i (.X(clknet_leaf_303_clk_i),
    .A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_304_clk_i (.X(clknet_leaf_304_clk_i),
    .A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_305_clk_i (.X(clknet_leaf_305_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_306_clk_i (.X(clknet_leaf_306_clk_i),
    .A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_307_clk_i (.X(clknet_leaf_307_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_308_clk_i (.X(clknet_leaf_308_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_309_clk_i (.X(clknet_leaf_309_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_310_clk_i (.X(clknet_leaf_310_clk_i),
    .A(clknet_6_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_311_clk_i (.X(clknet_leaf_311_clk_i),
    .A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_312_clk_i (.X(clknet_leaf_312_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_313_clk_i (.X(clknet_leaf_313_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_314_clk_i (.X(clknet_leaf_314_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_315_clk_i (.X(clknet_leaf_315_clk_i),
    .A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_316_clk_i (.X(clknet_leaf_316_clk_i),
    .A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_317_clk_i (.X(clknet_leaf_317_clk_i),
    .A(clknet_6_32_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_318_clk_i (.X(clknet_leaf_318_clk_i),
    .A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_319_clk_i (.X(clknet_leaf_319_clk_i),
    .A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_320_clk_i (.X(clknet_leaf_320_clk_i),
    .A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_321_clk_i (.X(clknet_leaf_321_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_322_clk_i (.X(clknet_leaf_322_clk_i),
    .A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_323_clk_i (.X(clknet_leaf_323_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_324_clk_i (.X(clknet_leaf_324_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_325_clk_i (.X(clknet_leaf_325_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_326_clk_i (.X(clknet_leaf_326_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_327_clk_i (.X(clknet_leaf_327_clk_i),
    .A(clknet_6_34_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_328_clk_i (.X(clknet_leaf_328_clk_i),
    .A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_329_clk_i (.X(clknet_leaf_329_clk_i),
    .A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_330_clk_i (.X(clknet_leaf_330_clk_i),
    .A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_331_clk_i (.X(clknet_leaf_331_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_332_clk_i (.X(clknet_leaf_332_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_333_clk_i (.X(clknet_leaf_333_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_334_clk_i (.X(clknet_leaf_334_clk_i),
    .A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_335_clk_i (.X(clknet_leaf_335_clk_i),
    .A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_336_clk_i (.X(clknet_leaf_336_clk_i),
    .A(clknet_6_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_337_clk_i (.X(clknet_leaf_337_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_338_clk_i (.X(clknet_leaf_338_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_339_clk_i (.X(clknet_leaf_339_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_340_clk_i (.X(clknet_leaf_340_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_341_clk_i (.X(clknet_leaf_341_clk_i),
    .A(clknet_6_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_342_clk_i (.X(clknet_leaf_342_clk_i),
    .A(clknet_6_0_0_clk_i));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_2_0_0_clk_i (.X(clknet_2_0_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_2_1_0_clk_i (.X(clknet_2_1_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_2_2_0_clk_i (.X(clknet_2_2_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_2_3_0_clk_i (.X(clknet_2_3_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_6_0_0_clk_i (.X(clknet_6_0_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_1_0_clk_i (.X(clknet_6_1_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_2_0_clk_i (.X(clknet_6_2_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_3_0_clk_i (.X(clknet_6_3_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_4_0_clk_i (.X(clknet_6_4_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_5_0_clk_i (.X(clknet_6_5_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_6_0_clk_i (.X(clknet_6_6_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_7_0_clk_i (.X(clknet_6_7_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_8_0_clk_i (.X(clknet_6_8_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_9_0_clk_i (.X(clknet_6_9_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_10_0_clk_i (.X(clknet_6_10_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_11_0_clk_i (.X(clknet_6_11_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_12_0_clk_i (.X(clknet_6_12_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_13_0_clk_i (.X(clknet_6_13_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_14_0_clk_i (.X(clknet_6_14_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_15_0_clk_i (.X(clknet_6_15_0_clk_i),
    .A(clknet_2_0_0_clk_i));
 sg13g2_buf_16 clkbuf_6_16_0_clk_i (.X(clknet_6_16_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_17_0_clk_i (.X(clknet_6_17_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_18_0_clk_i (.X(clknet_6_18_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_19_0_clk_i (.X(clknet_6_19_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_20_0_clk_i (.X(clknet_6_20_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_21_0_clk_i (.X(clknet_6_21_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_22_0_clk_i (.X(clknet_6_22_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_23_0_clk_i (.X(clknet_6_23_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_24_0_clk_i (.X(clknet_6_24_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_25_0_clk_i (.X(clknet_6_25_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_26_0_clk_i (.X(clknet_6_26_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_27_0_clk_i (.X(clknet_6_27_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_28_0_clk_i (.X(clknet_6_28_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_29_0_clk_i (.X(clknet_6_29_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_30_0_clk_i (.X(clknet_6_30_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_31_0_clk_i (.X(clknet_6_31_0_clk_i),
    .A(clknet_2_1_0_clk_i));
 sg13g2_buf_16 clkbuf_6_32_0_clk_i (.X(clknet_6_32_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_33_0_clk_i (.X(clknet_6_33_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_34_0_clk_i (.X(clknet_6_34_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_35_0_clk_i (.X(clknet_6_35_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_36_0_clk_i (.X(clknet_6_36_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_37_0_clk_i (.X(clknet_6_37_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_38_0_clk_i (.X(clknet_6_38_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_39_0_clk_i (.X(clknet_6_39_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_40_0_clk_i (.X(clknet_6_40_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_41_0_clk_i (.X(clknet_6_41_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_42_0_clk_i (.X(clknet_6_42_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_43_0_clk_i (.X(clknet_6_43_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_44_0_clk_i (.X(clknet_6_44_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_45_0_clk_i (.X(clknet_6_45_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_46_0_clk_i (.X(clknet_6_46_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_47_0_clk_i (.X(clknet_6_47_0_clk_i),
    .A(clknet_2_2_0_clk_i));
 sg13g2_buf_16 clkbuf_6_48_0_clk_i (.X(clknet_6_48_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_49_0_clk_i (.X(clknet_6_49_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_50_0_clk_i (.X(clknet_6_50_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_51_0_clk_i (.X(clknet_6_51_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_52_0_clk_i (.X(clknet_6_52_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_53_0_clk_i (.X(clknet_6_53_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_54_0_clk_i (.X(clknet_6_54_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_55_0_clk_i (.X(clknet_6_55_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_56_0_clk_i (.X(clknet_6_56_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_57_0_clk_i (.X(clknet_6_57_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_58_0_clk_i (.X(clknet_6_58_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_59_0_clk_i (.X(clknet_6_59_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_60_0_clk_i (.X(clknet_6_60_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_61_0_clk_i (.X(clknet_6_61_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_62_0_clk_i (.X(clknet_6_62_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkbuf_6_63_0_clk_i (.X(clknet_6_63_0_clk_i),
    .A(clknet_2_3_0_clk_i));
 sg13g2_buf_16 clkload0 (.A(clknet_6_1_0_clk_i));
 sg13g2_buf_16 clkload1 (.A(clknet_6_3_0_clk_i));
 sg13g2_inv_4 clkload2 (.A(clknet_6_4_0_clk_i));
 sg13g2_buf_16 clkload3 (.A(clknet_6_5_0_clk_i));
 sg13g2_buf_16 clkload4 (.A(clknet_6_6_0_clk_i));
 sg13g2_buf_16 clkload5 (.A(clknet_6_7_0_clk_i));
 sg13g2_buf_16 clkload6 (.A(clknet_6_9_0_clk_i));
 sg13g2_buf_16 clkload7 (.A(clknet_6_11_0_clk_i));
 sg13g2_buf_16 clkload8 (.A(clknet_6_13_0_clk_i));
 sg13g2_buf_16 clkload9 (.A(clknet_6_14_0_clk_i));
 sg13g2_buf_16 clkload10 (.A(clknet_6_15_0_clk_i));
 sg13g2_inv_4 clkload11 (.A(clknet_6_16_0_clk_i));
 sg13g2_buf_16 clkload12 (.A(clknet_6_17_0_clk_i));
 sg13g2_buf_16 clkload13 (.A(clknet_6_19_0_clk_i));
 sg13g2_buf_16 clkload14 (.A(clknet_6_21_0_clk_i));
 sg13g2_buf_16 clkload15 (.A(clknet_6_22_0_clk_i));
 sg13g2_buf_16 clkload16 (.A(clknet_6_23_0_clk_i));
 sg13g2_buf_16 clkload17 (.A(clknet_6_25_0_clk_i));
 sg13g2_inv_8 clkload18 (.A(clknet_6_27_0_clk_i));
 sg13g2_buf_16 clkload19 (.A(clknet_6_29_0_clk_i));
 sg13g2_buf_16 clkload20 (.A(clknet_6_30_0_clk_i));
 sg13g2_buf_16 clkload21 (.A(clknet_6_31_0_clk_i));
 sg13g2_buf_16 clkload22 (.A(clknet_6_33_0_clk_i));
 sg13g2_buf_16 clkload23 (.A(clknet_6_35_0_clk_i));
 sg13g2_buf_16 clkload24 (.A(clknet_6_37_0_clk_i));
 sg13g2_buf_16 clkload25 (.A(clknet_6_38_0_clk_i));
 sg13g2_buf_16 clkload26 (.A(clknet_6_39_0_clk_i));
 sg13g2_buf_16 clkload27 (.A(clknet_6_41_0_clk_i));
 sg13g2_buf_16 clkload28 (.A(clknet_6_43_0_clk_i));
 sg13g2_buf_16 clkload29 (.A(clknet_6_45_0_clk_i));
 sg13g2_buf_16 clkload30 (.A(clknet_6_46_0_clk_i));
 sg13g2_buf_16 clkload31 (.A(clknet_6_47_0_clk_i));
 sg13g2_buf_16 clkload32 (.A(clknet_6_49_0_clk_i));
 sg13g2_inv_4 clkload33 (.A(clknet_6_50_0_clk_i));
 sg13g2_buf_16 clkload34 (.A(clknet_6_51_0_clk_i));
 sg13g2_inv_8 clkload35 (.A(clknet_6_53_0_clk_i));
 sg13g2_buf_16 clkload36 (.A(clknet_6_54_0_clk_i));
 sg13g2_buf_16 clkload37 (.A(clknet_6_55_0_clk_i));
 sg13g2_inv_4 clkload38 (.A(clknet_6_56_0_clk_i));
 sg13g2_buf_16 clkload39 (.A(clknet_6_57_0_clk_i));
 sg13g2_buf_16 clkload40 (.A(clknet_6_58_0_clk_i));
 sg13g2_buf_16 clkload41 (.A(clknet_6_59_0_clk_i));
 sg13g2_buf_16 clkload42 (.A(clknet_6_61_0_clk_i));
 sg13g2_buf_16 clkload43 (.A(clknet_6_62_0_clk_i));
 sg13g2_buf_16 clkload44 (.A(clknet_6_63_0_clk_i));
 sg13g2_inv_4 clkload45 (.A(clknet_leaf_0_clk_i));
 sg13g2_inv_4 clkload46 (.A(clknet_leaf_2_clk_i));
 sg13g2_buf_8 clkload47 (.A(clknet_leaf_17_clk_i));
 sg13g2_inv_4 clkload48 (.A(clknet_leaf_342_clk_i));
 sg13g2_inv_2 clkload49 (.A(clknet_leaf_22_clk_i));
 sg13g2_inv_2 clkload50 (.A(clknet_leaf_23_clk_i));
 sg13g2_buf_8 clkload51 (.A(clknet_leaf_24_clk_i));
 sg13g2_inv_2 clkload52 (.A(clknet_leaf_3_clk_i));
 sg13g2_inv_1 clkload53 (.A(clknet_leaf_5_clk_i));
 sg13g2_buf_8 clkload54 (.A(clknet_leaf_14_clk_i));
 sg13g2_inv_1 clkload55 (.A(clknet_leaf_15_clk_i));
 sg13g2_inv_4 clkload56 (.A(clknet_leaf_21_clk_i));
 sg13g2_buf_8 clkload57 (.A(clknet_leaf_35_clk_i));
 sg13g2_inv_1 clkload58 (.A(clknet_leaf_36_clk_i));
 sg13g2_inv_1 clkload59 (.A(clknet_leaf_82_clk_i));
 sg13g2_inv_4 clkload60 (.A(clknet_leaf_83_clk_i));
 sg13g2_inv_1 clkload61 (.A(clknet_leaf_84_clk_i));
 sg13g2_buf_2 clkload62 (.A(clknet_leaf_81_clk_i));
 sg13g2_buf_8 clkload63 (.A(clknet_leaf_87_clk_i));
 sg13g2_inv_2 clkload64 (.A(clknet_leaf_88_clk_i));
 sg13g2_inv_2 clkload65 (.A(clknet_leaf_89_clk_i));
 sg13g2_buf_8 clkload66 (.A(clknet_leaf_30_clk_i));
 sg13g2_inv_2 clkload67 (.A(clknet_leaf_79_clk_i));
 sg13g2_inv_4 clkload68 (.A(clknet_leaf_73_clk_i));
 sg13g2_buf_8 clkload69 (.A(clknet_leaf_74_clk_i));
 sg13g2_inv_2 clkload70 (.A(clknet_leaf_75_clk_i));
 sg13g2_inv_1 clkload71 (.A(clknet_leaf_80_clk_i));
 sg13g2_inv_4 clkload72 (.A(clknet_leaf_6_clk_i));
 sg13g2_inv_4 clkload73 (.A(clknet_leaf_337_clk_i));
 sg13g2_inv_1 clkload74 (.A(clknet_leaf_338_clk_i));
 sg13g2_buf_8 clkload75 (.A(clknet_leaf_339_clk_i));
 sg13g2_inv_4 clkload76 (.A(clknet_leaf_341_clk_i));
 sg13g2_inv_2 clkload77 (.A(clknet_leaf_7_clk_i));
 sg13g2_buf_16 clkload78 (.A(clknet_leaf_8_clk_i));
 sg13g2_inv_4 clkload79 (.A(clknet_leaf_12_clk_i));
 sg13g2_inv_2 clkload80 (.A(clknet_leaf_311_clk_i));
 sg13g2_buf_8 clkload81 (.A(clknet_leaf_312_clk_i));
 sg13g2_buf_2 clkload82 (.A(clknet_leaf_314_clk_i));
 sg13g2_buf_8 clkload83 (.A(clknet_leaf_331_clk_i));
 sg13g2_buf_2 clkload84 (.A(clknet_leaf_333_clk_i));
 sg13g2_inv_2 clkload85 (.A(clknet_leaf_336_clk_i));
 sg13g2_inv_2 clkload86 (.A(clknet_leaf_328_clk_i));
 sg13g2_inv_2 clkload87 (.A(clknet_leaf_329_clk_i));
 sg13g2_inv_4 clkload88 (.A(clknet_leaf_334_clk_i));
 sg13g2_inv_4 clkload89 (.A(clknet_leaf_335_clk_i));
 sg13g2_inv_4 clkload90 (.A(clknet_leaf_10_clk_i));
 sg13g2_inv_1 clkload91 (.A(clknet_leaf_13_clk_i));
 sg13g2_buf_8 clkload92 (.A(clknet_leaf_39_clk_i));
 sg13g2_inv_2 clkload93 (.A(clknet_leaf_40_clk_i));
 sg13g2_inv_2 clkload94 (.A(clknet_leaf_32_clk_i));
 sg13g2_inv_2 clkload95 (.A(clknet_leaf_33_clk_i));
 sg13g2_buf_8 clkload96 (.A(clknet_leaf_38_clk_i));
 sg13g2_inv_4 clkload97 (.A(clknet_leaf_48_clk_i));
 sg13g2_inv_4 clkload98 (.A(clknet_leaf_61_clk_i));
 sg13g2_inv_4 clkload99 (.A(clknet_leaf_63_clk_i));
 sg13g2_inv_4 clkload100 (.A(clknet_leaf_65_clk_i));
 sg13g2_buf_8 clkload101 (.A(clknet_leaf_71_clk_i));
 sg13g2_inv_4 clkload102 (.A(clknet_leaf_72_clk_i));
 sg13g2_inv_1 clkload103 (.A(clknet_leaf_76_clk_i));
 sg13g2_inv_1 clkload104 (.A(clknet_leaf_77_clk_i));
 sg13g2_inv_4 clkload105 (.A(clknet_leaf_91_clk_i));
 sg13g2_buf_2 clkload106 (.A(clknet_leaf_93_clk_i));
 sg13g2_buf_2 clkload107 (.A(clknet_leaf_94_clk_i));
 sg13g2_buf_4 clkload108 (.A(clknet_leaf_106_clk_i));
 sg13g2_inv_1 clkload109 (.A(clknet_leaf_101_clk_i));
 sg13g2_buf_8 clkload110 (.A(clknet_leaf_104_clk_i));
 sg13g2_buf_8 clkload111 (.A(clknet_leaf_105_clk_i));
 sg13g2_inv_1 clkload112 (.A(clknet_leaf_108_clk_i));
 sg13g2_buf_8 clkload113 (.A(clknet_leaf_68_clk_i));
 sg13g2_inv_2 clkload114 (.A(clknet_leaf_70_clk_i));
 sg13g2_inv_2 clkload115 (.A(clknet_leaf_97_clk_i));
 sg13g2_buf_8 clkload116 (.A(clknet_leaf_100_clk_i));
 sg13g2_inv_1 clkload117 (.A(clknet_leaf_109_clk_i));
 sg13g2_inv_4 clkload118 (.A(clknet_leaf_110_clk_i));
 sg13g2_inv_4 clkload119 (.A(clknet_leaf_111_clk_i));
 sg13g2_inv_1 clkload120 (.A(clknet_leaf_112_clk_i));
 sg13g2_inv_4 clkload121 (.A(clknet_leaf_113_clk_i));
 sg13g2_inv_4 clkload122 (.A(clknet_leaf_114_clk_i));
 sg13g2_inv_4 clkload123 (.A(clknet_leaf_116_clk_i));
 sg13g2_inv_2 clkload124 (.A(clknet_leaf_117_clk_i));
 sg13g2_inv_1 clkload125 (.A(clknet_leaf_118_clk_i));
 sg13g2_buf_8 clkload126 (.A(clknet_leaf_124_clk_i));
 sg13g2_inv_2 clkload127 (.A(clknet_leaf_126_clk_i));
 sg13g2_inv_1 clkload128 (.A(clknet_leaf_120_clk_i));
 sg13g2_inv_1 clkload129 (.A(clknet_leaf_121_clk_i));
 sg13g2_inv_4 clkload130 (.A(clknet_leaf_122_clk_i));
 sg13g2_buf_8 clkload131 (.A(clknet_leaf_134_clk_i));
 sg13g2_inv_1 clkload132 (.A(clknet_leaf_66_clk_i));
 sg13g2_buf_8 clkload133 (.A(clknet_leaf_67_clk_i));
 sg13g2_inv_1 clkload134 (.A(clknet_leaf_162_clk_i));
 sg13g2_inv_4 clkload135 (.A(clknet_leaf_171_clk_i));
 sg13g2_inv_2 clkload136 (.A(clknet_leaf_157_clk_i));
 sg13g2_inv_1 clkload137 (.A(clknet_leaf_158_clk_i));
 sg13g2_inv_2 clkload138 (.A(clknet_leaf_159_clk_i));
 sg13g2_inv_2 clkload139 (.A(clknet_leaf_160_clk_i));
 sg13g2_buf_16 clkload140 (.A(clknet_leaf_164_clk_i));
 sg13g2_buf_2 clkload141 (.A(clknet_leaf_165_clk_i));
 sg13g2_inv_2 clkload142 (.A(clknet_leaf_166_clk_i));
 sg13g2_buf_4 clkload143 (.A(clknet_leaf_168_clk_i));
 sg13g2_buf_8 clkload144 (.A(clknet_leaf_170_clk_i));
 sg13g2_inv_4 clkload145 (.A(clknet_leaf_151_clk_i));
 sg13g2_inv_4 clkload146 (.A(clknet_leaf_153_clk_i));
 sg13g2_inv_1 clkload147 (.A(clknet_leaf_131_clk_i));
 sg13g2_inv_1 clkload148 (.A(clknet_leaf_155_clk_i));
 sg13g2_inv_1 clkload149 (.A(clknet_leaf_133_clk_i));
 sg13g2_inv_4 clkload150 (.A(clknet_leaf_135_clk_i));
 sg13g2_inv_4 clkload151 (.A(clknet_leaf_136_clk_i));
 sg13g2_buf_8 clkload152 (.A(clknet_leaf_137_clk_i));
 sg13g2_buf_8 clkload153 (.A(clknet_leaf_144_clk_i));
 sg13g2_inv_1 clkload154 (.A(clknet_leaf_145_clk_i));
 sg13g2_inv_2 clkload155 (.A(clknet_leaf_147_clk_i));
 sg13g2_inv_4 clkload156 (.A(clknet_leaf_149_clk_i));
 sg13g2_inv_2 clkload157 (.A(clknet_leaf_140_clk_i));
 sg13g2_inv_2 clkload158 (.A(clknet_leaf_141_clk_i));
 sg13g2_inv_1 clkload159 (.A(clknet_leaf_143_clk_i));
 sg13g2_inv_2 clkload160 (.A(clknet_leaf_188_clk_i));
 sg13g2_inv_4 clkload161 (.A(clknet_leaf_305_clk_i));
 sg13g2_inv_1 clkload162 (.A(clknet_leaf_308_clk_i));
 sg13g2_inv_4 clkload163 (.A(clknet_leaf_309_clk_i));
 sg13g2_inv_1 clkload164 (.A(clknet_leaf_313_clk_i));
 sg13g2_buf_16 clkload165 (.A(clknet_leaf_317_clk_i));
 sg13g2_buf_16 clkload166 (.A(clknet_leaf_302_clk_i));
 sg13g2_inv_2 clkload167 (.A(clknet_leaf_303_clk_i));
 sg13g2_buf_8 clkload168 (.A(clknet_leaf_304_clk_i));
 sg13g2_inv_2 clkload169 (.A(clknet_leaf_306_clk_i));
 sg13g2_inv_1 clkload170 (.A(clknet_leaf_321_clk_i));
 sg13g2_inv_4 clkload171 (.A(clknet_leaf_324_clk_i));
 sg13g2_inv_4 clkload172 (.A(clknet_leaf_326_clk_i));
 sg13g2_inv_1 clkload173 (.A(clknet_leaf_327_clk_i));
 sg13g2_inv_4 clkload174 (.A(clknet_leaf_315_clk_i));
 sg13g2_inv_2 clkload175 (.A(clknet_leaf_316_clk_i));
 sg13g2_inv_1 clkload176 (.A(clknet_leaf_320_clk_i));
 sg13g2_buf_8 clkload177 (.A(clknet_leaf_322_clk_i));
 sg13g2_buf_8 clkload178 (.A(clknet_leaf_34_clk_i));
 sg13g2_inv_4 clkload179 (.A(clknet_leaf_41_clk_i));
 sg13g2_buf_8 clkload180 (.A(clknet_leaf_42_clk_i));
 sg13g2_inv_1 clkload181 (.A(clknet_leaf_44_clk_i));
 sg13g2_inv_2 clkload182 (.A(clknet_leaf_50_clk_i));
 sg13g2_inv_2 clkload183 (.A(clknet_leaf_45_clk_i));
 sg13g2_buf_8 clkload184 (.A(clknet_leaf_46_clk_i));
 sg13g2_buf_8 clkload185 (.A(clknet_leaf_49_clk_i));
 sg13g2_inv_2 clkload186 (.A(clknet_leaf_51_clk_i));
 sg13g2_inv_2 clkload187 (.A(clknet_leaf_289_clk_i));
 sg13g2_inv_2 clkload188 (.A(clknet_leaf_290_clk_i));
 sg13g2_buf_8 clkload189 (.A(clknet_leaf_293_clk_i));
 sg13g2_buf_2 clkload190 (.A(clknet_leaf_294_clk_i));
 sg13g2_inv_2 clkload191 (.A(clknet_leaf_52_clk_i));
 sg13g2_inv_4 clkload192 (.A(clknet_leaf_53_clk_i));
 sg13g2_buf_2 clkload193 (.A(clknet_leaf_297_clk_i));
 sg13g2_buf_4 clkload194 (.A(clknet_leaf_298_clk_i));
 sg13g2_buf_2 clkload195 (.A(clknet_leaf_268_clk_i));
 sg13g2_buf_2 clkload196 (.A(clknet_leaf_270_clk_i));
 sg13g2_inv_1 clkload197 (.A(clknet_leaf_271_clk_i));
 sg13g2_buf_2 clkload198 (.A(clknet_leaf_272_clk_i));
 sg13g2_buf_2 clkload199 (.A(clknet_leaf_274_clk_i));
 sg13g2_buf_2 clkload200 (.A(clknet_leaf_273_clk_i));
 sg13g2_inv_4 clkload201 (.A(clknet_leaf_277_clk_i));
 sg13g2_inv_4 clkload202 (.A(clknet_leaf_280_clk_i));
 sg13g2_inv_2 clkload203 (.A(clknet_leaf_253_clk_i));
 sg13g2_buf_8 clkload204 (.A(clknet_leaf_254_clk_i));
 sg13g2_buf_8 clkload205 (.A(clknet_leaf_264_clk_i));
 sg13g2_inv_2 clkload206 (.A(clknet_leaf_265_clk_i));
 sg13g2_buf_8 clkload207 (.A(clknet_leaf_266_clk_i));
 sg13g2_buf_8 clkload208 (.A(clknet_leaf_260_clk_i));
 sg13g2_buf_2 clkload209 (.A(clknet_leaf_261_clk_i));
 sg13g2_buf_4 clkload210 (.A(clknet_leaf_262_clk_i));
 sg13g2_buf_2 clkload211 (.A(clknet_leaf_281_clk_i));
 sg13g2_buf_2 clkload212 (.A(clknet_leaf_259_clk_i));
 sg13g2_buf_16 clkload213 (.A(clknet_leaf_278_clk_i));
 sg13g2_inv_1 clkload214 (.A(clknet_leaf_279_clk_i));
 sg13g2_inv_4 clkload215 (.A(clknet_leaf_282_clk_i));
 sg13g2_buf_8 clkload216 (.A(clknet_leaf_284_clk_i));
 sg13g2_buf_8 clkload217 (.A(clknet_leaf_286_clk_i));
 sg13g2_inv_2 clkload218 (.A(clknet_leaf_288_clk_i));
 sg13g2_inv_2 clkload219 (.A(clknet_leaf_291_clk_i));
 sg13g2_buf_8 clkload220 (.A(clknet_leaf_319_clk_i));
 sg13g2_inv_2 clkload221 (.A(clknet_leaf_249_clk_i));
 sg13g2_inv_4 clkload222 (.A(clknet_leaf_250_clk_i));
 sg13g2_buf_2 clkload223 (.A(clknet_leaf_256_clk_i));
 sg13g2_buf_2 clkload224 (.A(clknet_leaf_257_clk_i));
 sg13g2_buf_8 clkload225 (.A(clknet_leaf_242_clk_i));
 sg13g2_inv_1 clkload226 (.A(clknet_leaf_243_clk_i));
 sg13g2_buf_8 clkload227 (.A(clknet_leaf_251_clk_i));
 sg13g2_inv_4 clkload228 (.A(clknet_leaf_252_clk_i));
 sg13g2_buf_8 clkload229 (.A(clknet_leaf_54_clk_i));
 sg13g2_inv_2 clkload230 (.A(clknet_leaf_55_clk_i));
 sg13g2_inv_2 clkload231 (.A(clknet_leaf_57_clk_i));
 sg13g2_buf_2 clkload232 (.A(clknet_leaf_174_clk_i));
 sg13g2_buf_2 clkload233 (.A(clknet_leaf_296_clk_i));
 sg13g2_inv_1 clkload234 (.A(clknet_leaf_58_clk_i));
 sg13g2_inv_4 clkload235 (.A(clknet_leaf_59_clk_i));
 sg13g2_buf_8 clkload236 (.A(clknet_leaf_175_clk_i));
 sg13g2_buf_8 clkload237 (.A(clknet_leaf_221_clk_i));
 sg13g2_buf_2 clkload238 (.A(clknet_leaf_226_clk_i));
 sg13g2_inv_2 clkload239 (.A(clknet_leaf_228_clk_i));
 sg13g2_inv_2 clkload240 (.A(clknet_leaf_285_clk_i));
 sg13g2_inv_2 clkload241 (.A(clknet_leaf_292_clk_i));
 sg13g2_inv_1 clkload242 (.A(clknet_leaf_222_clk_i));
 sg13g2_inv_4 clkload243 (.A(clknet_leaf_223_clk_i));
 sg13g2_inv_4 clkload244 (.A(clknet_leaf_225_clk_i));
 sg13g2_buf_2 clkload245 (.A(clknet_leaf_295_clk_i));
 sg13g2_buf_4 clkload246 (.A(clknet_leaf_172_clk_i));
 sg13g2_inv_4 clkload247 (.A(clknet_leaf_176_clk_i));
 sg13g2_buf_8 clkload248 (.A(clknet_leaf_177_clk_i));
 sg13g2_buf_8 clkload249 (.A(clknet_leaf_178_clk_i));
 sg13g2_inv_1 clkload250 (.A(clknet_leaf_179_clk_i));
 sg13g2_buf_4 clkload251 (.A(clknet_leaf_181_clk_i));
 sg13g2_inv_2 clkload252 (.A(clknet_leaf_186_clk_i));
 sg13g2_buf_8 clkload253 (.A(clknet_leaf_187_clk_i));
 sg13g2_buf_8 clkload254 (.A(clknet_leaf_213_clk_i));
 sg13g2_inv_2 clkload255 (.A(clknet_leaf_215_clk_i));
 sg13g2_buf_8 clkload256 (.A(clknet_leaf_216_clk_i));
 sg13g2_inv_4 clkload257 (.A(clknet_leaf_220_clk_i));
 sg13g2_inv_2 clkload258 (.A(clknet_leaf_183_clk_i));
 sg13g2_buf_2 clkload259 (.A(clknet_leaf_184_clk_i));
 sg13g2_inv_4 clkload260 (.A(clknet_leaf_185_clk_i));
 sg13g2_inv_2 clkload261 (.A(clknet_leaf_218_clk_i));
 sg13g2_buf_4 clkload262 (.A(clknet_leaf_230_clk_i));
 sg13g2_buf_4 clkload263 (.A(clknet_leaf_236_clk_i));
 sg13g2_inv_4 clkload264 (.A(clknet_leaf_246_clk_i));
 sg13g2_inv_4 clkload265 (.A(clknet_leaf_247_clk_i));
 sg13g2_buf_8 clkload266 (.A(clknet_leaf_235_clk_i));
 sg13g2_inv_2 clkload267 (.A(clknet_leaf_239_clk_i));
 sg13g2_inv_1 clkload268 (.A(clknet_leaf_244_clk_i));
 sg13g2_inv_2 clkload269 (.A(clknet_leaf_245_clk_i));
 sg13g2_buf_8 clkload270 (.A(clknet_leaf_231_clk_i));
 sg13g2_buf_2 clkload271 (.A(clknet_leaf_233_clk_i));
 sg13g2_inv_2 clkload272 (.A(clknet_leaf_237_clk_i));
 sg13g2_inv_4 clkload273 (.A(clknet_leaf_238_clk_i));
 sg13g2_inv_1 clkload274 (.A(clknet_leaf_208_clk_i));
 sg13g2_inv_2 clkload275 (.A(clknet_leaf_210_clk_i));
 sg13g2_buf_8 clkload276 (.A(clknet_leaf_211_clk_i));
 sg13g2_buf_4 clkload277 (.A(clknet_leaf_232_clk_i));
 sg13g2_inv_4 clkload278 (.A(clknet_leaf_195_clk_i));
 sg13g2_inv_4 clkload279 (.A(clknet_leaf_196_clk_i));
 sg13g2_buf_16 clkload280 (.A(clknet_leaf_204_clk_i));
 sg13g2_buf_4 clkload281 (.A(clknet_leaf_214_clk_i));
 sg13g2_inv_2 clkload282 (.A(clknet_leaf_217_clk_i));
 sg13g2_inv_4 clkload283 (.A(clknet_leaf_192_clk_i));
 sg13g2_buf_2 clkload284 (.A(clknet_leaf_193_clk_i));
 sg13g2_inv_2 clkload285 (.A(clknet_leaf_198_clk_i));
 sg13g2_buf_8 clkload286 (.A(clknet_leaf_201_clk_i));
 sg13g2_inv_1 clkload287 (.A(clknet_leaf_203_clk_i));
 sg13g2_buf_16 clkload288 (.A(clknet_leaf_205_clk_i));
 sg13g2_buf_8 clkload289 (.A(clknet_leaf_207_clk_i));
 sg13g2_buf_2 clkload290 (.A(clknet_leaf_212_clk_i));
 sg13g2_inv_4 clkload291 (.A(clknet_leaf_197_clk_i));
 sg13g2_buf_8 clkload292 (.A(clknet_leaf_199_clk_i));
 sg13g2_buf_8 clkload293 (.A(clknet_leaf_200_clk_i));
 sg13g2_xnor2_1 clone2490 (.Y(net2490),
    .A(_02290_),
    .B(_03016_));
 sg13g2_buf_4 rebuffer2491 (.X(net2491),
    .A(_03665_));
 sg13g2_xnor2_1 clone2494 (.Y(net2494),
    .A(_01877_),
    .B(_02869_));
 sg13g2_buf_4 rebuffer2495 (.X(net2495),
    .A(\cs_registers_i/_2287_ ));
 sg13g2_dlygate4sd3_1 hold2496 (.A(\cs_registers_i/_0000_ ),
    .X(net2496));
 sg13g2_dlygate4sd3_1 hold2497 (.A(\cs_registers_i/dcsr_q_0_ ),
    .X(net2497));
 sg13g2_dlygate4sd3_1 hold2498 (.A(\cs_registers_i/dcsr_q_26_ ),
    .X(net2498));
 sg13g2_dlygate4sd3_1 hold2499 (.A(\cs_registers_i/_0001_ ),
    .X(net2499));
 sg13g2_antennanp ANTENNA_1 (.A(_00602_));
 sg13g2_antennanp ANTENNA_2 (.A(_00620_));
 sg13g2_antennanp ANTENNA_3 (.A(_00638_));
 sg13g2_antennanp ANTENNA_4 (.A(_00654_));
 sg13g2_antennanp ANTENNA_5 (.A(_00713_));
 sg13g2_antennanp ANTENNA_6 (.A(_00735_));
 sg13g2_antennanp ANTENNA_7 (.A(_00753_));
 sg13g2_antennanp ANTENNA_8 (.A(_00780_));
 sg13g2_antennanp ANTENNA_9 (.A(_00785_));
 sg13g2_antennanp ANTENNA_10 (.A(_00834_));
 sg13g2_antennanp ANTENNA_11 (.A(_00857_));
 sg13g2_antennanp ANTENNA_12 (.A(_00878_));
 sg13g2_antennanp ANTENNA_13 (.A(_00904_));
 sg13g2_antennanp ANTENNA_14 (.A(_00941_));
 sg13g2_antennanp ANTENNA_15 (.A(_01002_));
 sg13g2_antennanp ANTENNA_16 (.A(_01031_));
 sg13g2_antennanp ANTENNA_17 (.A(_01085_));
 sg13g2_antennanp ANTENNA_18 (.A(_01173_));
 sg13g2_antennanp ANTENNA_19 (.A(_01306_));
 sg13g2_antennanp ANTENNA_20 (.A(_01475_));
 sg13g2_antennanp ANTENNA_21 (.A(_03318_));
 sg13g2_antennanp ANTENNA_22 (.A(_03550_));
 sg13g2_antennanp ANTENNA_23 (.A(_03564_));
 sg13g2_antennanp ANTENNA_24 (.A(_03564_));
 sg13g2_antennanp ANTENNA_25 (.A(_03564_));
 sg13g2_antennanp ANTENNA_26 (.A(_03564_));
 sg13g2_antennanp ANTENNA_27 (.A(_03605_));
 sg13g2_antennanp ANTENNA_28 (.A(_03605_));
 sg13g2_antennanp ANTENNA_29 (.A(_03605_));
 sg13g2_antennanp ANTENNA_30 (.A(_03610_));
 sg13g2_antennanp ANTENNA_31 (.A(_03610_));
 sg13g2_antennanp ANTENNA_32 (.A(_03684_));
 sg13g2_antennanp ANTENNA_33 (.A(_03684_));
 sg13g2_antennanp ANTENNA_34 (.A(_03695_));
 sg13g2_antennanp ANTENNA_35 (.A(_03712_));
 sg13g2_antennanp ANTENNA_36 (.A(_03719_));
 sg13g2_antennanp ANTENNA_37 (.A(_03724_));
 sg13g2_antennanp ANTENNA_38 (.A(_03730_));
 sg13g2_antennanp ANTENNA_39 (.A(_03797_));
 sg13g2_antennanp ANTENNA_40 (.A(_03838_));
 sg13g2_antennanp ANTENNA_41 (.A(net803));
 sg13g2_antennanp ANTENNA_42 (.A(net803));
 sg13g2_antennanp ANTENNA_43 (.A(net803));
 sg13g2_antennanp ANTENNA_44 (.A(net803));
 sg13g2_antennanp ANTENNA_45 (.A(_08337_));
 sg13g2_antennanp ANTENNA_46 (.A(_08375_));
 sg13g2_antennanp ANTENNA_47 (.A(_08414_));
 sg13g2_antennanp ANTENNA_48 (.A(_08614_));
 sg13g2_antennanp ANTENNA_49 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_50 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_51 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_52 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_53 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_54 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_55 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_56 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_57 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_58 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_59 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_60 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_61 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_62 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_63 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_64 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_65 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_66 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_67 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_68 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_69 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_70 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_71 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_72 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_73 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_74 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_75 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_76 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_77 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_78 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_79 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_80 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_81 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_82 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_83 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_84 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_85 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_86 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_87 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_88 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_89 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_90 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_91 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_92 (.A(boot_addr_i_21_));
 sg13g2_antennanp ANTENNA_93 (.A(boot_addr_i_21_));
 sg13g2_antennanp ANTENNA_94 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_95 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_96 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_97 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_98 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_99 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_100 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_101 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_102 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_103 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_104 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_105 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_106 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_107 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_108 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_109 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_110 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_111 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_112 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_113 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_114 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_115 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_116 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_117 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_118 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_119 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_120 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_121 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_122 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_123 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_124 (.A(crash_dump_o_32_));
 sg13g2_antennanp ANTENNA_125 (.A(crash_dump_o_32_));
 sg13g2_antennanp ANTENNA_126 (.A(crash_dump_o_32_));
 sg13g2_antennanp ANTENNA_127 (.A(crash_dump_o_65_));
 sg13g2_antennanp ANTENNA_128 (.A(crash_dump_o_65_));
 sg13g2_antennanp ANTENNA_129 (.A(crash_dump_o_65_));
 sg13g2_antennanp ANTENNA_130 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_131 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_132 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_133 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_134 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_135 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_136 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_137 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_138 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_139 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_140 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_141 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_142 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_143 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_144 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_145 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_146 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_147 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_148 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_149 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_150 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_151 (.A(crash_dump_o_97_));
 sg13g2_antennanp ANTENNA_152 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_153 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_154 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_155 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_156 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_157 (.A(csr_depc_5_));
 sg13g2_antennanp ANTENNA_158 (.A(csr_depc_5_));
 sg13g2_antennanp ANTENNA_159 (.A(csr_depc_5_));
 sg13g2_antennanp ANTENNA_160 (.A(csr_depc_9_));
 sg13g2_antennanp ANTENNA_161 (.A(csr_depc_9_));
 sg13g2_antennanp ANTENNA_162 (.A(csr_depc_9_));
 sg13g2_antennanp ANTENNA_163 (.A(csr_rdata_16_));
 sg13g2_antennanp ANTENNA_164 (.A(csr_rdata_21_));
 sg13g2_antennanp ANTENNA_165 (.A(data_addr_o_22_));
 sg13g2_antennanp ANTENNA_166 (.A(data_addr_o_22_));
 sg13g2_antennanp ANTENNA_167 (.A(data_addr_o_22_));
 sg13g2_antennanp ANTENNA_168 (.A(data_addr_o_23_));
 sg13g2_antennanp ANTENNA_169 (.A(data_addr_o_23_));
 sg13g2_antennanp ANTENNA_170 (.A(data_addr_o_23_));
 sg13g2_antennanp ANTENNA_171 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_172 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_173 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_174 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_175 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_176 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_177 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_178 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_179 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_180 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_181 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_182 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_183 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_184 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_185 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_186 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_187 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_188 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_189 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_190 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_191 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_192 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_193 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_194 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_195 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_196 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_197 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_198 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_199 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_200 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_201 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_202 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_203 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_204 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_205 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_206 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_207 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_208 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_209 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_210 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_211 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_212 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_antennanp ANTENNA_213 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_antennanp ANTENNA_214 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_antennanp ANTENNA_215 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_antennanp ANTENNA_216 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_13_ ));
 sg13g2_antennanp ANTENNA_217 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_218 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_219 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_220 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_221 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_222 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_223 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_224 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_225 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_226 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_227 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_228 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_229 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_230 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_231 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_232 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_233 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_234 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_235 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_236 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_237 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_238 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_239 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_240 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_241 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_242 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_25_ ));
 sg13g2_antennanp ANTENNA_243 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_244 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_245 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_246 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_247 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_248 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_249 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_250 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_251 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_252 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_253 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_254 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_255 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_256 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_257 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_258 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_259 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_260 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_261 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_262 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_263 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_264 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_265 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_266 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_267 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_268 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_269 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_270 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_271 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_272 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_273 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_274 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_275 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_276 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_277 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_278 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_279 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_280 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_281 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_282 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_283 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_284 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_285 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_286 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_287 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_288 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_289 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_290 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_291 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_292 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_293 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_294 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_295 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_296 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_297 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_298 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_299 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_300 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_301 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_302 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_303 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_304 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_305 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_306 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_307 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_308 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_309 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_310 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_311 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_312 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_313 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_314 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_315 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_316 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_317 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_318 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_319 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_320 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_321 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_322 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_323 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_324 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_325 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_326 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_327 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_328 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_329 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_330 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_331 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_332 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_333 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_334 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_335 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_336 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_337 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ));
 sg13g2_antennanp ANTENNA_338 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_11_ ));
 sg13g2_antennanp ANTENNA_339 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_340 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_341 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_342 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_343 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_344 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_345 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_346 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_347 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_348 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_antennanp ANTENNA_349 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_antennanp ANTENNA_350 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_antennanp ANTENNA_351 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_2_ ));
 sg13g2_antennanp ANTENNA_352 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ));
 sg13g2_antennanp ANTENNA_353 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_354 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_355 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_356 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_357 (.A(fetch_enable_i));
 sg13g2_antennanp ANTENNA_358 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_359 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_360 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_361 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_362 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_363 (.A(hart_id_i_12_));
 sg13g2_antennanp ANTENNA_364 (.A(hart_id_i_13_));
 sg13g2_antennanp ANTENNA_365 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_366 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_367 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_368 (.A(hart_id_i_16_));
 sg13g2_antennanp ANTENNA_369 (.A(hart_id_i_17_));
 sg13g2_antennanp ANTENNA_370 (.A(hart_id_i_18_));
 sg13g2_antennanp ANTENNA_371 (.A(hart_id_i_19_));
 sg13g2_antennanp ANTENNA_372 (.A(hart_id_i_1_));
 sg13g2_antennanp ANTENNA_373 (.A(hart_id_i_20_));
 sg13g2_antennanp ANTENNA_374 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_375 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_376 (.A(hart_id_i_23_));
 sg13g2_antennanp ANTENNA_377 (.A(hart_id_i_24_));
 sg13g2_antennanp ANTENNA_378 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_379 (.A(hart_id_i_26_));
 sg13g2_antennanp ANTENNA_380 (.A(hart_id_i_27_));
 sg13g2_antennanp ANTENNA_381 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_382 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_383 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_384 (.A(hart_id_i_30_));
 sg13g2_antennanp ANTENNA_385 (.A(hart_id_i_31_));
 sg13g2_antennanp ANTENNA_386 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_387 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_388 (.A(hart_id_i_4_));
 sg13g2_antennanp ANTENNA_389 (.A(hart_id_i_5_));
 sg13g2_antennanp ANTENNA_390 (.A(hart_id_i_6_));
 sg13g2_antennanp ANTENNA_391 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_392 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_393 (.A(hart_id_i_8_));
 sg13g2_antennanp ANTENNA_394 (.A(hart_id_i_8_));
 sg13g2_antennanp ANTENNA_395 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_396 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_397 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_398 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_399 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_400 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_401 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_402 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_403 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_404 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_405 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_406 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_407 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_408 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_409 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_410 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_411 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_412 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_413 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_414 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_415 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_416 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_417 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_418 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_419 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_420 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_421 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_422 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_423 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_424 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_425 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_426 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_427 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_428 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_429 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_430 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_431 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_432 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_433 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_434 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_435 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_436 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_437 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_438 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_439 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_440 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_441 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_442 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_443 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_444 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_445 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_446 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_447 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_448 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_449 (.A(irq_fast_i_4_));
 sg13g2_antennanp ANTENNA_450 (.A(irq_fast_i_4_));
 sg13g2_antennanp ANTENNA_451 (.A(irq_fast_i_4_));
 sg13g2_antennanp ANTENNA_452 (.A(irq_fast_i_4_));
 sg13g2_antennanp ANTENNA_453 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_454 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_455 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_456 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_457 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_458 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_459 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_460 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_461 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_462 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_463 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_464 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_465 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_466 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_467 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_468 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_469 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_470 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_471 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_472 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_473 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_474 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_475 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_476 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_477 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_478 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_479 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_480 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_481 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_482 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_483 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_484 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_485 (.A(perf_instr_ret_wb));
 sg13g2_antennanp ANTENNA_486 (.A(perf_instr_ret_wb));
 sg13g2_antennanp ANTENNA_487 (.A(perf_instr_ret_wb));
 sg13g2_antennanp ANTENNA_488 (.A(rf_wdata_wb_23_));
 sg13g2_antennanp ANTENNA_489 (.A(rf_wdata_wb_25_));
 sg13g2_antennanp ANTENNA_490 (.A(rf_wdata_wb_25_));
 sg13g2_antennanp ANTENNA_491 (.A(rf_wdata_wb_25_));
 sg13g2_antennanp ANTENNA_492 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_493 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_494 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_495 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_496 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_497 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_498 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_499 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_500 (.A(rf_wdata_wb_28_));
 sg13g2_antennanp ANTENNA_501 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_502 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_503 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_504 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_505 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_506 (.A(\cs_registers_i/_1034_ ));
 sg13g2_antennanp ANTENNA_507 (.A(\cs_registers_i/_1034_ ));
 sg13g2_antennanp ANTENNA_508 (.A(net513));
 sg13g2_antennanp ANTENNA_509 (.A(net513));
 sg13g2_antennanp ANTENNA_510 (.A(net513));
 sg13g2_antennanp ANTENNA_511 (.A(net513));
 sg13g2_antennanp ANTENNA_512 (.A(net513));
 sg13g2_antennanp ANTENNA_513 (.A(net513));
 sg13g2_antennanp ANTENNA_514 (.A(net513));
 sg13g2_antennanp ANTENNA_515 (.A(net513));
 sg13g2_antennanp ANTENNA_516 (.A(net513));
 sg13g2_antennanp ANTENNA_517 (.A(\cs_registers_i/_1694_ ));
 sg13g2_antennanp ANTENNA_518 (.A(\cs_registers_i/_1694_ ));
 sg13g2_antennanp ANTENNA_519 (.A(\cs_registers_i/_1694_ ));
 sg13g2_antennanp ANTENNA_520 (.A(\cs_registers_i/_1694_ ));
 sg13g2_antennanp ANTENNA_521 (.A(\register_file_i/_1893_ ));
 sg13g2_antennanp ANTENNA_522 (.A(\register_file_i/_2795_ ));
 sg13g2_antennanp ANTENNA_523 (.A(net149));
 sg13g2_antennanp ANTENNA_524 (.A(net149));
 sg13g2_antennanp ANTENNA_525 (.A(net149));
 sg13g2_antennanp ANTENNA_526 (.A(net149));
 sg13g2_antennanp ANTENNA_527 (.A(net149));
 sg13g2_antennanp ANTENNA_528 (.A(net149));
 sg13g2_antennanp ANTENNA_529 (.A(net149));
 sg13g2_antennanp ANTENNA_530 (.A(net149));
 sg13g2_antennanp ANTENNA_531 (.A(net86));
 sg13g2_antennanp ANTENNA_532 (.A(net86));
 sg13g2_antennanp ANTENNA_533 (.A(net86));
 sg13g2_antennanp ANTENNA_534 (.A(net86));
 sg13g2_antennanp ANTENNA_535 (.A(net86));
 sg13g2_antennanp ANTENNA_536 (.A(net86));
 sg13g2_antennanp ANTENNA_537 (.A(net86));
 sg13g2_antennanp ANTENNA_538 (.A(net86));
 sg13g2_antennanp ANTENNA_539 (.A(net1499));
 sg13g2_antennanp ANTENNA_540 (.A(net1499));
 sg13g2_antennanp ANTENNA_541 (.A(net1499));
 sg13g2_antennanp ANTENNA_542 (.A(net1499));
 sg13g2_antennanp ANTENNA_543 (.A(net1499));
 sg13g2_antennanp ANTENNA_544 (.A(net1499));
 sg13g2_antennanp ANTENNA_545 (.A(net1516));
 sg13g2_antennanp ANTENNA_546 (.A(net1516));
 sg13g2_antennanp ANTENNA_547 (.A(net1516));
 sg13g2_antennanp ANTENNA_548 (.A(net1516));
 sg13g2_antennanp ANTENNA_549 (.A(net1516));
 sg13g2_antennanp ANTENNA_550 (.A(net1516));
 sg13g2_antennanp ANTENNA_551 (.A(net1516));
 sg13g2_antennanp ANTENNA_552 (.A(net1516));
 sg13g2_antennanp ANTENNA_553 (.A(net1516));
 sg13g2_antennanp ANTENNA_554 (.A(net1516));
 sg13g2_antennanp ANTENNA_555 (.A(net1516));
 sg13g2_antennanp ANTENNA_556 (.A(net1651));
 sg13g2_antennanp ANTENNA_557 (.A(net1651));
 sg13g2_antennanp ANTENNA_558 (.A(net1651));
 sg13g2_antennanp ANTENNA_559 (.A(net1651));
 sg13g2_antennanp ANTENNA_560 (.A(net1651));
 sg13g2_antennanp ANTENNA_561 (.A(net1651));
 sg13g2_antennanp ANTENNA_562 (.A(net1651));
 sg13g2_antennanp ANTENNA_563 (.A(net1651));
 sg13g2_antennanp ANTENNA_564 (.A(net2006));
 sg13g2_antennanp ANTENNA_565 (.A(net2006));
 sg13g2_antennanp ANTENNA_566 (.A(net2006));
 sg13g2_antennanp ANTENNA_567 (.A(net2006));
 sg13g2_antennanp ANTENNA_568 (.A(net2465));
 sg13g2_antennanp ANTENNA_569 (.A(net2465));
 sg13g2_antennanp ANTENNA_570 (.A(net2465));
 sg13g2_antennanp ANTENNA_571 (.A(net2465));
 sg13g2_antennanp ANTENNA_572 (.A(net2465));
 sg13g2_antennanp ANTENNA_573 (.A(net2465));
 sg13g2_antennanp ANTENNA_574 (.A(net2490));
 sg13g2_antennanp ANTENNA_575 (.A(net2490));
 sg13g2_antennanp ANTENNA_576 (.A(net2490));
 sg13g2_antennanp ANTENNA_577 (.A(_00602_));
 sg13g2_antennanp ANTENNA_578 (.A(_00620_));
 sg13g2_antennanp ANTENNA_579 (.A(_00638_));
 sg13g2_antennanp ANTENNA_580 (.A(_00713_));
 sg13g2_antennanp ANTENNA_581 (.A(_00735_));
 sg13g2_antennanp ANTENNA_582 (.A(_00753_));
 sg13g2_antennanp ANTENNA_583 (.A(_00780_));
 sg13g2_antennanp ANTENNA_584 (.A(_00785_));
 sg13g2_antennanp ANTENNA_585 (.A(_00834_));
 sg13g2_antennanp ANTENNA_586 (.A(_00857_));
 sg13g2_antennanp ANTENNA_587 (.A(_00904_));
 sg13g2_antennanp ANTENNA_588 (.A(_00941_));
 sg13g2_antennanp ANTENNA_589 (.A(_01002_));
 sg13g2_antennanp ANTENNA_590 (.A(_01002_));
 sg13g2_antennanp ANTENNA_591 (.A(_01031_));
 sg13g2_antennanp ANTENNA_592 (.A(_01085_));
 sg13g2_antennanp ANTENNA_593 (.A(_01306_));
 sg13g2_antennanp ANTENNA_594 (.A(_01475_));
 sg13g2_antennanp ANTENNA_595 (.A(_03318_));
 sg13g2_antennanp ANTENNA_596 (.A(_03550_));
 sg13g2_antennanp ANTENNA_597 (.A(_03610_));
 sg13g2_antennanp ANTENNA_598 (.A(_03610_));
 sg13g2_antennanp ANTENNA_599 (.A(_03657_));
 sg13g2_antennanp ANTENNA_600 (.A(_03657_));
 sg13g2_antennanp ANTENNA_601 (.A(_03684_));
 sg13g2_antennanp ANTENNA_602 (.A(_03695_));
 sg13g2_antennanp ANTENNA_603 (.A(_03695_));
 sg13g2_antennanp ANTENNA_604 (.A(_03719_));
 sg13g2_antennanp ANTENNA_605 (.A(_03797_));
 sg13g2_antennanp ANTENNA_606 (.A(_03838_));
 sg13g2_antennanp ANTENNA_607 (.A(_08337_));
 sg13g2_antennanp ANTENNA_608 (.A(_08375_));
 sg13g2_antennanp ANTENNA_609 (.A(_08414_));
 sg13g2_antennanp ANTENNA_610 (.A(_08614_));
 sg13g2_antennanp ANTENNA_611 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_612 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_613 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_614 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_615 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_616 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_617 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_618 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_619 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_620 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_621 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_622 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_623 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_624 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_625 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_626 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_627 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_628 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_629 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_630 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_631 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_632 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_633 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_634 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_635 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_636 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_637 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_638 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_639 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_640 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_641 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_642 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_643 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_644 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_645 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_646 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_647 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_648 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_649 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_650 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_651 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_652 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_653 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_654 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_655 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_656 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_657 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_658 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_659 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_660 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_661 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_662 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_663 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_664 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_665 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_666 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_667 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_668 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_669 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_670 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_671 (.A(boot_addr_i_29_));
 sg13g2_antennanp ANTENNA_672 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_673 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_674 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_675 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_676 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_677 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_678 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_679 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_680 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_681 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_682 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_683 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_684 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_685 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_686 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_687 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_688 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_689 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_690 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_691 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_692 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_693 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_694 (.A(csr_rdata_16_));
 sg13g2_antennanp ANTENNA_695 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_696 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_697 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_698 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_699 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_700 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_701 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_702 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_703 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_704 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_705 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_706 (.A(data_addr_o_19_));
 sg13g2_antennanp ANTENNA_707 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_708 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_709 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_710 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_711 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_712 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_713 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_714 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_715 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_716 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_717 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_718 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_719 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_720 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_721 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_722 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_723 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_724 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_725 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_726 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_727 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_728 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_729 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_730 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_731 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_732 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_733 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_734 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_735 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_736 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_1_ ));
 sg13g2_antennanp ANTENNA_737 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_738 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_739 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_740 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_741 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_742 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_743 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_744 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_20_ ));
 sg13g2_antennanp ANTENNA_745 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_746 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_747 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_748 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_749 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_750 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_751 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_752 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_753 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_754 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_755 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_756 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_757 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_758 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_759 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_760 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_761 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_762 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_763 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_764 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_765 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_766 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_767 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_768 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_769 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_770 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_771 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_772 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_773 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_774 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_775 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_776 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_777 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_778 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_779 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_780 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_781 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_782 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_783 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_784 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_785 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_786 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_787 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_788 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_789 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_790 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_791 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_792 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_793 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_794 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_795 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_796 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_797 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_798 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_799 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_800 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_801 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_802 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_803 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_804 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_805 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_806 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_807 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_808 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_809 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_810 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_811 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_812 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_813 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_814 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_815 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_816 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_817 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_818 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_819 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_820 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_821 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_822 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_823 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_824 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_825 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_826 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_827 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_828 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_829 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_830 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_831 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_832 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_833 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_834 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_835 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_836 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_837 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_838 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_839 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_840 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_841 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_842 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_8_ ));
 sg13g2_antennanp ANTENNA_843 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_844 (.A(fetch_enable_i));
 sg13g2_antennanp ANTENNA_845 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_846 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_847 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_848 (.A(hart_id_i_12_));
 sg13g2_antennanp ANTENNA_849 (.A(hart_id_i_13_));
 sg13g2_antennanp ANTENNA_850 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_851 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_852 (.A(hart_id_i_16_));
 sg13g2_antennanp ANTENNA_853 (.A(hart_id_i_17_));
 sg13g2_antennanp ANTENNA_854 (.A(hart_id_i_18_));
 sg13g2_antennanp ANTENNA_855 (.A(hart_id_i_19_));
 sg13g2_antennanp ANTENNA_856 (.A(hart_id_i_1_));
 sg13g2_antennanp ANTENNA_857 (.A(hart_id_i_20_));
 sg13g2_antennanp ANTENNA_858 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_859 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_860 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_861 (.A(hart_id_i_23_));
 sg13g2_antennanp ANTENNA_862 (.A(hart_id_i_24_));
 sg13g2_antennanp ANTENNA_863 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_864 (.A(hart_id_i_26_));
 sg13g2_antennanp ANTENNA_865 (.A(hart_id_i_27_));
 sg13g2_antennanp ANTENNA_866 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_867 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_868 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_869 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_870 (.A(hart_id_i_30_));
 sg13g2_antennanp ANTENNA_871 (.A(hart_id_i_31_));
 sg13g2_antennanp ANTENNA_872 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_873 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_874 (.A(hart_id_i_4_));
 sg13g2_antennanp ANTENNA_875 (.A(hart_id_i_5_));
 sg13g2_antennanp ANTENNA_876 (.A(hart_id_i_5_));
 sg13g2_antennanp ANTENNA_877 (.A(hart_id_i_6_));
 sg13g2_antennanp ANTENNA_878 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_879 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_880 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_881 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_882 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_883 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_884 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_885 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_886 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_887 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_888 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_889 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_890 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_891 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_892 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_893 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_894 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_895 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_896 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_897 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_898 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_899 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_900 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_901 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_902 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_903 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_904 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_905 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_906 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_907 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_908 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_909 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_910 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_911 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_912 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_913 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_914 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_915 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_916 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_917 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_918 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_919 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_920 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_921 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_922 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_923 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_924 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_925 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_926 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_927 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_928 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_929 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_930 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_931 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_932 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_933 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_934 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_935 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_936 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_937 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_938 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_939 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_940 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_941 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_942 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_943 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_944 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_945 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_946 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_947 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_948 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_949 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_950 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_951 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_952 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_953 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_954 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_955 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_956 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_957 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_958 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_959 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_960 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_961 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_962 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_963 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_964 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_965 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_966 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_967 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_968 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_969 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_970 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_971 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_972 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_973 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_974 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_975 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_976 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_977 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_978 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_979 (.A(rf_wdata_wb_23_));
 sg13g2_antennanp ANTENNA_980 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_981 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_982 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_983 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_984 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_985 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_986 (.A(net513));
 sg13g2_antennanp ANTENNA_987 (.A(net513));
 sg13g2_antennanp ANTENNA_988 (.A(net513));
 sg13g2_antennanp ANTENNA_989 (.A(net513));
 sg13g2_antennanp ANTENNA_990 (.A(net513));
 sg13g2_antennanp ANTENNA_991 (.A(net513));
 sg13g2_antennanp ANTENNA_992 (.A(net513));
 sg13g2_antennanp ANTENNA_993 (.A(net513));
 sg13g2_antennanp ANTENNA_994 (.A(net1516));
 sg13g2_antennanp ANTENNA_995 (.A(net1516));
 sg13g2_antennanp ANTENNA_996 (.A(net1516));
 sg13g2_antennanp ANTENNA_997 (.A(net1516));
 sg13g2_antennanp ANTENNA_998 (.A(net2465));
 sg13g2_antennanp ANTENNA_999 (.A(net2465));
 sg13g2_antennanp ANTENNA_1000 (.A(net2465));
 sg13g2_antennanp ANTENNA_1001 (.A(net2465));
 sg13g2_antennanp ANTENNA_1002 (.A(net2465));
 sg13g2_antennanp ANTENNA_1003 (.A(net2465));
 sg13g2_antennanp ANTENNA_1004 (.A(_00602_));
 sg13g2_antennanp ANTENNA_1005 (.A(_00620_));
 sg13g2_antennanp ANTENNA_1006 (.A(_00638_));
 sg13g2_antennanp ANTENNA_1007 (.A(_00654_));
 sg13g2_antennanp ANTENNA_1008 (.A(_00713_));
 sg13g2_antennanp ANTENNA_1009 (.A(_00735_));
 sg13g2_antennanp ANTENNA_1010 (.A(_00780_));
 sg13g2_antennanp ANTENNA_1011 (.A(_00785_));
 sg13g2_antennanp ANTENNA_1012 (.A(_00834_));
 sg13g2_antennanp ANTENNA_1013 (.A(_00857_));
 sg13g2_antennanp ANTENNA_1014 (.A(_00904_));
 sg13g2_antennanp ANTENNA_1015 (.A(_01031_));
 sg13g2_antennanp ANTENNA_1016 (.A(_01306_));
 sg13g2_antennanp ANTENNA_1017 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1018 (.A(_03550_));
 sg13g2_antennanp ANTENNA_1019 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1020 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1021 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1022 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1023 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1024 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1025 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1026 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1027 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1028 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1029 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1030 (.A(_03719_));
 sg13g2_antennanp ANTENNA_1031 (.A(_03797_));
 sg13g2_antennanp ANTENNA_1032 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1033 (.A(_08337_));
 sg13g2_antennanp ANTENNA_1034 (.A(_08337_));
 sg13g2_antennanp ANTENNA_1035 (.A(_08375_));
 sg13g2_antennanp ANTENNA_1036 (.A(_08414_));
 sg13g2_antennanp ANTENNA_1037 (.A(_08614_));
 sg13g2_antennanp ANTENNA_1038 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1039 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1040 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1041 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1042 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1043 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1044 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1045 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1046 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1047 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1048 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1049 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1050 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1051 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1052 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1053 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1054 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1055 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1056 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1057 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1058 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1059 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1060 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1061 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1062 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1063 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1064 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1065 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1066 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1067 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1068 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1069 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1070 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1071 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1072 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1073 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1074 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1075 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1076 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1077 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1078 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1079 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1080 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1081 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1082 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1083 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1084 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1085 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1086 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1087 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1088 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1089 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1090 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1091 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_1092 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_1093 (.A(boot_addr_i_31_));
 sg13g2_antennanp ANTENNA_1094 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1095 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1096 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1097 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1098 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1099 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1100 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1101 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1102 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1103 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1104 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1105 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1106 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1107 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1108 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1109 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1110 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1111 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1112 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1113 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1114 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1115 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1116 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1117 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1118 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1119 (.A(data_addr_o_9_));
 sg13g2_antennanp ANTENNA_1120 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1121 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1122 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1123 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1124 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1125 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1126 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1127 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1128 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1129 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1130 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1131 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1132 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1133 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1134 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1135 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1136 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1137 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1138 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1139 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1140 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1141 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1142 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1143 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1144 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1145 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1146 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1147 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1148 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1149 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1150 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1151 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1152 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1153 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1154 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1155 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1156 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1157 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1158 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1159 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1160 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1161 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1162 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1163 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1164 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1165 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1166 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1167 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1168 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1169 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1170 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1171 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1172 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1173 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1174 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1175 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1176 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1177 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1178 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1179 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1180 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_1181 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_1182 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_8_ ));
 sg13g2_antennanp ANTENNA_1183 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1184 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1185 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1186 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1187 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1188 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1189 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1190 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1191 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1192 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1193 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1194 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1195 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1196 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1197 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1198 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1199 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1200 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1201 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1202 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1203 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1204 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1205 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1206 (.A(fetch_enable_i));
 sg13g2_antennanp ANTENNA_1207 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_1208 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_1209 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_1210 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_1211 (.A(hart_id_i_12_));
 sg13g2_antennanp ANTENNA_1212 (.A(hart_id_i_13_));
 sg13g2_antennanp ANTENNA_1213 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_1214 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_1215 (.A(hart_id_i_16_));
 sg13g2_antennanp ANTENNA_1216 (.A(hart_id_i_18_));
 sg13g2_antennanp ANTENNA_1217 (.A(hart_id_i_19_));
 sg13g2_antennanp ANTENNA_1218 (.A(hart_id_i_1_));
 sg13g2_antennanp ANTENNA_1219 (.A(hart_id_i_20_));
 sg13g2_antennanp ANTENNA_1220 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1221 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1222 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_1223 (.A(hart_id_i_23_));
 sg13g2_antennanp ANTENNA_1224 (.A(hart_id_i_24_));
 sg13g2_antennanp ANTENNA_1225 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_1226 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_1227 (.A(hart_id_i_27_));
 sg13g2_antennanp ANTENNA_1228 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_1229 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_1230 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1231 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1232 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1233 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1234 (.A(hart_id_i_30_));
 sg13g2_antennanp ANTENNA_1235 (.A(hart_id_i_31_));
 sg13g2_antennanp ANTENNA_1236 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1237 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1238 (.A(hart_id_i_4_));
 sg13g2_antennanp ANTENNA_1239 (.A(hart_id_i_5_));
 sg13g2_antennanp ANTENNA_1240 (.A(hart_id_i_5_));
 sg13g2_antennanp ANTENNA_1241 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_1242 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_1243 (.A(hart_id_i_8_));
 sg13g2_antennanp ANTENNA_1244 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_1245 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_1246 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1247 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1248 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1249 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1250 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1251 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1252 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1253 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_1254 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_1255 (.A(irq_fast_i_10_));
 sg13g2_antennanp ANTENNA_1256 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1257 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1258 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1259 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1260 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1261 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1262 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1263 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1264 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1265 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1266 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1267 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1268 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1269 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1270 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1271 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1272 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1273 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1274 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1275 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1276 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1277 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1278 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1279 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1280 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1281 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1282 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1283 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1284 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1285 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1286 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1287 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1288 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1289 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1290 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1291 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1292 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1293 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1294 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1295 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1296 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1297 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1298 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1299 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1300 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1301 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1302 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1303 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1304 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1305 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1306 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1307 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1308 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1309 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1310 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1311 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1312 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1313 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1314 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1315 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_1316 (.A(irq_pending_o));
 sg13g2_antennanp ANTENNA_1317 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1318 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1319 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1320 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1321 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1322 (.A(rf_wdata_wb_23_));
 sg13g2_antennanp ANTENNA_1323 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1324 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1325 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1326 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1327 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1328 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1329 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1330 (.A(net513));
 sg13g2_antennanp ANTENNA_1331 (.A(net513));
 sg13g2_antennanp ANTENNA_1332 (.A(net513));
 sg13g2_antennanp ANTENNA_1333 (.A(net513));
 sg13g2_antennanp ANTENNA_1334 (.A(net513));
 sg13g2_antennanp ANTENNA_1335 (.A(net513));
 sg13g2_antennanp ANTENNA_1336 (.A(net513));
 sg13g2_antennanp ANTENNA_1337 (.A(net513));
 sg13g2_antennanp ANTENNA_1338 (.A(net2465));
 sg13g2_antennanp ANTENNA_1339 (.A(net2465));
 sg13g2_antennanp ANTENNA_1340 (.A(net2465));
 sg13g2_antennanp ANTENNA_1341 (.A(net2465));
 sg13g2_antennanp ANTENNA_1342 (.A(net2465));
 sg13g2_antennanp ANTENNA_1343 (.A(net2465));
 sg13g2_antennanp ANTENNA_1344 (.A(net2465));
 sg13g2_antennanp ANTENNA_1345 (.A(net2465));
 sg13g2_antennanp ANTENNA_1346 (.A(net2465));
 sg13g2_antennanp ANTENNA_1347 (.A(net2465));
 sg13g2_antennanp ANTENNA_1348 (.A(_00602_));
 sg13g2_antennanp ANTENNA_1349 (.A(_00620_));
 sg13g2_antennanp ANTENNA_1350 (.A(_00638_));
 sg13g2_antennanp ANTENNA_1351 (.A(_00654_));
 sg13g2_antennanp ANTENNA_1352 (.A(_00713_));
 sg13g2_antennanp ANTENNA_1353 (.A(_00735_));
 sg13g2_antennanp ANTENNA_1354 (.A(_00780_));
 sg13g2_antennanp ANTENNA_1355 (.A(_00785_));
 sg13g2_antennanp ANTENNA_1356 (.A(_00834_));
 sg13g2_antennanp ANTENNA_1357 (.A(_00857_));
 sg13g2_antennanp ANTENNA_1358 (.A(_00904_));
 sg13g2_antennanp ANTENNA_1359 (.A(_01031_));
 sg13g2_antennanp ANTENNA_1360 (.A(_01306_));
 sg13g2_antennanp ANTENNA_1361 (.A(_03318_));
 sg13g2_antennanp ANTENNA_1362 (.A(_03550_));
 sg13g2_antennanp ANTENNA_1363 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1364 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1365 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1366 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1367 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1368 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1369 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1370 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1371 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1372 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1373 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1374 (.A(_03719_));
 sg13g2_antennanp ANTENNA_1375 (.A(_03797_));
 sg13g2_antennanp ANTENNA_1376 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1377 (.A(_08337_));
 sg13g2_antennanp ANTENNA_1378 (.A(_08375_));
 sg13g2_antennanp ANTENNA_1379 (.A(_08414_));
 sg13g2_antennanp ANTENNA_1380 (.A(_08614_));
 sg13g2_antennanp ANTENNA_1381 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1382 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1383 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1384 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1385 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1386 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1387 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1388 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1389 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1390 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1391 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1392 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1393 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1394 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1395 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1396 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1397 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1398 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1399 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1400 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1401 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1402 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1403 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1404 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1405 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1406 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1407 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1408 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1409 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1410 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1411 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1412 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1413 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1414 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1415 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1416 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1417 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1418 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1419 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1420 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1421 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1422 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1423 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1424 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1425 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1426 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1427 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1428 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1429 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1430 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1431 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1432 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1433 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1434 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1435 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1436 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1437 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1438 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1439 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1440 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1441 (.A(boot_addr_i_25_));
 sg13g2_antennanp ANTENNA_1442 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1443 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1444 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1445 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1446 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1447 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1448 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1449 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1450 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1451 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1452 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1453 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1454 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1455 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1456 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1457 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1458 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1459 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1460 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1461 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1462 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1463 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1464 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1465 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1466 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1467 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1468 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1469 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1470 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1471 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1472 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1473 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1474 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1475 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1476 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1477 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1478 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1479 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1480 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1481 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1482 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1483 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1484 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1485 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1486 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1487 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1488 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1489 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_27_ ));
 sg13g2_antennanp ANTENNA_1490 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1491 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1492 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1493 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1494 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1495 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1496 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1497 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1498 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1499 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1500 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1501 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1502 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1503 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_29_ ));
 sg13g2_antennanp ANTENNA_1504 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1505 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1506 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1507 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1508 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1509 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1510 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1511 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1512 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1513 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1514 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1515 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1516 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1517 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1518 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1519 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1520 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1521 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1522 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1523 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1524 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1525 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1526 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1527 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1528 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1529 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1530 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1531 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1532 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1533 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1534 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1535 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1536 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1537 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1538 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1539 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1540 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1541 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1542 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1543 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1544 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1545 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1546 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_9_ ));
 sg13g2_antennanp ANTENNA_1547 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1548 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1549 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1550 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1551 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1552 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1553 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1554 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1555 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1556 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_1557 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_1558 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_1559 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_1560 (.A(exc_cause_6_));
 sg13g2_antennanp ANTENNA_1561 (.A(fetch_enable_i));
 sg13g2_antennanp ANTENNA_1562 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_1563 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_1564 (.A(hart_id_i_10_));
 sg13g2_antennanp ANTENNA_1565 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_1566 (.A(hart_id_i_12_));
 sg13g2_antennanp ANTENNA_1567 (.A(hart_id_i_13_));
 sg13g2_antennanp ANTENNA_1568 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_1569 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_1570 (.A(hart_id_i_16_));
 sg13g2_antennanp ANTENNA_1571 (.A(hart_id_i_18_));
 sg13g2_antennanp ANTENNA_1572 (.A(hart_id_i_19_));
 sg13g2_antennanp ANTENNA_1573 (.A(hart_id_i_1_));
 sg13g2_antennanp ANTENNA_1574 (.A(hart_id_i_20_));
 sg13g2_antennanp ANTENNA_1575 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1576 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1577 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_1578 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_1579 (.A(hart_id_i_23_));
 sg13g2_antennanp ANTENNA_1580 (.A(hart_id_i_24_));
 sg13g2_antennanp ANTENNA_1581 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_1582 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_1583 (.A(hart_id_i_27_));
 sg13g2_antennanp ANTENNA_1584 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_1585 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_1586 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1587 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1588 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1589 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1590 (.A(hart_id_i_30_));
 sg13g2_antennanp ANTENNA_1591 (.A(hart_id_i_31_));
 sg13g2_antennanp ANTENNA_1592 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1593 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1594 (.A(hart_id_i_4_));
 sg13g2_antennanp ANTENNA_1595 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_1596 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_1597 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_1598 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_1599 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1600 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1601 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1602 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1603 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1604 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1605 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1606 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1607 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1608 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1609 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1610 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1611 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1612 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1613 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1614 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1615 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1616 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1617 (.A(irq_fast_i_12_));
 sg13g2_antennanp ANTENNA_1618 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1619 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1620 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1621 (.A(irq_fast_i_14_));
 sg13g2_antennanp ANTENNA_1622 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1623 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1624 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1625 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1626 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1627 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1628 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1629 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1630 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1631 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1632 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1633 (.A(irq_fast_i_3_));
 sg13g2_antennanp ANTENNA_1634 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1635 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1636 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1637 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1638 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1639 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1640 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1641 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1642 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1643 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1644 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1645 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1646 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1647 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1648 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1649 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1650 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1651 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1652 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1653 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1654 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1655 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1656 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1657 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1658 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1659 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1660 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1661 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1662 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1663 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1664 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1665 (.A(rf_wdata_wb_23_));
 sg13g2_antennanp ANTENNA_1666 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1667 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1668 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1669 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1670 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1671 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1672 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1673 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_1674 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_1675 (.A(net2465));
 sg13g2_antennanp ANTENNA_1676 (.A(net2465));
 sg13g2_antennanp ANTENNA_1677 (.A(net2465));
 sg13g2_antennanp ANTENNA_1678 (.A(net2465));
 sg13g2_antennanp ANTENNA_1679 (.A(net2465));
 sg13g2_antennanp ANTENNA_1680 (.A(net2465));
 sg13g2_antennanp ANTENNA_1681 (.A(net2465));
 sg13g2_antennanp ANTENNA_1682 (.A(_00602_));
 sg13g2_antennanp ANTENNA_1683 (.A(_00620_));
 sg13g2_antennanp ANTENNA_1684 (.A(_00638_));
 sg13g2_antennanp ANTENNA_1685 (.A(_00654_));
 sg13g2_antennanp ANTENNA_1686 (.A(_00713_));
 sg13g2_antennanp ANTENNA_1687 (.A(_00735_));
 sg13g2_antennanp ANTENNA_1688 (.A(_00780_));
 sg13g2_antennanp ANTENNA_1689 (.A(_00785_));
 sg13g2_antennanp ANTENNA_1690 (.A(_00834_));
 sg13g2_antennanp ANTENNA_1691 (.A(_00834_));
 sg13g2_antennanp ANTENNA_1692 (.A(_00857_));
 sg13g2_antennanp ANTENNA_1693 (.A(_00904_));
 sg13g2_antennanp ANTENNA_1694 (.A(_01031_));
 sg13g2_antennanp ANTENNA_1695 (.A(_01306_));
 sg13g2_antennanp ANTENNA_1696 (.A(_03550_));
 sg13g2_antennanp ANTENNA_1697 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1698 (.A(_03610_));
 sg13g2_antennanp ANTENNA_1699 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1700 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1701 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1702 (.A(_03630_));
 sg13g2_antennanp ANTENNA_1703 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1704 (.A(_03657_));
 sg13g2_antennanp ANTENNA_1705 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1706 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1707 (.A(_03695_));
 sg13g2_antennanp ANTENNA_1708 (.A(_03719_));
 sg13g2_antennanp ANTENNA_1709 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1710 (.A(_03838_));
 sg13g2_antennanp ANTENNA_1711 (.A(_08337_));
 sg13g2_antennanp ANTENNA_1712 (.A(_08375_));
 sg13g2_antennanp ANTENNA_1713 (.A(_08414_));
 sg13g2_antennanp ANTENNA_1714 (.A(_08614_));
 sg13g2_antennanp ANTENNA_1715 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1716 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1717 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1718 (.A(boot_addr_i_10_));
 sg13g2_antennanp ANTENNA_1719 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1720 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1721 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1722 (.A(boot_addr_i_11_));
 sg13g2_antennanp ANTENNA_1723 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1724 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1725 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1726 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1727 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1728 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1729 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1730 (.A(boot_addr_i_12_));
 sg13g2_antennanp ANTENNA_1731 (.A(boot_addr_i_13_));
 sg13g2_antennanp ANTENNA_1732 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1733 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1734 (.A(boot_addr_i_14_));
 sg13g2_antennanp ANTENNA_1735 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1736 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1737 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1738 (.A(boot_addr_i_15_));
 sg13g2_antennanp ANTENNA_1739 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1740 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1741 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1742 (.A(boot_addr_i_16_));
 sg13g2_antennanp ANTENNA_1743 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1744 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1745 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1746 (.A(boot_addr_i_17_));
 sg13g2_antennanp ANTENNA_1747 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1748 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1749 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1750 (.A(boot_addr_i_18_));
 sg13g2_antennanp ANTENNA_1751 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1752 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1753 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1754 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1755 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1756 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1757 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1758 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1759 (.A(boot_addr_i_20_));
 sg13g2_antennanp ANTENNA_1760 (.A(boot_addr_i_21_));
 sg13g2_antennanp ANTENNA_1761 (.A(boot_addr_i_21_));
 sg13g2_antennanp ANTENNA_1762 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1763 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1764 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1765 (.A(boot_addr_i_22_));
 sg13g2_antennanp ANTENNA_1766 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1767 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1768 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1769 (.A(boot_addr_i_23_));
 sg13g2_antennanp ANTENNA_1770 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1771 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1772 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1773 (.A(boot_addr_i_26_));
 sg13g2_antennanp ANTENNA_1774 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1775 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1776 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1777 (.A(boot_addr_i_27_));
 sg13g2_antennanp ANTENNA_1778 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1779 (.A(boot_addr_i_30_));
 sg13g2_antennanp ANTENNA_1780 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1781 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1782 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1783 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1784 (.A(boot_addr_i_9_));
 sg13g2_antennanp ANTENNA_1785 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1786 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1787 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1788 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1789 (.A(crash_dump_o_24_));
 sg13g2_antennanp ANTENNA_1790 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1791 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1792 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1793 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1794 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1795 (.A(crash_dump_o_8_));
 sg13g2_antennanp ANTENNA_1796 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1797 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1798 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1799 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1800 (.A(crash_dump_o_9_));
 sg13g2_antennanp ANTENNA_1801 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1802 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1803 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1804 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1805 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_10_ ));
 sg13g2_antennanp ANTENNA_1806 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1807 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1808 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1809 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1810 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1811 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_11_ ));
 sg13g2_antennanp ANTENNA_1812 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1813 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1814 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1815 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1816 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1817 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_15_ ));
 sg13g2_antennanp ANTENNA_1818 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1819 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1820 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1821 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1822 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1823 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_26_ ));
 sg13g2_antennanp ANTENNA_1824 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1825 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1826 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1827 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1828 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1829 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1830 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_2_ ));
 sg13g2_antennanp ANTENNA_1831 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_3_ ));
 sg13g2_antennanp ANTENNA_1832 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1833 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1834 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1835 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1836 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1837 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1838 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1839 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_4_ ));
 sg13g2_antennanp ANTENNA_1840 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1841 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1842 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1843 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1844 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1845 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1846 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1847 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1848 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1849 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1850 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1851 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_6_ ));
 sg13g2_antennanp ANTENNA_1852 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1853 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1854 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1855 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1856 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1857 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1858 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1859 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1860 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1861 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1862 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1863 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1864 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1865 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_a_i_7_ ));
 sg13g2_antennanp ANTENNA_1866 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1867 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1868 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1869 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_19_ ));
 sg13g2_antennanp ANTENNA_1870 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1871 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1872 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1873 (.A(\ex_block_i.gen_multdiv_fast.multdiv_i.op_b_i_20_ ));
 sg13g2_antennanp ANTENNA_1874 (.A(fetch_enable_i));
 sg13g2_antennanp ANTENNA_1875 (.A(hart_id_i_0_));
 sg13g2_antennanp ANTENNA_1876 (.A(hart_id_i_11_));
 sg13g2_antennanp ANTENNA_1877 (.A(hart_id_i_12_));
 sg13g2_antennanp ANTENNA_1878 (.A(hart_id_i_13_));
 sg13g2_antennanp ANTENNA_1879 (.A(hart_id_i_14_));
 sg13g2_antennanp ANTENNA_1880 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_1881 (.A(hart_id_i_15_));
 sg13g2_antennanp ANTENNA_1882 (.A(hart_id_i_16_));
 sg13g2_antennanp ANTENNA_1883 (.A(hart_id_i_18_));
 sg13g2_antennanp ANTENNA_1884 (.A(hart_id_i_19_));
 sg13g2_antennanp ANTENNA_1885 (.A(hart_id_i_20_));
 sg13g2_antennanp ANTENNA_1886 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1887 (.A(hart_id_i_21_));
 sg13g2_antennanp ANTENNA_1888 (.A(hart_id_i_22_));
 sg13g2_antennanp ANTENNA_1889 (.A(hart_id_i_23_));
 sg13g2_antennanp ANTENNA_1890 (.A(hart_id_i_24_));
 sg13g2_antennanp ANTENNA_1891 (.A(hart_id_i_25_));
 sg13g2_antennanp ANTENNA_1892 (.A(hart_id_i_27_));
 sg13g2_antennanp ANTENNA_1893 (.A(hart_id_i_28_));
 sg13g2_antennanp ANTENNA_1894 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1895 (.A(hart_id_i_29_));
 sg13g2_antennanp ANTENNA_1896 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1897 (.A(hart_id_i_2_));
 sg13g2_antennanp ANTENNA_1898 (.A(hart_id_i_31_));
 sg13g2_antennanp ANTENNA_1899 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1900 (.A(hart_id_i_3_));
 sg13g2_antennanp ANTENNA_1901 (.A(hart_id_i_4_));
 sg13g2_antennanp ANTENNA_1902 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_1903 (.A(hart_id_i_7_));
 sg13g2_antennanp ANTENNA_1904 (.A(hart_id_i_9_));
 sg13g2_antennanp ANTENNA_1905 (.A(instr_rvalid_i));
 sg13g2_antennanp ANTENNA_1906 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1907 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1908 (.A(irq_external_i));
 sg13g2_antennanp ANTENNA_1909 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1910 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1911 (.A(irq_fast_i_0_));
 sg13g2_antennanp ANTENNA_1912 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1913 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1914 (.A(irq_fast_i_11_));
 sg13g2_antennanp ANTENNA_1915 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1916 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1917 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1918 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1919 (.A(irq_fast_i_13_));
 sg13g2_antennanp ANTENNA_1920 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1921 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1922 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1923 (.A(irq_fast_i_15_));
 sg13g2_antennanp ANTENNA_1924 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1925 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1926 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1927 (.A(irq_fast_i_1_));
 sg13g2_antennanp ANTENNA_1928 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1929 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1930 (.A(irq_fast_i_2_));
 sg13g2_antennanp ANTENNA_1931 (.A(irq_fast_i_5_));
 sg13g2_antennanp ANTENNA_1932 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1933 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1934 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1935 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1936 (.A(irq_fast_i_6_));
 sg13g2_antennanp ANTENNA_1937 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1938 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1939 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1940 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1941 (.A(irq_fast_i_7_));
 sg13g2_antennanp ANTENNA_1942 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1943 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1944 (.A(irq_fast_i_8_));
 sg13g2_antennanp ANTENNA_1945 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1946 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1947 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1948 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1949 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1950 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1951 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1952 (.A(irq_fast_i_9_));
 sg13g2_antennanp ANTENNA_1953 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1954 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1955 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1956 (.A(irq_nm_i));
 sg13g2_antennanp ANTENNA_1957 (.A(irq_software_i));
 sg13g2_antennanp ANTENNA_1958 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1959 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1960 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1961 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1962 (.A(irq_timer_i));
 sg13g2_antennanp ANTENNA_1963 (.A(rf_wdata_wb_23_));
 sg13g2_antennanp ANTENNA_1964 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1965 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1966 (.A(rf_wdata_wb_27_));
 sg13g2_antennanp ANTENNA_1967 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1968 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1969 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1970 (.A(rf_wdata_wb_29_));
 sg13g2_antennanp ANTENNA_1971 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_1972 (.A(\cs_registers_i/_0702_ ));
 sg13g2_antennanp ANTENNA_1973 (.A(net1516));
 sg13g2_antennanp ANTENNA_1974 (.A(net1516));
 sg13g2_antennanp ANTENNA_1975 (.A(net1516));
 sg13g2_antennanp ANTENNA_1976 (.A(net1516));
 sg13g2_antennanp ANTENNA_1977 (.A(net1516));
 sg13g2_antennanp ANTENNA_1978 (.A(net2465));
 sg13g2_antennanp ANTENNA_1979 (.A(net2465));
 sg13g2_antennanp ANTENNA_1980 (.A(net2465));
 sg13g2_antennanp ANTENNA_1981 (.A(net2465));
 sg13g2_antennanp ANTENNA_1982 (.A(net2465));
 sg13g2_antennanp ANTENNA_1983 (.A(net2465));
 sg13g2_fill_8 FILLER_0_0 ();
 sg13g2_fill_8 FILLER_0_8 ();
 sg13g2_fill_8 FILLER_0_16 ();
 sg13g2_fill_8 FILLER_0_24 ();
 sg13g2_fill_8 FILLER_0_32 ();
 sg13g2_fill_8 FILLER_0_40 ();
 sg13g2_fill_8 FILLER_0_48 ();
 sg13g2_fill_8 FILLER_0_56 ();
 sg13g2_fill_8 FILLER_0_64 ();
 sg13g2_fill_8 FILLER_0_72 ();
 sg13g2_fill_8 FILLER_0_80 ();
 sg13g2_fill_8 FILLER_0_88 ();
 sg13g2_fill_8 FILLER_0_96 ();
 sg13g2_fill_8 FILLER_0_104 ();
 sg13g2_fill_8 FILLER_0_112 ();
 sg13g2_fill_8 FILLER_0_120 ();
 sg13g2_fill_8 FILLER_0_128 ();
 sg13g2_fill_8 FILLER_0_136 ();
 sg13g2_fill_8 FILLER_0_144 ();
 sg13g2_fill_8 FILLER_0_152 ();
 sg13g2_fill_8 FILLER_0_160 ();
 sg13g2_fill_8 FILLER_0_168 ();
 sg13g2_fill_8 FILLER_0_176 ();
 sg13g2_fill_8 FILLER_0_184 ();
 sg13g2_fill_8 FILLER_0_192 ();
 sg13g2_fill_8 FILLER_0_200 ();
 sg13g2_fill_8 FILLER_0_208 ();
 sg13g2_fill_8 FILLER_0_216 ();
 sg13g2_fill_8 FILLER_0_224 ();
 sg13g2_fill_8 FILLER_0_232 ();
 sg13g2_fill_8 FILLER_0_240 ();
 sg13g2_fill_8 FILLER_0_248 ();
 sg13g2_fill_8 FILLER_0_256 ();
 sg13g2_fill_8 FILLER_0_264 ();
 sg13g2_fill_8 FILLER_0_272 ();
 sg13g2_fill_8 FILLER_0_280 ();
 sg13g2_fill_8 FILLER_0_288 ();
 sg13g2_fill_8 FILLER_0_296 ();
 sg13g2_fill_8 FILLER_0_304 ();
 sg13g2_fill_8 FILLER_0_312 ();
 sg13g2_fill_8 FILLER_0_320 ();
 sg13g2_fill_8 FILLER_0_328 ();
 sg13g2_fill_8 FILLER_0_336 ();
 sg13g2_fill_8 FILLER_0_344 ();
 sg13g2_fill_8 FILLER_0_352 ();
 sg13g2_fill_8 FILLER_0_360 ();
 sg13g2_fill_8 FILLER_0_368 ();
 sg13g2_fill_8 FILLER_0_376 ();
 sg13g2_fill_8 FILLER_0_384 ();
 sg13g2_fill_8 FILLER_0_392 ();
 sg13g2_fill_8 FILLER_0_400 ();
 sg13g2_fill_8 FILLER_0_408 ();
 sg13g2_fill_8 FILLER_0_416 ();
 sg13g2_fill_8 FILLER_0_424 ();
 sg13g2_fill_8 FILLER_0_432 ();
 sg13g2_fill_8 FILLER_0_440 ();
 sg13g2_fill_8 FILLER_0_448 ();
 sg13g2_fill_8 FILLER_0_456 ();
 sg13g2_fill_8 FILLER_0_464 ();
 sg13g2_fill_8 FILLER_0_472 ();
 sg13g2_fill_8 FILLER_0_480 ();
 sg13g2_fill_8 FILLER_0_488 ();
 sg13g2_fill_8 FILLER_0_496 ();
 sg13g2_fill_8 FILLER_0_504 ();
 sg13g2_fill_8 FILLER_0_512 ();
 sg13g2_fill_8 FILLER_0_520 ();
 sg13g2_fill_8 FILLER_0_528 ();
 sg13g2_fill_8 FILLER_0_536 ();
 sg13g2_fill_8 FILLER_0_544 ();
 sg13g2_fill_8 FILLER_0_552 ();
 sg13g2_fill_8 FILLER_0_560 ();
 sg13g2_fill_8 FILLER_0_568 ();
 sg13g2_fill_8 FILLER_0_576 ();
 sg13g2_fill_8 FILLER_0_584 ();
 sg13g2_fill_8 FILLER_0_592 ();
 sg13g2_fill_8 FILLER_0_600 ();
 sg13g2_fill_8 FILLER_0_608 ();
 sg13g2_fill_8 FILLER_0_616 ();
 sg13g2_fill_8 FILLER_0_624 ();
 sg13g2_fill_8 FILLER_0_632 ();
 sg13g2_fill_8 FILLER_0_640 ();
 sg13g2_fill_8 FILLER_0_648 ();
 sg13g2_fill_8 FILLER_0_656 ();
 sg13g2_fill_8 FILLER_0_664 ();
 sg13g2_fill_8 FILLER_0_672 ();
 sg13g2_fill_8 FILLER_0_680 ();
 sg13g2_fill_8 FILLER_0_688 ();
 sg13g2_fill_8 FILLER_0_696 ();
 sg13g2_fill_8 FILLER_0_704 ();
 sg13g2_fill_8 FILLER_0_712 ();
 sg13g2_fill_8 FILLER_0_720 ();
 sg13g2_fill_8 FILLER_0_728 ();
 sg13g2_fill_8 FILLER_0_736 ();
 sg13g2_fill_8 FILLER_0_744 ();
 sg13g2_fill_8 FILLER_0_752 ();
 sg13g2_fill_8 FILLER_0_760 ();
 sg13g2_fill_8 FILLER_0_768 ();
 sg13g2_fill_8 FILLER_0_776 ();
 sg13g2_fill_8 FILLER_0_784 ();
 sg13g2_fill_8 FILLER_0_792 ();
 sg13g2_fill_8 FILLER_0_800 ();
 sg13g2_fill_8 FILLER_0_808 ();
 sg13g2_fill_2 FILLER_0_821 ();
 sg13g2_fill_1 FILLER_0_823 ();
 sg13g2_fill_8 FILLER_0_834 ();
 sg13g2_fill_8 FILLER_0_842 ();
 sg13g2_fill_8 FILLER_0_850 ();
 sg13g2_fill_8 FILLER_0_858 ();
 sg13g2_fill_8 FILLER_0_866 ();
 sg13g2_fill_8 FILLER_0_874 ();
 sg13g2_fill_8 FILLER_0_882 ();
 sg13g2_fill_8 FILLER_0_890 ();
 sg13g2_fill_8 FILLER_0_898 ();
 sg13g2_fill_8 FILLER_0_906 ();
 sg13g2_fill_8 FILLER_0_914 ();
 sg13g2_fill_8 FILLER_0_922 ();
 sg13g2_fill_8 FILLER_0_930 ();
 sg13g2_fill_8 FILLER_0_938 ();
 sg13g2_fill_8 FILLER_0_946 ();
 sg13g2_fill_8 FILLER_0_954 ();
 sg13g2_fill_8 FILLER_0_962 ();
 sg13g2_fill_8 FILLER_0_970 ();
 sg13g2_fill_8 FILLER_0_978 ();
 sg13g2_fill_8 FILLER_0_986 ();
 sg13g2_fill_8 FILLER_0_994 ();
 sg13g2_fill_8 FILLER_0_1002 ();
 sg13g2_fill_8 FILLER_0_1010 ();
 sg13g2_fill_8 FILLER_0_1018 ();
 sg13g2_fill_8 FILLER_0_1026 ();
 sg13g2_fill_8 FILLER_0_1034 ();
 sg13g2_fill_8 FILLER_0_1042 ();
 sg13g2_fill_8 FILLER_0_1050 ();
 sg13g2_fill_8 FILLER_0_1058 ();
 sg13g2_fill_8 FILLER_0_1066 ();
 sg13g2_fill_8 FILLER_0_1074 ();
 sg13g2_fill_8 FILLER_0_1082 ();
 sg13g2_fill_8 FILLER_0_1090 ();
 sg13g2_fill_8 FILLER_0_1098 ();
 sg13g2_fill_8 FILLER_0_1106 ();
 sg13g2_fill_8 FILLER_0_1114 ();
 sg13g2_fill_8 FILLER_0_1122 ();
 sg13g2_fill_8 FILLER_0_1130 ();
 sg13g2_fill_8 FILLER_0_1138 ();
 sg13g2_fill_8 FILLER_0_1146 ();
 sg13g2_fill_8 FILLER_0_1154 ();
 sg13g2_fill_8 FILLER_0_1162 ();
 sg13g2_fill_8 FILLER_0_1170 ();
 sg13g2_fill_8 FILLER_0_1178 ();
 sg13g2_fill_8 FILLER_0_1186 ();
 sg13g2_fill_8 FILLER_0_1194 ();
 sg13g2_fill_8 FILLER_0_1202 ();
 sg13g2_fill_8 FILLER_0_1210 ();
 sg13g2_fill_8 FILLER_0_1218 ();
 sg13g2_fill_8 FILLER_0_1226 ();
 sg13g2_fill_8 FILLER_0_1234 ();
 sg13g2_fill_8 FILLER_0_1242 ();
 sg13g2_fill_8 FILLER_0_1250 ();
 sg13g2_fill_8 FILLER_0_1258 ();
 sg13g2_fill_8 FILLER_0_1266 ();
 sg13g2_fill_8 FILLER_0_1274 ();
 sg13g2_fill_8 FILLER_0_1282 ();
 sg13g2_fill_8 FILLER_0_1290 ();
 sg13g2_fill_8 FILLER_0_1298 ();
 sg13g2_fill_8 FILLER_0_1306 ();
 sg13g2_fill_8 FILLER_0_1314 ();
 sg13g2_fill_8 FILLER_0_1322 ();
 sg13g2_fill_8 FILLER_0_1330 ();
 sg13g2_fill_8 FILLER_0_1338 ();
 sg13g2_fill_8 FILLER_0_1346 ();
 sg13g2_fill_8 FILLER_0_1354 ();
 sg13g2_fill_8 FILLER_0_1362 ();
 sg13g2_fill_8 FILLER_0_1370 ();
 sg13g2_fill_8 FILLER_0_1378 ();
 sg13g2_fill_8 FILLER_0_1386 ();
 sg13g2_fill_8 FILLER_0_1394 ();
 sg13g2_fill_8 FILLER_0_1402 ();
 sg13g2_fill_8 FILLER_0_1410 ();
 sg13g2_fill_8 FILLER_0_1418 ();
 sg13g2_fill_8 FILLER_0_1426 ();
 sg13g2_fill_8 FILLER_0_1434 ();
 sg13g2_fill_8 FILLER_0_1442 ();
 sg13g2_fill_8 FILLER_0_1450 ();
 sg13g2_fill_8 FILLER_0_1458 ();
 sg13g2_fill_8 FILLER_0_1466 ();
 sg13g2_fill_8 FILLER_0_1474 ();
 sg13g2_fill_8 FILLER_0_1482 ();
 sg13g2_fill_8 FILLER_0_1490 ();
 sg13g2_fill_8 FILLER_0_1498 ();
 sg13g2_fill_8 FILLER_0_1506 ();
 sg13g2_fill_8 FILLER_0_1514 ();
 sg13g2_fill_8 FILLER_0_1522 ();
 sg13g2_fill_8 FILLER_0_1530 ();
 sg13g2_fill_8 FILLER_0_1538 ();
 sg13g2_fill_8 FILLER_0_1546 ();
 sg13g2_fill_8 FILLER_0_1554 ();
 sg13g2_fill_8 FILLER_0_1562 ();
 sg13g2_fill_8 FILLER_0_1570 ();
 sg13g2_fill_2 FILLER_0_1578 ();
 sg13g2_fill_1 FILLER_0_1580 ();
 sg13g2_fill_4 FILLER_0_1585 ();
 sg13g2_fill_2 FILLER_0_1589 ();
 sg13g2_fill_1 FILLER_0_1591 ();
 sg13g2_fill_8 FILLER_1_0 ();
 sg13g2_fill_8 FILLER_1_8 ();
 sg13g2_fill_8 FILLER_1_16 ();
 sg13g2_fill_8 FILLER_1_24 ();
 sg13g2_fill_8 FILLER_1_32 ();
 sg13g2_fill_8 FILLER_1_40 ();
 sg13g2_fill_8 FILLER_1_48 ();
 sg13g2_fill_8 FILLER_1_56 ();
 sg13g2_fill_8 FILLER_1_64 ();
 sg13g2_fill_8 FILLER_1_72 ();
 sg13g2_fill_8 FILLER_1_80 ();
 sg13g2_fill_8 FILLER_1_88 ();
 sg13g2_fill_8 FILLER_1_96 ();
 sg13g2_fill_8 FILLER_1_104 ();
 sg13g2_fill_8 FILLER_1_112 ();
 sg13g2_fill_8 FILLER_1_120 ();
 sg13g2_fill_8 FILLER_1_128 ();
 sg13g2_fill_8 FILLER_1_136 ();
 sg13g2_fill_8 FILLER_1_144 ();
 sg13g2_fill_8 FILLER_1_152 ();
 sg13g2_fill_8 FILLER_1_160 ();
 sg13g2_fill_8 FILLER_1_168 ();
 sg13g2_fill_8 FILLER_1_176 ();
 sg13g2_fill_8 FILLER_1_184 ();
 sg13g2_fill_8 FILLER_1_192 ();
 sg13g2_fill_8 FILLER_1_200 ();
 sg13g2_fill_8 FILLER_1_208 ();
 sg13g2_fill_8 FILLER_1_216 ();
 sg13g2_fill_8 FILLER_1_224 ();
 sg13g2_fill_8 FILLER_1_232 ();
 sg13g2_fill_8 FILLER_1_240 ();
 sg13g2_fill_8 FILLER_1_248 ();
 sg13g2_fill_8 FILLER_1_256 ();
 sg13g2_fill_8 FILLER_1_264 ();
 sg13g2_fill_8 FILLER_1_272 ();
 sg13g2_fill_8 FILLER_1_280 ();
 sg13g2_fill_8 FILLER_1_288 ();
 sg13g2_fill_8 FILLER_1_296 ();
 sg13g2_fill_8 FILLER_1_304 ();
 sg13g2_fill_8 FILLER_1_312 ();
 sg13g2_fill_8 FILLER_1_320 ();
 sg13g2_fill_8 FILLER_1_328 ();
 sg13g2_fill_8 FILLER_1_336 ();
 sg13g2_fill_8 FILLER_1_344 ();
 sg13g2_fill_8 FILLER_1_352 ();
 sg13g2_fill_8 FILLER_1_360 ();
 sg13g2_fill_8 FILLER_1_368 ();
 sg13g2_fill_8 FILLER_1_376 ();
 sg13g2_fill_8 FILLER_1_384 ();
 sg13g2_fill_8 FILLER_1_392 ();
 sg13g2_fill_8 FILLER_1_400 ();
 sg13g2_fill_8 FILLER_1_408 ();
 sg13g2_fill_8 FILLER_1_416 ();
 sg13g2_fill_8 FILLER_1_424 ();
 sg13g2_fill_8 FILLER_1_432 ();
 sg13g2_fill_8 FILLER_1_440 ();
 sg13g2_fill_8 FILLER_1_448 ();
 sg13g2_fill_8 FILLER_1_456 ();
 sg13g2_fill_8 FILLER_1_464 ();
 sg13g2_fill_8 FILLER_1_472 ();
 sg13g2_fill_8 FILLER_1_480 ();
 sg13g2_fill_8 FILLER_1_488 ();
 sg13g2_fill_8 FILLER_1_496 ();
 sg13g2_fill_8 FILLER_1_504 ();
 sg13g2_fill_8 FILLER_1_512 ();
 sg13g2_fill_8 FILLER_1_520 ();
 sg13g2_fill_8 FILLER_1_528 ();
 sg13g2_fill_8 FILLER_1_536 ();
 sg13g2_fill_8 FILLER_1_544 ();
 sg13g2_fill_8 FILLER_1_552 ();
 sg13g2_fill_8 FILLER_1_560 ();
 sg13g2_fill_8 FILLER_1_568 ();
 sg13g2_fill_8 FILLER_1_576 ();
 sg13g2_fill_8 FILLER_1_584 ();
 sg13g2_fill_8 FILLER_1_592 ();
 sg13g2_fill_8 FILLER_1_600 ();
 sg13g2_fill_8 FILLER_1_608 ();
 sg13g2_fill_8 FILLER_1_616 ();
 sg13g2_fill_8 FILLER_1_624 ();
 sg13g2_fill_8 FILLER_1_632 ();
 sg13g2_fill_8 FILLER_1_640 ();
 sg13g2_fill_8 FILLER_1_648 ();
 sg13g2_fill_8 FILLER_1_656 ();
 sg13g2_fill_8 FILLER_1_664 ();
 sg13g2_fill_8 FILLER_1_672 ();
 sg13g2_fill_8 FILLER_1_680 ();
 sg13g2_fill_8 FILLER_1_688 ();
 sg13g2_fill_8 FILLER_1_696 ();
 sg13g2_fill_8 FILLER_1_704 ();
 sg13g2_fill_8 FILLER_1_712 ();
 sg13g2_fill_8 FILLER_1_720 ();
 sg13g2_fill_8 FILLER_1_728 ();
 sg13g2_fill_8 FILLER_1_736 ();
 sg13g2_fill_8 FILLER_1_744 ();
 sg13g2_fill_8 FILLER_1_752 ();
 sg13g2_fill_8 FILLER_1_760 ();
 sg13g2_fill_8 FILLER_1_768 ();
 sg13g2_fill_8 FILLER_1_776 ();
 sg13g2_fill_8 FILLER_1_784 ();
 sg13g2_fill_4 FILLER_1_792 ();
 sg13g2_fill_2 FILLER_1_796 ();
 sg13g2_fill_4 FILLER_1_824 ();
 sg13g2_fill_8 FILLER_1_854 ();
 sg13g2_fill_8 FILLER_1_862 ();
 sg13g2_fill_8 FILLER_1_870 ();
 sg13g2_fill_8 FILLER_1_878 ();
 sg13g2_fill_8 FILLER_1_886 ();
 sg13g2_fill_8 FILLER_1_894 ();
 sg13g2_fill_8 FILLER_1_902 ();
 sg13g2_fill_8 FILLER_1_910 ();
 sg13g2_fill_8 FILLER_1_918 ();
 sg13g2_fill_8 FILLER_1_926 ();
 sg13g2_fill_8 FILLER_1_934 ();
 sg13g2_fill_8 FILLER_1_942 ();
 sg13g2_fill_8 FILLER_1_950 ();
 sg13g2_fill_8 FILLER_1_958 ();
 sg13g2_fill_8 FILLER_1_966 ();
 sg13g2_fill_8 FILLER_1_974 ();
 sg13g2_fill_8 FILLER_1_982 ();
 sg13g2_fill_8 FILLER_1_990 ();
 sg13g2_fill_8 FILLER_1_998 ();
 sg13g2_fill_8 FILLER_1_1006 ();
 sg13g2_fill_8 FILLER_1_1014 ();
 sg13g2_fill_8 FILLER_1_1022 ();
 sg13g2_fill_8 FILLER_1_1030 ();
 sg13g2_fill_8 FILLER_1_1038 ();
 sg13g2_fill_8 FILLER_1_1046 ();
 sg13g2_fill_8 FILLER_1_1054 ();
 sg13g2_fill_8 FILLER_1_1062 ();
 sg13g2_fill_8 FILLER_1_1070 ();
 sg13g2_fill_8 FILLER_1_1078 ();
 sg13g2_fill_8 FILLER_1_1086 ();
 sg13g2_fill_8 FILLER_1_1094 ();
 sg13g2_fill_8 FILLER_1_1102 ();
 sg13g2_fill_8 FILLER_1_1110 ();
 sg13g2_fill_8 FILLER_1_1118 ();
 sg13g2_fill_8 FILLER_1_1126 ();
 sg13g2_fill_8 FILLER_1_1134 ();
 sg13g2_fill_8 FILLER_1_1142 ();
 sg13g2_fill_8 FILLER_1_1150 ();
 sg13g2_fill_8 FILLER_1_1158 ();
 sg13g2_fill_8 FILLER_1_1166 ();
 sg13g2_fill_8 FILLER_1_1174 ();
 sg13g2_fill_8 FILLER_1_1182 ();
 sg13g2_fill_8 FILLER_1_1190 ();
 sg13g2_fill_8 FILLER_1_1198 ();
 sg13g2_fill_8 FILLER_1_1206 ();
 sg13g2_fill_8 FILLER_1_1214 ();
 sg13g2_fill_8 FILLER_1_1222 ();
 sg13g2_fill_8 FILLER_1_1230 ();
 sg13g2_fill_8 FILLER_1_1238 ();
 sg13g2_fill_8 FILLER_1_1246 ();
 sg13g2_fill_8 FILLER_1_1254 ();
 sg13g2_fill_8 FILLER_1_1262 ();
 sg13g2_fill_8 FILLER_1_1270 ();
 sg13g2_fill_8 FILLER_1_1278 ();
 sg13g2_fill_8 FILLER_1_1286 ();
 sg13g2_fill_8 FILLER_1_1294 ();
 sg13g2_fill_8 FILLER_1_1302 ();
 sg13g2_fill_8 FILLER_1_1310 ();
 sg13g2_fill_8 FILLER_1_1318 ();
 sg13g2_fill_8 FILLER_1_1326 ();
 sg13g2_fill_8 FILLER_1_1334 ();
 sg13g2_fill_8 FILLER_1_1342 ();
 sg13g2_fill_8 FILLER_1_1350 ();
 sg13g2_fill_8 FILLER_1_1358 ();
 sg13g2_fill_8 FILLER_1_1366 ();
 sg13g2_fill_8 FILLER_1_1374 ();
 sg13g2_fill_8 FILLER_1_1382 ();
 sg13g2_fill_8 FILLER_1_1390 ();
 sg13g2_fill_8 FILLER_1_1398 ();
 sg13g2_fill_8 FILLER_1_1406 ();
 sg13g2_fill_8 FILLER_1_1414 ();
 sg13g2_fill_8 FILLER_1_1422 ();
 sg13g2_fill_8 FILLER_1_1430 ();
 sg13g2_fill_8 FILLER_1_1438 ();
 sg13g2_fill_8 FILLER_1_1446 ();
 sg13g2_fill_8 FILLER_1_1454 ();
 sg13g2_fill_8 FILLER_1_1462 ();
 sg13g2_fill_8 FILLER_1_1470 ();
 sg13g2_fill_8 FILLER_1_1478 ();
 sg13g2_fill_8 FILLER_1_1486 ();
 sg13g2_fill_8 FILLER_1_1494 ();
 sg13g2_fill_8 FILLER_1_1502 ();
 sg13g2_fill_8 FILLER_1_1510 ();
 sg13g2_fill_8 FILLER_1_1518 ();
 sg13g2_fill_8 FILLER_1_1526 ();
 sg13g2_fill_8 FILLER_1_1534 ();
 sg13g2_fill_8 FILLER_1_1542 ();
 sg13g2_fill_8 FILLER_1_1550 ();
 sg13g2_fill_8 FILLER_1_1558 ();
 sg13g2_fill_8 FILLER_1_1566 ();
 sg13g2_fill_2 FILLER_1_1574 ();
 sg13g2_fill_1 FILLER_1_1576 ();
 sg13g2_fill_2 FILLER_1_1589 ();
 sg13g2_fill_1 FILLER_1_1591 ();
 sg13g2_fill_8 FILLER_2_0 ();
 sg13g2_fill_8 FILLER_2_8 ();
 sg13g2_fill_8 FILLER_2_16 ();
 sg13g2_fill_8 FILLER_2_24 ();
 sg13g2_fill_8 FILLER_2_32 ();
 sg13g2_fill_8 FILLER_2_40 ();
 sg13g2_fill_8 FILLER_2_48 ();
 sg13g2_fill_8 FILLER_2_56 ();
 sg13g2_fill_8 FILLER_2_64 ();
 sg13g2_fill_8 FILLER_2_72 ();
 sg13g2_fill_8 FILLER_2_80 ();
 sg13g2_fill_8 FILLER_2_88 ();
 sg13g2_fill_8 FILLER_2_96 ();
 sg13g2_fill_8 FILLER_2_104 ();
 sg13g2_fill_8 FILLER_2_112 ();
 sg13g2_fill_8 FILLER_2_120 ();
 sg13g2_fill_8 FILLER_2_128 ();
 sg13g2_fill_8 FILLER_2_136 ();
 sg13g2_fill_8 FILLER_2_144 ();
 sg13g2_fill_8 FILLER_2_152 ();
 sg13g2_fill_8 FILLER_2_160 ();
 sg13g2_fill_8 FILLER_2_168 ();
 sg13g2_fill_8 FILLER_2_176 ();
 sg13g2_fill_8 FILLER_2_184 ();
 sg13g2_fill_8 FILLER_2_192 ();
 sg13g2_fill_8 FILLER_2_200 ();
 sg13g2_fill_8 FILLER_2_208 ();
 sg13g2_fill_8 FILLER_2_216 ();
 sg13g2_fill_8 FILLER_2_224 ();
 sg13g2_fill_8 FILLER_2_232 ();
 sg13g2_fill_8 FILLER_2_240 ();
 sg13g2_fill_8 FILLER_2_248 ();
 sg13g2_fill_8 FILLER_2_256 ();
 sg13g2_fill_8 FILLER_2_264 ();
 sg13g2_fill_8 FILLER_2_272 ();
 sg13g2_fill_8 FILLER_2_280 ();
 sg13g2_fill_8 FILLER_2_288 ();
 sg13g2_fill_8 FILLER_2_296 ();
 sg13g2_fill_8 FILLER_2_304 ();
 sg13g2_fill_8 FILLER_2_312 ();
 sg13g2_fill_8 FILLER_2_320 ();
 sg13g2_fill_8 FILLER_2_328 ();
 sg13g2_fill_8 FILLER_2_336 ();
 sg13g2_fill_8 FILLER_2_344 ();
 sg13g2_fill_8 FILLER_2_352 ();
 sg13g2_fill_8 FILLER_2_360 ();
 sg13g2_fill_8 FILLER_2_368 ();
 sg13g2_fill_8 FILLER_2_376 ();
 sg13g2_fill_8 FILLER_2_384 ();
 sg13g2_fill_8 FILLER_2_392 ();
 sg13g2_fill_8 FILLER_2_400 ();
 sg13g2_fill_8 FILLER_2_408 ();
 sg13g2_fill_8 FILLER_2_416 ();
 sg13g2_fill_8 FILLER_2_424 ();
 sg13g2_fill_8 FILLER_2_432 ();
 sg13g2_fill_8 FILLER_2_440 ();
 sg13g2_fill_8 FILLER_2_448 ();
 sg13g2_fill_8 FILLER_2_456 ();
 sg13g2_fill_8 FILLER_2_464 ();
 sg13g2_fill_8 FILLER_2_472 ();
 sg13g2_fill_8 FILLER_2_480 ();
 sg13g2_fill_8 FILLER_2_488 ();
 sg13g2_fill_8 FILLER_2_496 ();
 sg13g2_fill_8 FILLER_2_504 ();
 sg13g2_fill_8 FILLER_2_512 ();
 sg13g2_fill_8 FILLER_2_520 ();
 sg13g2_fill_8 FILLER_2_528 ();
 sg13g2_fill_8 FILLER_2_536 ();
 sg13g2_fill_8 FILLER_2_544 ();
 sg13g2_fill_8 FILLER_2_552 ();
 sg13g2_fill_8 FILLER_2_560 ();
 sg13g2_fill_8 FILLER_2_568 ();
 sg13g2_fill_8 FILLER_2_576 ();
 sg13g2_fill_8 FILLER_2_584 ();
 sg13g2_fill_8 FILLER_2_592 ();
 sg13g2_fill_8 FILLER_2_600 ();
 sg13g2_fill_8 FILLER_2_608 ();
 sg13g2_fill_8 FILLER_2_616 ();
 sg13g2_fill_8 FILLER_2_624 ();
 sg13g2_fill_8 FILLER_2_632 ();
 sg13g2_fill_8 FILLER_2_640 ();
 sg13g2_fill_8 FILLER_2_648 ();
 sg13g2_fill_8 FILLER_2_656 ();
 sg13g2_fill_8 FILLER_2_664 ();
 sg13g2_fill_8 FILLER_2_672 ();
 sg13g2_fill_8 FILLER_2_680 ();
 sg13g2_fill_8 FILLER_2_688 ();
 sg13g2_fill_8 FILLER_2_696 ();
 sg13g2_fill_8 FILLER_2_704 ();
 sg13g2_fill_8 FILLER_2_712 ();
 sg13g2_fill_8 FILLER_2_720 ();
 sg13g2_fill_8 FILLER_2_728 ();
 sg13g2_fill_8 FILLER_2_736 ();
 sg13g2_fill_8 FILLER_2_744 ();
 sg13g2_fill_8 FILLER_2_752 ();
 sg13g2_fill_8 FILLER_2_760 ();
 sg13g2_fill_8 FILLER_2_768 ();
 sg13g2_fill_8 FILLER_2_776 ();
 sg13g2_fill_8 FILLER_2_784 ();
 sg13g2_fill_8 FILLER_2_792 ();
 sg13g2_fill_1 FILLER_2_800 ();
 sg13g2_fill_8 FILLER_2_827 ();
 sg13g2_fill_2 FILLER_2_835 ();
 sg13g2_fill_1 FILLER_2_837 ();
 sg13g2_fill_8 FILLER_2_869 ();
 sg13g2_fill_2 FILLER_2_877 ();
 sg13g2_fill_1 FILLER_2_879 ();
 sg13g2_fill_8 FILLER_2_890 ();
 sg13g2_fill_4 FILLER_2_898 ();
 sg13g2_fill_1 FILLER_2_902 ();
 sg13g2_fill_8 FILLER_2_908 ();
 sg13g2_fill_8 FILLER_2_916 ();
 sg13g2_fill_8 FILLER_2_924 ();
 sg13g2_fill_8 FILLER_2_932 ();
 sg13g2_fill_8 FILLER_2_940 ();
 sg13g2_fill_8 FILLER_2_948 ();
 sg13g2_fill_8 FILLER_2_956 ();
 sg13g2_fill_8 FILLER_2_964 ();
 sg13g2_fill_8 FILLER_2_972 ();
 sg13g2_fill_8 FILLER_2_980 ();
 sg13g2_fill_8 FILLER_2_988 ();
 sg13g2_fill_8 FILLER_2_996 ();
 sg13g2_fill_8 FILLER_2_1004 ();
 sg13g2_fill_8 FILLER_2_1012 ();
 sg13g2_fill_8 FILLER_2_1020 ();
 sg13g2_fill_8 FILLER_2_1028 ();
 sg13g2_fill_8 FILLER_2_1036 ();
 sg13g2_fill_8 FILLER_2_1044 ();
 sg13g2_fill_8 FILLER_2_1052 ();
 sg13g2_fill_8 FILLER_2_1060 ();
 sg13g2_fill_8 FILLER_2_1068 ();
 sg13g2_fill_8 FILLER_2_1076 ();
 sg13g2_fill_8 FILLER_2_1084 ();
 sg13g2_fill_8 FILLER_2_1092 ();
 sg13g2_fill_8 FILLER_2_1100 ();
 sg13g2_fill_8 FILLER_2_1108 ();
 sg13g2_fill_8 FILLER_2_1116 ();
 sg13g2_fill_8 FILLER_2_1124 ();
 sg13g2_fill_8 FILLER_2_1132 ();
 sg13g2_fill_8 FILLER_2_1140 ();
 sg13g2_fill_8 FILLER_2_1148 ();
 sg13g2_fill_8 FILLER_2_1156 ();
 sg13g2_fill_8 FILLER_2_1164 ();
 sg13g2_fill_8 FILLER_2_1172 ();
 sg13g2_fill_8 FILLER_2_1180 ();
 sg13g2_fill_8 FILLER_2_1188 ();
 sg13g2_fill_8 FILLER_2_1196 ();
 sg13g2_fill_8 FILLER_2_1204 ();
 sg13g2_fill_8 FILLER_2_1212 ();
 sg13g2_fill_8 FILLER_2_1220 ();
 sg13g2_fill_8 FILLER_2_1228 ();
 sg13g2_fill_8 FILLER_2_1236 ();
 sg13g2_fill_8 FILLER_2_1244 ();
 sg13g2_fill_8 FILLER_2_1252 ();
 sg13g2_fill_8 FILLER_2_1260 ();
 sg13g2_fill_8 FILLER_2_1268 ();
 sg13g2_fill_8 FILLER_2_1276 ();
 sg13g2_fill_8 FILLER_2_1284 ();
 sg13g2_fill_8 FILLER_2_1292 ();
 sg13g2_fill_8 FILLER_2_1300 ();
 sg13g2_fill_8 FILLER_2_1308 ();
 sg13g2_fill_8 FILLER_2_1316 ();
 sg13g2_fill_8 FILLER_2_1324 ();
 sg13g2_fill_8 FILLER_2_1332 ();
 sg13g2_fill_8 FILLER_2_1340 ();
 sg13g2_fill_8 FILLER_2_1348 ();
 sg13g2_fill_8 FILLER_2_1356 ();
 sg13g2_fill_8 FILLER_2_1364 ();
 sg13g2_fill_8 FILLER_2_1372 ();
 sg13g2_fill_8 FILLER_2_1380 ();
 sg13g2_fill_8 FILLER_2_1388 ();
 sg13g2_fill_8 FILLER_2_1396 ();
 sg13g2_fill_8 FILLER_2_1404 ();
 sg13g2_fill_8 FILLER_2_1412 ();
 sg13g2_fill_8 FILLER_2_1420 ();
 sg13g2_fill_8 FILLER_2_1428 ();
 sg13g2_fill_8 FILLER_2_1436 ();
 sg13g2_fill_8 FILLER_2_1444 ();
 sg13g2_fill_8 FILLER_2_1452 ();
 sg13g2_fill_8 FILLER_2_1460 ();
 sg13g2_fill_8 FILLER_2_1468 ();
 sg13g2_fill_8 FILLER_2_1476 ();
 sg13g2_fill_8 FILLER_2_1484 ();
 sg13g2_fill_8 FILLER_2_1492 ();
 sg13g2_fill_8 FILLER_2_1500 ();
 sg13g2_fill_8 FILLER_2_1508 ();
 sg13g2_fill_8 FILLER_2_1516 ();
 sg13g2_fill_8 FILLER_2_1524 ();
 sg13g2_fill_8 FILLER_2_1532 ();
 sg13g2_fill_8 FILLER_2_1540 ();
 sg13g2_fill_8 FILLER_2_1548 ();
 sg13g2_fill_8 FILLER_2_1556 ();
 sg13g2_fill_8 FILLER_2_1564 ();
 sg13g2_fill_8 FILLER_2_1572 ();
 sg13g2_fill_1 FILLER_2_1580 ();
 sg13g2_fill_4 FILLER_2_1585 ();
 sg13g2_fill_2 FILLER_2_1589 ();
 sg13g2_fill_1 FILLER_2_1591 ();
 sg13g2_fill_8 FILLER_3_0 ();
 sg13g2_fill_8 FILLER_3_8 ();
 sg13g2_fill_8 FILLER_3_16 ();
 sg13g2_fill_8 FILLER_3_24 ();
 sg13g2_fill_8 FILLER_3_32 ();
 sg13g2_fill_8 FILLER_3_40 ();
 sg13g2_fill_8 FILLER_3_48 ();
 sg13g2_fill_8 FILLER_3_56 ();
 sg13g2_fill_8 FILLER_3_64 ();
 sg13g2_fill_8 FILLER_3_72 ();
 sg13g2_fill_8 FILLER_3_80 ();
 sg13g2_fill_8 FILLER_3_88 ();
 sg13g2_fill_8 FILLER_3_96 ();
 sg13g2_fill_8 FILLER_3_104 ();
 sg13g2_fill_8 FILLER_3_112 ();
 sg13g2_fill_8 FILLER_3_120 ();
 sg13g2_fill_8 FILLER_3_128 ();
 sg13g2_fill_8 FILLER_3_136 ();
 sg13g2_fill_8 FILLER_3_144 ();
 sg13g2_fill_8 FILLER_3_152 ();
 sg13g2_fill_8 FILLER_3_160 ();
 sg13g2_fill_8 FILLER_3_168 ();
 sg13g2_fill_8 FILLER_3_176 ();
 sg13g2_fill_8 FILLER_3_184 ();
 sg13g2_fill_8 FILLER_3_192 ();
 sg13g2_fill_8 FILLER_3_200 ();
 sg13g2_fill_8 FILLER_3_208 ();
 sg13g2_fill_8 FILLER_3_216 ();
 sg13g2_fill_8 FILLER_3_224 ();
 sg13g2_fill_8 FILLER_3_232 ();
 sg13g2_fill_8 FILLER_3_240 ();
 sg13g2_fill_8 FILLER_3_248 ();
 sg13g2_fill_8 FILLER_3_256 ();
 sg13g2_fill_8 FILLER_3_264 ();
 sg13g2_fill_8 FILLER_3_272 ();
 sg13g2_fill_8 FILLER_3_280 ();
 sg13g2_fill_8 FILLER_3_288 ();
 sg13g2_fill_8 FILLER_3_296 ();
 sg13g2_fill_8 FILLER_3_304 ();
 sg13g2_fill_8 FILLER_3_312 ();
 sg13g2_fill_8 FILLER_3_320 ();
 sg13g2_fill_8 FILLER_3_328 ();
 sg13g2_fill_8 FILLER_3_336 ();
 sg13g2_fill_8 FILLER_3_344 ();
 sg13g2_fill_8 FILLER_3_352 ();
 sg13g2_fill_8 FILLER_3_360 ();
 sg13g2_fill_8 FILLER_3_368 ();
 sg13g2_fill_8 FILLER_3_376 ();
 sg13g2_fill_8 FILLER_3_384 ();
 sg13g2_fill_8 FILLER_3_392 ();
 sg13g2_fill_8 FILLER_3_400 ();
 sg13g2_fill_8 FILLER_3_408 ();
 sg13g2_fill_8 FILLER_3_416 ();
 sg13g2_fill_8 FILLER_3_424 ();
 sg13g2_fill_8 FILLER_3_432 ();
 sg13g2_fill_8 FILLER_3_440 ();
 sg13g2_fill_8 FILLER_3_448 ();
 sg13g2_fill_8 FILLER_3_456 ();
 sg13g2_fill_8 FILLER_3_464 ();
 sg13g2_fill_8 FILLER_3_472 ();
 sg13g2_fill_8 FILLER_3_480 ();
 sg13g2_fill_8 FILLER_3_488 ();
 sg13g2_fill_8 FILLER_3_496 ();
 sg13g2_fill_8 FILLER_3_504 ();
 sg13g2_fill_8 FILLER_3_512 ();
 sg13g2_fill_8 FILLER_3_520 ();
 sg13g2_fill_8 FILLER_3_528 ();
 sg13g2_fill_8 FILLER_3_536 ();
 sg13g2_fill_8 FILLER_3_544 ();
 sg13g2_fill_8 FILLER_3_552 ();
 sg13g2_fill_8 FILLER_3_560 ();
 sg13g2_fill_8 FILLER_3_568 ();
 sg13g2_fill_8 FILLER_3_576 ();
 sg13g2_fill_8 FILLER_3_584 ();
 sg13g2_fill_8 FILLER_3_592 ();
 sg13g2_fill_8 FILLER_3_600 ();
 sg13g2_fill_8 FILLER_3_608 ();
 sg13g2_fill_8 FILLER_3_616 ();
 sg13g2_fill_8 FILLER_3_624 ();
 sg13g2_fill_8 FILLER_3_632 ();
 sg13g2_fill_8 FILLER_3_640 ();
 sg13g2_fill_8 FILLER_3_648 ();
 sg13g2_fill_8 FILLER_3_656 ();
 sg13g2_fill_8 FILLER_3_664 ();
 sg13g2_fill_8 FILLER_3_672 ();
 sg13g2_fill_8 FILLER_3_680 ();
 sg13g2_fill_8 FILLER_3_688 ();
 sg13g2_fill_8 FILLER_3_696 ();
 sg13g2_fill_8 FILLER_3_704 ();
 sg13g2_fill_8 FILLER_3_712 ();
 sg13g2_fill_8 FILLER_3_720 ();
 sg13g2_fill_8 FILLER_3_728 ();
 sg13g2_fill_8 FILLER_3_736 ();
 sg13g2_fill_8 FILLER_3_744 ();
 sg13g2_fill_8 FILLER_3_752 ();
 sg13g2_fill_8 FILLER_3_760 ();
 sg13g2_fill_8 FILLER_3_768 ();
 sg13g2_fill_8 FILLER_3_776 ();
 sg13g2_fill_2 FILLER_3_784 ();
 sg13g2_fill_8 FILLER_3_812 ();
 sg13g2_fill_1 FILLER_3_820 ();
 sg13g2_fill_2 FILLER_3_831 ();
 sg13g2_fill_4 FILLER_3_861 ();
 sg13g2_fill_2 FILLER_3_865 ();
 sg13g2_fill_2 FILLER_3_877 ();
 sg13g2_fill_8 FILLER_3_931 ();
 sg13g2_fill_8 FILLER_3_939 ();
 sg13g2_fill_8 FILLER_3_947 ();
 sg13g2_fill_8 FILLER_3_955 ();
 sg13g2_fill_8 FILLER_3_963 ();
 sg13g2_fill_8 FILLER_3_971 ();
 sg13g2_fill_8 FILLER_3_979 ();
 sg13g2_fill_8 FILLER_3_987 ();
 sg13g2_fill_8 FILLER_3_995 ();
 sg13g2_fill_8 FILLER_3_1003 ();
 sg13g2_fill_8 FILLER_3_1011 ();
 sg13g2_fill_8 FILLER_3_1019 ();
 sg13g2_fill_8 FILLER_3_1027 ();
 sg13g2_fill_8 FILLER_3_1035 ();
 sg13g2_fill_8 FILLER_3_1043 ();
 sg13g2_fill_8 FILLER_3_1051 ();
 sg13g2_fill_8 FILLER_3_1059 ();
 sg13g2_fill_8 FILLER_3_1067 ();
 sg13g2_fill_8 FILLER_3_1075 ();
 sg13g2_fill_8 FILLER_3_1083 ();
 sg13g2_fill_8 FILLER_3_1091 ();
 sg13g2_fill_8 FILLER_3_1099 ();
 sg13g2_fill_8 FILLER_3_1107 ();
 sg13g2_fill_8 FILLER_3_1115 ();
 sg13g2_fill_8 FILLER_3_1123 ();
 sg13g2_fill_8 FILLER_3_1131 ();
 sg13g2_fill_8 FILLER_3_1139 ();
 sg13g2_fill_8 FILLER_3_1147 ();
 sg13g2_fill_8 FILLER_3_1155 ();
 sg13g2_fill_8 FILLER_3_1163 ();
 sg13g2_fill_8 FILLER_3_1171 ();
 sg13g2_fill_8 FILLER_3_1179 ();
 sg13g2_fill_8 FILLER_3_1187 ();
 sg13g2_fill_8 FILLER_3_1195 ();
 sg13g2_fill_8 FILLER_3_1203 ();
 sg13g2_fill_8 FILLER_3_1211 ();
 sg13g2_fill_8 FILLER_3_1219 ();
 sg13g2_fill_8 FILLER_3_1227 ();
 sg13g2_fill_8 FILLER_3_1235 ();
 sg13g2_fill_8 FILLER_3_1243 ();
 sg13g2_fill_8 FILLER_3_1251 ();
 sg13g2_fill_8 FILLER_3_1259 ();
 sg13g2_fill_8 FILLER_3_1267 ();
 sg13g2_fill_8 FILLER_3_1275 ();
 sg13g2_fill_8 FILLER_3_1283 ();
 sg13g2_fill_8 FILLER_3_1291 ();
 sg13g2_fill_8 FILLER_3_1299 ();
 sg13g2_fill_8 FILLER_3_1307 ();
 sg13g2_fill_8 FILLER_3_1315 ();
 sg13g2_fill_8 FILLER_3_1323 ();
 sg13g2_fill_8 FILLER_3_1331 ();
 sg13g2_fill_8 FILLER_3_1339 ();
 sg13g2_fill_8 FILLER_3_1347 ();
 sg13g2_fill_8 FILLER_3_1355 ();
 sg13g2_fill_8 FILLER_3_1363 ();
 sg13g2_fill_8 FILLER_3_1371 ();
 sg13g2_fill_8 FILLER_3_1379 ();
 sg13g2_fill_8 FILLER_3_1387 ();
 sg13g2_fill_8 FILLER_3_1395 ();
 sg13g2_fill_8 FILLER_3_1403 ();
 sg13g2_fill_8 FILLER_3_1411 ();
 sg13g2_fill_8 FILLER_3_1419 ();
 sg13g2_fill_8 FILLER_3_1427 ();
 sg13g2_fill_8 FILLER_3_1435 ();
 sg13g2_fill_8 FILLER_3_1443 ();
 sg13g2_fill_8 FILLER_3_1451 ();
 sg13g2_fill_8 FILLER_3_1459 ();
 sg13g2_fill_8 FILLER_3_1467 ();
 sg13g2_fill_8 FILLER_3_1475 ();
 sg13g2_fill_8 FILLER_3_1483 ();
 sg13g2_fill_8 FILLER_3_1491 ();
 sg13g2_fill_8 FILLER_3_1499 ();
 sg13g2_fill_8 FILLER_3_1507 ();
 sg13g2_fill_8 FILLER_3_1515 ();
 sg13g2_fill_8 FILLER_3_1523 ();
 sg13g2_fill_8 FILLER_3_1531 ();
 sg13g2_fill_8 FILLER_3_1539 ();
 sg13g2_fill_8 FILLER_3_1547 ();
 sg13g2_fill_8 FILLER_3_1555 ();
 sg13g2_fill_8 FILLER_3_1563 ();
 sg13g2_fill_8 FILLER_3_1571 ();
 sg13g2_fill_8 FILLER_3_1579 ();
 sg13g2_fill_4 FILLER_3_1587 ();
 sg13g2_fill_1 FILLER_3_1591 ();
 sg13g2_fill_8 FILLER_4_0 ();
 sg13g2_fill_8 FILLER_4_8 ();
 sg13g2_fill_8 FILLER_4_16 ();
 sg13g2_fill_8 FILLER_4_24 ();
 sg13g2_fill_8 FILLER_4_32 ();
 sg13g2_fill_8 FILLER_4_40 ();
 sg13g2_fill_8 FILLER_4_48 ();
 sg13g2_fill_8 FILLER_4_56 ();
 sg13g2_fill_8 FILLER_4_64 ();
 sg13g2_fill_8 FILLER_4_72 ();
 sg13g2_fill_8 FILLER_4_80 ();
 sg13g2_fill_8 FILLER_4_88 ();
 sg13g2_fill_8 FILLER_4_96 ();
 sg13g2_fill_8 FILLER_4_104 ();
 sg13g2_fill_8 FILLER_4_112 ();
 sg13g2_fill_8 FILLER_4_120 ();
 sg13g2_fill_8 FILLER_4_128 ();
 sg13g2_fill_8 FILLER_4_136 ();
 sg13g2_fill_8 FILLER_4_144 ();
 sg13g2_fill_8 FILLER_4_152 ();
 sg13g2_fill_8 FILLER_4_160 ();
 sg13g2_fill_8 FILLER_4_168 ();
 sg13g2_fill_8 FILLER_4_176 ();
 sg13g2_fill_8 FILLER_4_184 ();
 sg13g2_fill_8 FILLER_4_192 ();
 sg13g2_fill_8 FILLER_4_200 ();
 sg13g2_fill_8 FILLER_4_208 ();
 sg13g2_fill_8 FILLER_4_216 ();
 sg13g2_fill_8 FILLER_4_224 ();
 sg13g2_fill_8 FILLER_4_232 ();
 sg13g2_fill_8 FILLER_4_240 ();
 sg13g2_fill_8 FILLER_4_248 ();
 sg13g2_fill_8 FILLER_4_256 ();
 sg13g2_fill_8 FILLER_4_264 ();
 sg13g2_fill_8 FILLER_4_272 ();
 sg13g2_fill_8 FILLER_4_280 ();
 sg13g2_fill_8 FILLER_4_288 ();
 sg13g2_fill_8 FILLER_4_296 ();
 sg13g2_fill_8 FILLER_4_304 ();
 sg13g2_fill_8 FILLER_4_312 ();
 sg13g2_fill_8 FILLER_4_320 ();
 sg13g2_fill_8 FILLER_4_328 ();
 sg13g2_fill_8 FILLER_4_336 ();
 sg13g2_fill_8 FILLER_4_344 ();
 sg13g2_fill_8 FILLER_4_352 ();
 sg13g2_fill_8 FILLER_4_360 ();
 sg13g2_fill_8 FILLER_4_368 ();
 sg13g2_fill_8 FILLER_4_376 ();
 sg13g2_fill_8 FILLER_4_384 ();
 sg13g2_fill_8 FILLER_4_392 ();
 sg13g2_fill_8 FILLER_4_400 ();
 sg13g2_fill_8 FILLER_4_408 ();
 sg13g2_fill_8 FILLER_4_416 ();
 sg13g2_fill_8 FILLER_4_424 ();
 sg13g2_fill_8 FILLER_4_432 ();
 sg13g2_fill_8 FILLER_4_440 ();
 sg13g2_fill_8 FILLER_4_448 ();
 sg13g2_fill_8 FILLER_4_456 ();
 sg13g2_fill_8 FILLER_4_464 ();
 sg13g2_fill_8 FILLER_4_472 ();
 sg13g2_fill_8 FILLER_4_480 ();
 sg13g2_fill_8 FILLER_4_488 ();
 sg13g2_fill_8 FILLER_4_496 ();
 sg13g2_fill_8 FILLER_4_504 ();
 sg13g2_fill_8 FILLER_4_512 ();
 sg13g2_fill_8 FILLER_4_520 ();
 sg13g2_fill_8 FILLER_4_528 ();
 sg13g2_fill_8 FILLER_4_536 ();
 sg13g2_fill_8 FILLER_4_544 ();
 sg13g2_fill_8 FILLER_4_552 ();
 sg13g2_fill_8 FILLER_4_560 ();
 sg13g2_fill_8 FILLER_4_568 ();
 sg13g2_fill_8 FILLER_4_576 ();
 sg13g2_fill_8 FILLER_4_584 ();
 sg13g2_fill_8 FILLER_4_592 ();
 sg13g2_fill_8 FILLER_4_600 ();
 sg13g2_fill_8 FILLER_4_608 ();
 sg13g2_fill_8 FILLER_4_616 ();
 sg13g2_fill_8 FILLER_4_624 ();
 sg13g2_fill_8 FILLER_4_632 ();
 sg13g2_fill_8 FILLER_4_640 ();
 sg13g2_fill_8 FILLER_4_648 ();
 sg13g2_fill_8 FILLER_4_656 ();
 sg13g2_fill_8 FILLER_4_664 ();
 sg13g2_fill_8 FILLER_4_672 ();
 sg13g2_fill_8 FILLER_4_680 ();
 sg13g2_fill_8 FILLER_4_688 ();
 sg13g2_fill_8 FILLER_4_696 ();
 sg13g2_fill_8 FILLER_4_704 ();
 sg13g2_fill_8 FILLER_4_712 ();
 sg13g2_fill_8 FILLER_4_720 ();
 sg13g2_fill_8 FILLER_4_728 ();
 sg13g2_fill_8 FILLER_4_736 ();
 sg13g2_fill_8 FILLER_4_744 ();
 sg13g2_fill_8 FILLER_4_752 ();
 sg13g2_fill_8 FILLER_4_760 ();
 sg13g2_fill_8 FILLER_4_768 ();
 sg13g2_fill_4 FILLER_4_776 ();
 sg13g2_fill_1 FILLER_4_780 ();
 sg13g2_fill_8 FILLER_4_791 ();
 sg13g2_fill_8 FILLER_4_799 ();
 sg13g2_fill_8 FILLER_4_807 ();
 sg13g2_fill_8 FILLER_4_815 ();
 sg13g2_fill_8 FILLER_4_823 ();
 sg13g2_fill_8 FILLER_4_831 ();
 sg13g2_fill_4 FILLER_4_865 ();
 sg13g2_fill_8 FILLER_4_895 ();
 sg13g2_fill_8 FILLER_4_903 ();
 sg13g2_fill_8 FILLER_4_911 ();
 sg13g2_fill_8 FILLER_4_919 ();
 sg13g2_fill_8 FILLER_4_927 ();
 sg13g2_fill_8 FILLER_4_935 ();
 sg13g2_fill_8 FILLER_4_943 ();
 sg13g2_fill_8 FILLER_4_951 ();
 sg13g2_fill_8 FILLER_4_959 ();
 sg13g2_fill_8 FILLER_4_967 ();
 sg13g2_fill_8 FILLER_4_975 ();
 sg13g2_fill_8 FILLER_4_983 ();
 sg13g2_fill_8 FILLER_4_991 ();
 sg13g2_fill_8 FILLER_4_999 ();
 sg13g2_fill_8 FILLER_4_1007 ();
 sg13g2_fill_8 FILLER_4_1015 ();
 sg13g2_fill_8 FILLER_4_1023 ();
 sg13g2_fill_8 FILLER_4_1031 ();
 sg13g2_fill_8 FILLER_4_1039 ();
 sg13g2_fill_8 FILLER_4_1047 ();
 sg13g2_fill_8 FILLER_4_1055 ();
 sg13g2_fill_8 FILLER_4_1063 ();
 sg13g2_fill_8 FILLER_4_1071 ();
 sg13g2_fill_8 FILLER_4_1079 ();
 sg13g2_fill_8 FILLER_4_1087 ();
 sg13g2_fill_8 FILLER_4_1095 ();
 sg13g2_fill_8 FILLER_4_1103 ();
 sg13g2_fill_8 FILLER_4_1111 ();
 sg13g2_fill_8 FILLER_4_1119 ();
 sg13g2_fill_8 FILLER_4_1127 ();
 sg13g2_fill_8 FILLER_4_1135 ();
 sg13g2_fill_8 FILLER_4_1143 ();
 sg13g2_fill_8 FILLER_4_1151 ();
 sg13g2_fill_8 FILLER_4_1159 ();
 sg13g2_fill_8 FILLER_4_1167 ();
 sg13g2_fill_8 FILLER_4_1175 ();
 sg13g2_fill_8 FILLER_4_1183 ();
 sg13g2_fill_8 FILLER_4_1191 ();
 sg13g2_fill_8 FILLER_4_1199 ();
 sg13g2_fill_8 FILLER_4_1207 ();
 sg13g2_fill_8 FILLER_4_1215 ();
 sg13g2_fill_8 FILLER_4_1223 ();
 sg13g2_fill_8 FILLER_4_1231 ();
 sg13g2_fill_8 FILLER_4_1239 ();
 sg13g2_fill_8 FILLER_4_1247 ();
 sg13g2_fill_8 FILLER_4_1255 ();
 sg13g2_fill_8 FILLER_4_1263 ();
 sg13g2_fill_8 FILLER_4_1271 ();
 sg13g2_fill_8 FILLER_4_1279 ();
 sg13g2_fill_8 FILLER_4_1287 ();
 sg13g2_fill_8 FILLER_4_1295 ();
 sg13g2_fill_8 FILLER_4_1303 ();
 sg13g2_fill_8 FILLER_4_1311 ();
 sg13g2_fill_8 FILLER_4_1319 ();
 sg13g2_fill_8 FILLER_4_1327 ();
 sg13g2_fill_8 FILLER_4_1335 ();
 sg13g2_fill_8 FILLER_4_1343 ();
 sg13g2_fill_8 FILLER_4_1351 ();
 sg13g2_fill_8 FILLER_4_1359 ();
 sg13g2_fill_8 FILLER_4_1367 ();
 sg13g2_fill_8 FILLER_4_1375 ();
 sg13g2_fill_8 FILLER_4_1383 ();
 sg13g2_fill_8 FILLER_4_1391 ();
 sg13g2_fill_8 FILLER_4_1399 ();
 sg13g2_fill_8 FILLER_4_1407 ();
 sg13g2_fill_8 FILLER_4_1415 ();
 sg13g2_fill_8 FILLER_4_1423 ();
 sg13g2_fill_8 FILLER_4_1431 ();
 sg13g2_fill_8 FILLER_4_1439 ();
 sg13g2_fill_8 FILLER_4_1447 ();
 sg13g2_fill_8 FILLER_4_1455 ();
 sg13g2_fill_8 FILLER_4_1463 ();
 sg13g2_fill_8 FILLER_4_1471 ();
 sg13g2_fill_8 FILLER_4_1479 ();
 sg13g2_fill_8 FILLER_4_1487 ();
 sg13g2_fill_8 FILLER_4_1495 ();
 sg13g2_fill_8 FILLER_4_1503 ();
 sg13g2_fill_8 FILLER_4_1511 ();
 sg13g2_fill_8 FILLER_4_1519 ();
 sg13g2_fill_8 FILLER_4_1527 ();
 sg13g2_fill_8 FILLER_4_1535 ();
 sg13g2_fill_8 FILLER_4_1543 ();
 sg13g2_fill_8 FILLER_4_1551 ();
 sg13g2_fill_8 FILLER_4_1559 ();
 sg13g2_fill_8 FILLER_4_1567 ();
 sg13g2_fill_8 FILLER_4_1575 ();
 sg13g2_fill_8 FILLER_4_1583 ();
 sg13g2_fill_1 FILLER_4_1591 ();
 sg13g2_fill_8 FILLER_5_0 ();
 sg13g2_fill_8 FILLER_5_8 ();
 sg13g2_fill_8 FILLER_5_16 ();
 sg13g2_fill_8 FILLER_5_24 ();
 sg13g2_fill_8 FILLER_5_32 ();
 sg13g2_fill_8 FILLER_5_40 ();
 sg13g2_fill_8 FILLER_5_48 ();
 sg13g2_fill_8 FILLER_5_56 ();
 sg13g2_fill_8 FILLER_5_64 ();
 sg13g2_fill_8 FILLER_5_72 ();
 sg13g2_fill_8 FILLER_5_80 ();
 sg13g2_fill_8 FILLER_5_88 ();
 sg13g2_fill_8 FILLER_5_96 ();
 sg13g2_fill_8 FILLER_5_104 ();
 sg13g2_fill_8 FILLER_5_112 ();
 sg13g2_fill_8 FILLER_5_120 ();
 sg13g2_fill_8 FILLER_5_128 ();
 sg13g2_fill_8 FILLER_5_136 ();
 sg13g2_fill_8 FILLER_5_144 ();
 sg13g2_fill_8 FILLER_5_152 ();
 sg13g2_fill_8 FILLER_5_160 ();
 sg13g2_fill_8 FILLER_5_168 ();
 sg13g2_fill_8 FILLER_5_176 ();
 sg13g2_fill_8 FILLER_5_184 ();
 sg13g2_fill_8 FILLER_5_192 ();
 sg13g2_fill_8 FILLER_5_200 ();
 sg13g2_fill_8 FILLER_5_208 ();
 sg13g2_fill_8 FILLER_5_216 ();
 sg13g2_fill_8 FILLER_5_224 ();
 sg13g2_fill_8 FILLER_5_232 ();
 sg13g2_fill_8 FILLER_5_240 ();
 sg13g2_fill_8 FILLER_5_248 ();
 sg13g2_fill_8 FILLER_5_256 ();
 sg13g2_fill_8 FILLER_5_264 ();
 sg13g2_fill_8 FILLER_5_272 ();
 sg13g2_fill_8 FILLER_5_280 ();
 sg13g2_fill_8 FILLER_5_288 ();
 sg13g2_fill_8 FILLER_5_296 ();
 sg13g2_fill_8 FILLER_5_304 ();
 sg13g2_fill_8 FILLER_5_312 ();
 sg13g2_fill_8 FILLER_5_320 ();
 sg13g2_fill_8 FILLER_5_328 ();
 sg13g2_fill_8 FILLER_5_336 ();
 sg13g2_fill_8 FILLER_5_344 ();
 sg13g2_fill_8 FILLER_5_352 ();
 sg13g2_fill_8 FILLER_5_360 ();
 sg13g2_fill_8 FILLER_5_368 ();
 sg13g2_fill_8 FILLER_5_376 ();
 sg13g2_fill_8 FILLER_5_384 ();
 sg13g2_fill_8 FILLER_5_392 ();
 sg13g2_fill_8 FILLER_5_400 ();
 sg13g2_fill_8 FILLER_5_408 ();
 sg13g2_fill_8 FILLER_5_416 ();
 sg13g2_fill_8 FILLER_5_424 ();
 sg13g2_fill_8 FILLER_5_432 ();
 sg13g2_fill_8 FILLER_5_440 ();
 sg13g2_fill_8 FILLER_5_448 ();
 sg13g2_fill_8 FILLER_5_456 ();
 sg13g2_fill_8 FILLER_5_464 ();
 sg13g2_fill_8 FILLER_5_472 ();
 sg13g2_fill_8 FILLER_5_480 ();
 sg13g2_fill_8 FILLER_5_488 ();
 sg13g2_fill_8 FILLER_5_496 ();
 sg13g2_fill_8 FILLER_5_504 ();
 sg13g2_fill_8 FILLER_5_512 ();
 sg13g2_fill_8 FILLER_5_520 ();
 sg13g2_fill_8 FILLER_5_528 ();
 sg13g2_fill_8 FILLER_5_536 ();
 sg13g2_fill_8 FILLER_5_544 ();
 sg13g2_fill_8 FILLER_5_552 ();
 sg13g2_fill_8 FILLER_5_560 ();
 sg13g2_fill_8 FILLER_5_568 ();
 sg13g2_fill_8 FILLER_5_576 ();
 sg13g2_fill_8 FILLER_5_584 ();
 sg13g2_fill_8 FILLER_5_592 ();
 sg13g2_fill_8 FILLER_5_600 ();
 sg13g2_fill_8 FILLER_5_608 ();
 sg13g2_fill_8 FILLER_5_616 ();
 sg13g2_fill_8 FILLER_5_624 ();
 sg13g2_fill_8 FILLER_5_632 ();
 sg13g2_fill_8 FILLER_5_640 ();
 sg13g2_fill_8 FILLER_5_648 ();
 sg13g2_fill_8 FILLER_5_656 ();
 sg13g2_fill_8 FILLER_5_664 ();
 sg13g2_fill_8 FILLER_5_672 ();
 sg13g2_fill_8 FILLER_5_680 ();
 sg13g2_fill_8 FILLER_5_688 ();
 sg13g2_fill_8 FILLER_5_696 ();
 sg13g2_fill_8 FILLER_5_704 ();
 sg13g2_fill_8 FILLER_5_712 ();
 sg13g2_fill_8 FILLER_5_720 ();
 sg13g2_fill_8 FILLER_5_728 ();
 sg13g2_fill_8 FILLER_5_736 ();
 sg13g2_fill_8 FILLER_5_744 ();
 sg13g2_fill_8 FILLER_5_752 ();
 sg13g2_fill_8 FILLER_5_760 ();
 sg13g2_fill_8 FILLER_5_768 ();
 sg13g2_fill_2 FILLER_5_776 ();
 sg13g2_fill_4 FILLER_5_791 ();
 sg13g2_fill_2 FILLER_5_795 ();
 sg13g2_fill_1 FILLER_5_797 ();
 sg13g2_fill_8 FILLER_5_824 ();
 sg13g2_fill_8 FILLER_5_868 ();
 sg13g2_fill_8 FILLER_5_876 ();
 sg13g2_fill_8 FILLER_5_884 ();
 sg13g2_fill_8 FILLER_5_892 ();
 sg13g2_fill_8 FILLER_5_900 ();
 sg13g2_fill_8 FILLER_5_908 ();
 sg13g2_fill_2 FILLER_5_916 ();
 sg13g2_fill_1 FILLER_5_918 ();
 sg13g2_fill_8 FILLER_5_945 ();
 sg13g2_fill_8 FILLER_5_953 ();
 sg13g2_fill_8 FILLER_5_961 ();
 sg13g2_fill_8 FILLER_5_969 ();
 sg13g2_fill_8 FILLER_5_977 ();
 sg13g2_fill_8 FILLER_5_985 ();
 sg13g2_fill_8 FILLER_5_993 ();
 sg13g2_fill_8 FILLER_5_1001 ();
 sg13g2_fill_8 FILLER_5_1009 ();
 sg13g2_fill_8 FILLER_5_1017 ();
 sg13g2_fill_8 FILLER_5_1025 ();
 sg13g2_fill_8 FILLER_5_1033 ();
 sg13g2_fill_8 FILLER_5_1041 ();
 sg13g2_fill_8 FILLER_5_1049 ();
 sg13g2_fill_2 FILLER_5_1057 ();
 sg13g2_fill_1 FILLER_5_1109 ();
 sg13g2_fill_8 FILLER_5_1135 ();
 sg13g2_fill_8 FILLER_5_1143 ();
 sg13g2_fill_8 FILLER_5_1151 ();
 sg13g2_fill_8 FILLER_5_1159 ();
 sg13g2_fill_8 FILLER_5_1167 ();
 sg13g2_fill_8 FILLER_5_1175 ();
 sg13g2_fill_8 FILLER_5_1183 ();
 sg13g2_fill_8 FILLER_5_1191 ();
 sg13g2_fill_8 FILLER_5_1199 ();
 sg13g2_fill_8 FILLER_5_1207 ();
 sg13g2_fill_8 FILLER_5_1215 ();
 sg13g2_fill_8 FILLER_5_1223 ();
 sg13g2_fill_8 FILLER_5_1231 ();
 sg13g2_fill_8 FILLER_5_1239 ();
 sg13g2_fill_8 FILLER_5_1247 ();
 sg13g2_fill_8 FILLER_5_1255 ();
 sg13g2_fill_8 FILLER_5_1263 ();
 sg13g2_fill_8 FILLER_5_1271 ();
 sg13g2_fill_8 FILLER_5_1279 ();
 sg13g2_fill_8 FILLER_5_1287 ();
 sg13g2_fill_8 FILLER_5_1295 ();
 sg13g2_fill_8 FILLER_5_1303 ();
 sg13g2_fill_8 FILLER_5_1311 ();
 sg13g2_fill_8 FILLER_5_1319 ();
 sg13g2_fill_8 FILLER_5_1327 ();
 sg13g2_fill_8 FILLER_5_1335 ();
 sg13g2_fill_8 FILLER_5_1343 ();
 sg13g2_fill_8 FILLER_5_1351 ();
 sg13g2_fill_8 FILLER_5_1359 ();
 sg13g2_fill_8 FILLER_5_1367 ();
 sg13g2_fill_8 FILLER_5_1375 ();
 sg13g2_fill_8 FILLER_5_1383 ();
 sg13g2_fill_8 FILLER_5_1391 ();
 sg13g2_fill_8 FILLER_5_1399 ();
 sg13g2_fill_8 FILLER_5_1407 ();
 sg13g2_fill_8 FILLER_5_1415 ();
 sg13g2_fill_8 FILLER_5_1423 ();
 sg13g2_fill_8 FILLER_5_1431 ();
 sg13g2_fill_8 FILLER_5_1439 ();
 sg13g2_fill_8 FILLER_5_1447 ();
 sg13g2_fill_8 FILLER_5_1455 ();
 sg13g2_fill_8 FILLER_5_1463 ();
 sg13g2_fill_8 FILLER_5_1471 ();
 sg13g2_fill_8 FILLER_5_1479 ();
 sg13g2_fill_8 FILLER_5_1487 ();
 sg13g2_fill_8 FILLER_5_1495 ();
 sg13g2_fill_8 FILLER_5_1503 ();
 sg13g2_fill_8 FILLER_5_1511 ();
 sg13g2_fill_8 FILLER_5_1519 ();
 sg13g2_fill_8 FILLER_5_1527 ();
 sg13g2_fill_8 FILLER_5_1535 ();
 sg13g2_fill_8 FILLER_5_1543 ();
 sg13g2_fill_8 FILLER_5_1551 ();
 sg13g2_fill_8 FILLER_5_1559 ();
 sg13g2_fill_8 FILLER_5_1567 ();
 sg13g2_fill_8 FILLER_5_1575 ();
 sg13g2_fill_8 FILLER_5_1583 ();
 sg13g2_fill_1 FILLER_5_1591 ();
 sg13g2_fill_8 FILLER_6_0 ();
 sg13g2_fill_8 FILLER_6_8 ();
 sg13g2_fill_8 FILLER_6_16 ();
 sg13g2_fill_8 FILLER_6_24 ();
 sg13g2_fill_8 FILLER_6_32 ();
 sg13g2_fill_8 FILLER_6_40 ();
 sg13g2_fill_8 FILLER_6_48 ();
 sg13g2_fill_8 FILLER_6_56 ();
 sg13g2_fill_8 FILLER_6_64 ();
 sg13g2_fill_8 FILLER_6_72 ();
 sg13g2_fill_8 FILLER_6_80 ();
 sg13g2_fill_8 FILLER_6_88 ();
 sg13g2_fill_8 FILLER_6_96 ();
 sg13g2_fill_8 FILLER_6_104 ();
 sg13g2_fill_8 FILLER_6_112 ();
 sg13g2_fill_8 FILLER_6_120 ();
 sg13g2_fill_8 FILLER_6_128 ();
 sg13g2_fill_8 FILLER_6_136 ();
 sg13g2_fill_8 FILLER_6_144 ();
 sg13g2_fill_8 FILLER_6_152 ();
 sg13g2_fill_8 FILLER_6_160 ();
 sg13g2_fill_8 FILLER_6_168 ();
 sg13g2_fill_8 FILLER_6_176 ();
 sg13g2_fill_8 FILLER_6_184 ();
 sg13g2_fill_8 FILLER_6_192 ();
 sg13g2_fill_8 FILLER_6_200 ();
 sg13g2_fill_8 FILLER_6_208 ();
 sg13g2_fill_8 FILLER_6_216 ();
 sg13g2_fill_8 FILLER_6_224 ();
 sg13g2_fill_8 FILLER_6_232 ();
 sg13g2_fill_8 FILLER_6_240 ();
 sg13g2_fill_8 FILLER_6_248 ();
 sg13g2_fill_8 FILLER_6_256 ();
 sg13g2_fill_8 FILLER_6_264 ();
 sg13g2_fill_8 FILLER_6_272 ();
 sg13g2_fill_8 FILLER_6_280 ();
 sg13g2_fill_8 FILLER_6_288 ();
 sg13g2_fill_8 FILLER_6_296 ();
 sg13g2_fill_8 FILLER_6_304 ();
 sg13g2_fill_8 FILLER_6_312 ();
 sg13g2_fill_8 FILLER_6_320 ();
 sg13g2_fill_8 FILLER_6_328 ();
 sg13g2_fill_8 FILLER_6_336 ();
 sg13g2_fill_8 FILLER_6_344 ();
 sg13g2_fill_8 FILLER_6_352 ();
 sg13g2_fill_8 FILLER_6_360 ();
 sg13g2_fill_8 FILLER_6_368 ();
 sg13g2_fill_8 FILLER_6_376 ();
 sg13g2_fill_8 FILLER_6_384 ();
 sg13g2_fill_8 FILLER_6_392 ();
 sg13g2_fill_8 FILLER_6_400 ();
 sg13g2_fill_8 FILLER_6_408 ();
 sg13g2_fill_8 FILLER_6_416 ();
 sg13g2_fill_8 FILLER_6_424 ();
 sg13g2_fill_8 FILLER_6_432 ();
 sg13g2_fill_8 FILLER_6_440 ();
 sg13g2_fill_8 FILLER_6_448 ();
 sg13g2_fill_8 FILLER_6_456 ();
 sg13g2_fill_8 FILLER_6_464 ();
 sg13g2_fill_8 FILLER_6_472 ();
 sg13g2_fill_8 FILLER_6_480 ();
 sg13g2_fill_8 FILLER_6_488 ();
 sg13g2_fill_8 FILLER_6_496 ();
 sg13g2_fill_8 FILLER_6_504 ();
 sg13g2_fill_8 FILLER_6_512 ();
 sg13g2_fill_8 FILLER_6_520 ();
 sg13g2_fill_8 FILLER_6_528 ();
 sg13g2_fill_8 FILLER_6_536 ();
 sg13g2_fill_8 FILLER_6_544 ();
 sg13g2_fill_8 FILLER_6_552 ();
 sg13g2_fill_8 FILLER_6_560 ();
 sg13g2_fill_8 FILLER_6_568 ();
 sg13g2_fill_8 FILLER_6_576 ();
 sg13g2_fill_8 FILLER_6_584 ();
 sg13g2_fill_8 FILLER_6_592 ();
 sg13g2_fill_8 FILLER_6_600 ();
 sg13g2_fill_8 FILLER_6_608 ();
 sg13g2_fill_8 FILLER_6_616 ();
 sg13g2_fill_8 FILLER_6_624 ();
 sg13g2_fill_8 FILLER_6_632 ();
 sg13g2_fill_8 FILLER_6_640 ();
 sg13g2_fill_8 FILLER_6_648 ();
 sg13g2_fill_8 FILLER_6_656 ();
 sg13g2_fill_8 FILLER_6_664 ();
 sg13g2_fill_8 FILLER_6_672 ();
 sg13g2_fill_8 FILLER_6_680 ();
 sg13g2_fill_8 FILLER_6_688 ();
 sg13g2_fill_8 FILLER_6_696 ();
 sg13g2_fill_8 FILLER_6_704 ();
 sg13g2_fill_8 FILLER_6_712 ();
 sg13g2_fill_8 FILLER_6_720 ();
 sg13g2_fill_8 FILLER_6_728 ();
 sg13g2_fill_8 FILLER_6_736 ();
 sg13g2_fill_4 FILLER_6_744 ();
 sg13g2_fill_2 FILLER_6_748 ();
 sg13g2_fill_1 FILLER_6_750 ();
 sg13g2_fill_4 FILLER_6_777 ();
 sg13g2_fill_1 FILLER_6_781 ();
 sg13g2_fill_4 FILLER_6_795 ();
 sg13g2_fill_2 FILLER_6_799 ();
 sg13g2_fill_4 FILLER_6_809 ();
 sg13g2_fill_1 FILLER_6_813 ();
 sg13g2_fill_2 FILLER_6_819 ();
 sg13g2_fill_8 FILLER_6_855 ();
 sg13g2_fill_8 FILLER_6_863 ();
 sg13g2_fill_8 FILLER_6_871 ();
 sg13g2_fill_1 FILLER_6_879 ();
 sg13g2_fill_1 FILLER_6_921 ();
 sg13g2_fill_8 FILLER_6_948 ();
 sg13g2_fill_8 FILLER_6_956 ();
 sg13g2_fill_8 FILLER_6_964 ();
 sg13g2_fill_8 FILLER_6_972 ();
 sg13g2_fill_8 FILLER_6_980 ();
 sg13g2_fill_8 FILLER_6_988 ();
 sg13g2_fill_8 FILLER_6_996 ();
 sg13g2_fill_8 FILLER_6_1004 ();
 sg13g2_fill_8 FILLER_6_1012 ();
 sg13g2_fill_8 FILLER_6_1020 ();
 sg13g2_fill_8 FILLER_6_1028 ();
 sg13g2_fill_8 FILLER_6_1036 ();
 sg13g2_fill_8 FILLER_6_1044 ();
 sg13g2_fill_8 FILLER_6_1052 ();
 sg13g2_fill_8 FILLER_6_1060 ();
 sg13g2_fill_8 FILLER_6_1068 ();
 sg13g2_fill_8 FILLER_6_1076 ();
 sg13g2_fill_8 FILLER_6_1084 ();
 sg13g2_fill_1 FILLER_6_1092 ();
 sg13g2_fill_2 FILLER_6_1107 ();
 sg13g2_fill_1 FILLER_6_1109 ();
 sg13g2_fill_8 FILLER_6_1140 ();
 sg13g2_fill_8 FILLER_6_1148 ();
 sg13g2_fill_8 FILLER_6_1156 ();
 sg13g2_fill_8 FILLER_6_1164 ();
 sg13g2_fill_8 FILLER_6_1172 ();
 sg13g2_fill_8 FILLER_6_1180 ();
 sg13g2_fill_8 FILLER_6_1188 ();
 sg13g2_fill_8 FILLER_6_1196 ();
 sg13g2_fill_8 FILLER_6_1204 ();
 sg13g2_fill_8 FILLER_6_1212 ();
 sg13g2_fill_8 FILLER_6_1220 ();
 sg13g2_fill_8 FILLER_6_1228 ();
 sg13g2_fill_8 FILLER_6_1236 ();
 sg13g2_fill_8 FILLER_6_1244 ();
 sg13g2_fill_8 FILLER_6_1252 ();
 sg13g2_fill_8 FILLER_6_1260 ();
 sg13g2_fill_8 FILLER_6_1268 ();
 sg13g2_fill_8 FILLER_6_1276 ();
 sg13g2_fill_8 FILLER_6_1284 ();
 sg13g2_fill_8 FILLER_6_1292 ();
 sg13g2_fill_8 FILLER_6_1300 ();
 sg13g2_fill_8 FILLER_6_1308 ();
 sg13g2_fill_8 FILLER_6_1316 ();
 sg13g2_fill_8 FILLER_6_1324 ();
 sg13g2_fill_8 FILLER_6_1332 ();
 sg13g2_fill_8 FILLER_6_1340 ();
 sg13g2_fill_8 FILLER_6_1348 ();
 sg13g2_fill_8 FILLER_6_1356 ();
 sg13g2_fill_8 FILLER_6_1364 ();
 sg13g2_fill_8 FILLER_6_1372 ();
 sg13g2_fill_8 FILLER_6_1380 ();
 sg13g2_fill_8 FILLER_6_1388 ();
 sg13g2_fill_8 FILLER_6_1396 ();
 sg13g2_fill_8 FILLER_6_1404 ();
 sg13g2_fill_8 FILLER_6_1412 ();
 sg13g2_fill_8 FILLER_6_1420 ();
 sg13g2_fill_8 FILLER_6_1428 ();
 sg13g2_fill_8 FILLER_6_1436 ();
 sg13g2_fill_8 FILLER_6_1444 ();
 sg13g2_fill_8 FILLER_6_1452 ();
 sg13g2_fill_8 FILLER_6_1460 ();
 sg13g2_fill_8 FILLER_6_1468 ();
 sg13g2_fill_8 FILLER_6_1476 ();
 sg13g2_fill_8 FILLER_6_1484 ();
 sg13g2_fill_8 FILLER_6_1492 ();
 sg13g2_fill_8 FILLER_6_1500 ();
 sg13g2_fill_8 FILLER_6_1508 ();
 sg13g2_fill_8 FILLER_6_1516 ();
 sg13g2_fill_8 FILLER_6_1524 ();
 sg13g2_fill_8 FILLER_6_1532 ();
 sg13g2_fill_8 FILLER_6_1540 ();
 sg13g2_fill_8 FILLER_6_1548 ();
 sg13g2_fill_8 FILLER_6_1556 ();
 sg13g2_fill_8 FILLER_6_1564 ();
 sg13g2_fill_8 FILLER_6_1572 ();
 sg13g2_fill_8 FILLER_6_1580 ();
 sg13g2_fill_4 FILLER_6_1588 ();
 sg13g2_fill_8 FILLER_7_0 ();
 sg13g2_fill_8 FILLER_7_8 ();
 sg13g2_fill_8 FILLER_7_16 ();
 sg13g2_fill_8 FILLER_7_24 ();
 sg13g2_fill_8 FILLER_7_32 ();
 sg13g2_fill_8 FILLER_7_40 ();
 sg13g2_fill_8 FILLER_7_48 ();
 sg13g2_fill_8 FILLER_7_56 ();
 sg13g2_fill_8 FILLER_7_64 ();
 sg13g2_fill_8 FILLER_7_72 ();
 sg13g2_fill_8 FILLER_7_80 ();
 sg13g2_fill_8 FILLER_7_88 ();
 sg13g2_fill_8 FILLER_7_96 ();
 sg13g2_fill_8 FILLER_7_104 ();
 sg13g2_fill_8 FILLER_7_112 ();
 sg13g2_fill_8 FILLER_7_120 ();
 sg13g2_fill_8 FILLER_7_128 ();
 sg13g2_fill_8 FILLER_7_136 ();
 sg13g2_fill_8 FILLER_7_144 ();
 sg13g2_fill_8 FILLER_7_152 ();
 sg13g2_fill_8 FILLER_7_160 ();
 sg13g2_fill_8 FILLER_7_168 ();
 sg13g2_fill_8 FILLER_7_176 ();
 sg13g2_fill_8 FILLER_7_184 ();
 sg13g2_fill_8 FILLER_7_192 ();
 sg13g2_fill_8 FILLER_7_200 ();
 sg13g2_fill_8 FILLER_7_208 ();
 sg13g2_fill_8 FILLER_7_216 ();
 sg13g2_fill_8 FILLER_7_224 ();
 sg13g2_fill_8 FILLER_7_232 ();
 sg13g2_fill_8 FILLER_7_240 ();
 sg13g2_fill_8 FILLER_7_248 ();
 sg13g2_fill_8 FILLER_7_256 ();
 sg13g2_fill_8 FILLER_7_264 ();
 sg13g2_fill_8 FILLER_7_272 ();
 sg13g2_fill_8 FILLER_7_280 ();
 sg13g2_fill_8 FILLER_7_288 ();
 sg13g2_fill_8 FILLER_7_296 ();
 sg13g2_fill_8 FILLER_7_304 ();
 sg13g2_fill_8 FILLER_7_312 ();
 sg13g2_fill_8 FILLER_7_320 ();
 sg13g2_fill_8 FILLER_7_328 ();
 sg13g2_fill_8 FILLER_7_336 ();
 sg13g2_fill_8 FILLER_7_344 ();
 sg13g2_fill_8 FILLER_7_352 ();
 sg13g2_fill_8 FILLER_7_360 ();
 sg13g2_fill_8 FILLER_7_368 ();
 sg13g2_fill_8 FILLER_7_376 ();
 sg13g2_fill_8 FILLER_7_384 ();
 sg13g2_fill_8 FILLER_7_392 ();
 sg13g2_fill_8 FILLER_7_400 ();
 sg13g2_fill_8 FILLER_7_408 ();
 sg13g2_fill_8 FILLER_7_416 ();
 sg13g2_fill_8 FILLER_7_424 ();
 sg13g2_fill_8 FILLER_7_432 ();
 sg13g2_fill_8 FILLER_7_440 ();
 sg13g2_fill_8 FILLER_7_448 ();
 sg13g2_fill_8 FILLER_7_456 ();
 sg13g2_fill_8 FILLER_7_464 ();
 sg13g2_fill_8 FILLER_7_472 ();
 sg13g2_fill_8 FILLER_7_480 ();
 sg13g2_fill_8 FILLER_7_488 ();
 sg13g2_fill_8 FILLER_7_496 ();
 sg13g2_fill_8 FILLER_7_504 ();
 sg13g2_fill_8 FILLER_7_512 ();
 sg13g2_fill_8 FILLER_7_520 ();
 sg13g2_fill_8 FILLER_7_528 ();
 sg13g2_fill_8 FILLER_7_536 ();
 sg13g2_fill_8 FILLER_7_544 ();
 sg13g2_fill_8 FILLER_7_552 ();
 sg13g2_fill_8 FILLER_7_560 ();
 sg13g2_fill_8 FILLER_7_568 ();
 sg13g2_fill_8 FILLER_7_576 ();
 sg13g2_fill_8 FILLER_7_584 ();
 sg13g2_fill_8 FILLER_7_592 ();
 sg13g2_fill_8 FILLER_7_600 ();
 sg13g2_fill_8 FILLER_7_608 ();
 sg13g2_fill_8 FILLER_7_616 ();
 sg13g2_fill_8 FILLER_7_624 ();
 sg13g2_fill_8 FILLER_7_632 ();
 sg13g2_fill_8 FILLER_7_640 ();
 sg13g2_fill_8 FILLER_7_648 ();
 sg13g2_fill_8 FILLER_7_656 ();
 sg13g2_fill_8 FILLER_7_664 ();
 sg13g2_fill_8 FILLER_7_672 ();
 sg13g2_fill_8 FILLER_7_680 ();
 sg13g2_fill_8 FILLER_7_688 ();
 sg13g2_fill_8 FILLER_7_696 ();
 sg13g2_fill_8 FILLER_7_704 ();
 sg13g2_fill_8 FILLER_7_712 ();
 sg13g2_fill_8 FILLER_7_720 ();
 sg13g2_fill_8 FILLER_7_728 ();
 sg13g2_fill_8 FILLER_7_736 ();
 sg13g2_fill_8 FILLER_7_744 ();
 sg13g2_fill_8 FILLER_7_752 ();
 sg13g2_fill_2 FILLER_7_760 ();
 sg13g2_fill_2 FILLER_7_818 ();
 sg13g2_fill_1 FILLER_7_820 ();
 sg13g2_fill_8 FILLER_7_842 ();
 sg13g2_fill_8 FILLER_7_850 ();
 sg13g2_fill_2 FILLER_7_858 ();
 sg13g2_fill_1 FILLER_7_860 ();
 sg13g2_fill_1 FILLER_7_877 ();
 sg13g2_fill_8 FILLER_7_929 ();
 sg13g2_fill_8 FILLER_7_937 ();
 sg13g2_fill_1 FILLER_7_945 ();
 sg13g2_fill_8 FILLER_7_951 ();
 sg13g2_fill_4 FILLER_7_959 ();
 sg13g2_fill_1 FILLER_7_963 ();
 sg13g2_fill_8 FILLER_7_990 ();
 sg13g2_fill_8 FILLER_7_998 ();
 sg13g2_fill_8 FILLER_7_1006 ();
 sg13g2_fill_8 FILLER_7_1014 ();
 sg13g2_fill_8 FILLER_7_1022 ();
 sg13g2_fill_8 FILLER_7_1030 ();
 sg13g2_fill_8 FILLER_7_1038 ();
 sg13g2_fill_8 FILLER_7_1046 ();
 sg13g2_fill_8 FILLER_7_1054 ();
 sg13g2_fill_8 FILLER_7_1062 ();
 sg13g2_fill_8 FILLER_7_1070 ();
 sg13g2_fill_4 FILLER_7_1078 ();
 sg13g2_fill_4 FILLER_7_1108 ();
 sg13g2_fill_1 FILLER_7_1112 ();
 sg13g2_fill_8 FILLER_7_1138 ();
 sg13g2_fill_8 FILLER_7_1146 ();
 sg13g2_fill_8 FILLER_7_1154 ();
 sg13g2_fill_8 FILLER_7_1162 ();
 sg13g2_fill_8 FILLER_7_1170 ();
 sg13g2_fill_8 FILLER_7_1178 ();
 sg13g2_fill_8 FILLER_7_1186 ();
 sg13g2_fill_8 FILLER_7_1194 ();
 sg13g2_fill_8 FILLER_7_1202 ();
 sg13g2_fill_8 FILLER_7_1210 ();
 sg13g2_fill_8 FILLER_7_1218 ();
 sg13g2_fill_8 FILLER_7_1226 ();
 sg13g2_fill_8 FILLER_7_1234 ();
 sg13g2_fill_8 FILLER_7_1242 ();
 sg13g2_fill_8 FILLER_7_1250 ();
 sg13g2_fill_8 FILLER_7_1258 ();
 sg13g2_fill_8 FILLER_7_1266 ();
 sg13g2_fill_8 FILLER_7_1274 ();
 sg13g2_fill_8 FILLER_7_1282 ();
 sg13g2_fill_8 FILLER_7_1290 ();
 sg13g2_fill_8 FILLER_7_1298 ();
 sg13g2_fill_8 FILLER_7_1306 ();
 sg13g2_fill_8 FILLER_7_1314 ();
 sg13g2_fill_8 FILLER_7_1322 ();
 sg13g2_fill_8 FILLER_7_1330 ();
 sg13g2_fill_8 FILLER_7_1338 ();
 sg13g2_fill_8 FILLER_7_1346 ();
 sg13g2_fill_8 FILLER_7_1354 ();
 sg13g2_fill_8 FILLER_7_1362 ();
 sg13g2_fill_8 FILLER_7_1370 ();
 sg13g2_fill_8 FILLER_7_1378 ();
 sg13g2_fill_8 FILLER_7_1386 ();
 sg13g2_fill_8 FILLER_7_1394 ();
 sg13g2_fill_8 FILLER_7_1402 ();
 sg13g2_fill_8 FILLER_7_1410 ();
 sg13g2_fill_8 FILLER_7_1418 ();
 sg13g2_fill_8 FILLER_7_1426 ();
 sg13g2_fill_8 FILLER_7_1434 ();
 sg13g2_fill_8 FILLER_7_1442 ();
 sg13g2_fill_8 FILLER_7_1450 ();
 sg13g2_fill_8 FILLER_7_1458 ();
 sg13g2_fill_8 FILLER_7_1466 ();
 sg13g2_fill_8 FILLER_7_1474 ();
 sg13g2_fill_8 FILLER_7_1482 ();
 sg13g2_fill_8 FILLER_7_1490 ();
 sg13g2_fill_8 FILLER_7_1498 ();
 sg13g2_fill_8 FILLER_7_1506 ();
 sg13g2_fill_8 FILLER_7_1514 ();
 sg13g2_fill_8 FILLER_7_1522 ();
 sg13g2_fill_8 FILLER_7_1530 ();
 sg13g2_fill_8 FILLER_7_1538 ();
 sg13g2_fill_8 FILLER_7_1546 ();
 sg13g2_fill_8 FILLER_7_1554 ();
 sg13g2_fill_8 FILLER_7_1562 ();
 sg13g2_fill_8 FILLER_7_1570 ();
 sg13g2_fill_8 FILLER_7_1578 ();
 sg13g2_fill_4 FILLER_7_1586 ();
 sg13g2_fill_2 FILLER_7_1590 ();
 sg13g2_fill_8 FILLER_8_0 ();
 sg13g2_fill_8 FILLER_8_8 ();
 sg13g2_fill_8 FILLER_8_16 ();
 sg13g2_fill_8 FILLER_8_24 ();
 sg13g2_fill_8 FILLER_8_32 ();
 sg13g2_fill_8 FILLER_8_40 ();
 sg13g2_fill_8 FILLER_8_48 ();
 sg13g2_fill_8 FILLER_8_56 ();
 sg13g2_fill_8 FILLER_8_64 ();
 sg13g2_fill_8 FILLER_8_72 ();
 sg13g2_fill_8 FILLER_8_80 ();
 sg13g2_fill_8 FILLER_8_88 ();
 sg13g2_fill_8 FILLER_8_96 ();
 sg13g2_fill_8 FILLER_8_104 ();
 sg13g2_fill_8 FILLER_8_112 ();
 sg13g2_fill_8 FILLER_8_120 ();
 sg13g2_fill_8 FILLER_8_128 ();
 sg13g2_fill_8 FILLER_8_136 ();
 sg13g2_fill_8 FILLER_8_144 ();
 sg13g2_fill_8 FILLER_8_152 ();
 sg13g2_fill_8 FILLER_8_160 ();
 sg13g2_fill_8 FILLER_8_168 ();
 sg13g2_fill_8 FILLER_8_176 ();
 sg13g2_fill_8 FILLER_8_184 ();
 sg13g2_fill_8 FILLER_8_192 ();
 sg13g2_fill_8 FILLER_8_200 ();
 sg13g2_fill_8 FILLER_8_208 ();
 sg13g2_fill_8 FILLER_8_216 ();
 sg13g2_fill_8 FILLER_8_224 ();
 sg13g2_fill_8 FILLER_8_232 ();
 sg13g2_fill_8 FILLER_8_240 ();
 sg13g2_fill_8 FILLER_8_248 ();
 sg13g2_fill_8 FILLER_8_256 ();
 sg13g2_fill_8 FILLER_8_264 ();
 sg13g2_fill_8 FILLER_8_272 ();
 sg13g2_fill_8 FILLER_8_280 ();
 sg13g2_fill_8 FILLER_8_288 ();
 sg13g2_fill_8 FILLER_8_296 ();
 sg13g2_fill_8 FILLER_8_304 ();
 sg13g2_fill_8 FILLER_8_312 ();
 sg13g2_fill_8 FILLER_8_320 ();
 sg13g2_fill_8 FILLER_8_328 ();
 sg13g2_fill_8 FILLER_8_336 ();
 sg13g2_fill_8 FILLER_8_344 ();
 sg13g2_fill_8 FILLER_8_352 ();
 sg13g2_fill_8 FILLER_8_360 ();
 sg13g2_fill_8 FILLER_8_368 ();
 sg13g2_fill_8 FILLER_8_376 ();
 sg13g2_fill_8 FILLER_8_384 ();
 sg13g2_fill_8 FILLER_8_392 ();
 sg13g2_fill_8 FILLER_8_400 ();
 sg13g2_fill_8 FILLER_8_408 ();
 sg13g2_fill_8 FILLER_8_416 ();
 sg13g2_fill_8 FILLER_8_424 ();
 sg13g2_fill_8 FILLER_8_432 ();
 sg13g2_fill_8 FILLER_8_440 ();
 sg13g2_fill_8 FILLER_8_448 ();
 sg13g2_fill_8 FILLER_8_456 ();
 sg13g2_fill_8 FILLER_8_464 ();
 sg13g2_fill_8 FILLER_8_472 ();
 sg13g2_fill_8 FILLER_8_480 ();
 sg13g2_fill_8 FILLER_8_488 ();
 sg13g2_fill_8 FILLER_8_496 ();
 sg13g2_fill_8 FILLER_8_504 ();
 sg13g2_fill_8 FILLER_8_512 ();
 sg13g2_fill_8 FILLER_8_520 ();
 sg13g2_fill_8 FILLER_8_528 ();
 sg13g2_fill_8 FILLER_8_536 ();
 sg13g2_fill_8 FILLER_8_544 ();
 sg13g2_fill_8 FILLER_8_552 ();
 sg13g2_fill_8 FILLER_8_560 ();
 sg13g2_fill_8 FILLER_8_568 ();
 sg13g2_fill_8 FILLER_8_576 ();
 sg13g2_fill_8 FILLER_8_584 ();
 sg13g2_fill_8 FILLER_8_592 ();
 sg13g2_fill_8 FILLER_8_600 ();
 sg13g2_fill_8 FILLER_8_608 ();
 sg13g2_fill_8 FILLER_8_616 ();
 sg13g2_fill_8 FILLER_8_624 ();
 sg13g2_fill_8 FILLER_8_632 ();
 sg13g2_fill_8 FILLER_8_640 ();
 sg13g2_fill_2 FILLER_8_648 ();
 sg13g2_fill_8 FILLER_8_660 ();
 sg13g2_fill_8 FILLER_8_668 ();
 sg13g2_fill_8 FILLER_8_676 ();
 sg13g2_fill_8 FILLER_8_684 ();
 sg13g2_fill_8 FILLER_8_692 ();
 sg13g2_fill_8 FILLER_8_700 ();
 sg13g2_fill_8 FILLER_8_708 ();
 sg13g2_fill_8 FILLER_8_716 ();
 sg13g2_fill_8 FILLER_8_724 ();
 sg13g2_fill_8 FILLER_8_732 ();
 sg13g2_fill_8 FILLER_8_740 ();
 sg13g2_fill_8 FILLER_8_748 ();
 sg13g2_fill_8 FILLER_8_756 ();
 sg13g2_fill_4 FILLER_8_764 ();
 sg13g2_fill_2 FILLER_8_768 ();
 sg13g2_fill_2 FILLER_8_806 ();
 sg13g2_fill_1 FILLER_8_808 ();
 sg13g2_fill_4 FILLER_8_830 ();
 sg13g2_fill_2 FILLER_8_834 ();
 sg13g2_fill_1 FILLER_8_836 ();
 sg13g2_fill_2 FILLER_8_873 ();
 sg13g2_fill_8 FILLER_8_886 ();
 sg13g2_fill_2 FILLER_8_894 ();
 sg13g2_fill_4 FILLER_8_901 ();
 sg13g2_fill_4 FILLER_8_936 ();
 sg13g2_fill_1 FILLER_8_940 ();
 sg13g2_fill_8 FILLER_8_977 ();
 sg13g2_fill_8 FILLER_8_985 ();
 sg13g2_fill_8 FILLER_8_993 ();
 sg13g2_fill_8 FILLER_8_1001 ();
 sg13g2_fill_8 FILLER_8_1009 ();
 sg13g2_fill_8 FILLER_8_1017 ();
 sg13g2_fill_8 FILLER_8_1025 ();
 sg13g2_fill_4 FILLER_8_1033 ();
 sg13g2_fill_2 FILLER_8_1037 ();
 sg13g2_fill_8 FILLER_8_1047 ();
 sg13g2_fill_4 FILLER_8_1055 ();
 sg13g2_fill_8 FILLER_8_1095 ();
 sg13g2_fill_8 FILLER_8_1139 ();
 sg13g2_fill_1 FILLER_8_1147 ();
 sg13g2_fill_8 FILLER_8_1174 ();
 sg13g2_fill_8 FILLER_8_1182 ();
 sg13g2_fill_8 FILLER_8_1190 ();
 sg13g2_fill_8 FILLER_8_1198 ();
 sg13g2_fill_8 FILLER_8_1206 ();
 sg13g2_fill_8 FILLER_8_1214 ();
 sg13g2_fill_8 FILLER_8_1222 ();
 sg13g2_fill_8 FILLER_8_1230 ();
 sg13g2_fill_8 FILLER_8_1238 ();
 sg13g2_fill_8 FILLER_8_1246 ();
 sg13g2_fill_8 FILLER_8_1254 ();
 sg13g2_fill_8 FILLER_8_1262 ();
 sg13g2_fill_8 FILLER_8_1270 ();
 sg13g2_fill_8 FILLER_8_1278 ();
 sg13g2_fill_8 FILLER_8_1286 ();
 sg13g2_fill_8 FILLER_8_1294 ();
 sg13g2_fill_8 FILLER_8_1302 ();
 sg13g2_fill_8 FILLER_8_1310 ();
 sg13g2_fill_8 FILLER_8_1318 ();
 sg13g2_fill_8 FILLER_8_1326 ();
 sg13g2_fill_8 FILLER_8_1334 ();
 sg13g2_fill_8 FILLER_8_1342 ();
 sg13g2_fill_8 FILLER_8_1350 ();
 sg13g2_fill_8 FILLER_8_1358 ();
 sg13g2_fill_8 FILLER_8_1366 ();
 sg13g2_fill_8 FILLER_8_1374 ();
 sg13g2_fill_8 FILLER_8_1382 ();
 sg13g2_fill_8 FILLER_8_1390 ();
 sg13g2_fill_8 FILLER_8_1398 ();
 sg13g2_fill_8 FILLER_8_1406 ();
 sg13g2_fill_8 FILLER_8_1414 ();
 sg13g2_fill_8 FILLER_8_1422 ();
 sg13g2_fill_8 FILLER_8_1430 ();
 sg13g2_fill_8 FILLER_8_1438 ();
 sg13g2_fill_8 FILLER_8_1446 ();
 sg13g2_fill_8 FILLER_8_1454 ();
 sg13g2_fill_8 FILLER_8_1462 ();
 sg13g2_fill_8 FILLER_8_1470 ();
 sg13g2_fill_8 FILLER_8_1478 ();
 sg13g2_fill_8 FILLER_8_1486 ();
 sg13g2_fill_8 FILLER_8_1494 ();
 sg13g2_fill_8 FILLER_8_1502 ();
 sg13g2_fill_8 FILLER_8_1510 ();
 sg13g2_fill_8 FILLER_8_1518 ();
 sg13g2_fill_8 FILLER_8_1526 ();
 sg13g2_fill_8 FILLER_8_1534 ();
 sg13g2_fill_8 FILLER_8_1542 ();
 sg13g2_fill_8 FILLER_8_1550 ();
 sg13g2_fill_8 FILLER_8_1558 ();
 sg13g2_fill_8 FILLER_8_1566 ();
 sg13g2_fill_8 FILLER_8_1574 ();
 sg13g2_fill_8 FILLER_8_1582 ();
 sg13g2_fill_2 FILLER_8_1590 ();
 sg13g2_fill_8 FILLER_9_0 ();
 sg13g2_fill_8 FILLER_9_8 ();
 sg13g2_fill_8 FILLER_9_16 ();
 sg13g2_fill_8 FILLER_9_24 ();
 sg13g2_fill_8 FILLER_9_32 ();
 sg13g2_fill_8 FILLER_9_40 ();
 sg13g2_fill_8 FILLER_9_48 ();
 sg13g2_fill_8 FILLER_9_56 ();
 sg13g2_fill_8 FILLER_9_64 ();
 sg13g2_fill_8 FILLER_9_72 ();
 sg13g2_fill_8 FILLER_9_80 ();
 sg13g2_fill_8 FILLER_9_88 ();
 sg13g2_fill_8 FILLER_9_96 ();
 sg13g2_fill_8 FILLER_9_104 ();
 sg13g2_fill_8 FILLER_9_112 ();
 sg13g2_fill_8 FILLER_9_120 ();
 sg13g2_fill_8 FILLER_9_128 ();
 sg13g2_fill_8 FILLER_9_136 ();
 sg13g2_fill_8 FILLER_9_144 ();
 sg13g2_fill_8 FILLER_9_152 ();
 sg13g2_fill_8 FILLER_9_160 ();
 sg13g2_fill_8 FILLER_9_168 ();
 sg13g2_fill_8 FILLER_9_176 ();
 sg13g2_fill_8 FILLER_9_184 ();
 sg13g2_fill_8 FILLER_9_192 ();
 sg13g2_fill_8 FILLER_9_200 ();
 sg13g2_fill_8 FILLER_9_208 ();
 sg13g2_fill_8 FILLER_9_216 ();
 sg13g2_fill_8 FILLER_9_224 ();
 sg13g2_fill_8 FILLER_9_232 ();
 sg13g2_fill_8 FILLER_9_240 ();
 sg13g2_fill_8 FILLER_9_248 ();
 sg13g2_fill_8 FILLER_9_256 ();
 sg13g2_fill_8 FILLER_9_264 ();
 sg13g2_fill_8 FILLER_9_272 ();
 sg13g2_fill_8 FILLER_9_280 ();
 sg13g2_fill_8 FILLER_9_288 ();
 sg13g2_fill_8 FILLER_9_296 ();
 sg13g2_fill_8 FILLER_9_304 ();
 sg13g2_fill_8 FILLER_9_312 ();
 sg13g2_fill_8 FILLER_9_320 ();
 sg13g2_fill_8 FILLER_9_328 ();
 sg13g2_fill_8 FILLER_9_336 ();
 sg13g2_fill_8 FILLER_9_344 ();
 sg13g2_fill_8 FILLER_9_352 ();
 sg13g2_fill_8 FILLER_9_360 ();
 sg13g2_fill_8 FILLER_9_368 ();
 sg13g2_fill_8 FILLER_9_376 ();
 sg13g2_fill_8 FILLER_9_384 ();
 sg13g2_fill_8 FILLER_9_392 ();
 sg13g2_fill_8 FILLER_9_400 ();
 sg13g2_fill_8 FILLER_9_408 ();
 sg13g2_fill_8 FILLER_9_416 ();
 sg13g2_fill_8 FILLER_9_424 ();
 sg13g2_fill_8 FILLER_9_432 ();
 sg13g2_fill_8 FILLER_9_440 ();
 sg13g2_fill_8 FILLER_9_448 ();
 sg13g2_fill_8 FILLER_9_456 ();
 sg13g2_fill_8 FILLER_9_464 ();
 sg13g2_fill_8 FILLER_9_472 ();
 sg13g2_fill_8 FILLER_9_480 ();
 sg13g2_fill_8 FILLER_9_488 ();
 sg13g2_fill_8 FILLER_9_496 ();
 sg13g2_fill_8 FILLER_9_504 ();
 sg13g2_fill_8 FILLER_9_512 ();
 sg13g2_fill_8 FILLER_9_520 ();
 sg13g2_fill_8 FILLER_9_528 ();
 sg13g2_fill_8 FILLER_9_536 ();
 sg13g2_fill_8 FILLER_9_544 ();
 sg13g2_fill_8 FILLER_9_552 ();
 sg13g2_fill_8 FILLER_9_560 ();
 sg13g2_fill_8 FILLER_9_568 ();
 sg13g2_fill_8 FILLER_9_576 ();
 sg13g2_fill_8 FILLER_9_584 ();
 sg13g2_fill_8 FILLER_9_592 ();
 sg13g2_fill_8 FILLER_9_600 ();
 sg13g2_fill_8 FILLER_9_608 ();
 sg13g2_fill_8 FILLER_9_616 ();
 sg13g2_fill_8 FILLER_9_624 ();
 sg13g2_fill_8 FILLER_9_632 ();
 sg13g2_fill_8 FILLER_9_640 ();
 sg13g2_fill_4 FILLER_9_648 ();
 sg13g2_fill_4 FILLER_9_655 ();
 sg13g2_fill_1 FILLER_9_659 ();
 sg13g2_fill_2 FILLER_9_694 ();
 sg13g2_fill_1 FILLER_9_696 ();
 sg13g2_fill_2 FILLER_9_710 ();
 sg13g2_fill_8 FILLER_9_715 ();
 sg13g2_fill_8 FILLER_9_723 ();
 sg13g2_fill_8 FILLER_9_731 ();
 sg13g2_fill_8 FILLER_9_739 ();
 sg13g2_fill_4 FILLER_9_747 ();
 sg13g2_fill_2 FILLER_9_751 ();
 sg13g2_fill_8 FILLER_9_820 ();
 sg13g2_fill_2 FILLER_9_828 ();
 sg13g2_fill_1 FILLER_9_830 ();
 sg13g2_fill_8 FILLER_9_852 ();
 sg13g2_fill_8 FILLER_9_860 ();
 sg13g2_fill_4 FILLER_9_868 ();
 sg13g2_fill_2 FILLER_9_872 ();
 sg13g2_fill_1 FILLER_9_874 ();
 sg13g2_fill_8 FILLER_9_896 ();
 sg13g2_fill_8 FILLER_9_904 ();
 sg13g2_fill_1 FILLER_9_912 ();
 sg13g2_fill_8 FILLER_9_923 ();
 sg13g2_fill_8 FILLER_9_931 ();
 sg13g2_fill_8 FILLER_9_939 ();
 sg13g2_fill_4 FILLER_9_947 ();
 sg13g2_fill_2 FILLER_9_951 ();
 sg13g2_fill_8 FILLER_9_993 ();
 sg13g2_fill_8 FILLER_9_1001 ();
 sg13g2_fill_4 FILLER_9_1009 ();
 sg13g2_fill_1 FILLER_9_1013 ();
 sg13g2_fill_2 FILLER_9_1048 ();
 sg13g2_fill_1 FILLER_9_1050 ();
 sg13g2_fill_8 FILLER_9_1061 ();
 sg13g2_fill_4 FILLER_9_1069 ();
 sg13g2_fill_2 FILLER_9_1073 ();
 sg13g2_fill_8 FILLER_9_1090 ();
 sg13g2_fill_8 FILLER_9_1098 ();
 sg13g2_fill_2 FILLER_9_1111 ();
 sg13g2_fill_1 FILLER_9_1129 ();
 sg13g2_fill_8 FILLER_9_1160 ();
 sg13g2_fill_8 FILLER_9_1168 ();
 sg13g2_fill_8 FILLER_9_1176 ();
 sg13g2_fill_8 FILLER_9_1184 ();
 sg13g2_fill_8 FILLER_9_1192 ();
 sg13g2_fill_8 FILLER_9_1200 ();
 sg13g2_fill_8 FILLER_9_1208 ();
 sg13g2_fill_8 FILLER_9_1216 ();
 sg13g2_fill_8 FILLER_9_1224 ();
 sg13g2_fill_8 FILLER_9_1232 ();
 sg13g2_fill_8 FILLER_9_1240 ();
 sg13g2_fill_8 FILLER_9_1248 ();
 sg13g2_fill_8 FILLER_9_1256 ();
 sg13g2_fill_8 FILLER_9_1264 ();
 sg13g2_fill_8 FILLER_9_1272 ();
 sg13g2_fill_8 FILLER_9_1280 ();
 sg13g2_fill_8 FILLER_9_1288 ();
 sg13g2_fill_8 FILLER_9_1296 ();
 sg13g2_fill_8 FILLER_9_1304 ();
 sg13g2_fill_8 FILLER_9_1312 ();
 sg13g2_fill_8 FILLER_9_1320 ();
 sg13g2_fill_8 FILLER_9_1328 ();
 sg13g2_fill_8 FILLER_9_1336 ();
 sg13g2_fill_8 FILLER_9_1344 ();
 sg13g2_fill_8 FILLER_9_1352 ();
 sg13g2_fill_8 FILLER_9_1360 ();
 sg13g2_fill_8 FILLER_9_1368 ();
 sg13g2_fill_8 FILLER_9_1376 ();
 sg13g2_fill_8 FILLER_9_1384 ();
 sg13g2_fill_8 FILLER_9_1392 ();
 sg13g2_fill_8 FILLER_9_1400 ();
 sg13g2_fill_8 FILLER_9_1408 ();
 sg13g2_fill_8 FILLER_9_1416 ();
 sg13g2_fill_8 FILLER_9_1424 ();
 sg13g2_fill_8 FILLER_9_1432 ();
 sg13g2_fill_8 FILLER_9_1440 ();
 sg13g2_fill_8 FILLER_9_1448 ();
 sg13g2_fill_8 FILLER_9_1456 ();
 sg13g2_fill_8 FILLER_9_1464 ();
 sg13g2_fill_8 FILLER_9_1472 ();
 sg13g2_fill_8 FILLER_9_1480 ();
 sg13g2_fill_8 FILLER_9_1488 ();
 sg13g2_fill_8 FILLER_9_1496 ();
 sg13g2_fill_8 FILLER_9_1504 ();
 sg13g2_fill_8 FILLER_9_1512 ();
 sg13g2_fill_8 FILLER_9_1520 ();
 sg13g2_fill_8 FILLER_9_1528 ();
 sg13g2_fill_8 FILLER_9_1536 ();
 sg13g2_fill_8 FILLER_9_1544 ();
 sg13g2_fill_8 FILLER_9_1552 ();
 sg13g2_fill_8 FILLER_9_1560 ();
 sg13g2_fill_8 FILLER_9_1568 ();
 sg13g2_fill_8 FILLER_9_1576 ();
 sg13g2_fill_8 FILLER_9_1584 ();
 sg13g2_fill_8 FILLER_10_0 ();
 sg13g2_fill_8 FILLER_10_8 ();
 sg13g2_fill_8 FILLER_10_16 ();
 sg13g2_fill_8 FILLER_10_24 ();
 sg13g2_fill_8 FILLER_10_32 ();
 sg13g2_fill_8 FILLER_10_40 ();
 sg13g2_fill_8 FILLER_10_48 ();
 sg13g2_fill_8 FILLER_10_56 ();
 sg13g2_fill_8 FILLER_10_64 ();
 sg13g2_fill_8 FILLER_10_72 ();
 sg13g2_fill_8 FILLER_10_80 ();
 sg13g2_fill_8 FILLER_10_88 ();
 sg13g2_fill_8 FILLER_10_96 ();
 sg13g2_fill_8 FILLER_10_104 ();
 sg13g2_fill_8 FILLER_10_112 ();
 sg13g2_fill_8 FILLER_10_120 ();
 sg13g2_fill_8 FILLER_10_128 ();
 sg13g2_fill_8 FILLER_10_136 ();
 sg13g2_fill_8 FILLER_10_144 ();
 sg13g2_fill_8 FILLER_10_152 ();
 sg13g2_fill_8 FILLER_10_160 ();
 sg13g2_fill_8 FILLER_10_168 ();
 sg13g2_fill_8 FILLER_10_176 ();
 sg13g2_fill_8 FILLER_10_184 ();
 sg13g2_fill_8 FILLER_10_192 ();
 sg13g2_fill_8 FILLER_10_200 ();
 sg13g2_fill_8 FILLER_10_208 ();
 sg13g2_fill_8 FILLER_10_216 ();
 sg13g2_fill_8 FILLER_10_224 ();
 sg13g2_fill_8 FILLER_10_232 ();
 sg13g2_fill_8 FILLER_10_240 ();
 sg13g2_fill_8 FILLER_10_248 ();
 sg13g2_fill_8 FILLER_10_256 ();
 sg13g2_fill_8 FILLER_10_264 ();
 sg13g2_fill_8 FILLER_10_272 ();
 sg13g2_fill_8 FILLER_10_280 ();
 sg13g2_fill_8 FILLER_10_288 ();
 sg13g2_fill_8 FILLER_10_296 ();
 sg13g2_fill_8 FILLER_10_304 ();
 sg13g2_fill_8 FILLER_10_312 ();
 sg13g2_fill_8 FILLER_10_320 ();
 sg13g2_fill_8 FILLER_10_328 ();
 sg13g2_fill_8 FILLER_10_336 ();
 sg13g2_fill_8 FILLER_10_344 ();
 sg13g2_fill_8 FILLER_10_352 ();
 sg13g2_fill_8 FILLER_10_360 ();
 sg13g2_fill_8 FILLER_10_368 ();
 sg13g2_fill_8 FILLER_10_376 ();
 sg13g2_fill_8 FILLER_10_384 ();
 sg13g2_fill_8 FILLER_10_392 ();
 sg13g2_fill_8 FILLER_10_400 ();
 sg13g2_fill_8 FILLER_10_408 ();
 sg13g2_fill_8 FILLER_10_416 ();
 sg13g2_fill_8 FILLER_10_424 ();
 sg13g2_fill_8 FILLER_10_432 ();
 sg13g2_fill_8 FILLER_10_440 ();
 sg13g2_fill_8 FILLER_10_448 ();
 sg13g2_fill_8 FILLER_10_456 ();
 sg13g2_fill_8 FILLER_10_464 ();
 sg13g2_fill_8 FILLER_10_472 ();
 sg13g2_fill_8 FILLER_10_480 ();
 sg13g2_fill_8 FILLER_10_488 ();
 sg13g2_fill_8 FILLER_10_496 ();
 sg13g2_fill_8 FILLER_10_504 ();
 sg13g2_fill_8 FILLER_10_512 ();
 sg13g2_fill_8 FILLER_10_520 ();
 sg13g2_fill_8 FILLER_10_528 ();
 sg13g2_fill_8 FILLER_10_536 ();
 sg13g2_fill_8 FILLER_10_544 ();
 sg13g2_fill_8 FILLER_10_552 ();
 sg13g2_fill_8 FILLER_10_560 ();
 sg13g2_fill_8 FILLER_10_568 ();
 sg13g2_fill_8 FILLER_10_576 ();
 sg13g2_fill_8 FILLER_10_584 ();
 sg13g2_fill_8 FILLER_10_592 ();
 sg13g2_fill_8 FILLER_10_600 ();
 sg13g2_fill_8 FILLER_10_608 ();
 sg13g2_fill_8 FILLER_10_616 ();
 sg13g2_fill_8 FILLER_10_624 ();
 sg13g2_fill_8 FILLER_10_632 ();
 sg13g2_fill_4 FILLER_10_645 ();
 sg13g2_fill_2 FILLER_10_649 ();
 sg13g2_fill_1 FILLER_10_651 ();
 sg13g2_fill_8 FILLER_10_662 ();
 sg13g2_fill_1 FILLER_10_670 ();
 sg13g2_fill_8 FILLER_10_677 ();
 sg13g2_fill_8 FILLER_10_685 ();
 sg13g2_fill_4 FILLER_10_693 ();
 sg13g2_fill_1 FILLER_10_697 ();
 sg13g2_fill_1 FILLER_10_711 ();
 sg13g2_fill_1 FILLER_10_772 ();
 sg13g2_fill_8 FILLER_10_783 ();
 sg13g2_fill_8 FILLER_10_791 ();
 sg13g2_fill_8 FILLER_10_799 ();
 sg13g2_fill_8 FILLER_10_807 ();
 sg13g2_fill_8 FILLER_10_815 ();
 sg13g2_fill_8 FILLER_10_836 ();
 sg13g2_fill_8 FILLER_10_844 ();
 sg13g2_fill_4 FILLER_10_852 ();
 sg13g2_fill_1 FILLER_10_856 ();
 sg13g2_fill_8 FILLER_10_883 ();
 sg13g2_fill_1 FILLER_10_917 ();
 sg13g2_fill_8 FILLER_10_944 ();
 sg13g2_fill_8 FILLER_10_952 ();
 sg13g2_fill_2 FILLER_10_960 ();
 sg13g2_fill_2 FILLER_10_992 ();
 sg13g2_fill_1 FILLER_10_994 ();
 sg13g2_fill_8 FILLER_10_1025 ();
 sg13g2_fill_4 FILLER_10_1033 ();
 sg13g2_fill_2 FILLER_10_1037 ();
 sg13g2_fill_1 FILLER_10_1039 ();
 sg13g2_fill_4 FILLER_10_1076 ();
 sg13g2_fill_2 FILLER_10_1080 ();
 sg13g2_fill_1 FILLER_10_1082 ();
 sg13g2_fill_1 FILLER_10_1091 ();
 sg13g2_fill_2 FILLER_10_1114 ();
 sg13g2_fill_1 FILLER_10_1141 ();
 sg13g2_fill_8 FILLER_10_1152 ();
 sg13g2_fill_4 FILLER_10_1160 ();
 sg13g2_fill_1 FILLER_10_1164 ();
 sg13g2_fill_8 FILLER_10_1173 ();
 sg13g2_fill_8 FILLER_10_1181 ();
 sg13g2_fill_8 FILLER_10_1189 ();
 sg13g2_fill_8 FILLER_10_1197 ();
 sg13g2_fill_8 FILLER_10_1205 ();
 sg13g2_fill_8 FILLER_10_1213 ();
 sg13g2_fill_8 FILLER_10_1221 ();
 sg13g2_fill_8 FILLER_10_1229 ();
 sg13g2_fill_8 FILLER_10_1237 ();
 sg13g2_fill_8 FILLER_10_1245 ();
 sg13g2_fill_8 FILLER_10_1253 ();
 sg13g2_fill_8 FILLER_10_1261 ();
 sg13g2_fill_8 FILLER_10_1269 ();
 sg13g2_fill_8 FILLER_10_1277 ();
 sg13g2_fill_8 FILLER_10_1285 ();
 sg13g2_fill_8 FILLER_10_1293 ();
 sg13g2_fill_8 FILLER_10_1301 ();
 sg13g2_fill_8 FILLER_10_1309 ();
 sg13g2_fill_8 FILLER_10_1317 ();
 sg13g2_fill_8 FILLER_10_1325 ();
 sg13g2_fill_8 FILLER_10_1333 ();
 sg13g2_fill_8 FILLER_10_1341 ();
 sg13g2_fill_8 FILLER_10_1349 ();
 sg13g2_fill_8 FILLER_10_1357 ();
 sg13g2_fill_8 FILLER_10_1365 ();
 sg13g2_fill_8 FILLER_10_1373 ();
 sg13g2_fill_8 FILLER_10_1381 ();
 sg13g2_fill_8 FILLER_10_1389 ();
 sg13g2_fill_8 FILLER_10_1397 ();
 sg13g2_fill_8 FILLER_10_1405 ();
 sg13g2_fill_8 FILLER_10_1413 ();
 sg13g2_fill_8 FILLER_10_1421 ();
 sg13g2_fill_8 FILLER_10_1429 ();
 sg13g2_fill_8 FILLER_10_1437 ();
 sg13g2_fill_8 FILLER_10_1445 ();
 sg13g2_fill_8 FILLER_10_1453 ();
 sg13g2_fill_8 FILLER_10_1461 ();
 sg13g2_fill_8 FILLER_10_1469 ();
 sg13g2_fill_8 FILLER_10_1477 ();
 sg13g2_fill_8 FILLER_10_1485 ();
 sg13g2_fill_8 FILLER_10_1493 ();
 sg13g2_fill_8 FILLER_10_1501 ();
 sg13g2_fill_8 FILLER_10_1509 ();
 sg13g2_fill_8 FILLER_10_1517 ();
 sg13g2_fill_8 FILLER_10_1525 ();
 sg13g2_fill_8 FILLER_10_1533 ();
 sg13g2_fill_8 FILLER_10_1541 ();
 sg13g2_fill_8 FILLER_10_1549 ();
 sg13g2_fill_8 FILLER_10_1557 ();
 sg13g2_fill_8 FILLER_10_1565 ();
 sg13g2_fill_8 FILLER_10_1573 ();
 sg13g2_fill_8 FILLER_10_1581 ();
 sg13g2_fill_2 FILLER_10_1589 ();
 sg13g2_fill_1 FILLER_10_1591 ();
 sg13g2_fill_8 FILLER_11_0 ();
 sg13g2_fill_8 FILLER_11_8 ();
 sg13g2_fill_8 FILLER_11_16 ();
 sg13g2_fill_8 FILLER_11_24 ();
 sg13g2_fill_8 FILLER_11_32 ();
 sg13g2_fill_8 FILLER_11_40 ();
 sg13g2_fill_8 FILLER_11_48 ();
 sg13g2_fill_8 FILLER_11_56 ();
 sg13g2_fill_8 FILLER_11_64 ();
 sg13g2_fill_8 FILLER_11_72 ();
 sg13g2_fill_8 FILLER_11_80 ();
 sg13g2_fill_8 FILLER_11_88 ();
 sg13g2_fill_8 FILLER_11_96 ();
 sg13g2_fill_8 FILLER_11_104 ();
 sg13g2_fill_8 FILLER_11_112 ();
 sg13g2_fill_8 FILLER_11_120 ();
 sg13g2_fill_8 FILLER_11_128 ();
 sg13g2_fill_8 FILLER_11_136 ();
 sg13g2_fill_8 FILLER_11_144 ();
 sg13g2_fill_8 FILLER_11_152 ();
 sg13g2_fill_8 FILLER_11_160 ();
 sg13g2_fill_8 FILLER_11_168 ();
 sg13g2_fill_8 FILLER_11_176 ();
 sg13g2_fill_8 FILLER_11_184 ();
 sg13g2_fill_8 FILLER_11_192 ();
 sg13g2_fill_8 FILLER_11_200 ();
 sg13g2_fill_8 FILLER_11_208 ();
 sg13g2_fill_8 FILLER_11_216 ();
 sg13g2_fill_8 FILLER_11_224 ();
 sg13g2_fill_8 FILLER_11_232 ();
 sg13g2_fill_8 FILLER_11_240 ();
 sg13g2_fill_8 FILLER_11_248 ();
 sg13g2_fill_8 FILLER_11_256 ();
 sg13g2_fill_8 FILLER_11_264 ();
 sg13g2_fill_8 FILLER_11_272 ();
 sg13g2_fill_8 FILLER_11_280 ();
 sg13g2_fill_8 FILLER_11_288 ();
 sg13g2_fill_8 FILLER_11_296 ();
 sg13g2_fill_8 FILLER_11_304 ();
 sg13g2_fill_8 FILLER_11_312 ();
 sg13g2_fill_8 FILLER_11_320 ();
 sg13g2_fill_8 FILLER_11_328 ();
 sg13g2_fill_8 FILLER_11_336 ();
 sg13g2_fill_8 FILLER_11_344 ();
 sg13g2_fill_8 FILLER_11_352 ();
 sg13g2_fill_8 FILLER_11_360 ();
 sg13g2_fill_8 FILLER_11_368 ();
 sg13g2_fill_8 FILLER_11_376 ();
 sg13g2_fill_8 FILLER_11_384 ();
 sg13g2_fill_8 FILLER_11_392 ();
 sg13g2_fill_8 FILLER_11_400 ();
 sg13g2_fill_8 FILLER_11_408 ();
 sg13g2_fill_8 FILLER_11_416 ();
 sg13g2_fill_8 FILLER_11_424 ();
 sg13g2_fill_8 FILLER_11_432 ();
 sg13g2_fill_8 FILLER_11_440 ();
 sg13g2_fill_8 FILLER_11_448 ();
 sg13g2_fill_8 FILLER_11_456 ();
 sg13g2_fill_8 FILLER_11_464 ();
 sg13g2_fill_8 FILLER_11_472 ();
 sg13g2_fill_8 FILLER_11_480 ();
 sg13g2_fill_8 FILLER_11_488 ();
 sg13g2_fill_8 FILLER_11_496 ();
 sg13g2_fill_8 FILLER_11_504 ();
 sg13g2_fill_8 FILLER_11_512 ();
 sg13g2_fill_8 FILLER_11_520 ();
 sg13g2_fill_8 FILLER_11_528 ();
 sg13g2_fill_8 FILLER_11_536 ();
 sg13g2_fill_8 FILLER_11_544 ();
 sg13g2_fill_8 FILLER_11_552 ();
 sg13g2_fill_8 FILLER_11_560 ();
 sg13g2_fill_8 FILLER_11_568 ();
 sg13g2_fill_8 FILLER_11_576 ();
 sg13g2_fill_8 FILLER_11_584 ();
 sg13g2_fill_8 FILLER_11_592 ();
 sg13g2_fill_8 FILLER_11_600 ();
 sg13g2_fill_8 FILLER_11_608 ();
 sg13g2_fill_2 FILLER_11_616 ();
 sg13g2_fill_2 FILLER_11_644 ();
 sg13g2_fill_1 FILLER_11_646 ();
 sg13g2_fill_1 FILLER_11_663 ();
 sg13g2_fill_1 FILLER_11_677 ();
 sg13g2_fill_1 FILLER_11_708 ();
 sg13g2_fill_8 FILLER_11_739 ();
 sg13g2_fill_1 FILLER_11_747 ();
 sg13g2_fill_8 FILLER_11_774 ();
 sg13g2_fill_2 FILLER_11_782 ();
 sg13g2_fill_8 FILLER_11_809 ();
 sg13g2_fill_4 FILLER_11_843 ();
 sg13g2_fill_2 FILLER_11_847 ();
 sg13g2_fill_8 FILLER_11_854 ();
 sg13g2_fill_8 FILLER_11_862 ();
 sg13g2_fill_4 FILLER_11_870 ();
 sg13g2_fill_2 FILLER_11_874 ();
 sg13g2_fill_1 FILLER_11_876 ();
 sg13g2_fill_2 FILLER_11_897 ();
 sg13g2_fill_8 FILLER_11_909 ();
 sg13g2_fill_8 FILLER_11_917 ();
 sg13g2_fill_4 FILLER_11_925 ();
 sg13g2_fill_4 FILLER_11_980 ();
 sg13g2_fill_4 FILLER_11_989 ();
 sg13g2_fill_2 FILLER_11_993 ();
 sg13g2_fill_8 FILLER_11_1005 ();
 sg13g2_fill_2 FILLER_11_1013 ();
 sg13g2_fill_1 FILLER_11_1015 ();
 sg13g2_fill_8 FILLER_11_1024 ();
 sg13g2_fill_8 FILLER_11_1032 ();
 sg13g2_fill_8 FILLER_11_1040 ();
 sg13g2_fill_8 FILLER_11_1048 ();
 sg13g2_fill_4 FILLER_11_1056 ();
 sg13g2_fill_2 FILLER_11_1060 ();
 sg13g2_fill_2 FILLER_11_1086 ();
 sg13g2_fill_1 FILLER_11_1094 ();
 sg13g2_fill_2 FILLER_11_1100 ();
 sg13g2_fill_1 FILLER_11_1102 ();
 sg13g2_fill_1 FILLER_11_1111 ();
 sg13g2_fill_8 FILLER_11_1183 ();
 sg13g2_fill_8 FILLER_11_1191 ();
 sg13g2_fill_8 FILLER_11_1199 ();
 sg13g2_fill_8 FILLER_11_1207 ();
 sg13g2_fill_8 FILLER_11_1215 ();
 sg13g2_fill_8 FILLER_11_1223 ();
 sg13g2_fill_8 FILLER_11_1231 ();
 sg13g2_fill_8 FILLER_11_1239 ();
 sg13g2_fill_8 FILLER_11_1247 ();
 sg13g2_fill_8 FILLER_11_1255 ();
 sg13g2_fill_8 FILLER_11_1263 ();
 sg13g2_fill_8 FILLER_11_1271 ();
 sg13g2_fill_8 FILLER_11_1279 ();
 sg13g2_fill_8 FILLER_11_1287 ();
 sg13g2_fill_8 FILLER_11_1295 ();
 sg13g2_fill_8 FILLER_11_1303 ();
 sg13g2_fill_8 FILLER_11_1311 ();
 sg13g2_fill_8 FILLER_11_1319 ();
 sg13g2_fill_8 FILLER_11_1327 ();
 sg13g2_fill_8 FILLER_11_1335 ();
 sg13g2_fill_8 FILLER_11_1343 ();
 sg13g2_fill_8 FILLER_11_1351 ();
 sg13g2_fill_8 FILLER_11_1359 ();
 sg13g2_fill_8 FILLER_11_1367 ();
 sg13g2_fill_8 FILLER_11_1375 ();
 sg13g2_fill_8 FILLER_11_1383 ();
 sg13g2_fill_8 FILLER_11_1391 ();
 sg13g2_fill_8 FILLER_11_1399 ();
 sg13g2_fill_8 FILLER_11_1407 ();
 sg13g2_fill_8 FILLER_11_1415 ();
 sg13g2_fill_8 FILLER_11_1423 ();
 sg13g2_fill_8 FILLER_11_1431 ();
 sg13g2_fill_8 FILLER_11_1439 ();
 sg13g2_fill_8 FILLER_11_1447 ();
 sg13g2_fill_8 FILLER_11_1455 ();
 sg13g2_fill_8 FILLER_11_1463 ();
 sg13g2_fill_8 FILLER_11_1471 ();
 sg13g2_fill_8 FILLER_11_1479 ();
 sg13g2_fill_8 FILLER_11_1487 ();
 sg13g2_fill_8 FILLER_11_1495 ();
 sg13g2_fill_8 FILLER_11_1503 ();
 sg13g2_fill_8 FILLER_11_1511 ();
 sg13g2_fill_8 FILLER_11_1519 ();
 sg13g2_fill_8 FILLER_11_1527 ();
 sg13g2_fill_8 FILLER_11_1535 ();
 sg13g2_fill_8 FILLER_11_1543 ();
 sg13g2_fill_8 FILLER_11_1551 ();
 sg13g2_fill_8 FILLER_11_1559 ();
 sg13g2_fill_8 FILLER_11_1567 ();
 sg13g2_fill_8 FILLER_11_1575 ();
 sg13g2_fill_8 FILLER_11_1583 ();
 sg13g2_fill_1 FILLER_11_1591 ();
 sg13g2_fill_8 FILLER_12_0 ();
 sg13g2_fill_8 FILLER_12_8 ();
 sg13g2_fill_8 FILLER_12_16 ();
 sg13g2_fill_8 FILLER_12_24 ();
 sg13g2_fill_8 FILLER_12_32 ();
 sg13g2_fill_8 FILLER_12_40 ();
 sg13g2_fill_8 FILLER_12_48 ();
 sg13g2_fill_8 FILLER_12_56 ();
 sg13g2_fill_8 FILLER_12_64 ();
 sg13g2_fill_8 FILLER_12_72 ();
 sg13g2_fill_8 FILLER_12_80 ();
 sg13g2_fill_8 FILLER_12_88 ();
 sg13g2_fill_8 FILLER_12_96 ();
 sg13g2_fill_8 FILLER_12_104 ();
 sg13g2_fill_8 FILLER_12_112 ();
 sg13g2_fill_8 FILLER_12_120 ();
 sg13g2_fill_8 FILLER_12_128 ();
 sg13g2_fill_8 FILLER_12_136 ();
 sg13g2_fill_8 FILLER_12_144 ();
 sg13g2_fill_8 FILLER_12_152 ();
 sg13g2_fill_8 FILLER_12_160 ();
 sg13g2_fill_8 FILLER_12_168 ();
 sg13g2_fill_8 FILLER_12_176 ();
 sg13g2_fill_8 FILLER_12_184 ();
 sg13g2_fill_8 FILLER_12_192 ();
 sg13g2_fill_8 FILLER_12_200 ();
 sg13g2_fill_8 FILLER_12_208 ();
 sg13g2_fill_8 FILLER_12_216 ();
 sg13g2_fill_8 FILLER_12_224 ();
 sg13g2_fill_8 FILLER_12_232 ();
 sg13g2_fill_8 FILLER_12_240 ();
 sg13g2_fill_8 FILLER_12_248 ();
 sg13g2_fill_8 FILLER_12_256 ();
 sg13g2_fill_8 FILLER_12_264 ();
 sg13g2_fill_8 FILLER_12_272 ();
 sg13g2_fill_8 FILLER_12_280 ();
 sg13g2_fill_8 FILLER_12_288 ();
 sg13g2_fill_8 FILLER_12_296 ();
 sg13g2_fill_8 FILLER_12_304 ();
 sg13g2_fill_8 FILLER_12_312 ();
 sg13g2_fill_8 FILLER_12_320 ();
 sg13g2_fill_8 FILLER_12_328 ();
 sg13g2_fill_8 FILLER_12_336 ();
 sg13g2_fill_8 FILLER_12_344 ();
 sg13g2_fill_8 FILLER_12_352 ();
 sg13g2_fill_8 FILLER_12_360 ();
 sg13g2_fill_8 FILLER_12_368 ();
 sg13g2_fill_8 FILLER_12_376 ();
 sg13g2_fill_8 FILLER_12_384 ();
 sg13g2_fill_8 FILLER_12_392 ();
 sg13g2_fill_8 FILLER_12_400 ();
 sg13g2_fill_8 FILLER_12_408 ();
 sg13g2_fill_8 FILLER_12_416 ();
 sg13g2_fill_8 FILLER_12_424 ();
 sg13g2_fill_8 FILLER_12_432 ();
 sg13g2_fill_8 FILLER_12_440 ();
 sg13g2_fill_8 FILLER_12_448 ();
 sg13g2_fill_8 FILLER_12_456 ();
 sg13g2_fill_8 FILLER_12_464 ();
 sg13g2_fill_8 FILLER_12_472 ();
 sg13g2_fill_8 FILLER_12_480 ();
 sg13g2_fill_8 FILLER_12_488 ();
 sg13g2_fill_8 FILLER_12_496 ();
 sg13g2_fill_8 FILLER_12_504 ();
 sg13g2_fill_8 FILLER_12_512 ();
 sg13g2_fill_8 FILLER_12_520 ();
 sg13g2_fill_8 FILLER_12_528 ();
 sg13g2_fill_8 FILLER_12_536 ();
 sg13g2_fill_8 FILLER_12_544 ();
 sg13g2_fill_8 FILLER_12_552 ();
 sg13g2_fill_8 FILLER_12_560 ();
 sg13g2_fill_8 FILLER_12_568 ();
 sg13g2_fill_8 FILLER_12_576 ();
 sg13g2_fill_8 FILLER_12_584 ();
 sg13g2_fill_8 FILLER_12_608 ();
 sg13g2_fill_8 FILLER_12_616 ();
 sg13g2_fill_4 FILLER_12_624 ();
 sg13g2_fill_2 FILLER_12_628 ();
 sg13g2_fill_2 FILLER_12_659 ();
 sg13g2_fill_1 FILLER_12_661 ();
 sg13g2_fill_8 FILLER_12_703 ();
 sg13g2_fill_1 FILLER_12_711 ();
 sg13g2_fill_8 FILLER_12_715 ();
 sg13g2_fill_8 FILLER_12_723 ();
 sg13g2_fill_8 FILLER_12_731 ();
 sg13g2_fill_8 FILLER_12_739 ();
 sg13g2_fill_4 FILLER_12_747 ();
 sg13g2_fill_8 FILLER_12_776 ();
 sg13g2_fill_1 FILLER_12_815 ();
 sg13g2_fill_8 FILLER_12_826 ();
 sg13g2_fill_8 FILLER_12_834 ();
 sg13g2_fill_2 FILLER_12_842 ();
 sg13g2_fill_8 FILLER_12_870 ();
 sg13g2_fill_8 FILLER_12_878 ();
 sg13g2_fill_4 FILLER_12_886 ();
 sg13g2_fill_2 FILLER_12_890 ();
 sg13g2_fill_1 FILLER_12_892 ();
 sg13g2_fill_1 FILLER_12_940 ();
 sg13g2_fill_8 FILLER_12_951 ();
 sg13g2_fill_4 FILLER_12_965 ();
 sg13g2_fill_1 FILLER_12_978 ();
 sg13g2_fill_4 FILLER_12_1005 ();
 sg13g2_fill_2 FILLER_12_1009 ();
 sg13g2_fill_1 FILLER_12_1011 ();
 sg13g2_fill_4 FILLER_12_1022 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_8 FILLER_12_1062 ();
 sg13g2_fill_2 FILLER_12_1070 ();
 sg13g2_fill_2 FILLER_12_1080 ();
 sg13g2_fill_1 FILLER_12_1082 ();
 sg13g2_fill_2 FILLER_12_1127 ();
 sg13g2_fill_1 FILLER_12_1163 ();
 sg13g2_fill_8 FILLER_12_1196 ();
 sg13g2_fill_8 FILLER_12_1204 ();
 sg13g2_fill_8 FILLER_12_1212 ();
 sg13g2_fill_8 FILLER_12_1220 ();
 sg13g2_fill_8 FILLER_12_1228 ();
 sg13g2_fill_8 FILLER_12_1236 ();
 sg13g2_fill_8 FILLER_12_1244 ();
 sg13g2_fill_8 FILLER_12_1252 ();
 sg13g2_fill_8 FILLER_12_1260 ();
 sg13g2_fill_8 FILLER_12_1268 ();
 sg13g2_fill_8 FILLER_12_1276 ();
 sg13g2_fill_8 FILLER_12_1284 ();
 sg13g2_fill_8 FILLER_12_1292 ();
 sg13g2_fill_8 FILLER_12_1300 ();
 sg13g2_fill_8 FILLER_12_1308 ();
 sg13g2_fill_8 FILLER_12_1316 ();
 sg13g2_fill_8 FILLER_12_1324 ();
 sg13g2_fill_8 FILLER_12_1332 ();
 sg13g2_fill_8 FILLER_12_1340 ();
 sg13g2_fill_8 FILLER_12_1348 ();
 sg13g2_fill_8 FILLER_12_1356 ();
 sg13g2_fill_8 FILLER_12_1364 ();
 sg13g2_fill_8 FILLER_12_1372 ();
 sg13g2_fill_8 FILLER_12_1380 ();
 sg13g2_fill_8 FILLER_12_1388 ();
 sg13g2_fill_8 FILLER_12_1396 ();
 sg13g2_fill_8 FILLER_12_1404 ();
 sg13g2_fill_8 FILLER_12_1412 ();
 sg13g2_fill_8 FILLER_12_1420 ();
 sg13g2_fill_8 FILLER_12_1428 ();
 sg13g2_fill_8 FILLER_12_1436 ();
 sg13g2_fill_8 FILLER_12_1444 ();
 sg13g2_fill_8 FILLER_12_1452 ();
 sg13g2_fill_8 FILLER_12_1460 ();
 sg13g2_fill_8 FILLER_12_1468 ();
 sg13g2_fill_8 FILLER_12_1476 ();
 sg13g2_fill_8 FILLER_12_1484 ();
 sg13g2_fill_8 FILLER_12_1492 ();
 sg13g2_fill_8 FILLER_12_1500 ();
 sg13g2_fill_8 FILLER_12_1508 ();
 sg13g2_fill_8 FILLER_12_1516 ();
 sg13g2_fill_8 FILLER_12_1524 ();
 sg13g2_fill_8 FILLER_12_1532 ();
 sg13g2_fill_8 FILLER_12_1540 ();
 sg13g2_fill_8 FILLER_12_1548 ();
 sg13g2_fill_8 FILLER_12_1556 ();
 sg13g2_fill_8 FILLER_12_1564 ();
 sg13g2_fill_8 FILLER_12_1572 ();
 sg13g2_fill_8 FILLER_12_1580 ();
 sg13g2_fill_4 FILLER_12_1588 ();
 sg13g2_fill_8 FILLER_13_0 ();
 sg13g2_fill_8 FILLER_13_8 ();
 sg13g2_fill_8 FILLER_13_16 ();
 sg13g2_fill_8 FILLER_13_24 ();
 sg13g2_fill_8 FILLER_13_32 ();
 sg13g2_fill_8 FILLER_13_40 ();
 sg13g2_fill_8 FILLER_13_48 ();
 sg13g2_fill_8 FILLER_13_56 ();
 sg13g2_fill_8 FILLER_13_64 ();
 sg13g2_fill_8 FILLER_13_72 ();
 sg13g2_fill_8 FILLER_13_80 ();
 sg13g2_fill_8 FILLER_13_88 ();
 sg13g2_fill_8 FILLER_13_96 ();
 sg13g2_fill_8 FILLER_13_104 ();
 sg13g2_fill_8 FILLER_13_112 ();
 sg13g2_fill_8 FILLER_13_120 ();
 sg13g2_fill_8 FILLER_13_128 ();
 sg13g2_fill_8 FILLER_13_136 ();
 sg13g2_fill_8 FILLER_13_144 ();
 sg13g2_fill_8 FILLER_13_152 ();
 sg13g2_fill_8 FILLER_13_160 ();
 sg13g2_fill_8 FILLER_13_168 ();
 sg13g2_fill_8 FILLER_13_176 ();
 sg13g2_fill_8 FILLER_13_184 ();
 sg13g2_fill_8 FILLER_13_192 ();
 sg13g2_fill_8 FILLER_13_200 ();
 sg13g2_fill_8 FILLER_13_208 ();
 sg13g2_fill_8 FILLER_13_216 ();
 sg13g2_fill_8 FILLER_13_224 ();
 sg13g2_fill_8 FILLER_13_232 ();
 sg13g2_fill_8 FILLER_13_240 ();
 sg13g2_fill_8 FILLER_13_248 ();
 sg13g2_fill_8 FILLER_13_256 ();
 sg13g2_fill_8 FILLER_13_264 ();
 sg13g2_fill_8 FILLER_13_272 ();
 sg13g2_fill_8 FILLER_13_280 ();
 sg13g2_fill_8 FILLER_13_288 ();
 sg13g2_fill_8 FILLER_13_296 ();
 sg13g2_fill_8 FILLER_13_304 ();
 sg13g2_fill_8 FILLER_13_312 ();
 sg13g2_fill_8 FILLER_13_320 ();
 sg13g2_fill_8 FILLER_13_328 ();
 sg13g2_fill_8 FILLER_13_336 ();
 sg13g2_fill_8 FILLER_13_344 ();
 sg13g2_fill_8 FILLER_13_352 ();
 sg13g2_fill_8 FILLER_13_360 ();
 sg13g2_fill_8 FILLER_13_368 ();
 sg13g2_fill_8 FILLER_13_376 ();
 sg13g2_fill_8 FILLER_13_384 ();
 sg13g2_fill_8 FILLER_13_392 ();
 sg13g2_fill_8 FILLER_13_400 ();
 sg13g2_fill_8 FILLER_13_408 ();
 sg13g2_fill_8 FILLER_13_416 ();
 sg13g2_fill_4 FILLER_13_424 ();
 sg13g2_fill_1 FILLER_13_428 ();
 sg13g2_fill_4 FILLER_13_439 ();
 sg13g2_fill_8 FILLER_13_453 ();
 sg13g2_fill_8 FILLER_13_461 ();
 sg13g2_fill_8 FILLER_13_469 ();
 sg13g2_fill_8 FILLER_13_477 ();
 sg13g2_fill_8 FILLER_13_485 ();
 sg13g2_fill_8 FILLER_13_493 ();
 sg13g2_fill_8 FILLER_13_537 ();
 sg13g2_fill_8 FILLER_13_545 ();
 sg13g2_fill_8 FILLER_13_553 ();
 sg13g2_fill_8 FILLER_13_561 ();
 sg13g2_fill_8 FILLER_13_569 ();
 sg13g2_fill_8 FILLER_13_577 ();
 sg13g2_fill_8 FILLER_13_585 ();
 sg13g2_fill_8 FILLER_13_623 ();
 sg13g2_fill_8 FILLER_13_631 ();
 sg13g2_fill_4 FILLER_13_639 ();
 sg13g2_fill_2 FILLER_13_643 ();
 sg13g2_fill_8 FILLER_13_679 ();
 sg13g2_fill_8 FILLER_13_687 ();
 sg13g2_fill_8 FILLER_13_695 ();
 sg13g2_fill_8 FILLER_13_703 ();
 sg13g2_fill_2 FILLER_13_732 ();
 sg13g2_fill_1 FILLER_13_739 ();
 sg13g2_fill_8 FILLER_13_786 ();
 sg13g2_fill_8 FILLER_13_794 ();
 sg13g2_fill_8 FILLER_13_802 ();
 sg13g2_fill_1 FILLER_13_810 ();
 sg13g2_fill_1 FILLER_13_837 ();
 sg13g2_fill_4 FILLER_13_863 ();
 sg13g2_fill_8 FILLER_13_893 ();
 sg13g2_fill_8 FILLER_13_901 ();
 sg13g2_fill_2 FILLER_13_909 ();
 sg13g2_fill_1 FILLER_13_911 ();
 sg13g2_fill_2 FILLER_13_940 ();
 sg13g2_fill_1 FILLER_13_942 ();
 sg13g2_fill_1 FILLER_13_953 ();
 sg13g2_fill_1 FILLER_13_974 ();
 sg13g2_fill_8 FILLER_13_994 ();
 sg13g2_fill_8 FILLER_13_1002 ();
 sg13g2_fill_2 FILLER_13_1010 ();
 sg13g2_fill_1 FILLER_13_1063 ();
 sg13g2_fill_8 FILLER_13_1069 ();
 sg13g2_fill_8 FILLER_13_1077 ();
 sg13g2_fill_8 FILLER_13_1085 ();
 sg13g2_fill_8 FILLER_13_1093 ();
 sg13g2_fill_8 FILLER_13_1101 ();
 sg13g2_fill_8 FILLER_13_1109 ();
 sg13g2_fill_1 FILLER_13_1117 ();
 sg13g2_fill_8 FILLER_13_1183 ();
 sg13g2_fill_8 FILLER_13_1191 ();
 sg13g2_fill_8 FILLER_13_1199 ();
 sg13g2_fill_8 FILLER_13_1207 ();
 sg13g2_fill_8 FILLER_13_1215 ();
 sg13g2_fill_8 FILLER_13_1223 ();
 sg13g2_fill_8 FILLER_13_1231 ();
 sg13g2_fill_8 FILLER_13_1239 ();
 sg13g2_fill_8 FILLER_13_1247 ();
 sg13g2_fill_8 FILLER_13_1255 ();
 sg13g2_fill_8 FILLER_13_1263 ();
 sg13g2_fill_8 FILLER_13_1271 ();
 sg13g2_fill_8 FILLER_13_1279 ();
 sg13g2_fill_8 FILLER_13_1287 ();
 sg13g2_fill_8 FILLER_13_1295 ();
 sg13g2_fill_8 FILLER_13_1303 ();
 sg13g2_fill_8 FILLER_13_1311 ();
 sg13g2_fill_8 FILLER_13_1319 ();
 sg13g2_fill_8 FILLER_13_1327 ();
 sg13g2_fill_8 FILLER_13_1335 ();
 sg13g2_fill_8 FILLER_13_1343 ();
 sg13g2_fill_8 FILLER_13_1351 ();
 sg13g2_fill_8 FILLER_13_1359 ();
 sg13g2_fill_8 FILLER_13_1367 ();
 sg13g2_fill_8 FILLER_13_1375 ();
 sg13g2_fill_8 FILLER_13_1383 ();
 sg13g2_fill_8 FILLER_13_1391 ();
 sg13g2_fill_8 FILLER_13_1399 ();
 sg13g2_fill_8 FILLER_13_1407 ();
 sg13g2_fill_8 FILLER_13_1415 ();
 sg13g2_fill_8 FILLER_13_1423 ();
 sg13g2_fill_8 FILLER_13_1431 ();
 sg13g2_fill_8 FILLER_13_1439 ();
 sg13g2_fill_8 FILLER_13_1447 ();
 sg13g2_fill_8 FILLER_13_1455 ();
 sg13g2_fill_8 FILLER_13_1463 ();
 sg13g2_fill_8 FILLER_13_1471 ();
 sg13g2_fill_8 FILLER_13_1479 ();
 sg13g2_fill_8 FILLER_13_1487 ();
 sg13g2_fill_8 FILLER_13_1495 ();
 sg13g2_fill_8 FILLER_13_1503 ();
 sg13g2_fill_8 FILLER_13_1511 ();
 sg13g2_fill_8 FILLER_13_1519 ();
 sg13g2_fill_8 FILLER_13_1527 ();
 sg13g2_fill_8 FILLER_13_1535 ();
 sg13g2_fill_8 FILLER_13_1543 ();
 sg13g2_fill_8 FILLER_13_1551 ();
 sg13g2_fill_8 FILLER_13_1559 ();
 sg13g2_fill_8 FILLER_13_1567 ();
 sg13g2_fill_8 FILLER_13_1575 ();
 sg13g2_fill_8 FILLER_13_1583 ();
 sg13g2_fill_1 FILLER_13_1591 ();
 sg13g2_fill_8 FILLER_14_0 ();
 sg13g2_fill_8 FILLER_14_8 ();
 sg13g2_fill_8 FILLER_14_16 ();
 sg13g2_fill_8 FILLER_14_24 ();
 sg13g2_fill_8 FILLER_14_32 ();
 sg13g2_fill_8 FILLER_14_40 ();
 sg13g2_fill_8 FILLER_14_48 ();
 sg13g2_fill_8 FILLER_14_56 ();
 sg13g2_fill_8 FILLER_14_64 ();
 sg13g2_fill_8 FILLER_14_72 ();
 sg13g2_fill_8 FILLER_14_80 ();
 sg13g2_fill_8 FILLER_14_88 ();
 sg13g2_fill_8 FILLER_14_96 ();
 sg13g2_fill_8 FILLER_14_104 ();
 sg13g2_fill_8 FILLER_14_112 ();
 sg13g2_fill_8 FILLER_14_120 ();
 sg13g2_fill_8 FILLER_14_128 ();
 sg13g2_fill_8 FILLER_14_136 ();
 sg13g2_fill_8 FILLER_14_144 ();
 sg13g2_fill_8 FILLER_14_152 ();
 sg13g2_fill_8 FILLER_14_160 ();
 sg13g2_fill_8 FILLER_14_168 ();
 sg13g2_fill_8 FILLER_14_176 ();
 sg13g2_fill_8 FILLER_14_184 ();
 sg13g2_fill_8 FILLER_14_192 ();
 sg13g2_fill_8 FILLER_14_200 ();
 sg13g2_fill_8 FILLER_14_208 ();
 sg13g2_fill_8 FILLER_14_216 ();
 sg13g2_fill_8 FILLER_14_224 ();
 sg13g2_fill_8 FILLER_14_232 ();
 sg13g2_fill_8 FILLER_14_240 ();
 sg13g2_fill_8 FILLER_14_248 ();
 sg13g2_fill_8 FILLER_14_256 ();
 sg13g2_fill_8 FILLER_14_264 ();
 sg13g2_fill_8 FILLER_14_272 ();
 sg13g2_fill_8 FILLER_14_280 ();
 sg13g2_fill_8 FILLER_14_288 ();
 sg13g2_fill_8 FILLER_14_296 ();
 sg13g2_fill_8 FILLER_14_304 ();
 sg13g2_fill_8 FILLER_14_312 ();
 sg13g2_fill_8 FILLER_14_320 ();
 sg13g2_fill_8 FILLER_14_328 ();
 sg13g2_fill_8 FILLER_14_336 ();
 sg13g2_fill_8 FILLER_14_344 ();
 sg13g2_fill_8 FILLER_14_352 ();
 sg13g2_fill_8 FILLER_14_360 ();
 sg13g2_fill_8 FILLER_14_368 ();
 sg13g2_fill_8 FILLER_14_376 ();
 sg13g2_fill_8 FILLER_14_384 ();
 sg13g2_fill_8 FILLER_14_392 ();
 sg13g2_fill_8 FILLER_14_400 ();
 sg13g2_fill_8 FILLER_14_408 ();
 sg13g2_fill_8 FILLER_14_416 ();
 sg13g2_fill_8 FILLER_14_476 ();
 sg13g2_fill_4 FILLER_14_519 ();
 sg13g2_fill_8 FILLER_14_549 ();
 sg13g2_fill_8 FILLER_14_557 ();
 sg13g2_fill_8 FILLER_14_565 ();
 sg13g2_fill_8 FILLER_14_573 ();
 sg13g2_fill_8 FILLER_14_581 ();
 sg13g2_fill_8 FILLER_14_589 ();
 sg13g2_fill_8 FILLER_14_597 ();
 sg13g2_fill_8 FILLER_14_605 ();
 sg13g2_fill_4 FILLER_14_613 ();
 sg13g2_fill_2 FILLER_14_617 ();
 sg13g2_fill_1 FILLER_14_619 ();
 sg13g2_fill_2 FILLER_14_646 ();
 sg13g2_fill_2 FILLER_14_651 ();
 sg13g2_fill_4 FILLER_14_672 ();
 sg13g2_fill_2 FILLER_14_676 ();
 sg13g2_fill_1 FILLER_14_678 ();
 sg13g2_fill_4 FILLER_14_705 ();
 sg13g2_fill_2 FILLER_14_722 ();
 sg13g2_fill_1 FILLER_14_724 ();
 sg13g2_fill_2 FILLER_14_769 ();
 sg13g2_fill_2 FILLER_14_807 ();
 sg13g2_fill_1 FILLER_14_827 ();
 sg13g2_fill_2 FILLER_14_869 ();
 sg13g2_fill_8 FILLER_14_892 ();
 sg13g2_fill_1 FILLER_14_900 ();
 sg13g2_fill_8 FILLER_14_908 ();
 sg13g2_fill_8 FILLER_14_960 ();
 sg13g2_fill_1 FILLER_14_968 ();
 sg13g2_fill_2 FILLER_14_974 ();
 sg13g2_fill_8 FILLER_14_986 ();
 sg13g2_fill_4 FILLER_14_994 ();
 sg13g2_fill_1 FILLER_14_998 ();
 sg13g2_fill_8 FILLER_14_1008 ();
 sg13g2_fill_8 FILLER_14_1016 ();
 sg13g2_fill_8 FILLER_14_1024 ();
 sg13g2_fill_4 FILLER_14_1032 ();
 sg13g2_fill_2 FILLER_14_1036 ();
 sg13g2_fill_1 FILLER_14_1058 ();
 sg13g2_fill_4 FILLER_14_1095 ();
 sg13g2_fill_2 FILLER_14_1099 ();
 sg13g2_fill_1 FILLER_14_1135 ();
 sg13g2_fill_8 FILLER_14_1141 ();
 sg13g2_fill_8 FILLER_14_1149 ();
 sg13g2_fill_2 FILLER_14_1157 ();
 sg13g2_fill_2 FILLER_14_1173 ();
 sg13g2_fill_1 FILLER_14_1175 ();
 sg13g2_fill_8 FILLER_14_1202 ();
 sg13g2_fill_1 FILLER_14_1210 ();
 sg13g2_fill_8 FILLER_14_1244 ();
 sg13g2_fill_8 FILLER_14_1252 ();
 sg13g2_fill_8 FILLER_14_1260 ();
 sg13g2_fill_8 FILLER_14_1268 ();
 sg13g2_fill_8 FILLER_14_1276 ();
 sg13g2_fill_8 FILLER_14_1284 ();
 sg13g2_fill_8 FILLER_14_1292 ();
 sg13g2_fill_8 FILLER_14_1300 ();
 sg13g2_fill_8 FILLER_14_1308 ();
 sg13g2_fill_8 FILLER_14_1316 ();
 sg13g2_fill_8 FILLER_14_1324 ();
 sg13g2_fill_8 FILLER_14_1332 ();
 sg13g2_fill_8 FILLER_14_1340 ();
 sg13g2_fill_8 FILLER_14_1348 ();
 sg13g2_fill_8 FILLER_14_1356 ();
 sg13g2_fill_8 FILLER_14_1364 ();
 sg13g2_fill_8 FILLER_14_1372 ();
 sg13g2_fill_8 FILLER_14_1380 ();
 sg13g2_fill_8 FILLER_14_1388 ();
 sg13g2_fill_8 FILLER_14_1396 ();
 sg13g2_fill_8 FILLER_14_1404 ();
 sg13g2_fill_8 FILLER_14_1412 ();
 sg13g2_fill_8 FILLER_14_1420 ();
 sg13g2_fill_8 FILLER_14_1428 ();
 sg13g2_fill_8 FILLER_14_1436 ();
 sg13g2_fill_8 FILLER_14_1444 ();
 sg13g2_fill_8 FILLER_14_1452 ();
 sg13g2_fill_8 FILLER_14_1460 ();
 sg13g2_fill_8 FILLER_14_1468 ();
 sg13g2_fill_8 FILLER_14_1476 ();
 sg13g2_fill_8 FILLER_14_1484 ();
 sg13g2_fill_8 FILLER_14_1492 ();
 sg13g2_fill_8 FILLER_14_1500 ();
 sg13g2_fill_8 FILLER_14_1508 ();
 sg13g2_fill_8 FILLER_14_1516 ();
 sg13g2_fill_8 FILLER_14_1524 ();
 sg13g2_fill_8 FILLER_14_1532 ();
 sg13g2_fill_8 FILLER_14_1540 ();
 sg13g2_fill_8 FILLER_14_1548 ();
 sg13g2_fill_8 FILLER_14_1556 ();
 sg13g2_fill_8 FILLER_14_1564 ();
 sg13g2_fill_8 FILLER_14_1572 ();
 sg13g2_fill_8 FILLER_14_1580 ();
 sg13g2_fill_4 FILLER_14_1588 ();
 sg13g2_fill_8 FILLER_15_0 ();
 sg13g2_fill_8 FILLER_15_8 ();
 sg13g2_fill_8 FILLER_15_16 ();
 sg13g2_fill_8 FILLER_15_24 ();
 sg13g2_fill_8 FILLER_15_32 ();
 sg13g2_fill_8 FILLER_15_40 ();
 sg13g2_fill_8 FILLER_15_48 ();
 sg13g2_fill_8 FILLER_15_56 ();
 sg13g2_fill_8 FILLER_15_64 ();
 sg13g2_fill_8 FILLER_15_72 ();
 sg13g2_fill_8 FILLER_15_80 ();
 sg13g2_fill_8 FILLER_15_88 ();
 sg13g2_fill_8 FILLER_15_96 ();
 sg13g2_fill_8 FILLER_15_104 ();
 sg13g2_fill_8 FILLER_15_112 ();
 sg13g2_fill_8 FILLER_15_120 ();
 sg13g2_fill_8 FILLER_15_128 ();
 sg13g2_fill_8 FILLER_15_136 ();
 sg13g2_fill_8 FILLER_15_144 ();
 sg13g2_fill_8 FILLER_15_152 ();
 sg13g2_fill_8 FILLER_15_160 ();
 sg13g2_fill_8 FILLER_15_168 ();
 sg13g2_fill_8 FILLER_15_176 ();
 sg13g2_fill_8 FILLER_15_184 ();
 sg13g2_fill_8 FILLER_15_192 ();
 sg13g2_fill_8 FILLER_15_200 ();
 sg13g2_fill_8 FILLER_15_208 ();
 sg13g2_fill_8 FILLER_15_216 ();
 sg13g2_fill_8 FILLER_15_224 ();
 sg13g2_fill_8 FILLER_15_232 ();
 sg13g2_fill_8 FILLER_15_240 ();
 sg13g2_fill_8 FILLER_15_248 ();
 sg13g2_fill_8 FILLER_15_256 ();
 sg13g2_fill_8 FILLER_15_264 ();
 sg13g2_fill_8 FILLER_15_272 ();
 sg13g2_fill_8 FILLER_15_280 ();
 sg13g2_fill_8 FILLER_15_288 ();
 sg13g2_fill_8 FILLER_15_296 ();
 sg13g2_fill_8 FILLER_15_304 ();
 sg13g2_fill_8 FILLER_15_312 ();
 sg13g2_fill_8 FILLER_15_320 ();
 sg13g2_fill_8 FILLER_15_328 ();
 sg13g2_fill_8 FILLER_15_336 ();
 sg13g2_fill_8 FILLER_15_344 ();
 sg13g2_fill_8 FILLER_15_352 ();
 sg13g2_fill_8 FILLER_15_360 ();
 sg13g2_fill_8 FILLER_15_368 ();
 sg13g2_fill_8 FILLER_15_376 ();
 sg13g2_fill_8 FILLER_15_384 ();
 sg13g2_fill_8 FILLER_15_392 ();
 sg13g2_fill_8 FILLER_15_400 ();
 sg13g2_fill_8 FILLER_15_408 ();
 sg13g2_fill_8 FILLER_15_416 ();
 sg13g2_fill_8 FILLER_15_424 ();
 sg13g2_fill_8 FILLER_15_432 ();
 sg13g2_fill_8 FILLER_15_440 ();
 sg13g2_fill_8 FILLER_15_448 ();
 sg13g2_fill_8 FILLER_15_526 ();
 sg13g2_fill_8 FILLER_15_534 ();
 sg13g2_fill_8 FILLER_15_552 ();
 sg13g2_fill_8 FILLER_15_560 ();
 sg13g2_fill_4 FILLER_15_568 ();
 sg13g2_fill_1 FILLER_15_572 ();
 sg13g2_fill_8 FILLER_15_603 ();
 sg13g2_fill_8 FILLER_15_611 ();
 sg13g2_fill_4 FILLER_15_619 ();
 sg13g2_fill_2 FILLER_15_623 ();
 sg13g2_fill_1 FILLER_15_635 ();
 sg13g2_fill_1 FILLER_15_641 ();
 sg13g2_fill_1 FILLER_15_666 ();
 sg13g2_fill_8 FILLER_15_677 ();
 sg13g2_fill_2 FILLER_15_685 ();
 sg13g2_fill_1 FILLER_15_687 ();
 sg13g2_fill_8 FILLER_15_696 ();
 sg13g2_fill_4 FILLER_15_704 ();
 sg13g2_fill_2 FILLER_15_745 ();
 sg13g2_fill_1 FILLER_15_747 ();
 sg13g2_fill_2 FILLER_15_753 ();
 sg13g2_fill_8 FILLER_15_773 ();
 sg13g2_fill_1 FILLER_15_781 ();
 sg13g2_fill_8 FILLER_15_808 ();
 sg13g2_fill_8 FILLER_15_816 ();
 sg13g2_fill_8 FILLER_15_824 ();
 sg13g2_fill_4 FILLER_15_832 ();
 sg13g2_fill_1 FILLER_15_836 ();
 sg13g2_fill_4 FILLER_15_858 ();
 sg13g2_fill_1 FILLER_15_862 ();
 sg13g2_fill_8 FILLER_15_873 ();
 sg13g2_fill_8 FILLER_15_881 ();
 sg13g2_fill_4 FILLER_15_889 ();
 sg13g2_fill_2 FILLER_15_919 ();
 sg13g2_fill_1 FILLER_15_925 ();
 sg13g2_fill_8 FILLER_15_930 ();
 sg13g2_fill_4 FILLER_15_938 ();
 sg13g2_fill_1 FILLER_15_942 ();
 sg13g2_fill_8 FILLER_15_948 ();
 sg13g2_fill_4 FILLER_15_956 ();
 sg13g2_fill_1 FILLER_15_960 ();
 sg13g2_fill_8 FILLER_15_975 ();
 sg13g2_fill_8 FILLER_15_983 ();
 sg13g2_fill_1 FILLER_15_991 ();
 sg13g2_fill_1 FILLER_15_1018 ();
 sg13g2_fill_4 FILLER_15_1070 ();
 sg13g2_fill_8 FILLER_15_1110 ();
 sg13g2_fill_1 FILLER_15_1118 ();
 sg13g2_fill_2 FILLER_15_1127 ();
 sg13g2_fill_2 FILLER_15_1165 ();
 sg13g2_fill_1 FILLER_15_1167 ();
 sg13g2_fill_8 FILLER_15_1233 ();
 sg13g2_fill_1 FILLER_15_1241 ();
 sg13g2_fill_8 FILLER_15_1267 ();
 sg13g2_fill_8 FILLER_15_1275 ();
 sg13g2_fill_8 FILLER_15_1283 ();
 sg13g2_fill_8 FILLER_15_1291 ();
 sg13g2_fill_8 FILLER_15_1299 ();
 sg13g2_fill_8 FILLER_15_1307 ();
 sg13g2_fill_8 FILLER_15_1315 ();
 sg13g2_fill_8 FILLER_15_1323 ();
 sg13g2_fill_8 FILLER_15_1331 ();
 sg13g2_fill_8 FILLER_15_1339 ();
 sg13g2_fill_8 FILLER_15_1347 ();
 sg13g2_fill_8 FILLER_15_1355 ();
 sg13g2_fill_8 FILLER_15_1363 ();
 sg13g2_fill_8 FILLER_15_1371 ();
 sg13g2_fill_8 FILLER_15_1379 ();
 sg13g2_fill_8 FILLER_15_1387 ();
 sg13g2_fill_8 FILLER_15_1395 ();
 sg13g2_fill_8 FILLER_15_1403 ();
 sg13g2_fill_8 FILLER_15_1411 ();
 sg13g2_fill_8 FILLER_15_1419 ();
 sg13g2_fill_8 FILLER_15_1427 ();
 sg13g2_fill_8 FILLER_15_1435 ();
 sg13g2_fill_8 FILLER_15_1443 ();
 sg13g2_fill_8 FILLER_15_1451 ();
 sg13g2_fill_8 FILLER_15_1459 ();
 sg13g2_fill_8 FILLER_15_1467 ();
 sg13g2_fill_8 FILLER_15_1475 ();
 sg13g2_fill_8 FILLER_15_1483 ();
 sg13g2_fill_8 FILLER_15_1491 ();
 sg13g2_fill_8 FILLER_15_1499 ();
 sg13g2_fill_8 FILLER_15_1507 ();
 sg13g2_fill_8 FILLER_15_1515 ();
 sg13g2_fill_8 FILLER_15_1523 ();
 sg13g2_fill_8 FILLER_15_1531 ();
 sg13g2_fill_8 FILLER_15_1539 ();
 sg13g2_fill_8 FILLER_15_1547 ();
 sg13g2_fill_8 FILLER_15_1555 ();
 sg13g2_fill_8 FILLER_15_1563 ();
 sg13g2_fill_8 FILLER_15_1571 ();
 sg13g2_fill_8 FILLER_15_1579 ();
 sg13g2_fill_4 FILLER_15_1587 ();
 sg13g2_fill_1 FILLER_15_1591 ();
 sg13g2_fill_8 FILLER_16_0 ();
 sg13g2_fill_8 FILLER_16_8 ();
 sg13g2_fill_8 FILLER_16_16 ();
 sg13g2_fill_8 FILLER_16_24 ();
 sg13g2_fill_8 FILLER_16_32 ();
 sg13g2_fill_8 FILLER_16_40 ();
 sg13g2_fill_8 FILLER_16_48 ();
 sg13g2_fill_8 FILLER_16_56 ();
 sg13g2_fill_8 FILLER_16_64 ();
 sg13g2_fill_8 FILLER_16_72 ();
 sg13g2_fill_8 FILLER_16_80 ();
 sg13g2_fill_8 FILLER_16_88 ();
 sg13g2_fill_8 FILLER_16_96 ();
 sg13g2_fill_8 FILLER_16_104 ();
 sg13g2_fill_8 FILLER_16_112 ();
 sg13g2_fill_8 FILLER_16_120 ();
 sg13g2_fill_8 FILLER_16_128 ();
 sg13g2_fill_8 FILLER_16_136 ();
 sg13g2_fill_8 FILLER_16_144 ();
 sg13g2_fill_8 FILLER_16_152 ();
 sg13g2_fill_8 FILLER_16_160 ();
 sg13g2_fill_8 FILLER_16_168 ();
 sg13g2_fill_8 FILLER_16_176 ();
 sg13g2_fill_8 FILLER_16_184 ();
 sg13g2_fill_8 FILLER_16_192 ();
 sg13g2_fill_8 FILLER_16_200 ();
 sg13g2_fill_8 FILLER_16_208 ();
 sg13g2_fill_8 FILLER_16_216 ();
 sg13g2_fill_8 FILLER_16_224 ();
 sg13g2_fill_8 FILLER_16_232 ();
 sg13g2_fill_8 FILLER_16_240 ();
 sg13g2_fill_8 FILLER_16_248 ();
 sg13g2_fill_8 FILLER_16_256 ();
 sg13g2_fill_8 FILLER_16_264 ();
 sg13g2_fill_8 FILLER_16_272 ();
 sg13g2_fill_8 FILLER_16_280 ();
 sg13g2_fill_8 FILLER_16_288 ();
 sg13g2_fill_8 FILLER_16_296 ();
 sg13g2_fill_8 FILLER_16_304 ();
 sg13g2_fill_8 FILLER_16_312 ();
 sg13g2_fill_8 FILLER_16_320 ();
 sg13g2_fill_8 FILLER_16_328 ();
 sg13g2_fill_8 FILLER_16_336 ();
 sg13g2_fill_8 FILLER_16_344 ();
 sg13g2_fill_8 FILLER_16_352 ();
 sg13g2_fill_8 FILLER_16_360 ();
 sg13g2_fill_8 FILLER_16_368 ();
 sg13g2_fill_8 FILLER_16_376 ();
 sg13g2_fill_8 FILLER_16_384 ();
 sg13g2_fill_8 FILLER_16_392 ();
 sg13g2_fill_8 FILLER_16_400 ();
 sg13g2_fill_4 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_16_438 ();
 sg13g2_fill_1 FILLER_16_440 ();
 sg13g2_fill_8 FILLER_16_451 ();
 sg13g2_fill_1 FILLER_16_459 ();
 sg13g2_fill_2 FILLER_16_468 ();
 sg13g2_fill_8 FILLER_16_480 ();
 sg13g2_fill_4 FILLER_16_488 ();
 sg13g2_fill_2 FILLER_16_492 ();
 sg13g2_fill_8 FILLER_16_498 ();
 sg13g2_fill_8 FILLER_16_506 ();
 sg13g2_fill_1 FILLER_16_514 ();
 sg13g2_fill_8 FILLER_16_525 ();
 sg13g2_fill_8 FILLER_16_533 ();
 sg13g2_fill_4 FILLER_16_567 ();
 sg13g2_fill_1 FILLER_16_571 ();
 sg13g2_fill_1 FILLER_16_629 ();
 sg13g2_fill_8 FILLER_16_637 ();
 sg13g2_fill_4 FILLER_16_645 ();
 sg13g2_fill_2 FILLER_16_649 ();
 sg13g2_fill_2 FILLER_16_666 ();
 sg13g2_fill_1 FILLER_16_668 ();
 sg13g2_fill_4 FILLER_16_674 ();
 sg13g2_fill_8 FILLER_16_704 ();
 sg13g2_fill_4 FILLER_16_712 ();
 sg13g2_fill_1 FILLER_16_716 ();
 sg13g2_fill_4 FILLER_16_724 ();
 sg13g2_fill_4 FILLER_16_733 ();
 sg13g2_fill_1 FILLER_16_737 ();
 sg13g2_fill_4 FILLER_16_742 ();
 sg13g2_fill_2 FILLER_16_746 ();
 sg13g2_fill_1 FILLER_16_753 ();
 sg13g2_fill_8 FILLER_16_776 ();
 sg13g2_fill_8 FILLER_16_784 ();
 sg13g2_fill_2 FILLER_16_792 ();
 sg13g2_fill_1 FILLER_16_794 ();
 sg13g2_fill_4 FILLER_16_815 ();
 sg13g2_fill_2 FILLER_16_819 ();
 sg13g2_fill_8 FILLER_16_839 ();
 sg13g2_fill_4 FILLER_16_847 ();
 sg13g2_fill_2 FILLER_16_851 ();
 sg13g2_fill_4 FILLER_16_861 ();
 sg13g2_fill_2 FILLER_16_865 ();
 sg13g2_fill_1 FILLER_16_867 ();
 sg13g2_fill_4 FILLER_16_894 ();
 sg13g2_fill_2 FILLER_16_903 ();
 sg13g2_fill_2 FILLER_16_914 ();
 sg13g2_fill_8 FILLER_16_925 ();
 sg13g2_fill_8 FILLER_16_933 ();
 sg13g2_fill_8 FILLER_16_941 ();
 sg13g2_fill_4 FILLER_16_949 ();
 sg13g2_fill_1 FILLER_16_953 ();
 sg13g2_fill_2 FILLER_16_974 ();
 sg13g2_fill_1 FILLER_16_976 ();
 sg13g2_fill_8 FILLER_16_1013 ();
 sg13g2_fill_8 FILLER_16_1021 ();
 sg13g2_fill_4 FILLER_16_1029 ();
 sg13g2_fill_1 FILLER_16_1033 ();
 sg13g2_fill_1 FILLER_16_1078 ();
 sg13g2_fill_4 FILLER_16_1095 ();
 sg13g2_fill_2 FILLER_16_1099 ();
 sg13g2_fill_1 FILLER_16_1101 ();
 sg13g2_fill_8 FILLER_16_1113 ();
 sg13g2_fill_8 FILLER_16_1121 ();
 sg13g2_fill_4 FILLER_16_1129 ();
 sg13g2_fill_8 FILLER_16_1190 ();
 sg13g2_fill_8 FILLER_16_1198 ();
 sg13g2_fill_4 FILLER_16_1206 ();
 sg13g2_fill_8 FILLER_16_1215 ();
 sg13g2_fill_8 FILLER_16_1223 ();
 sg13g2_fill_4 FILLER_16_1231 ();
 sg13g2_fill_2 FILLER_16_1235 ();
 sg13g2_fill_1 FILLER_16_1237 ();
 sg13g2_fill_8 FILLER_16_1263 ();
 sg13g2_fill_8 FILLER_16_1271 ();
 sg13g2_fill_8 FILLER_16_1279 ();
 sg13g2_fill_8 FILLER_16_1287 ();
 sg13g2_fill_8 FILLER_16_1295 ();
 sg13g2_fill_8 FILLER_16_1303 ();
 sg13g2_fill_8 FILLER_16_1311 ();
 sg13g2_fill_8 FILLER_16_1319 ();
 sg13g2_fill_8 FILLER_16_1327 ();
 sg13g2_fill_8 FILLER_16_1335 ();
 sg13g2_fill_8 FILLER_16_1343 ();
 sg13g2_fill_8 FILLER_16_1351 ();
 sg13g2_fill_8 FILLER_16_1359 ();
 sg13g2_fill_8 FILLER_16_1367 ();
 sg13g2_fill_8 FILLER_16_1375 ();
 sg13g2_fill_8 FILLER_16_1383 ();
 sg13g2_fill_8 FILLER_16_1391 ();
 sg13g2_fill_8 FILLER_16_1399 ();
 sg13g2_fill_8 FILLER_16_1407 ();
 sg13g2_fill_8 FILLER_16_1415 ();
 sg13g2_fill_8 FILLER_16_1423 ();
 sg13g2_fill_8 FILLER_16_1431 ();
 sg13g2_fill_8 FILLER_16_1439 ();
 sg13g2_fill_8 FILLER_16_1447 ();
 sg13g2_fill_8 FILLER_16_1455 ();
 sg13g2_fill_8 FILLER_16_1463 ();
 sg13g2_fill_8 FILLER_16_1471 ();
 sg13g2_fill_8 FILLER_16_1479 ();
 sg13g2_fill_8 FILLER_16_1487 ();
 sg13g2_fill_8 FILLER_16_1495 ();
 sg13g2_fill_8 FILLER_16_1503 ();
 sg13g2_fill_8 FILLER_16_1511 ();
 sg13g2_fill_8 FILLER_16_1519 ();
 sg13g2_fill_8 FILLER_16_1527 ();
 sg13g2_fill_8 FILLER_16_1535 ();
 sg13g2_fill_8 FILLER_16_1543 ();
 sg13g2_fill_8 FILLER_16_1551 ();
 sg13g2_fill_8 FILLER_16_1559 ();
 sg13g2_fill_8 FILLER_16_1567 ();
 sg13g2_fill_8 FILLER_16_1575 ();
 sg13g2_fill_8 FILLER_16_1583 ();
 sg13g2_fill_1 FILLER_16_1591 ();
 sg13g2_fill_8 FILLER_17_0 ();
 sg13g2_fill_8 FILLER_17_8 ();
 sg13g2_fill_8 FILLER_17_16 ();
 sg13g2_fill_8 FILLER_17_24 ();
 sg13g2_fill_8 FILLER_17_32 ();
 sg13g2_fill_8 FILLER_17_40 ();
 sg13g2_fill_8 FILLER_17_48 ();
 sg13g2_fill_8 FILLER_17_56 ();
 sg13g2_fill_8 FILLER_17_64 ();
 sg13g2_fill_8 FILLER_17_72 ();
 sg13g2_fill_8 FILLER_17_80 ();
 sg13g2_fill_8 FILLER_17_88 ();
 sg13g2_fill_8 FILLER_17_96 ();
 sg13g2_fill_8 FILLER_17_104 ();
 sg13g2_fill_8 FILLER_17_112 ();
 sg13g2_fill_8 FILLER_17_120 ();
 sg13g2_fill_8 FILLER_17_128 ();
 sg13g2_fill_8 FILLER_17_136 ();
 sg13g2_fill_8 FILLER_17_144 ();
 sg13g2_fill_8 FILLER_17_152 ();
 sg13g2_fill_8 FILLER_17_160 ();
 sg13g2_fill_8 FILLER_17_168 ();
 sg13g2_fill_8 FILLER_17_176 ();
 sg13g2_fill_8 FILLER_17_184 ();
 sg13g2_fill_8 FILLER_17_192 ();
 sg13g2_fill_8 FILLER_17_200 ();
 sg13g2_fill_8 FILLER_17_208 ();
 sg13g2_fill_8 FILLER_17_216 ();
 sg13g2_fill_8 FILLER_17_224 ();
 sg13g2_fill_8 FILLER_17_232 ();
 sg13g2_fill_8 FILLER_17_240 ();
 sg13g2_fill_8 FILLER_17_248 ();
 sg13g2_fill_8 FILLER_17_256 ();
 sg13g2_fill_8 FILLER_17_264 ();
 sg13g2_fill_8 FILLER_17_272 ();
 sg13g2_fill_8 FILLER_17_280 ();
 sg13g2_fill_8 FILLER_17_288 ();
 sg13g2_fill_8 FILLER_17_296 ();
 sg13g2_fill_8 FILLER_17_304 ();
 sg13g2_fill_8 FILLER_17_312 ();
 sg13g2_fill_8 FILLER_17_320 ();
 sg13g2_fill_8 FILLER_17_328 ();
 sg13g2_fill_8 FILLER_17_336 ();
 sg13g2_fill_8 FILLER_17_344 ();
 sg13g2_fill_8 FILLER_17_352 ();
 sg13g2_fill_8 FILLER_17_360 ();
 sg13g2_fill_8 FILLER_17_368 ();
 sg13g2_fill_8 FILLER_17_376 ();
 sg13g2_fill_8 FILLER_17_384 ();
 sg13g2_fill_8 FILLER_17_392 ();
 sg13g2_fill_8 FILLER_17_400 ();
 sg13g2_fill_4 FILLER_17_485 ();
 sg13g2_fill_2 FILLER_17_489 ();
 sg13g2_fill_4 FILLER_17_543 ();
 sg13g2_fill_8 FILLER_17_555 ();
 sg13g2_fill_8 FILLER_17_563 ();
 sg13g2_fill_8 FILLER_17_571 ();
 sg13g2_fill_8 FILLER_17_579 ();
 sg13g2_fill_8 FILLER_17_587 ();
 sg13g2_fill_8 FILLER_17_595 ();
 sg13g2_fill_1 FILLER_17_603 ();
 sg13g2_fill_8 FILLER_17_622 ();
 sg13g2_fill_4 FILLER_17_630 ();
 sg13g2_fill_2 FILLER_17_634 ();
 sg13g2_fill_1 FILLER_17_636 ();
 sg13g2_fill_2 FILLER_17_661 ();
 sg13g2_fill_1 FILLER_17_673 ();
 sg13g2_fill_8 FILLER_17_679 ();
 sg13g2_fill_4 FILLER_17_708 ();
 sg13g2_fill_2 FILLER_17_712 ();
 sg13g2_fill_2 FILLER_17_724 ();
 sg13g2_fill_1 FILLER_17_731 ();
 sg13g2_fill_1 FILLER_17_754 ();
 sg13g2_fill_2 FILLER_17_768 ();
 sg13g2_fill_1 FILLER_17_770 ();
 sg13g2_fill_8 FILLER_17_792 ();
 sg13g2_fill_4 FILLER_17_800 ();
 sg13g2_fill_2 FILLER_17_804 ();
 sg13g2_fill_1 FILLER_17_806 ();
 sg13g2_fill_8 FILLER_17_817 ();
 sg13g2_fill_4 FILLER_17_825 ();
 sg13g2_fill_1 FILLER_17_829 ();
 sg13g2_fill_4 FILLER_17_892 ();
 sg13g2_fill_2 FILLER_17_896 ();
 sg13g2_fill_1 FILLER_17_898 ();
 sg13g2_fill_8 FILLER_17_903 ();
 sg13g2_fill_1 FILLER_17_911 ();
 sg13g2_fill_4 FILLER_17_920 ();
 sg13g2_fill_1 FILLER_17_924 ();
 sg13g2_fill_1 FILLER_17_957 ();
 sg13g2_fill_2 FILLER_17_964 ();
 sg13g2_fill_1 FILLER_17_1004 ();
 sg13g2_fill_8 FILLER_17_1034 ();
 sg13g2_fill_8 FILLER_17_1048 ();
 sg13g2_fill_2 FILLER_17_1056 ();
 sg13g2_fill_8 FILLER_17_1062 ();
 sg13g2_fill_4 FILLER_17_1070 ();
 sg13g2_fill_1 FILLER_17_1074 ();
 sg13g2_fill_1 FILLER_17_1085 ();
 sg13g2_fill_8 FILLER_17_1091 ();
 sg13g2_fill_8 FILLER_17_1099 ();
 sg13g2_fill_8 FILLER_17_1107 ();
 sg13g2_fill_1 FILLER_17_1115 ();
 sg13g2_fill_4 FILLER_17_1154 ();
 sg13g2_fill_1 FILLER_17_1158 ();
 sg13g2_fill_4 FILLER_17_1167 ();
 sg13g2_fill_8 FILLER_17_1196 ();
 sg13g2_fill_1 FILLER_17_1204 ();
 sg13g2_fill_8 FILLER_17_1241 ();
 sg13g2_fill_8 FILLER_17_1249 ();
 sg13g2_fill_8 FILLER_17_1257 ();
 sg13g2_fill_8 FILLER_17_1265 ();
 sg13g2_fill_8 FILLER_17_1273 ();
 sg13g2_fill_8 FILLER_17_1281 ();
 sg13g2_fill_8 FILLER_17_1289 ();
 sg13g2_fill_8 FILLER_17_1297 ();
 sg13g2_fill_8 FILLER_17_1305 ();
 sg13g2_fill_8 FILLER_17_1313 ();
 sg13g2_fill_8 FILLER_17_1321 ();
 sg13g2_fill_8 FILLER_17_1329 ();
 sg13g2_fill_8 FILLER_17_1337 ();
 sg13g2_fill_8 FILLER_17_1345 ();
 sg13g2_fill_8 FILLER_17_1353 ();
 sg13g2_fill_8 FILLER_17_1361 ();
 sg13g2_fill_8 FILLER_17_1369 ();
 sg13g2_fill_8 FILLER_17_1377 ();
 sg13g2_fill_8 FILLER_17_1385 ();
 sg13g2_fill_8 FILLER_17_1393 ();
 sg13g2_fill_8 FILLER_17_1401 ();
 sg13g2_fill_8 FILLER_17_1409 ();
 sg13g2_fill_8 FILLER_17_1417 ();
 sg13g2_fill_8 FILLER_17_1425 ();
 sg13g2_fill_8 FILLER_17_1433 ();
 sg13g2_fill_8 FILLER_17_1441 ();
 sg13g2_fill_8 FILLER_17_1449 ();
 sg13g2_fill_8 FILLER_17_1457 ();
 sg13g2_fill_8 FILLER_17_1465 ();
 sg13g2_fill_8 FILLER_17_1473 ();
 sg13g2_fill_8 FILLER_17_1481 ();
 sg13g2_fill_8 FILLER_17_1489 ();
 sg13g2_fill_8 FILLER_17_1497 ();
 sg13g2_fill_8 FILLER_17_1505 ();
 sg13g2_fill_8 FILLER_17_1513 ();
 sg13g2_fill_8 FILLER_17_1521 ();
 sg13g2_fill_8 FILLER_17_1529 ();
 sg13g2_fill_8 FILLER_17_1537 ();
 sg13g2_fill_8 FILLER_17_1545 ();
 sg13g2_fill_8 FILLER_17_1553 ();
 sg13g2_fill_8 FILLER_17_1561 ();
 sg13g2_fill_8 FILLER_17_1569 ();
 sg13g2_fill_8 FILLER_17_1577 ();
 sg13g2_fill_4 FILLER_17_1585 ();
 sg13g2_fill_2 FILLER_17_1589 ();
 sg13g2_fill_1 FILLER_17_1591 ();
 sg13g2_fill_8 FILLER_18_0 ();
 sg13g2_fill_8 FILLER_18_8 ();
 sg13g2_fill_8 FILLER_18_16 ();
 sg13g2_fill_8 FILLER_18_24 ();
 sg13g2_fill_8 FILLER_18_32 ();
 sg13g2_fill_8 FILLER_18_40 ();
 sg13g2_fill_8 FILLER_18_48 ();
 sg13g2_fill_8 FILLER_18_56 ();
 sg13g2_fill_8 FILLER_18_64 ();
 sg13g2_fill_8 FILLER_18_72 ();
 sg13g2_fill_8 FILLER_18_80 ();
 sg13g2_fill_8 FILLER_18_88 ();
 sg13g2_fill_8 FILLER_18_96 ();
 sg13g2_fill_8 FILLER_18_104 ();
 sg13g2_fill_8 FILLER_18_112 ();
 sg13g2_fill_8 FILLER_18_120 ();
 sg13g2_fill_8 FILLER_18_128 ();
 sg13g2_fill_8 FILLER_18_136 ();
 sg13g2_fill_8 FILLER_18_144 ();
 sg13g2_fill_8 FILLER_18_152 ();
 sg13g2_fill_8 FILLER_18_160 ();
 sg13g2_fill_8 FILLER_18_168 ();
 sg13g2_fill_8 FILLER_18_176 ();
 sg13g2_fill_8 FILLER_18_184 ();
 sg13g2_fill_8 FILLER_18_192 ();
 sg13g2_fill_8 FILLER_18_200 ();
 sg13g2_fill_8 FILLER_18_208 ();
 sg13g2_fill_8 FILLER_18_216 ();
 sg13g2_fill_8 FILLER_18_224 ();
 sg13g2_fill_8 FILLER_18_232 ();
 sg13g2_fill_8 FILLER_18_240 ();
 sg13g2_fill_8 FILLER_18_248 ();
 sg13g2_fill_8 FILLER_18_256 ();
 sg13g2_fill_8 FILLER_18_264 ();
 sg13g2_fill_8 FILLER_18_272 ();
 sg13g2_fill_8 FILLER_18_280 ();
 sg13g2_fill_8 FILLER_18_288 ();
 sg13g2_fill_8 FILLER_18_296 ();
 sg13g2_fill_8 FILLER_18_304 ();
 sg13g2_fill_8 FILLER_18_312 ();
 sg13g2_fill_8 FILLER_18_320 ();
 sg13g2_fill_8 FILLER_18_328 ();
 sg13g2_fill_8 FILLER_18_336 ();
 sg13g2_fill_8 FILLER_18_344 ();
 sg13g2_fill_8 FILLER_18_352 ();
 sg13g2_fill_8 FILLER_18_360 ();
 sg13g2_fill_8 FILLER_18_368 ();
 sg13g2_fill_8 FILLER_18_376 ();
 sg13g2_fill_8 FILLER_18_384 ();
 sg13g2_fill_8 FILLER_18_392 ();
 sg13g2_fill_4 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_406 ();
 sg13g2_fill_8 FILLER_18_417 ();
 sg13g2_fill_8 FILLER_18_425 ();
 sg13g2_fill_4 FILLER_18_433 ();
 sg13g2_fill_2 FILLER_18_437 ();
 sg13g2_fill_1 FILLER_18_439 ();
 sg13g2_fill_8 FILLER_18_450 ();
 sg13g2_fill_8 FILLER_18_458 ();
 sg13g2_fill_1 FILLER_18_492 ();
 sg13g2_fill_8 FILLER_18_503 ();
 sg13g2_fill_8 FILLER_18_511 ();
 sg13g2_fill_8 FILLER_18_519 ();
 sg13g2_fill_8 FILLER_18_527 ();
 sg13g2_fill_2 FILLER_18_535 ();
 sg13g2_fill_8 FILLER_18_547 ();
 sg13g2_fill_4 FILLER_18_563 ();
 sg13g2_fill_2 FILLER_18_567 ();
 sg13g2_fill_8 FILLER_18_598 ();
 sg13g2_fill_4 FILLER_18_622 ();
 sg13g2_fill_1 FILLER_18_626 ();
 sg13g2_fill_4 FILLER_18_633 ();
 sg13g2_fill_1 FILLER_18_642 ();
 sg13g2_fill_2 FILLER_18_647 ();
 sg13g2_fill_1 FILLER_18_649 ();
 sg13g2_fill_8 FILLER_18_664 ();
 sg13g2_fill_8 FILLER_18_672 ();
 sg13g2_fill_2 FILLER_18_706 ();
 sg13g2_fill_1 FILLER_18_708 ();
 sg13g2_fill_4 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_743 ();
 sg13g2_fill_4 FILLER_18_793 ();
 sg13g2_fill_2 FILLER_18_797 ();
 sg13g2_fill_4 FILLER_18_861 ();
 sg13g2_fill_2 FILLER_18_865 ();
 sg13g2_fill_1 FILLER_18_867 ();
 sg13g2_fill_4 FILLER_18_883 ();
 sg13g2_fill_8 FILLER_18_958 ();
 sg13g2_fill_8 FILLER_18_966 ();
 sg13g2_fill_8 FILLER_18_974 ();
 sg13g2_fill_1 FILLER_18_982 ();
 sg13g2_fill_2 FILLER_18_988 ();
 sg13g2_fill_1 FILLER_18_990 ();
 sg13g2_fill_4 FILLER_18_996 ();
 sg13g2_fill_2 FILLER_18_1020 ();
 sg13g2_fill_4 FILLER_18_1048 ();
 sg13g2_fill_2 FILLER_18_1052 ();
 sg13g2_fill_1 FILLER_18_1054 ();
 sg13g2_fill_2 FILLER_18_1081 ();
 sg13g2_fill_1 FILLER_18_1083 ();
 sg13g2_fill_8 FILLER_18_1120 ();
 sg13g2_fill_4 FILLER_18_1128 ();
 sg13g2_fill_4 FILLER_18_1142 ();
 sg13g2_fill_2 FILLER_18_1146 ();
 sg13g2_fill_1 FILLER_18_1148 ();
 sg13g2_fill_2 FILLER_18_1159 ();
 sg13g2_fill_4 FILLER_18_1220 ();
 sg13g2_fill_2 FILLER_18_1224 ();
 sg13g2_fill_1 FILLER_18_1226 ();
 sg13g2_fill_8 FILLER_18_1235 ();
 sg13g2_fill_1 FILLER_18_1243 ();
 sg13g2_fill_2 FILLER_18_1249 ();
 sg13g2_fill_8 FILLER_18_1281 ();
 sg13g2_fill_8 FILLER_18_1289 ();
 sg13g2_fill_8 FILLER_18_1297 ();
 sg13g2_fill_8 FILLER_18_1305 ();
 sg13g2_fill_8 FILLER_18_1313 ();
 sg13g2_fill_8 FILLER_18_1321 ();
 sg13g2_fill_8 FILLER_18_1329 ();
 sg13g2_fill_8 FILLER_18_1337 ();
 sg13g2_fill_8 FILLER_18_1345 ();
 sg13g2_fill_8 FILLER_18_1353 ();
 sg13g2_fill_8 FILLER_18_1361 ();
 sg13g2_fill_8 FILLER_18_1369 ();
 sg13g2_fill_8 FILLER_18_1377 ();
 sg13g2_fill_8 FILLER_18_1385 ();
 sg13g2_fill_8 FILLER_18_1393 ();
 sg13g2_fill_8 FILLER_18_1401 ();
 sg13g2_fill_8 FILLER_18_1409 ();
 sg13g2_fill_8 FILLER_18_1417 ();
 sg13g2_fill_8 FILLER_18_1425 ();
 sg13g2_fill_8 FILLER_18_1433 ();
 sg13g2_fill_8 FILLER_18_1441 ();
 sg13g2_fill_8 FILLER_18_1449 ();
 sg13g2_fill_8 FILLER_18_1457 ();
 sg13g2_fill_8 FILLER_18_1465 ();
 sg13g2_fill_8 FILLER_18_1473 ();
 sg13g2_fill_8 FILLER_18_1481 ();
 sg13g2_fill_8 FILLER_18_1489 ();
 sg13g2_fill_8 FILLER_18_1497 ();
 sg13g2_fill_8 FILLER_18_1505 ();
 sg13g2_fill_8 FILLER_18_1513 ();
 sg13g2_fill_8 FILLER_18_1521 ();
 sg13g2_fill_8 FILLER_18_1529 ();
 sg13g2_fill_8 FILLER_18_1537 ();
 sg13g2_fill_8 FILLER_18_1545 ();
 sg13g2_fill_8 FILLER_18_1553 ();
 sg13g2_fill_8 FILLER_18_1561 ();
 sg13g2_fill_8 FILLER_18_1569 ();
 sg13g2_fill_8 FILLER_18_1577 ();
 sg13g2_fill_4 FILLER_18_1585 ();
 sg13g2_fill_2 FILLER_18_1589 ();
 sg13g2_fill_1 FILLER_18_1591 ();
 sg13g2_fill_8 FILLER_19_0 ();
 sg13g2_fill_8 FILLER_19_8 ();
 sg13g2_fill_8 FILLER_19_16 ();
 sg13g2_fill_8 FILLER_19_24 ();
 sg13g2_fill_8 FILLER_19_32 ();
 sg13g2_fill_8 FILLER_19_40 ();
 sg13g2_fill_8 FILLER_19_48 ();
 sg13g2_fill_8 FILLER_19_56 ();
 sg13g2_fill_8 FILLER_19_64 ();
 sg13g2_fill_8 FILLER_19_72 ();
 sg13g2_fill_8 FILLER_19_80 ();
 sg13g2_fill_8 FILLER_19_88 ();
 sg13g2_fill_8 FILLER_19_96 ();
 sg13g2_fill_8 FILLER_19_104 ();
 sg13g2_fill_8 FILLER_19_112 ();
 sg13g2_fill_8 FILLER_19_120 ();
 sg13g2_fill_8 FILLER_19_128 ();
 sg13g2_fill_8 FILLER_19_136 ();
 sg13g2_fill_8 FILLER_19_144 ();
 sg13g2_fill_8 FILLER_19_152 ();
 sg13g2_fill_8 FILLER_19_160 ();
 sg13g2_fill_8 FILLER_19_168 ();
 sg13g2_fill_8 FILLER_19_176 ();
 sg13g2_fill_8 FILLER_19_184 ();
 sg13g2_fill_8 FILLER_19_192 ();
 sg13g2_fill_8 FILLER_19_200 ();
 sg13g2_fill_8 FILLER_19_208 ();
 sg13g2_fill_8 FILLER_19_216 ();
 sg13g2_fill_8 FILLER_19_224 ();
 sg13g2_fill_8 FILLER_19_232 ();
 sg13g2_fill_8 FILLER_19_240 ();
 sg13g2_fill_8 FILLER_19_248 ();
 sg13g2_fill_8 FILLER_19_256 ();
 sg13g2_fill_8 FILLER_19_264 ();
 sg13g2_fill_8 FILLER_19_272 ();
 sg13g2_fill_8 FILLER_19_280 ();
 sg13g2_fill_8 FILLER_19_288 ();
 sg13g2_fill_8 FILLER_19_296 ();
 sg13g2_fill_8 FILLER_19_304 ();
 sg13g2_fill_8 FILLER_19_312 ();
 sg13g2_fill_8 FILLER_19_320 ();
 sg13g2_fill_8 FILLER_19_328 ();
 sg13g2_fill_8 FILLER_19_336 ();
 sg13g2_fill_8 FILLER_19_344 ();
 sg13g2_fill_8 FILLER_19_352 ();
 sg13g2_fill_8 FILLER_19_360 ();
 sg13g2_fill_8 FILLER_19_368 ();
 sg13g2_fill_8 FILLER_19_376 ();
 sg13g2_fill_8 FILLER_19_384 ();
 sg13g2_fill_8 FILLER_19_392 ();
 sg13g2_fill_8 FILLER_19_400 ();
 sg13g2_fill_4 FILLER_19_408 ();
 sg13g2_fill_1 FILLER_19_412 ();
 sg13g2_fill_8 FILLER_19_423 ();
 sg13g2_fill_1 FILLER_19_431 ();
 sg13g2_fill_8 FILLER_19_457 ();
 sg13g2_fill_8 FILLER_19_465 ();
 sg13g2_fill_8 FILLER_19_473 ();
 sg13g2_fill_8 FILLER_19_481 ();
 sg13g2_fill_1 FILLER_19_489 ();
 sg13g2_fill_8 FILLER_19_516 ();
 sg13g2_fill_4 FILLER_19_524 ();
 sg13g2_fill_2 FILLER_19_528 ();
 sg13g2_fill_4 FILLER_19_540 ();
 sg13g2_fill_1 FILLER_19_544 ();
 sg13g2_fill_2 FILLER_19_571 ();
 sg13g2_fill_1 FILLER_19_573 ();
 sg13g2_fill_2 FILLER_19_600 ();
 sg13g2_fill_1 FILLER_19_602 ();
 sg13g2_fill_4 FILLER_19_618 ();
 sg13g2_fill_1 FILLER_19_630 ();
 sg13g2_fill_8 FILLER_19_644 ();
 sg13g2_fill_2 FILLER_19_652 ();
 sg13g2_fill_8 FILLER_19_680 ();
 sg13g2_fill_8 FILLER_19_688 ();
 sg13g2_fill_8 FILLER_19_704 ();
 sg13g2_fill_8 FILLER_19_712 ();
 sg13g2_fill_4 FILLER_19_725 ();
 sg13g2_fill_2 FILLER_19_729 ();
 sg13g2_fill_1 FILLER_19_731 ();
 sg13g2_fill_4 FILLER_19_736 ();
 sg13g2_fill_1 FILLER_19_740 ();
 sg13g2_fill_8 FILLER_19_774 ();
 sg13g2_fill_2 FILLER_19_782 ();
 sg13g2_fill_1 FILLER_19_784 ();
 sg13g2_fill_2 FILLER_19_798 ();
 sg13g2_fill_1 FILLER_19_800 ();
 sg13g2_fill_8 FILLER_19_809 ();
 sg13g2_fill_4 FILLER_19_817 ();
 sg13g2_fill_2 FILLER_19_821 ();
 sg13g2_fill_8 FILLER_19_833 ();
 sg13g2_fill_1 FILLER_19_841 ();
 sg13g2_fill_2 FILLER_19_867 ();
 sg13g2_fill_2 FILLER_19_894 ();
 sg13g2_fill_1 FILLER_19_896 ();
 sg13g2_fill_1 FILLER_19_922 ();
 sg13g2_fill_8 FILLER_19_936 ();
 sg13g2_fill_8 FILLER_19_944 ();
 sg13g2_fill_4 FILLER_19_982 ();
 sg13g2_fill_2 FILLER_19_986 ();
 sg13g2_fill_1 FILLER_19_988 ();
 sg13g2_fill_4 FILLER_19_1070 ();
 sg13g2_fill_1 FILLER_19_1074 ();
 sg13g2_fill_1 FILLER_19_1080 ();
 sg13g2_fill_8 FILLER_19_1107 ();
 sg13g2_fill_4 FILLER_19_1161 ();
 sg13g2_fill_8 FILLER_19_1195 ();
 sg13g2_fill_4 FILLER_19_1203 ();
 sg13g2_fill_2 FILLER_19_1248 ();
 sg13g2_fill_8 FILLER_19_1280 ();
 sg13g2_fill_8 FILLER_19_1288 ();
 sg13g2_fill_8 FILLER_19_1296 ();
 sg13g2_fill_8 FILLER_19_1304 ();
 sg13g2_fill_8 FILLER_19_1312 ();
 sg13g2_fill_8 FILLER_19_1320 ();
 sg13g2_fill_8 FILLER_19_1328 ();
 sg13g2_fill_8 FILLER_19_1336 ();
 sg13g2_fill_8 FILLER_19_1344 ();
 sg13g2_fill_8 FILLER_19_1352 ();
 sg13g2_fill_8 FILLER_19_1360 ();
 sg13g2_fill_8 FILLER_19_1368 ();
 sg13g2_fill_8 FILLER_19_1376 ();
 sg13g2_fill_8 FILLER_19_1384 ();
 sg13g2_fill_8 FILLER_19_1392 ();
 sg13g2_fill_8 FILLER_19_1400 ();
 sg13g2_fill_8 FILLER_19_1408 ();
 sg13g2_fill_8 FILLER_19_1416 ();
 sg13g2_fill_8 FILLER_19_1424 ();
 sg13g2_fill_8 FILLER_19_1432 ();
 sg13g2_fill_8 FILLER_19_1440 ();
 sg13g2_fill_8 FILLER_19_1448 ();
 sg13g2_fill_8 FILLER_19_1456 ();
 sg13g2_fill_8 FILLER_19_1464 ();
 sg13g2_fill_8 FILLER_19_1472 ();
 sg13g2_fill_8 FILLER_19_1480 ();
 sg13g2_fill_8 FILLER_19_1488 ();
 sg13g2_fill_8 FILLER_19_1496 ();
 sg13g2_fill_8 FILLER_19_1504 ();
 sg13g2_fill_8 FILLER_19_1512 ();
 sg13g2_fill_8 FILLER_19_1520 ();
 sg13g2_fill_8 FILLER_19_1528 ();
 sg13g2_fill_8 FILLER_19_1536 ();
 sg13g2_fill_8 FILLER_19_1544 ();
 sg13g2_fill_8 FILLER_19_1552 ();
 sg13g2_fill_8 FILLER_19_1560 ();
 sg13g2_fill_8 FILLER_19_1568 ();
 sg13g2_fill_8 FILLER_19_1576 ();
 sg13g2_fill_8 FILLER_19_1584 ();
 sg13g2_fill_8 FILLER_20_0 ();
 sg13g2_fill_8 FILLER_20_8 ();
 sg13g2_fill_8 FILLER_20_16 ();
 sg13g2_fill_8 FILLER_20_24 ();
 sg13g2_fill_8 FILLER_20_32 ();
 sg13g2_fill_8 FILLER_20_40 ();
 sg13g2_fill_8 FILLER_20_48 ();
 sg13g2_fill_8 FILLER_20_56 ();
 sg13g2_fill_8 FILLER_20_64 ();
 sg13g2_fill_8 FILLER_20_72 ();
 sg13g2_fill_8 FILLER_20_80 ();
 sg13g2_fill_8 FILLER_20_88 ();
 sg13g2_fill_8 FILLER_20_96 ();
 sg13g2_fill_8 FILLER_20_104 ();
 sg13g2_fill_8 FILLER_20_112 ();
 sg13g2_fill_8 FILLER_20_120 ();
 sg13g2_fill_8 FILLER_20_128 ();
 sg13g2_fill_8 FILLER_20_136 ();
 sg13g2_fill_8 FILLER_20_144 ();
 sg13g2_fill_8 FILLER_20_152 ();
 sg13g2_fill_8 FILLER_20_160 ();
 sg13g2_fill_8 FILLER_20_168 ();
 sg13g2_fill_8 FILLER_20_176 ();
 sg13g2_fill_8 FILLER_20_184 ();
 sg13g2_fill_8 FILLER_20_192 ();
 sg13g2_fill_8 FILLER_20_200 ();
 sg13g2_fill_8 FILLER_20_208 ();
 sg13g2_fill_8 FILLER_20_216 ();
 sg13g2_fill_8 FILLER_20_224 ();
 sg13g2_fill_8 FILLER_20_232 ();
 sg13g2_fill_8 FILLER_20_240 ();
 sg13g2_fill_8 FILLER_20_248 ();
 sg13g2_fill_8 FILLER_20_256 ();
 sg13g2_fill_8 FILLER_20_264 ();
 sg13g2_fill_8 FILLER_20_272 ();
 sg13g2_fill_8 FILLER_20_280 ();
 sg13g2_fill_8 FILLER_20_288 ();
 sg13g2_fill_8 FILLER_20_296 ();
 sg13g2_fill_8 FILLER_20_304 ();
 sg13g2_fill_8 FILLER_20_312 ();
 sg13g2_fill_8 FILLER_20_320 ();
 sg13g2_fill_8 FILLER_20_328 ();
 sg13g2_fill_8 FILLER_20_336 ();
 sg13g2_fill_8 FILLER_20_344 ();
 sg13g2_fill_8 FILLER_20_352 ();
 sg13g2_fill_8 FILLER_20_360 ();
 sg13g2_fill_8 FILLER_20_368 ();
 sg13g2_fill_4 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_fill_4 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_413 ();
 sg13g2_fill_2 FILLER_20_477 ();
 sg13g2_fill_1 FILLER_20_479 ();
 sg13g2_fill_8 FILLER_20_500 ();
 sg13g2_fill_2 FILLER_20_508 ();
 sg13g2_fill_8 FILLER_20_562 ();
 sg13g2_fill_4 FILLER_20_570 ();
 sg13g2_fill_2 FILLER_20_574 ();
 sg13g2_fill_4 FILLER_20_579 ();
 sg13g2_fill_1 FILLER_20_627 ();
 sg13g2_fill_8 FILLER_20_633 ();
 sg13g2_fill_4 FILLER_20_641 ();
 sg13g2_fill_2 FILLER_20_645 ();
 sg13g2_fill_1 FILLER_20_647 ();
 sg13g2_fill_8 FILLER_20_658 ();
 sg13g2_fill_8 FILLER_20_666 ();
 sg13g2_fill_8 FILLER_20_674 ();
 sg13g2_fill_4 FILLER_20_682 ();
 sg13g2_fill_2 FILLER_20_686 ();
 sg13g2_fill_8 FILLER_20_713 ();
 sg13g2_fill_8 FILLER_20_768 ();
 sg13g2_fill_8 FILLER_20_776 ();
 sg13g2_fill_2 FILLER_20_784 ();
 sg13g2_fill_4 FILLER_20_799 ();
 sg13g2_fill_8 FILLER_20_839 ();
 sg13g2_fill_2 FILLER_20_873 ();
 sg13g2_fill_8 FILLER_20_924 ();
 sg13g2_fill_8 FILLER_20_932 ();
 sg13g2_fill_8 FILLER_20_940 ();
 sg13g2_fill_4 FILLER_20_948 ();
 sg13g2_fill_2 FILLER_20_952 ();
 sg13g2_fill_8 FILLER_20_964 ();
 sg13g2_fill_8 FILLER_20_972 ();
 sg13g2_fill_2 FILLER_20_980 ();
 sg13g2_fill_1 FILLER_20_982 ();
 sg13g2_fill_8 FILLER_20_993 ();
 sg13g2_fill_8 FILLER_20_1001 ();
 sg13g2_fill_4 FILLER_20_1009 ();
 sg13g2_fill_2 FILLER_20_1013 ();
 sg13g2_fill_1 FILLER_20_1015 ();
 sg13g2_fill_8 FILLER_20_1047 ();
 sg13g2_fill_4 FILLER_20_1055 ();
 sg13g2_fill_2 FILLER_20_1059 ();
 sg13g2_fill_1 FILLER_20_1061 ();
 sg13g2_fill_8 FILLER_20_1070 ();
 sg13g2_fill_4 FILLER_20_1078 ();
 sg13g2_fill_2 FILLER_20_1082 ();
 sg13g2_fill_2 FILLER_20_1090 ();
 sg13g2_fill_1 FILLER_20_1092 ();
 sg13g2_fill_8 FILLER_20_1158 ();
 sg13g2_fill_8 FILLER_20_1166 ();
 sg13g2_fill_8 FILLER_20_1236 ();
 sg13g2_fill_1 FILLER_20_1244 ();
 sg13g2_fill_8 FILLER_20_1253 ();
 sg13g2_fill_8 FILLER_20_1261 ();
 sg13g2_fill_2 FILLER_20_1269 ();
 sg13g2_fill_8 FILLER_20_1284 ();
 sg13g2_fill_8 FILLER_20_1292 ();
 sg13g2_fill_8 FILLER_20_1300 ();
 sg13g2_fill_8 FILLER_20_1308 ();
 sg13g2_fill_8 FILLER_20_1316 ();
 sg13g2_fill_8 FILLER_20_1324 ();
 sg13g2_fill_8 FILLER_20_1332 ();
 sg13g2_fill_8 FILLER_20_1340 ();
 sg13g2_fill_8 FILLER_20_1348 ();
 sg13g2_fill_8 FILLER_20_1356 ();
 sg13g2_fill_8 FILLER_20_1364 ();
 sg13g2_fill_8 FILLER_20_1372 ();
 sg13g2_fill_8 FILLER_20_1380 ();
 sg13g2_fill_8 FILLER_20_1388 ();
 sg13g2_fill_8 FILLER_20_1396 ();
 sg13g2_fill_8 FILLER_20_1404 ();
 sg13g2_fill_8 FILLER_20_1412 ();
 sg13g2_fill_8 FILLER_20_1420 ();
 sg13g2_fill_8 FILLER_20_1428 ();
 sg13g2_fill_8 FILLER_20_1436 ();
 sg13g2_fill_8 FILLER_20_1444 ();
 sg13g2_fill_8 FILLER_20_1452 ();
 sg13g2_fill_8 FILLER_20_1460 ();
 sg13g2_fill_8 FILLER_20_1468 ();
 sg13g2_fill_8 FILLER_20_1476 ();
 sg13g2_fill_8 FILLER_20_1484 ();
 sg13g2_fill_8 FILLER_20_1492 ();
 sg13g2_fill_8 FILLER_20_1500 ();
 sg13g2_fill_8 FILLER_20_1508 ();
 sg13g2_fill_8 FILLER_20_1516 ();
 sg13g2_fill_8 FILLER_20_1524 ();
 sg13g2_fill_8 FILLER_20_1532 ();
 sg13g2_fill_8 FILLER_20_1540 ();
 sg13g2_fill_8 FILLER_20_1548 ();
 sg13g2_fill_8 FILLER_20_1556 ();
 sg13g2_fill_8 FILLER_20_1564 ();
 sg13g2_fill_8 FILLER_20_1572 ();
 sg13g2_fill_8 FILLER_20_1580 ();
 sg13g2_fill_4 FILLER_20_1588 ();
 sg13g2_fill_8 FILLER_21_0 ();
 sg13g2_fill_8 FILLER_21_8 ();
 sg13g2_fill_8 FILLER_21_16 ();
 sg13g2_fill_8 FILLER_21_24 ();
 sg13g2_fill_8 FILLER_21_32 ();
 sg13g2_fill_8 FILLER_21_40 ();
 sg13g2_fill_8 FILLER_21_48 ();
 sg13g2_fill_8 FILLER_21_56 ();
 sg13g2_fill_8 FILLER_21_64 ();
 sg13g2_fill_8 FILLER_21_72 ();
 sg13g2_fill_8 FILLER_21_80 ();
 sg13g2_fill_8 FILLER_21_88 ();
 sg13g2_fill_8 FILLER_21_96 ();
 sg13g2_fill_8 FILLER_21_104 ();
 sg13g2_fill_8 FILLER_21_112 ();
 sg13g2_fill_8 FILLER_21_120 ();
 sg13g2_fill_8 FILLER_21_128 ();
 sg13g2_fill_8 FILLER_21_136 ();
 sg13g2_fill_8 FILLER_21_144 ();
 sg13g2_fill_8 FILLER_21_152 ();
 sg13g2_fill_8 FILLER_21_160 ();
 sg13g2_fill_8 FILLER_21_168 ();
 sg13g2_fill_8 FILLER_21_176 ();
 sg13g2_fill_8 FILLER_21_184 ();
 sg13g2_fill_8 FILLER_21_192 ();
 sg13g2_fill_8 FILLER_21_200 ();
 sg13g2_fill_8 FILLER_21_208 ();
 sg13g2_fill_8 FILLER_21_216 ();
 sg13g2_fill_8 FILLER_21_224 ();
 sg13g2_fill_8 FILLER_21_232 ();
 sg13g2_fill_8 FILLER_21_240 ();
 sg13g2_fill_8 FILLER_21_248 ();
 sg13g2_fill_8 FILLER_21_256 ();
 sg13g2_fill_8 FILLER_21_264 ();
 sg13g2_fill_8 FILLER_21_272 ();
 sg13g2_fill_8 FILLER_21_280 ();
 sg13g2_fill_8 FILLER_21_288 ();
 sg13g2_fill_8 FILLER_21_296 ();
 sg13g2_fill_8 FILLER_21_304 ();
 sg13g2_fill_8 FILLER_21_312 ();
 sg13g2_fill_8 FILLER_21_320 ();
 sg13g2_fill_8 FILLER_21_328 ();
 sg13g2_fill_8 FILLER_21_336 ();
 sg13g2_fill_8 FILLER_21_344 ();
 sg13g2_fill_8 FILLER_21_352 ();
 sg13g2_fill_8 FILLER_21_360 ();
 sg13g2_fill_8 FILLER_21_368 ();
 sg13g2_fill_8 FILLER_21_376 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_fill_8 FILLER_21_423 ();
 sg13g2_fill_8 FILLER_21_431 ();
 sg13g2_fill_8 FILLER_21_439 ();
 sg13g2_fill_4 FILLER_21_447 ();
 sg13g2_fill_2 FILLER_21_451 ();
 sg13g2_fill_8 FILLER_21_505 ();
 sg13g2_fill_8 FILLER_21_548 ();
 sg13g2_fill_8 FILLER_21_556 ();
 sg13g2_fill_4 FILLER_21_564 ();
 sg13g2_fill_2 FILLER_21_568 ();
 sg13g2_fill_1 FILLER_21_570 ();
 sg13g2_fill_8 FILLER_21_606 ();
 sg13g2_fill_4 FILLER_21_614 ();
 sg13g2_fill_2 FILLER_21_618 ();
 sg13g2_fill_4 FILLER_21_632 ();
 sg13g2_fill_2 FILLER_21_666 ();
 sg13g2_fill_4 FILLER_21_748 ();
 sg13g2_fill_8 FILLER_21_788 ();
 sg13g2_fill_8 FILLER_21_796 ();
 sg13g2_fill_8 FILLER_21_804 ();
 sg13g2_fill_8 FILLER_21_812 ();
 sg13g2_fill_8 FILLER_21_820 ();
 sg13g2_fill_2 FILLER_21_828 ();
 sg13g2_fill_8 FILLER_21_885 ();
 sg13g2_fill_8 FILLER_21_893 ();
 sg13g2_fill_1 FILLER_21_901 ();
 sg13g2_fill_4 FILLER_21_928 ();
 sg13g2_fill_2 FILLER_21_932 ();
 sg13g2_fill_2 FILLER_21_964 ();
 sg13g2_fill_1 FILLER_21_966 ();
 sg13g2_fill_8 FILLER_21_1003 ();
 sg13g2_fill_4 FILLER_21_1011 ();
 sg13g2_fill_1 FILLER_21_1025 ();
 sg13g2_fill_8 FILLER_21_1030 ();
 sg13g2_fill_2 FILLER_21_1038 ();
 sg13g2_fill_1 FILLER_21_1040 ();
 sg13g2_fill_4 FILLER_21_1088 ();
 sg13g2_fill_1 FILLER_21_1092 ();
 sg13g2_fill_8 FILLER_21_1123 ();
 sg13g2_fill_8 FILLER_21_1131 ();
 sg13g2_fill_2 FILLER_21_1139 ();
 sg13g2_fill_1 FILLER_21_1157 ();
 sg13g2_fill_8 FILLER_21_1170 ();
 sg13g2_fill_8 FILLER_21_1178 ();
 sg13g2_fill_8 FILLER_21_1186 ();
 sg13g2_fill_1 FILLER_21_1194 ();
 sg13g2_fill_8 FILLER_21_1203 ();
 sg13g2_fill_8 FILLER_21_1211 ();
 sg13g2_fill_2 FILLER_21_1219 ();
 sg13g2_fill_1 FILLER_21_1221 ();
 sg13g2_fill_8 FILLER_21_1243 ();
 sg13g2_fill_4 FILLER_21_1251 ();
 sg13g2_fill_1 FILLER_21_1255 ();
 sg13g2_fill_1 FILLER_21_1270 ();
 sg13g2_fill_8 FILLER_21_1296 ();
 sg13g2_fill_8 FILLER_21_1304 ();
 sg13g2_fill_8 FILLER_21_1312 ();
 sg13g2_fill_8 FILLER_21_1320 ();
 sg13g2_fill_8 FILLER_21_1328 ();
 sg13g2_fill_8 FILLER_21_1336 ();
 sg13g2_fill_8 FILLER_21_1344 ();
 sg13g2_fill_8 FILLER_21_1352 ();
 sg13g2_fill_8 FILLER_21_1360 ();
 sg13g2_fill_8 FILLER_21_1368 ();
 sg13g2_fill_8 FILLER_21_1376 ();
 sg13g2_fill_8 FILLER_21_1384 ();
 sg13g2_fill_8 FILLER_21_1392 ();
 sg13g2_fill_8 FILLER_21_1400 ();
 sg13g2_fill_8 FILLER_21_1408 ();
 sg13g2_fill_8 FILLER_21_1416 ();
 sg13g2_fill_8 FILLER_21_1424 ();
 sg13g2_fill_8 FILLER_21_1432 ();
 sg13g2_fill_8 FILLER_21_1440 ();
 sg13g2_fill_8 FILLER_21_1448 ();
 sg13g2_fill_8 FILLER_21_1456 ();
 sg13g2_fill_8 FILLER_21_1464 ();
 sg13g2_fill_8 FILLER_21_1472 ();
 sg13g2_fill_8 FILLER_21_1480 ();
 sg13g2_fill_8 FILLER_21_1488 ();
 sg13g2_fill_8 FILLER_21_1496 ();
 sg13g2_fill_8 FILLER_21_1504 ();
 sg13g2_fill_8 FILLER_21_1512 ();
 sg13g2_fill_8 FILLER_21_1520 ();
 sg13g2_fill_8 FILLER_21_1528 ();
 sg13g2_fill_8 FILLER_21_1536 ();
 sg13g2_fill_8 FILLER_21_1544 ();
 sg13g2_fill_8 FILLER_21_1552 ();
 sg13g2_fill_8 FILLER_21_1560 ();
 sg13g2_fill_8 FILLER_21_1568 ();
 sg13g2_fill_8 FILLER_21_1576 ();
 sg13g2_fill_8 FILLER_21_1584 ();
 sg13g2_fill_8 FILLER_22_0 ();
 sg13g2_fill_8 FILLER_22_8 ();
 sg13g2_fill_8 FILLER_22_16 ();
 sg13g2_fill_8 FILLER_22_24 ();
 sg13g2_fill_8 FILLER_22_32 ();
 sg13g2_fill_8 FILLER_22_40 ();
 sg13g2_fill_8 FILLER_22_48 ();
 sg13g2_fill_8 FILLER_22_56 ();
 sg13g2_fill_8 FILLER_22_64 ();
 sg13g2_fill_8 FILLER_22_72 ();
 sg13g2_fill_8 FILLER_22_80 ();
 sg13g2_fill_8 FILLER_22_88 ();
 sg13g2_fill_8 FILLER_22_96 ();
 sg13g2_fill_8 FILLER_22_104 ();
 sg13g2_fill_8 FILLER_22_112 ();
 sg13g2_fill_8 FILLER_22_120 ();
 sg13g2_fill_8 FILLER_22_128 ();
 sg13g2_fill_8 FILLER_22_136 ();
 sg13g2_fill_8 FILLER_22_144 ();
 sg13g2_fill_8 FILLER_22_152 ();
 sg13g2_fill_8 FILLER_22_160 ();
 sg13g2_fill_8 FILLER_22_168 ();
 sg13g2_fill_8 FILLER_22_176 ();
 sg13g2_fill_8 FILLER_22_184 ();
 sg13g2_fill_8 FILLER_22_192 ();
 sg13g2_fill_8 FILLER_22_200 ();
 sg13g2_fill_8 FILLER_22_208 ();
 sg13g2_fill_8 FILLER_22_216 ();
 sg13g2_fill_8 FILLER_22_224 ();
 sg13g2_fill_8 FILLER_22_232 ();
 sg13g2_fill_8 FILLER_22_240 ();
 sg13g2_fill_8 FILLER_22_248 ();
 sg13g2_fill_8 FILLER_22_256 ();
 sg13g2_fill_8 FILLER_22_264 ();
 sg13g2_fill_8 FILLER_22_272 ();
 sg13g2_fill_8 FILLER_22_280 ();
 sg13g2_fill_8 FILLER_22_288 ();
 sg13g2_fill_8 FILLER_22_296 ();
 sg13g2_fill_8 FILLER_22_304 ();
 sg13g2_fill_8 FILLER_22_312 ();
 sg13g2_fill_8 FILLER_22_320 ();
 sg13g2_fill_8 FILLER_22_328 ();
 sg13g2_fill_8 FILLER_22_336 ();
 sg13g2_fill_8 FILLER_22_344 ();
 sg13g2_fill_8 FILLER_22_352 ();
 sg13g2_fill_8 FILLER_22_360 ();
 sg13g2_fill_8 FILLER_22_368 ();
 sg13g2_fill_8 FILLER_22_376 ();
 sg13g2_fill_8 FILLER_22_390 ();
 sg13g2_fill_8 FILLER_22_398 ();
 sg13g2_fill_4 FILLER_22_416 ();
 sg13g2_fill_2 FILLER_22_420 ();
 sg13g2_fill_4 FILLER_22_458 ();
 sg13g2_fill_2 FILLER_22_462 ();
 sg13g2_fill_1 FILLER_22_464 ();
 sg13g2_fill_8 FILLER_22_513 ();
 sg13g2_fill_8 FILLER_22_521 ();
 sg13g2_fill_8 FILLER_22_529 ();
 sg13g2_fill_1 FILLER_22_537 ();
 sg13g2_fill_8 FILLER_22_564 ();
 sg13g2_fill_8 FILLER_22_572 ();
 sg13g2_fill_8 FILLER_22_580 ();
 sg13g2_fill_8 FILLER_22_588 ();
 sg13g2_fill_8 FILLER_22_596 ();
 sg13g2_fill_2 FILLER_22_604 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_fill_8 FILLER_22_634 ();
 sg13g2_fill_8 FILLER_22_642 ();
 sg13g2_fill_8 FILLER_22_650 ();
 sg13g2_fill_8 FILLER_22_658 ();
 sg13g2_fill_8 FILLER_22_666 ();
 sg13g2_fill_2 FILLER_22_674 ();
 sg13g2_fill_1 FILLER_22_681 ();
 sg13g2_fill_4 FILLER_22_689 ();
 sg13g2_fill_2 FILLER_22_693 ();
 sg13g2_fill_1 FILLER_22_695 ();
 sg13g2_fill_8 FILLER_22_722 ();
 sg13g2_fill_1 FILLER_22_730 ();
 sg13g2_fill_8 FILLER_22_736 ();
 sg13g2_fill_2 FILLER_22_744 ();
 sg13g2_fill_2 FILLER_22_790 ();
 sg13g2_fill_4 FILLER_22_836 ();
 sg13g2_fill_4 FILLER_22_866 ();
 sg13g2_fill_1 FILLER_22_870 ();
 sg13g2_fill_1 FILLER_22_922 ();
 sg13g2_fill_8 FILLER_22_949 ();
 sg13g2_fill_4 FILLER_22_957 ();
 sg13g2_fill_1 FILLER_22_961 ();
 sg13g2_fill_2 FILLER_22_967 ();
 sg13g2_fill_8 FILLER_22_979 ();
 sg13g2_fill_8 FILLER_22_987 ();
 sg13g2_fill_4 FILLER_22_995 ();
 sg13g2_fill_2 FILLER_22_999 ();
 sg13g2_fill_4 FILLER_22_1027 ();
 sg13g2_fill_2 FILLER_22_1031 ();
 sg13g2_fill_1 FILLER_22_1033 ();
 sg13g2_fill_1 FILLER_22_1083 ();
 sg13g2_fill_8 FILLER_22_1094 ();
 sg13g2_fill_8 FILLER_22_1102 ();
 sg13g2_fill_8 FILLER_22_1110 ();
 sg13g2_fill_8 FILLER_22_1118 ();
 sg13g2_fill_1 FILLER_22_1126 ();
 sg13g2_fill_2 FILLER_22_1166 ();
 sg13g2_fill_8 FILLER_22_1182 ();
 sg13g2_fill_2 FILLER_22_1190 ();
 sg13g2_fill_1 FILLER_22_1192 ();
 sg13g2_fill_8 FILLER_22_1201 ();
 sg13g2_fill_1 FILLER_22_1209 ();
 sg13g2_fill_4 FILLER_22_1220 ();
 sg13g2_fill_1 FILLER_22_1224 ();
 sg13g2_fill_8 FILLER_22_1297 ();
 sg13g2_fill_8 FILLER_22_1305 ();
 sg13g2_fill_8 FILLER_22_1313 ();
 sg13g2_fill_8 FILLER_22_1321 ();
 sg13g2_fill_8 FILLER_22_1329 ();
 sg13g2_fill_8 FILLER_22_1337 ();
 sg13g2_fill_8 FILLER_22_1345 ();
 sg13g2_fill_8 FILLER_22_1353 ();
 sg13g2_fill_8 FILLER_22_1361 ();
 sg13g2_fill_8 FILLER_22_1369 ();
 sg13g2_fill_8 FILLER_22_1377 ();
 sg13g2_fill_8 FILLER_22_1385 ();
 sg13g2_fill_8 FILLER_22_1393 ();
 sg13g2_fill_8 FILLER_22_1401 ();
 sg13g2_fill_8 FILLER_22_1409 ();
 sg13g2_fill_8 FILLER_22_1417 ();
 sg13g2_fill_8 FILLER_22_1425 ();
 sg13g2_fill_8 FILLER_22_1433 ();
 sg13g2_fill_8 FILLER_22_1441 ();
 sg13g2_fill_8 FILLER_22_1449 ();
 sg13g2_fill_8 FILLER_22_1457 ();
 sg13g2_fill_8 FILLER_22_1465 ();
 sg13g2_fill_8 FILLER_22_1473 ();
 sg13g2_fill_8 FILLER_22_1481 ();
 sg13g2_fill_8 FILLER_22_1489 ();
 sg13g2_fill_8 FILLER_22_1497 ();
 sg13g2_fill_8 FILLER_22_1505 ();
 sg13g2_fill_8 FILLER_22_1513 ();
 sg13g2_fill_8 FILLER_22_1521 ();
 sg13g2_fill_8 FILLER_22_1529 ();
 sg13g2_fill_8 FILLER_22_1537 ();
 sg13g2_fill_8 FILLER_22_1545 ();
 sg13g2_fill_8 FILLER_22_1553 ();
 sg13g2_fill_8 FILLER_22_1561 ();
 sg13g2_fill_8 FILLER_22_1569 ();
 sg13g2_fill_8 FILLER_22_1577 ();
 sg13g2_fill_4 FILLER_22_1585 ();
 sg13g2_fill_2 FILLER_22_1589 ();
 sg13g2_fill_1 FILLER_22_1591 ();
 sg13g2_fill_8 FILLER_23_0 ();
 sg13g2_fill_8 FILLER_23_8 ();
 sg13g2_fill_8 FILLER_23_16 ();
 sg13g2_fill_8 FILLER_23_24 ();
 sg13g2_fill_8 FILLER_23_32 ();
 sg13g2_fill_8 FILLER_23_40 ();
 sg13g2_fill_8 FILLER_23_48 ();
 sg13g2_fill_8 FILLER_23_56 ();
 sg13g2_fill_8 FILLER_23_64 ();
 sg13g2_fill_8 FILLER_23_72 ();
 sg13g2_fill_8 FILLER_23_80 ();
 sg13g2_fill_8 FILLER_23_88 ();
 sg13g2_fill_8 FILLER_23_96 ();
 sg13g2_fill_8 FILLER_23_104 ();
 sg13g2_fill_8 FILLER_23_112 ();
 sg13g2_fill_8 FILLER_23_120 ();
 sg13g2_fill_8 FILLER_23_128 ();
 sg13g2_fill_8 FILLER_23_136 ();
 sg13g2_fill_8 FILLER_23_144 ();
 sg13g2_fill_8 FILLER_23_152 ();
 sg13g2_fill_8 FILLER_23_160 ();
 sg13g2_fill_8 FILLER_23_168 ();
 sg13g2_fill_8 FILLER_23_176 ();
 sg13g2_fill_8 FILLER_23_184 ();
 sg13g2_fill_8 FILLER_23_192 ();
 sg13g2_fill_8 FILLER_23_200 ();
 sg13g2_fill_8 FILLER_23_208 ();
 sg13g2_fill_8 FILLER_23_216 ();
 sg13g2_fill_8 FILLER_23_224 ();
 sg13g2_fill_8 FILLER_23_232 ();
 sg13g2_fill_8 FILLER_23_240 ();
 sg13g2_fill_8 FILLER_23_248 ();
 sg13g2_fill_8 FILLER_23_256 ();
 sg13g2_fill_8 FILLER_23_264 ();
 sg13g2_fill_8 FILLER_23_272 ();
 sg13g2_fill_8 FILLER_23_280 ();
 sg13g2_fill_8 FILLER_23_288 ();
 sg13g2_fill_8 FILLER_23_296 ();
 sg13g2_fill_8 FILLER_23_304 ();
 sg13g2_fill_8 FILLER_23_312 ();
 sg13g2_fill_8 FILLER_23_320 ();
 sg13g2_fill_8 FILLER_23_328 ();
 sg13g2_fill_8 FILLER_23_336 ();
 sg13g2_fill_8 FILLER_23_344 ();
 sg13g2_fill_8 FILLER_23_352 ();
 sg13g2_fill_8 FILLER_23_360 ();
 sg13g2_fill_4 FILLER_23_368 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_fill_8 FILLER_23_419 ();
 sg13g2_fill_4 FILLER_23_427 ();
 sg13g2_fill_8 FILLER_23_441 ();
 sg13g2_fill_8 FILLER_23_449 ();
 sg13g2_fill_2 FILLER_23_457 ();
 sg13g2_fill_1 FILLER_23_459 ();
 sg13g2_fill_8 FILLER_23_470 ();
 sg13g2_fill_4 FILLER_23_504 ();
 sg13g2_fill_2 FILLER_23_600 ();
 sg13g2_fill_1 FILLER_23_607 ();
 sg13g2_fill_8 FILLER_23_617 ();
 sg13g2_fill_1 FILLER_23_630 ();
 sg13g2_fill_2 FILLER_23_659 ();
 sg13g2_fill_1 FILLER_23_661 ();
 sg13g2_fill_8 FILLER_23_690 ();
 sg13g2_fill_8 FILLER_23_698 ();
 sg13g2_fill_2 FILLER_23_706 ();
 sg13g2_fill_1 FILLER_23_708 ();
 sg13g2_fill_2 FILLER_23_719 ();
 sg13g2_fill_8 FILLER_23_727 ();
 sg13g2_fill_8 FILLER_23_735 ();
 sg13g2_fill_1 FILLER_23_743 ();
 sg13g2_fill_2 FILLER_23_754 ();
 sg13g2_fill_8 FILLER_23_802 ();
 sg13g2_fill_8 FILLER_23_810 ();
 sg13g2_fill_8 FILLER_23_818 ();
 sg13g2_fill_8 FILLER_23_826 ();
 sg13g2_fill_4 FILLER_23_834 ();
 sg13g2_fill_2 FILLER_23_838 ();
 sg13g2_fill_8 FILLER_23_850 ();
 sg13g2_fill_4 FILLER_23_858 ();
 sg13g2_fill_4 FILLER_23_888 ();
 sg13g2_fill_2 FILLER_23_892 ();
 sg13g2_fill_1 FILLER_23_894 ();
 sg13g2_fill_4 FILLER_23_935 ();
 sg13g2_fill_2 FILLER_23_970 ();
 sg13g2_fill_1 FILLER_23_972 ();
 sg13g2_fill_2 FILLER_23_999 ();
 sg13g2_fill_8 FILLER_23_1011 ();
 sg13g2_fill_8 FILLER_23_1019 ();
 sg13g2_fill_1 FILLER_23_1027 ();
 sg13g2_fill_1 FILLER_23_1064 ();
 sg13g2_fill_4 FILLER_23_1069 ();
 sg13g2_fill_4 FILLER_23_1099 ();
 sg13g2_fill_2 FILLER_23_1103 ();
 sg13g2_fill_8 FILLER_23_1145 ();
 sg13g2_fill_8 FILLER_23_1153 ();
 sg13g2_fill_2 FILLER_23_1161 ();
 sg13g2_fill_1 FILLER_23_1203 ();
 sg13g2_fill_8 FILLER_23_1238 ();
 sg13g2_fill_8 FILLER_23_1246 ();
 sg13g2_fill_4 FILLER_23_1254 ();
 sg13g2_fill_2 FILLER_23_1258 ();
 sg13g2_fill_1 FILLER_23_1268 ();
 sg13g2_fill_8 FILLER_23_1299 ();
 sg13g2_fill_8 FILLER_23_1307 ();
 sg13g2_fill_8 FILLER_23_1315 ();
 sg13g2_fill_8 FILLER_23_1323 ();
 sg13g2_fill_8 FILLER_23_1331 ();
 sg13g2_fill_8 FILLER_23_1339 ();
 sg13g2_fill_8 FILLER_23_1347 ();
 sg13g2_fill_8 FILLER_23_1355 ();
 sg13g2_fill_8 FILLER_23_1363 ();
 sg13g2_fill_8 FILLER_23_1371 ();
 sg13g2_fill_8 FILLER_23_1379 ();
 sg13g2_fill_8 FILLER_23_1387 ();
 sg13g2_fill_8 FILLER_23_1395 ();
 sg13g2_fill_8 FILLER_23_1403 ();
 sg13g2_fill_8 FILLER_23_1411 ();
 sg13g2_fill_8 FILLER_23_1419 ();
 sg13g2_fill_8 FILLER_23_1427 ();
 sg13g2_fill_8 FILLER_23_1435 ();
 sg13g2_fill_8 FILLER_23_1443 ();
 sg13g2_fill_8 FILLER_23_1451 ();
 sg13g2_fill_8 FILLER_23_1459 ();
 sg13g2_fill_8 FILLER_23_1467 ();
 sg13g2_fill_8 FILLER_23_1475 ();
 sg13g2_fill_8 FILLER_23_1483 ();
 sg13g2_fill_8 FILLER_23_1491 ();
 sg13g2_fill_8 FILLER_23_1499 ();
 sg13g2_fill_8 FILLER_23_1507 ();
 sg13g2_fill_8 FILLER_23_1515 ();
 sg13g2_fill_8 FILLER_23_1523 ();
 sg13g2_fill_8 FILLER_23_1531 ();
 sg13g2_fill_8 FILLER_23_1539 ();
 sg13g2_fill_8 FILLER_23_1547 ();
 sg13g2_fill_8 FILLER_23_1555 ();
 sg13g2_fill_8 FILLER_23_1563 ();
 sg13g2_fill_8 FILLER_23_1571 ();
 sg13g2_fill_8 FILLER_23_1579 ();
 sg13g2_fill_4 FILLER_23_1587 ();
 sg13g2_fill_1 FILLER_23_1591 ();
 sg13g2_fill_8 FILLER_24_0 ();
 sg13g2_fill_8 FILLER_24_8 ();
 sg13g2_fill_8 FILLER_24_16 ();
 sg13g2_fill_8 FILLER_24_24 ();
 sg13g2_fill_8 FILLER_24_32 ();
 sg13g2_fill_8 FILLER_24_40 ();
 sg13g2_fill_8 FILLER_24_48 ();
 sg13g2_fill_8 FILLER_24_56 ();
 sg13g2_fill_8 FILLER_24_64 ();
 sg13g2_fill_8 FILLER_24_72 ();
 sg13g2_fill_8 FILLER_24_80 ();
 sg13g2_fill_8 FILLER_24_88 ();
 sg13g2_fill_8 FILLER_24_96 ();
 sg13g2_fill_8 FILLER_24_104 ();
 sg13g2_fill_8 FILLER_24_112 ();
 sg13g2_fill_8 FILLER_24_120 ();
 sg13g2_fill_8 FILLER_24_128 ();
 sg13g2_fill_8 FILLER_24_136 ();
 sg13g2_fill_8 FILLER_24_144 ();
 sg13g2_fill_8 FILLER_24_152 ();
 sg13g2_fill_8 FILLER_24_160 ();
 sg13g2_fill_8 FILLER_24_168 ();
 sg13g2_fill_8 FILLER_24_176 ();
 sg13g2_fill_8 FILLER_24_184 ();
 sg13g2_fill_8 FILLER_24_192 ();
 sg13g2_fill_8 FILLER_24_200 ();
 sg13g2_fill_8 FILLER_24_208 ();
 sg13g2_fill_8 FILLER_24_216 ();
 sg13g2_fill_8 FILLER_24_224 ();
 sg13g2_fill_8 FILLER_24_232 ();
 sg13g2_fill_8 FILLER_24_240 ();
 sg13g2_fill_8 FILLER_24_248 ();
 sg13g2_fill_8 FILLER_24_256 ();
 sg13g2_fill_8 FILLER_24_264 ();
 sg13g2_fill_8 FILLER_24_272 ();
 sg13g2_fill_8 FILLER_24_280 ();
 sg13g2_fill_8 FILLER_24_288 ();
 sg13g2_fill_8 FILLER_24_296 ();
 sg13g2_fill_8 FILLER_24_304 ();
 sg13g2_fill_8 FILLER_24_312 ();
 sg13g2_fill_8 FILLER_24_320 ();
 sg13g2_fill_8 FILLER_24_328 ();
 sg13g2_fill_8 FILLER_24_336 ();
 sg13g2_fill_8 FILLER_24_344 ();
 sg13g2_fill_8 FILLER_24_352 ();
 sg13g2_fill_1 FILLER_24_360 ();
 sg13g2_fill_1 FILLER_24_413 ();
 sg13g2_fill_2 FILLER_24_424 ();
 sg13g2_fill_8 FILLER_24_488 ();
 sg13g2_fill_4 FILLER_24_496 ();
 sg13g2_fill_4 FILLER_24_536 ();
 sg13g2_fill_2 FILLER_24_540 ();
 sg13g2_fill_1 FILLER_24_542 ();
 sg13g2_fill_8 FILLER_24_553 ();
 sg13g2_fill_1 FILLER_24_561 ();
 sg13g2_fill_8 FILLER_24_567 ();
 sg13g2_fill_4 FILLER_24_575 ();
 sg13g2_fill_1 FILLER_24_579 ();
 sg13g2_fill_1 FILLER_24_625 ();
 sg13g2_fill_2 FILLER_24_631 ();
 sg13g2_fill_1 FILLER_24_633 ();
 sg13g2_fill_4 FILLER_24_644 ();
 sg13g2_fill_2 FILLER_24_687 ();
 sg13g2_fill_4 FILLER_24_719 ();
 sg13g2_fill_1 FILLER_24_723 ();
 sg13g2_fill_8 FILLER_24_782 ();
 sg13g2_fill_8 FILLER_24_790 ();
 sg13g2_fill_2 FILLER_24_798 ();
 sg13g2_fill_1 FILLER_24_800 ();
 sg13g2_fill_8 FILLER_24_837 ();
 sg13g2_fill_8 FILLER_24_845 ();
 sg13g2_fill_4 FILLER_24_853 ();
 sg13g2_fill_2 FILLER_24_857 ();
 sg13g2_fill_8 FILLER_24_869 ();
 sg13g2_fill_8 FILLER_24_877 ();
 sg13g2_fill_2 FILLER_24_890 ();
 sg13g2_fill_8 FILLER_24_927 ();
 sg13g2_fill_8 FILLER_24_935 ();
 sg13g2_fill_4 FILLER_24_943 ();
 sg13g2_fill_2 FILLER_24_947 ();
 sg13g2_fill_1 FILLER_24_949 ();
 sg13g2_fill_8 FILLER_24_975 ();
 sg13g2_fill_8 FILLER_24_983 ();
 sg13g2_fill_8 FILLER_24_991 ();
 sg13g2_fill_4 FILLER_24_999 ();
 sg13g2_fill_2 FILLER_24_1003 ();
 sg13g2_fill_1 FILLER_24_1005 ();
 sg13g2_fill_8 FILLER_24_1057 ();
 sg13g2_fill_8 FILLER_24_1065 ();
 sg13g2_fill_2 FILLER_24_1081 ();
 sg13g2_fill_1 FILLER_24_1083 ();
 sg13g2_fill_4 FILLER_24_1087 ();
 sg13g2_fill_2 FILLER_24_1091 ();
 sg13g2_fill_4 FILLER_24_1098 ();
 sg13g2_fill_1 FILLER_24_1102 ();
 sg13g2_fill_8 FILLER_24_1114 ();
 sg13g2_fill_8 FILLER_24_1122 ();
 sg13g2_fill_8 FILLER_24_1130 ();
 sg13g2_fill_4 FILLER_24_1138 ();
 sg13g2_fill_1 FILLER_24_1142 ();
 sg13g2_fill_8 FILLER_24_1153 ();
 sg13g2_fill_4 FILLER_24_1161 ();
 sg13g2_fill_2 FILLER_24_1165 ();
 sg13g2_fill_1 FILLER_24_1167 ();
 sg13g2_fill_8 FILLER_24_1172 ();
 sg13g2_fill_4 FILLER_24_1180 ();
 sg13g2_fill_4 FILLER_24_1189 ();
 sg13g2_fill_1 FILLER_24_1193 ();
 sg13g2_fill_8 FILLER_24_1199 ();
 sg13g2_fill_8 FILLER_24_1207 ();
 sg13g2_fill_8 FILLER_24_1215 ();
 sg13g2_fill_1 FILLER_24_1223 ();
 sg13g2_fill_8 FILLER_24_1229 ();
 sg13g2_fill_8 FILLER_24_1237 ();
 sg13g2_fill_8 FILLER_24_1245 ();
 sg13g2_fill_4 FILLER_24_1253 ();
 sg13g2_fill_8 FILLER_24_1263 ();
 sg13g2_fill_8 FILLER_24_1271 ();
 sg13g2_fill_8 FILLER_24_1279 ();
 sg13g2_fill_8 FILLER_24_1287 ();
 sg13g2_fill_8 FILLER_24_1295 ();
 sg13g2_fill_8 FILLER_24_1303 ();
 sg13g2_fill_8 FILLER_24_1311 ();
 sg13g2_fill_8 FILLER_24_1319 ();
 sg13g2_fill_8 FILLER_24_1327 ();
 sg13g2_fill_8 FILLER_24_1335 ();
 sg13g2_fill_8 FILLER_24_1343 ();
 sg13g2_fill_8 FILLER_24_1351 ();
 sg13g2_fill_8 FILLER_24_1359 ();
 sg13g2_fill_8 FILLER_24_1367 ();
 sg13g2_fill_8 FILLER_24_1375 ();
 sg13g2_fill_8 FILLER_24_1383 ();
 sg13g2_fill_8 FILLER_24_1391 ();
 sg13g2_fill_8 FILLER_24_1399 ();
 sg13g2_fill_8 FILLER_24_1407 ();
 sg13g2_fill_8 FILLER_24_1415 ();
 sg13g2_fill_8 FILLER_24_1423 ();
 sg13g2_fill_8 FILLER_24_1431 ();
 sg13g2_fill_8 FILLER_24_1439 ();
 sg13g2_fill_8 FILLER_24_1447 ();
 sg13g2_fill_8 FILLER_24_1455 ();
 sg13g2_fill_8 FILLER_24_1463 ();
 sg13g2_fill_8 FILLER_24_1471 ();
 sg13g2_fill_8 FILLER_24_1479 ();
 sg13g2_fill_8 FILLER_24_1487 ();
 sg13g2_fill_8 FILLER_24_1495 ();
 sg13g2_fill_8 FILLER_24_1503 ();
 sg13g2_fill_8 FILLER_24_1511 ();
 sg13g2_fill_8 FILLER_24_1519 ();
 sg13g2_fill_8 FILLER_24_1527 ();
 sg13g2_fill_8 FILLER_24_1535 ();
 sg13g2_fill_8 FILLER_24_1543 ();
 sg13g2_fill_8 FILLER_24_1551 ();
 sg13g2_fill_8 FILLER_24_1559 ();
 sg13g2_fill_8 FILLER_24_1567 ();
 sg13g2_fill_8 FILLER_24_1575 ();
 sg13g2_fill_8 FILLER_24_1583 ();
 sg13g2_fill_1 FILLER_24_1591 ();
 sg13g2_fill_8 FILLER_25_0 ();
 sg13g2_fill_8 FILLER_25_8 ();
 sg13g2_fill_8 FILLER_25_16 ();
 sg13g2_fill_8 FILLER_25_24 ();
 sg13g2_fill_8 FILLER_25_32 ();
 sg13g2_fill_8 FILLER_25_40 ();
 sg13g2_fill_8 FILLER_25_48 ();
 sg13g2_fill_8 FILLER_25_56 ();
 sg13g2_fill_8 FILLER_25_64 ();
 sg13g2_fill_8 FILLER_25_72 ();
 sg13g2_fill_8 FILLER_25_80 ();
 sg13g2_fill_8 FILLER_25_88 ();
 sg13g2_fill_8 FILLER_25_96 ();
 sg13g2_fill_8 FILLER_25_104 ();
 sg13g2_fill_8 FILLER_25_112 ();
 sg13g2_fill_8 FILLER_25_120 ();
 sg13g2_fill_8 FILLER_25_128 ();
 sg13g2_fill_8 FILLER_25_136 ();
 sg13g2_fill_8 FILLER_25_144 ();
 sg13g2_fill_8 FILLER_25_152 ();
 sg13g2_fill_8 FILLER_25_160 ();
 sg13g2_fill_8 FILLER_25_168 ();
 sg13g2_fill_8 FILLER_25_176 ();
 sg13g2_fill_8 FILLER_25_184 ();
 sg13g2_fill_8 FILLER_25_192 ();
 sg13g2_fill_8 FILLER_25_200 ();
 sg13g2_fill_8 FILLER_25_208 ();
 sg13g2_fill_8 FILLER_25_216 ();
 sg13g2_fill_8 FILLER_25_224 ();
 sg13g2_fill_8 FILLER_25_232 ();
 sg13g2_fill_8 FILLER_25_240 ();
 sg13g2_fill_8 FILLER_25_248 ();
 sg13g2_fill_8 FILLER_25_256 ();
 sg13g2_fill_8 FILLER_25_264 ();
 sg13g2_fill_8 FILLER_25_272 ();
 sg13g2_fill_8 FILLER_25_280 ();
 sg13g2_fill_8 FILLER_25_288 ();
 sg13g2_fill_8 FILLER_25_296 ();
 sg13g2_fill_8 FILLER_25_304 ();
 sg13g2_fill_8 FILLER_25_312 ();
 sg13g2_fill_8 FILLER_25_320 ();
 sg13g2_fill_8 FILLER_25_328 ();
 sg13g2_fill_8 FILLER_25_336 ();
 sg13g2_fill_8 FILLER_25_344 ();
 sg13g2_fill_4 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_356 ();
 sg13g2_fill_8 FILLER_25_384 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_fill_1 FILLER_25_419 ();
 sg13g2_fill_8 FILLER_25_430 ();
 sg13g2_fill_8 FILLER_25_438 ();
 sg13g2_fill_8 FILLER_25_446 ();
 sg13g2_fill_8 FILLER_25_454 ();
 sg13g2_fill_8 FILLER_25_467 ();
 sg13g2_fill_4 FILLER_25_475 ();
 sg13g2_fill_8 FILLER_25_489 ();
 sg13g2_fill_8 FILLER_25_497 ();
 sg13g2_fill_1 FILLER_25_505 ();
 sg13g2_fill_8 FILLER_25_516 ();
 sg13g2_fill_8 FILLER_25_524 ();
 sg13g2_fill_8 FILLER_25_532 ();
 sg13g2_fill_2 FILLER_25_540 ();
 sg13g2_fill_1 FILLER_25_542 ();
 sg13g2_fill_8 FILLER_25_594 ();
 sg13g2_fill_8 FILLER_25_602 ();
 sg13g2_fill_2 FILLER_25_610 ();
 sg13g2_fill_8 FILLER_25_616 ();
 sg13g2_fill_4 FILLER_25_624 ();
 sg13g2_fill_2 FILLER_25_633 ();
 sg13g2_fill_8 FILLER_25_639 ();
 sg13g2_fill_4 FILLER_25_647 ();
 sg13g2_fill_2 FILLER_25_651 ();
 sg13g2_fill_8 FILLER_25_657 ();
 sg13g2_fill_8 FILLER_25_665 ();
 sg13g2_fill_4 FILLER_25_673 ();
 sg13g2_fill_1 FILLER_25_677 ();
 sg13g2_fill_8 FILLER_25_703 ();
 sg13g2_fill_8 FILLER_25_711 ();
 sg13g2_fill_8 FILLER_25_719 ();
 sg13g2_fill_8 FILLER_25_727 ();
 sg13g2_fill_8 FILLER_25_735 ();
 sg13g2_fill_2 FILLER_25_743 ();
 sg13g2_fill_4 FILLER_25_754 ();
 sg13g2_fill_2 FILLER_25_758 ();
 sg13g2_fill_4 FILLER_25_764 ();
 sg13g2_fill_2 FILLER_25_802 ();
 sg13g2_fill_2 FILLER_25_830 ();
 sg13g2_fill_8 FILLER_25_862 ();
 sg13g2_fill_8 FILLER_25_870 ();
 sg13g2_fill_2 FILLER_25_878 ();
 sg13g2_fill_8 FILLER_25_944 ();
 sg13g2_fill_2 FILLER_25_952 ();
 sg13g2_fill_1 FILLER_25_954 ();
 sg13g2_fill_1 FILLER_25_970 ();
 sg13g2_fill_8 FILLER_25_1007 ();
 sg13g2_fill_8 FILLER_25_1015 ();
 sg13g2_fill_8 FILLER_25_1023 ();
 sg13g2_fill_1 FILLER_25_1031 ();
 sg13g2_fill_2 FILLER_25_1052 ();
 sg13g2_fill_4 FILLER_25_1058 ();
 sg13g2_fill_2 FILLER_25_1062 ();
 sg13g2_fill_4 FILLER_25_1070 ();
 sg13g2_fill_2 FILLER_25_1074 ();
 sg13g2_fill_2 FILLER_25_1081 ();
 sg13g2_fill_1 FILLER_25_1083 ();
 sg13g2_fill_8 FILLER_25_1088 ();
 sg13g2_fill_1 FILLER_25_1096 ();
 sg13g2_fill_1 FILLER_25_1105 ();
 sg13g2_fill_4 FILLER_25_1110 ();
 sg13g2_fill_1 FILLER_25_1114 ();
 sg13g2_fill_2 FILLER_25_1207 ();
 sg13g2_fill_1 FILLER_25_1209 ();
 sg13g2_fill_8 FILLER_25_1215 ();
 sg13g2_fill_1 FILLER_25_1223 ();
 sg13g2_fill_1 FILLER_25_1266 ();
 sg13g2_fill_8 FILLER_25_1297 ();
 sg13g2_fill_8 FILLER_25_1305 ();
 sg13g2_fill_8 FILLER_25_1313 ();
 sg13g2_fill_8 FILLER_25_1321 ();
 sg13g2_fill_8 FILLER_25_1329 ();
 sg13g2_fill_8 FILLER_25_1337 ();
 sg13g2_fill_8 FILLER_25_1345 ();
 sg13g2_fill_8 FILLER_25_1353 ();
 sg13g2_fill_8 FILLER_25_1361 ();
 sg13g2_fill_8 FILLER_25_1369 ();
 sg13g2_fill_8 FILLER_25_1377 ();
 sg13g2_fill_8 FILLER_25_1385 ();
 sg13g2_fill_8 FILLER_25_1393 ();
 sg13g2_fill_8 FILLER_25_1401 ();
 sg13g2_fill_8 FILLER_25_1409 ();
 sg13g2_fill_8 FILLER_25_1417 ();
 sg13g2_fill_8 FILLER_25_1425 ();
 sg13g2_fill_8 FILLER_25_1433 ();
 sg13g2_fill_8 FILLER_25_1441 ();
 sg13g2_fill_8 FILLER_25_1449 ();
 sg13g2_fill_8 FILLER_25_1457 ();
 sg13g2_fill_8 FILLER_25_1465 ();
 sg13g2_fill_8 FILLER_25_1473 ();
 sg13g2_fill_8 FILLER_25_1481 ();
 sg13g2_fill_8 FILLER_25_1489 ();
 sg13g2_fill_8 FILLER_25_1497 ();
 sg13g2_fill_8 FILLER_25_1505 ();
 sg13g2_fill_8 FILLER_25_1513 ();
 sg13g2_fill_8 FILLER_25_1521 ();
 sg13g2_fill_8 FILLER_25_1529 ();
 sg13g2_fill_8 FILLER_25_1537 ();
 sg13g2_fill_8 FILLER_25_1545 ();
 sg13g2_fill_8 FILLER_25_1553 ();
 sg13g2_fill_8 FILLER_25_1561 ();
 sg13g2_fill_8 FILLER_25_1569 ();
 sg13g2_fill_8 FILLER_25_1577 ();
 sg13g2_fill_4 FILLER_25_1585 ();
 sg13g2_fill_2 FILLER_25_1589 ();
 sg13g2_fill_1 FILLER_25_1591 ();
 sg13g2_fill_8 FILLER_26_0 ();
 sg13g2_fill_8 FILLER_26_8 ();
 sg13g2_fill_8 FILLER_26_16 ();
 sg13g2_fill_8 FILLER_26_24 ();
 sg13g2_fill_8 FILLER_26_32 ();
 sg13g2_fill_8 FILLER_26_40 ();
 sg13g2_fill_8 FILLER_26_48 ();
 sg13g2_fill_8 FILLER_26_56 ();
 sg13g2_fill_8 FILLER_26_64 ();
 sg13g2_fill_8 FILLER_26_72 ();
 sg13g2_fill_8 FILLER_26_80 ();
 sg13g2_fill_8 FILLER_26_88 ();
 sg13g2_fill_8 FILLER_26_96 ();
 sg13g2_fill_8 FILLER_26_104 ();
 sg13g2_fill_8 FILLER_26_112 ();
 sg13g2_fill_8 FILLER_26_120 ();
 sg13g2_fill_8 FILLER_26_128 ();
 sg13g2_fill_8 FILLER_26_136 ();
 sg13g2_fill_8 FILLER_26_144 ();
 sg13g2_fill_8 FILLER_26_152 ();
 sg13g2_fill_8 FILLER_26_160 ();
 sg13g2_fill_8 FILLER_26_168 ();
 sg13g2_fill_8 FILLER_26_176 ();
 sg13g2_fill_8 FILLER_26_184 ();
 sg13g2_fill_8 FILLER_26_192 ();
 sg13g2_fill_8 FILLER_26_200 ();
 sg13g2_fill_8 FILLER_26_208 ();
 sg13g2_fill_8 FILLER_26_216 ();
 sg13g2_fill_8 FILLER_26_224 ();
 sg13g2_fill_8 FILLER_26_232 ();
 sg13g2_fill_8 FILLER_26_240 ();
 sg13g2_fill_8 FILLER_26_248 ();
 sg13g2_fill_8 FILLER_26_256 ();
 sg13g2_fill_8 FILLER_26_264 ();
 sg13g2_fill_8 FILLER_26_272 ();
 sg13g2_fill_8 FILLER_26_280 ();
 sg13g2_fill_8 FILLER_26_288 ();
 sg13g2_fill_8 FILLER_26_296 ();
 sg13g2_fill_8 FILLER_26_304 ();
 sg13g2_fill_8 FILLER_26_312 ();
 sg13g2_fill_8 FILLER_26_320 ();
 sg13g2_fill_8 FILLER_26_328 ();
 sg13g2_fill_8 FILLER_26_336 ();
 sg13g2_fill_8 FILLER_26_344 ();
 sg13g2_fill_8 FILLER_26_352 ();
 sg13g2_fill_4 FILLER_26_395 ();
 sg13g2_fill_1 FILLER_26_399 ();
 sg13g2_fill_8 FILLER_26_410 ();
 sg13g2_fill_2 FILLER_26_418 ();
 sg13g2_fill_1 FILLER_26_420 ();
 sg13g2_fill_8 FILLER_26_457 ();
 sg13g2_fill_4 FILLER_26_465 ();
 sg13g2_fill_2 FILLER_26_469 ();
 sg13g2_fill_4 FILLER_26_491 ();
 sg13g2_fill_1 FILLER_26_495 ();
 sg13g2_fill_8 FILLER_26_516 ();
 sg13g2_fill_1 FILLER_26_524 ();
 sg13g2_fill_1 FILLER_26_545 ();
 sg13g2_fill_8 FILLER_26_572 ();
 sg13g2_fill_8 FILLER_26_580 ();
 sg13g2_fill_8 FILLER_26_614 ();
 sg13g2_fill_8 FILLER_26_622 ();
 sg13g2_fill_4 FILLER_26_630 ();
 sg13g2_fill_1 FILLER_26_634 ();
 sg13g2_fill_8 FILLER_26_642 ();
 sg13g2_fill_1 FILLER_26_650 ();
 sg13g2_fill_2 FILLER_26_659 ();
 sg13g2_fill_1 FILLER_26_661 ();
 sg13g2_fill_8 FILLER_26_672 ();
 sg13g2_fill_8 FILLER_26_680 ();
 sg13g2_fill_8 FILLER_26_688 ();
 sg13g2_fill_4 FILLER_26_696 ();
 sg13g2_fill_2 FILLER_26_700 ();
 sg13g2_fill_1 FILLER_26_702 ();
 sg13g2_fill_2 FILLER_26_710 ();
 sg13g2_fill_1 FILLER_26_712 ();
 sg13g2_fill_4 FILLER_26_738 ();
 sg13g2_fill_2 FILLER_26_742 ();
 sg13g2_fill_8 FILLER_26_755 ();
 sg13g2_fill_4 FILLER_26_763 ();
 sg13g2_fill_1 FILLER_26_767 ();
 sg13g2_fill_4 FILLER_26_778 ();
 sg13g2_fill_2 FILLER_26_782 ();
 sg13g2_fill_1 FILLER_26_784 ();
 sg13g2_fill_4 FILLER_26_811 ();
 sg13g2_fill_8 FILLER_26_835 ();
 sg13g2_fill_1 FILLER_26_843 ();
 sg13g2_fill_8 FILLER_26_854 ();
 sg13g2_fill_8 FILLER_26_862 ();
 sg13g2_fill_8 FILLER_26_870 ();
 sg13g2_fill_2 FILLER_26_878 ();
 sg13g2_fill_1 FILLER_26_880 ();
 sg13g2_fill_8 FILLER_26_907 ();
 sg13g2_fill_2 FILLER_26_915 ();
 sg13g2_fill_4 FILLER_26_985 ();
 sg13g2_fill_4 FILLER_26_994 ();
 sg13g2_fill_1 FILLER_26_998 ();
 sg13g2_fill_8 FILLER_26_1009 ();
 sg13g2_fill_4 FILLER_26_1017 ();
 sg13g2_fill_2 FILLER_26_1021 ();
 sg13g2_fill_4 FILLER_26_1060 ();
 sg13g2_fill_1 FILLER_26_1064 ();
 sg13g2_fill_2 FILLER_26_1075 ();
 sg13g2_fill_8 FILLER_26_1162 ();
 sg13g2_fill_4 FILLER_26_1170 ();
 sg13g2_fill_8 FILLER_26_1184 ();
 sg13g2_fill_4 FILLER_26_1192 ();
 sg13g2_fill_2 FILLER_26_1196 ();
 sg13g2_fill_1 FILLER_26_1198 ();
 sg13g2_fill_4 FILLER_26_1243 ();
 sg13g2_fill_2 FILLER_26_1247 ();
 sg13g2_fill_1 FILLER_26_1249 ();
 sg13g2_fill_4 FILLER_26_1258 ();
 sg13g2_fill_8 FILLER_26_1270 ();
 sg13g2_fill_8 FILLER_26_1278 ();
 sg13g2_fill_8 FILLER_26_1286 ();
 sg13g2_fill_8 FILLER_26_1294 ();
 sg13g2_fill_8 FILLER_26_1302 ();
 sg13g2_fill_8 FILLER_26_1310 ();
 sg13g2_fill_8 FILLER_26_1318 ();
 sg13g2_fill_8 FILLER_26_1326 ();
 sg13g2_fill_8 FILLER_26_1334 ();
 sg13g2_fill_8 FILLER_26_1342 ();
 sg13g2_fill_8 FILLER_26_1350 ();
 sg13g2_fill_8 FILLER_26_1358 ();
 sg13g2_fill_8 FILLER_26_1366 ();
 sg13g2_fill_8 FILLER_26_1374 ();
 sg13g2_fill_8 FILLER_26_1382 ();
 sg13g2_fill_8 FILLER_26_1390 ();
 sg13g2_fill_8 FILLER_26_1398 ();
 sg13g2_fill_8 FILLER_26_1406 ();
 sg13g2_fill_8 FILLER_26_1414 ();
 sg13g2_fill_8 FILLER_26_1422 ();
 sg13g2_fill_8 FILLER_26_1430 ();
 sg13g2_fill_8 FILLER_26_1438 ();
 sg13g2_fill_8 FILLER_26_1446 ();
 sg13g2_fill_8 FILLER_26_1454 ();
 sg13g2_fill_8 FILLER_26_1462 ();
 sg13g2_fill_8 FILLER_26_1470 ();
 sg13g2_fill_8 FILLER_26_1478 ();
 sg13g2_fill_8 FILLER_26_1486 ();
 sg13g2_fill_8 FILLER_26_1494 ();
 sg13g2_fill_8 FILLER_26_1502 ();
 sg13g2_fill_8 FILLER_26_1510 ();
 sg13g2_fill_8 FILLER_26_1518 ();
 sg13g2_fill_8 FILLER_26_1526 ();
 sg13g2_fill_8 FILLER_26_1534 ();
 sg13g2_fill_8 FILLER_26_1542 ();
 sg13g2_fill_8 FILLER_26_1550 ();
 sg13g2_fill_8 FILLER_26_1558 ();
 sg13g2_fill_8 FILLER_26_1566 ();
 sg13g2_fill_8 FILLER_26_1574 ();
 sg13g2_fill_8 FILLER_26_1582 ();
 sg13g2_fill_2 FILLER_26_1590 ();
 sg13g2_fill_8 FILLER_27_0 ();
 sg13g2_fill_8 FILLER_27_8 ();
 sg13g2_fill_8 FILLER_27_16 ();
 sg13g2_fill_8 FILLER_27_24 ();
 sg13g2_fill_8 FILLER_27_32 ();
 sg13g2_fill_8 FILLER_27_40 ();
 sg13g2_fill_8 FILLER_27_48 ();
 sg13g2_fill_8 FILLER_27_56 ();
 sg13g2_fill_8 FILLER_27_64 ();
 sg13g2_fill_8 FILLER_27_72 ();
 sg13g2_fill_8 FILLER_27_80 ();
 sg13g2_fill_8 FILLER_27_88 ();
 sg13g2_fill_8 FILLER_27_96 ();
 sg13g2_fill_8 FILLER_27_104 ();
 sg13g2_fill_8 FILLER_27_112 ();
 sg13g2_fill_8 FILLER_27_120 ();
 sg13g2_fill_8 FILLER_27_128 ();
 sg13g2_fill_8 FILLER_27_136 ();
 sg13g2_fill_8 FILLER_27_144 ();
 sg13g2_fill_8 FILLER_27_152 ();
 sg13g2_fill_8 FILLER_27_160 ();
 sg13g2_fill_8 FILLER_27_168 ();
 sg13g2_fill_8 FILLER_27_176 ();
 sg13g2_fill_8 FILLER_27_184 ();
 sg13g2_fill_8 FILLER_27_192 ();
 sg13g2_fill_8 FILLER_27_200 ();
 sg13g2_fill_8 FILLER_27_208 ();
 sg13g2_fill_8 FILLER_27_216 ();
 sg13g2_fill_8 FILLER_27_224 ();
 sg13g2_fill_8 FILLER_27_232 ();
 sg13g2_fill_8 FILLER_27_240 ();
 sg13g2_fill_8 FILLER_27_248 ();
 sg13g2_fill_8 FILLER_27_256 ();
 sg13g2_fill_8 FILLER_27_264 ();
 sg13g2_fill_8 FILLER_27_272 ();
 sg13g2_fill_8 FILLER_27_280 ();
 sg13g2_fill_8 FILLER_27_288 ();
 sg13g2_fill_8 FILLER_27_296 ();
 sg13g2_fill_8 FILLER_27_304 ();
 sg13g2_fill_8 FILLER_27_312 ();
 sg13g2_fill_8 FILLER_27_320 ();
 sg13g2_fill_8 FILLER_27_328 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_8 FILLER_27_346 ();
 sg13g2_fill_8 FILLER_27_354 ();
 sg13g2_fill_8 FILLER_27_362 ();
 sg13g2_fill_4 FILLER_27_383 ();
 sg13g2_fill_8 FILLER_27_413 ();
 sg13g2_fill_4 FILLER_27_421 ();
 sg13g2_fill_1 FILLER_27_425 ();
 sg13g2_fill_1 FILLER_27_436 ();
 sg13g2_fill_8 FILLER_27_447 ();
 sg13g2_fill_4 FILLER_27_465 ();
 sg13g2_fill_2 FILLER_27_469 ();
 sg13g2_fill_1 FILLER_27_471 ();
 sg13g2_fill_4 FILLER_27_482 ();
 sg13g2_fill_4 FILLER_27_492 ();
 sg13g2_fill_1 FILLER_27_496 ();
 sg13g2_fill_4 FILLER_27_507 ();
 sg13g2_fill_8 FILLER_27_533 ();
 sg13g2_fill_8 FILLER_27_541 ();
 sg13g2_fill_8 FILLER_27_549 ();
 sg13g2_fill_8 FILLER_27_557 ();
 sg13g2_fill_4 FILLER_27_565 ();
 sg13g2_fill_2 FILLER_27_569 ();
 sg13g2_fill_8 FILLER_27_597 ();
 sg13g2_fill_2 FILLER_27_605 ();
 sg13g2_fill_1 FILLER_27_607 ();
 sg13g2_fill_1 FILLER_27_671 ();
 sg13g2_fill_2 FILLER_27_685 ();
 sg13g2_fill_1 FILLER_27_687 ();
 sg13g2_fill_2 FILLER_27_697 ();
 sg13g2_fill_4 FILLER_27_706 ();
 sg13g2_fill_1 FILLER_27_756 ();
 sg13g2_fill_1 FILLER_27_766 ();
 sg13g2_fill_8 FILLER_27_776 ();
 sg13g2_fill_8 FILLER_27_784 ();
 sg13g2_fill_8 FILLER_27_792 ();
 sg13g2_fill_4 FILLER_27_800 ();
 sg13g2_fill_8 FILLER_27_809 ();
 sg13g2_fill_8 FILLER_27_817 ();
 sg13g2_fill_4 FILLER_27_825 ();
 sg13g2_fill_2 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_831 ();
 sg13g2_fill_2 FILLER_27_838 ();
 sg13g2_fill_1 FILLER_27_840 ();
 sg13g2_fill_2 FILLER_27_898 ();
 sg13g2_fill_8 FILLER_27_931 ();
 sg13g2_fill_1 FILLER_27_939 ();
 sg13g2_fill_8 FILLER_27_945 ();
 sg13g2_fill_2 FILLER_27_953 ();
 sg13g2_fill_2 FILLER_27_1037 ();
 sg13g2_fill_8 FILLER_27_1095 ();
 sg13g2_fill_2 FILLER_27_1103 ();
 sg13g2_fill_1 FILLER_27_1130 ();
 sg13g2_fill_1 FILLER_27_1144 ();
 sg13g2_fill_8 FILLER_27_1166 ();
 sg13g2_fill_8 FILLER_27_1174 ();
 sg13g2_fill_8 FILLER_27_1182 ();
 sg13g2_fill_8 FILLER_27_1190 ();
 sg13g2_fill_2 FILLER_27_1198 ();
 sg13g2_fill_1 FILLER_27_1200 ();
 sg13g2_fill_2 FILLER_27_1210 ();
 sg13g2_fill_1 FILLER_27_1212 ();
 sg13g2_fill_4 FILLER_27_1227 ();
 sg13g2_fill_4 FILLER_27_1242 ();
 sg13g2_fill_1 FILLER_27_1246 ();
 sg13g2_fill_8 FILLER_27_1283 ();
 sg13g2_fill_8 FILLER_27_1291 ();
 sg13g2_fill_8 FILLER_27_1299 ();
 sg13g2_fill_8 FILLER_27_1307 ();
 sg13g2_fill_8 FILLER_27_1315 ();
 sg13g2_fill_8 FILLER_27_1323 ();
 sg13g2_fill_8 FILLER_27_1331 ();
 sg13g2_fill_8 FILLER_27_1339 ();
 sg13g2_fill_8 FILLER_27_1347 ();
 sg13g2_fill_8 FILLER_27_1355 ();
 sg13g2_fill_8 FILLER_27_1363 ();
 sg13g2_fill_8 FILLER_27_1371 ();
 sg13g2_fill_8 FILLER_27_1379 ();
 sg13g2_fill_8 FILLER_27_1387 ();
 sg13g2_fill_8 FILLER_27_1395 ();
 sg13g2_fill_8 FILLER_27_1403 ();
 sg13g2_fill_8 FILLER_27_1411 ();
 sg13g2_fill_8 FILLER_27_1419 ();
 sg13g2_fill_8 FILLER_27_1427 ();
 sg13g2_fill_8 FILLER_27_1435 ();
 sg13g2_fill_8 FILLER_27_1443 ();
 sg13g2_fill_8 FILLER_27_1451 ();
 sg13g2_fill_8 FILLER_27_1459 ();
 sg13g2_fill_8 FILLER_27_1467 ();
 sg13g2_fill_8 FILLER_27_1475 ();
 sg13g2_fill_8 FILLER_27_1483 ();
 sg13g2_fill_8 FILLER_27_1491 ();
 sg13g2_fill_8 FILLER_27_1499 ();
 sg13g2_fill_8 FILLER_27_1507 ();
 sg13g2_fill_8 FILLER_27_1515 ();
 sg13g2_fill_8 FILLER_27_1523 ();
 sg13g2_fill_8 FILLER_27_1531 ();
 sg13g2_fill_8 FILLER_27_1539 ();
 sg13g2_fill_8 FILLER_27_1547 ();
 sg13g2_fill_8 FILLER_27_1555 ();
 sg13g2_fill_8 FILLER_27_1563 ();
 sg13g2_fill_8 FILLER_27_1571 ();
 sg13g2_fill_8 FILLER_27_1579 ();
 sg13g2_fill_4 FILLER_27_1587 ();
 sg13g2_fill_1 FILLER_27_1591 ();
 sg13g2_fill_8 FILLER_28_0 ();
 sg13g2_fill_8 FILLER_28_8 ();
 sg13g2_fill_8 FILLER_28_16 ();
 sg13g2_fill_8 FILLER_28_24 ();
 sg13g2_fill_8 FILLER_28_32 ();
 sg13g2_fill_8 FILLER_28_40 ();
 sg13g2_fill_8 FILLER_28_48 ();
 sg13g2_fill_8 FILLER_28_56 ();
 sg13g2_fill_8 FILLER_28_64 ();
 sg13g2_fill_8 FILLER_28_72 ();
 sg13g2_fill_8 FILLER_28_80 ();
 sg13g2_fill_8 FILLER_28_88 ();
 sg13g2_fill_8 FILLER_28_96 ();
 sg13g2_fill_8 FILLER_28_104 ();
 sg13g2_fill_8 FILLER_28_112 ();
 sg13g2_fill_8 FILLER_28_120 ();
 sg13g2_fill_8 FILLER_28_128 ();
 sg13g2_fill_8 FILLER_28_136 ();
 sg13g2_fill_8 FILLER_28_144 ();
 sg13g2_fill_8 FILLER_28_152 ();
 sg13g2_fill_8 FILLER_28_160 ();
 sg13g2_fill_8 FILLER_28_168 ();
 sg13g2_fill_8 FILLER_28_176 ();
 sg13g2_fill_8 FILLER_28_184 ();
 sg13g2_fill_8 FILLER_28_192 ();
 sg13g2_fill_8 FILLER_28_200 ();
 sg13g2_fill_8 FILLER_28_208 ();
 sg13g2_fill_8 FILLER_28_216 ();
 sg13g2_fill_8 FILLER_28_224 ();
 sg13g2_fill_8 FILLER_28_232 ();
 sg13g2_fill_8 FILLER_28_240 ();
 sg13g2_fill_8 FILLER_28_248 ();
 sg13g2_fill_8 FILLER_28_256 ();
 sg13g2_fill_8 FILLER_28_264 ();
 sg13g2_fill_8 FILLER_28_272 ();
 sg13g2_fill_8 FILLER_28_280 ();
 sg13g2_fill_8 FILLER_28_288 ();
 sg13g2_fill_8 FILLER_28_296 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_8 FILLER_28_393 ();
 sg13g2_fill_4 FILLER_28_401 ();
 sg13g2_fill_2 FILLER_28_425 ();
 sg13g2_fill_1 FILLER_28_447 ();
 sg13g2_fill_4 FILLER_28_458 ();
 sg13g2_fill_1 FILLER_28_462 ();
 sg13g2_fill_8 FILLER_28_473 ();
 sg13g2_fill_2 FILLER_28_481 ();
 sg13g2_fill_1 FILLER_28_483 ();
 sg13g2_fill_8 FILLER_28_490 ();
 sg13g2_fill_4 FILLER_28_498 ();
 sg13g2_fill_8 FILLER_28_512 ();
 sg13g2_fill_1 FILLER_28_520 ();
 sg13g2_fill_2 FILLER_28_541 ();
 sg13g2_fill_1 FILLER_28_543 ();
 sg13g2_fill_8 FILLER_28_564 ();
 sg13g2_fill_2 FILLER_28_572 ();
 sg13g2_fill_1 FILLER_28_574 ();
 sg13g2_fill_1 FILLER_28_578 ();
 sg13g2_fill_8 FILLER_28_626 ();
 sg13g2_fill_8 FILLER_28_634 ();
 sg13g2_fill_4 FILLER_28_642 ();
 sg13g2_fill_2 FILLER_28_646 ();
 sg13g2_fill_1 FILLER_28_648 ();
 sg13g2_fill_2 FILLER_28_663 ();
 sg13g2_fill_1 FILLER_28_726 ();
 sg13g2_fill_4 FILLER_28_737 ();
 sg13g2_fill_2 FILLER_28_741 ();
 sg13g2_fill_1 FILLER_28_743 ();
 sg13g2_fill_2 FILLER_28_751 ();
 sg13g2_fill_1 FILLER_28_753 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_fill_8 FILLER_28_796 ();
 sg13g2_fill_4 FILLER_28_804 ();
 sg13g2_fill_4 FILLER_28_820 ();
 sg13g2_fill_2 FILLER_28_824 ();
 sg13g2_fill_2 FILLER_28_845 ();
 sg13g2_fill_4 FILLER_28_887 ();
 sg13g2_fill_2 FILLER_28_927 ();
 sg13g2_fill_1 FILLER_28_929 ();
 sg13g2_fill_1 FILLER_28_981 ();
 sg13g2_fill_8 FILLER_28_995 ();
 sg13g2_fill_8 FILLER_28_1003 ();
 sg13g2_fill_4 FILLER_28_1011 ();
 sg13g2_fill_8 FILLER_28_1019 ();
 sg13g2_fill_8 FILLER_28_1027 ();
 sg13g2_fill_2 FILLER_28_1035 ();
 sg13g2_fill_1 FILLER_28_1042 ();
 sg13g2_fill_8 FILLER_28_1058 ();
 sg13g2_fill_4 FILLER_28_1066 ();
 sg13g2_fill_2 FILLER_28_1074 ();
 sg13g2_fill_2 FILLER_28_1080 ();
 sg13g2_fill_2 FILLER_28_1107 ();
 sg13g2_fill_1 FILLER_28_1109 ();
 sg13g2_fill_2 FILLER_28_1146 ();
 sg13g2_fill_1 FILLER_28_1148 ();
 sg13g2_fill_8 FILLER_28_1155 ();
 sg13g2_fill_8 FILLER_28_1163 ();
 sg13g2_fill_4 FILLER_28_1171 ();
 sg13g2_fill_2 FILLER_28_1201 ();
 sg13g2_fill_1 FILLER_28_1203 ();
 sg13g2_fill_4 FILLER_28_1209 ();
 sg13g2_fill_8 FILLER_28_1248 ();
 sg13g2_fill_8 FILLER_28_1256 ();
 sg13g2_fill_4 FILLER_28_1264 ();
 sg13g2_fill_2 FILLER_28_1268 ();
 sg13g2_fill_8 FILLER_28_1295 ();
 sg13g2_fill_8 FILLER_28_1303 ();
 sg13g2_fill_8 FILLER_28_1311 ();
 sg13g2_fill_8 FILLER_28_1319 ();
 sg13g2_fill_8 FILLER_28_1327 ();
 sg13g2_fill_8 FILLER_28_1335 ();
 sg13g2_fill_8 FILLER_28_1343 ();
 sg13g2_fill_8 FILLER_28_1351 ();
 sg13g2_fill_8 FILLER_28_1359 ();
 sg13g2_fill_8 FILLER_28_1367 ();
 sg13g2_fill_8 FILLER_28_1375 ();
 sg13g2_fill_8 FILLER_28_1383 ();
 sg13g2_fill_8 FILLER_28_1391 ();
 sg13g2_fill_8 FILLER_28_1399 ();
 sg13g2_fill_8 FILLER_28_1407 ();
 sg13g2_fill_8 FILLER_28_1415 ();
 sg13g2_fill_8 FILLER_28_1423 ();
 sg13g2_fill_8 FILLER_28_1431 ();
 sg13g2_fill_8 FILLER_28_1439 ();
 sg13g2_fill_8 FILLER_28_1447 ();
 sg13g2_fill_8 FILLER_28_1455 ();
 sg13g2_fill_8 FILLER_28_1463 ();
 sg13g2_fill_8 FILLER_28_1471 ();
 sg13g2_fill_8 FILLER_28_1479 ();
 sg13g2_fill_8 FILLER_28_1487 ();
 sg13g2_fill_8 FILLER_28_1495 ();
 sg13g2_fill_8 FILLER_28_1503 ();
 sg13g2_fill_8 FILLER_28_1511 ();
 sg13g2_fill_8 FILLER_28_1519 ();
 sg13g2_fill_8 FILLER_28_1527 ();
 sg13g2_fill_8 FILLER_28_1535 ();
 sg13g2_fill_8 FILLER_28_1543 ();
 sg13g2_fill_8 FILLER_28_1551 ();
 sg13g2_fill_8 FILLER_28_1559 ();
 sg13g2_fill_8 FILLER_28_1567 ();
 sg13g2_fill_8 FILLER_28_1575 ();
 sg13g2_fill_8 FILLER_28_1583 ();
 sg13g2_fill_1 FILLER_28_1591 ();
 sg13g2_fill_8 FILLER_29_0 ();
 sg13g2_fill_8 FILLER_29_8 ();
 sg13g2_fill_8 FILLER_29_16 ();
 sg13g2_fill_8 FILLER_29_24 ();
 sg13g2_fill_8 FILLER_29_32 ();
 sg13g2_fill_8 FILLER_29_40 ();
 sg13g2_fill_8 FILLER_29_48 ();
 sg13g2_fill_8 FILLER_29_56 ();
 sg13g2_fill_8 FILLER_29_64 ();
 sg13g2_fill_8 FILLER_29_72 ();
 sg13g2_fill_8 FILLER_29_80 ();
 sg13g2_fill_8 FILLER_29_88 ();
 sg13g2_fill_8 FILLER_29_96 ();
 sg13g2_fill_8 FILLER_29_104 ();
 sg13g2_fill_8 FILLER_29_112 ();
 sg13g2_fill_8 FILLER_29_120 ();
 sg13g2_fill_8 FILLER_29_128 ();
 sg13g2_fill_8 FILLER_29_136 ();
 sg13g2_fill_8 FILLER_29_144 ();
 sg13g2_fill_8 FILLER_29_152 ();
 sg13g2_fill_8 FILLER_29_160 ();
 sg13g2_fill_8 FILLER_29_168 ();
 sg13g2_fill_8 FILLER_29_176 ();
 sg13g2_fill_8 FILLER_29_184 ();
 sg13g2_fill_8 FILLER_29_192 ();
 sg13g2_fill_8 FILLER_29_200 ();
 sg13g2_fill_8 FILLER_29_208 ();
 sg13g2_fill_8 FILLER_29_216 ();
 sg13g2_fill_8 FILLER_29_224 ();
 sg13g2_fill_8 FILLER_29_232 ();
 sg13g2_fill_8 FILLER_29_240 ();
 sg13g2_fill_8 FILLER_29_248 ();
 sg13g2_fill_4 FILLER_29_256 ();
 sg13g2_fill_8 FILLER_29_286 ();
 sg13g2_fill_4 FILLER_29_294 ();
 sg13g2_fill_4 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_338 ();
 sg13g2_fill_8 FILLER_29_376 ();
 sg13g2_fill_4 FILLER_29_384 ();
 sg13g2_fill_1 FILLER_29_388 ();
 sg13g2_fill_8 FILLER_29_415 ();
 sg13g2_fill_8 FILLER_29_423 ();
 sg13g2_fill_8 FILLER_29_431 ();
 sg13g2_fill_8 FILLER_29_439 ();
 sg13g2_fill_8 FILLER_29_447 ();
 sg13g2_fill_8 FILLER_29_473 ();
 sg13g2_fill_8 FILLER_29_481 ();
 sg13g2_fill_8 FILLER_29_489 ();
 sg13g2_fill_4 FILLER_29_497 ();
 sg13g2_fill_1 FILLER_29_501 ();
 sg13g2_fill_8 FILLER_29_512 ();
 sg13g2_fill_8 FILLER_29_520 ();
 sg13g2_fill_2 FILLER_29_528 ();
 sg13g2_fill_1 FILLER_29_530 ();
 sg13g2_fill_8 FILLER_29_577 ();
 sg13g2_fill_8 FILLER_29_585 ();
 sg13g2_fill_8 FILLER_29_593 ();
 sg13g2_fill_8 FILLER_29_601 ();
 sg13g2_fill_8 FILLER_29_609 ();
 sg13g2_fill_1 FILLER_29_628 ();
 sg13g2_fill_8 FILLER_29_637 ();
 sg13g2_fill_8 FILLER_29_645 ();
 sg13g2_fill_8 FILLER_29_664 ();
 sg13g2_fill_2 FILLER_29_672 ();
 sg13g2_fill_1 FILLER_29_674 ();
 sg13g2_fill_1 FILLER_29_680 ();
 sg13g2_fill_4 FILLER_29_685 ();
 sg13g2_fill_4 FILLER_29_694 ();
 sg13g2_fill_8 FILLER_29_708 ();
 sg13g2_fill_8 FILLER_29_716 ();
 sg13g2_fill_1 FILLER_29_724 ();
 sg13g2_fill_4 FILLER_29_752 ();
 sg13g2_fill_8 FILLER_29_792 ();
 sg13g2_fill_4 FILLER_29_800 ();
 sg13g2_fill_1 FILLER_29_804 ();
 sg13g2_fill_8 FILLER_29_829 ();
 sg13g2_fill_2 FILLER_29_837 ();
 sg13g2_fill_1 FILLER_29_839 ();
 sg13g2_fill_8 FILLER_29_848 ();
 sg13g2_fill_4 FILLER_29_856 ();
 sg13g2_fill_8 FILLER_29_864 ();
 sg13g2_fill_8 FILLER_29_872 ();
 sg13g2_fill_2 FILLER_29_880 ();
 sg13g2_fill_1 FILLER_29_882 ();
 sg13g2_fill_2 FILLER_29_898 ();
 sg13g2_fill_8 FILLER_29_928 ();
 sg13g2_fill_8 FILLER_29_936 ();
 sg13g2_fill_8 FILLER_29_944 ();
 sg13g2_fill_8 FILLER_29_952 ();
 sg13g2_fill_1 FILLER_29_970 ();
 sg13g2_fill_2 FILLER_29_985 ();
 sg13g2_fill_1 FILLER_29_987 ();
 sg13g2_fill_8 FILLER_29_993 ();
 sg13g2_fill_4 FILLER_29_1001 ();
 sg13g2_fill_8 FILLER_29_1021 ();
 sg13g2_fill_2 FILLER_29_1029 ();
 sg13g2_fill_1 FILLER_29_1031 ();
 sg13g2_fill_2 FILLER_29_1052 ();
 sg13g2_fill_1 FILLER_29_1054 ();
 sg13g2_fill_8 FILLER_29_1059 ();
 sg13g2_fill_8 FILLER_29_1067 ();
 sg13g2_fill_2 FILLER_29_1075 ();
 sg13g2_fill_2 FILLER_29_1107 ();
 sg13g2_fill_1 FILLER_29_1109 ();
 sg13g2_fill_4 FILLER_29_1167 ();
 sg13g2_fill_2 FILLER_29_1171 ();
 sg13g2_fill_1 FILLER_29_1199 ();
 sg13g2_fill_2 FILLER_29_1236 ();
 sg13g2_fill_1 FILLER_29_1238 ();
 sg13g2_fill_4 FILLER_29_1264 ();
 sg13g2_fill_2 FILLER_29_1268 ();
 sg13g2_fill_1 FILLER_29_1270 ();
 sg13g2_fill_8 FILLER_29_1315 ();
 sg13g2_fill_8 FILLER_29_1323 ();
 sg13g2_fill_8 FILLER_29_1331 ();
 sg13g2_fill_8 FILLER_29_1339 ();
 sg13g2_fill_8 FILLER_29_1347 ();
 sg13g2_fill_8 FILLER_29_1355 ();
 sg13g2_fill_8 FILLER_29_1363 ();
 sg13g2_fill_8 FILLER_29_1371 ();
 sg13g2_fill_8 FILLER_29_1379 ();
 sg13g2_fill_8 FILLER_29_1387 ();
 sg13g2_fill_8 FILLER_29_1395 ();
 sg13g2_fill_8 FILLER_29_1403 ();
 sg13g2_fill_8 FILLER_29_1411 ();
 sg13g2_fill_8 FILLER_29_1419 ();
 sg13g2_fill_8 FILLER_29_1427 ();
 sg13g2_fill_8 FILLER_29_1435 ();
 sg13g2_fill_8 FILLER_29_1443 ();
 sg13g2_fill_8 FILLER_29_1451 ();
 sg13g2_fill_8 FILLER_29_1459 ();
 sg13g2_fill_8 FILLER_29_1467 ();
 sg13g2_fill_8 FILLER_29_1475 ();
 sg13g2_fill_8 FILLER_29_1483 ();
 sg13g2_fill_8 FILLER_29_1491 ();
 sg13g2_fill_8 FILLER_29_1499 ();
 sg13g2_fill_8 FILLER_29_1507 ();
 sg13g2_fill_8 FILLER_29_1515 ();
 sg13g2_fill_8 FILLER_29_1523 ();
 sg13g2_fill_8 FILLER_29_1531 ();
 sg13g2_fill_8 FILLER_29_1539 ();
 sg13g2_fill_8 FILLER_29_1547 ();
 sg13g2_fill_8 FILLER_29_1555 ();
 sg13g2_fill_8 FILLER_29_1563 ();
 sg13g2_fill_8 FILLER_29_1571 ();
 sg13g2_fill_8 FILLER_29_1579 ();
 sg13g2_fill_4 FILLER_29_1587 ();
 sg13g2_fill_1 FILLER_29_1591 ();
 sg13g2_fill_8 FILLER_30_0 ();
 sg13g2_fill_8 FILLER_30_8 ();
 sg13g2_fill_8 FILLER_30_16 ();
 sg13g2_fill_8 FILLER_30_24 ();
 sg13g2_fill_8 FILLER_30_32 ();
 sg13g2_fill_8 FILLER_30_40 ();
 sg13g2_fill_8 FILLER_30_48 ();
 sg13g2_fill_8 FILLER_30_56 ();
 sg13g2_fill_8 FILLER_30_64 ();
 sg13g2_fill_8 FILLER_30_72 ();
 sg13g2_fill_8 FILLER_30_80 ();
 sg13g2_fill_8 FILLER_30_88 ();
 sg13g2_fill_8 FILLER_30_96 ();
 sg13g2_fill_8 FILLER_30_104 ();
 sg13g2_fill_8 FILLER_30_112 ();
 sg13g2_fill_8 FILLER_30_120 ();
 sg13g2_fill_8 FILLER_30_128 ();
 sg13g2_fill_8 FILLER_30_136 ();
 sg13g2_fill_8 FILLER_30_144 ();
 sg13g2_fill_8 FILLER_30_152 ();
 sg13g2_fill_8 FILLER_30_160 ();
 sg13g2_fill_8 FILLER_30_168 ();
 sg13g2_fill_8 FILLER_30_176 ();
 sg13g2_fill_8 FILLER_30_184 ();
 sg13g2_fill_8 FILLER_30_192 ();
 sg13g2_fill_8 FILLER_30_200 ();
 sg13g2_fill_8 FILLER_30_208 ();
 sg13g2_fill_8 FILLER_30_216 ();
 sg13g2_fill_8 FILLER_30_224 ();
 sg13g2_fill_4 FILLER_30_232 ();
 sg13g2_fill_8 FILLER_30_246 ();
 sg13g2_fill_8 FILLER_30_254 ();
 sg13g2_fill_4 FILLER_30_262 ();
 sg13g2_fill_8 FILLER_30_292 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_8 FILLER_30_322 ();
 sg13g2_fill_8 FILLER_30_330 ();
 sg13g2_fill_8 FILLER_30_338 ();
 sg13g2_fill_4 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_350 ();
 sg13g2_fill_4 FILLER_30_377 ();
 sg13g2_fill_8 FILLER_30_391 ();
 sg13g2_fill_4 FILLER_30_399 ();
 sg13g2_fill_8 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_421 ();
 sg13g2_fill_4 FILLER_30_441 ();
 sg13g2_fill_2 FILLER_30_445 ();
 sg13g2_fill_1 FILLER_30_447 ();
 sg13g2_fill_8 FILLER_30_458 ();
 sg13g2_fill_4 FILLER_30_466 ();
 sg13g2_fill_2 FILLER_30_470 ();
 sg13g2_fill_8 FILLER_30_498 ();
 sg13g2_fill_8 FILLER_30_506 ();
 sg13g2_fill_4 FILLER_30_514 ();
 sg13g2_fill_2 FILLER_30_518 ();
 sg13g2_fill_8 FILLER_30_540 ();
 sg13g2_fill_4 FILLER_30_548 ();
 sg13g2_fill_8 FILLER_30_562 ();
 sg13g2_fill_4 FILLER_30_570 ();
 sg13g2_fill_1 FILLER_30_574 ();
 sg13g2_fill_8 FILLER_30_586 ();
 sg13g2_fill_8 FILLER_30_594 ();
 sg13g2_fill_1 FILLER_30_609 ();
 sg13g2_fill_4 FILLER_30_621 ();
 sg13g2_fill_1 FILLER_30_625 ();
 sg13g2_fill_2 FILLER_30_639 ();
 sg13g2_fill_2 FILLER_30_651 ();
 sg13g2_fill_1 FILLER_30_653 ();
 sg13g2_fill_2 FILLER_30_662 ();
 sg13g2_fill_1 FILLER_30_668 ();
 sg13g2_fill_2 FILLER_30_682 ();
 sg13g2_fill_1 FILLER_30_684 ();
 sg13g2_fill_2 FILLER_30_692 ();
 sg13g2_fill_1 FILLER_30_694 ();
 sg13g2_fill_4 FILLER_30_711 ();
 sg13g2_fill_1 FILLER_30_740 ();
 sg13g2_fill_2 FILLER_30_746 ();
 sg13g2_fill_4 FILLER_30_778 ();
 sg13g2_fill_2 FILLER_30_782 ();
 sg13g2_fill_8 FILLER_30_792 ();
 sg13g2_fill_8 FILLER_30_800 ();
 sg13g2_fill_4 FILLER_30_808 ();
 sg13g2_fill_2 FILLER_30_848 ();
 sg13g2_fill_4 FILLER_30_868 ();
 sg13g2_fill_8 FILLER_30_895 ();
 sg13g2_fill_2 FILLER_30_933 ();
 sg13g2_fill_1 FILLER_30_935 ();
 sg13g2_fill_8 FILLER_30_942 ();
 sg13g2_fill_4 FILLER_30_950 ();
 sg13g2_fill_2 FILLER_30_954 ();
 sg13g2_fill_1 FILLER_30_956 ();
 sg13g2_fill_4 FILLER_30_962 ();
 sg13g2_fill_2 FILLER_30_966 ();
 sg13g2_fill_1 FILLER_30_968 ();
 sg13g2_fill_1 FILLER_30_974 ();
 sg13g2_fill_1 FILLER_30_988 ();
 sg13g2_fill_2 FILLER_30_1008 ();
 sg13g2_fill_2 FILLER_30_1046 ();
 sg13g2_fill_4 FILLER_30_1074 ();
 sg13g2_fill_2 FILLER_30_1078 ();
 sg13g2_fill_8 FILLER_30_1114 ();
 sg13g2_fill_8 FILLER_30_1122 ();
 sg13g2_fill_8 FILLER_30_1130 ();
 sg13g2_fill_4 FILLER_30_1138 ();
 sg13g2_fill_2 FILLER_30_1142 ();
 sg13g2_fill_1 FILLER_30_1144 ();
 sg13g2_fill_2 FILLER_30_1166 ();
 sg13g2_fill_1 FILLER_30_1168 ();
 sg13g2_fill_8 FILLER_30_1189 ();
 sg13g2_fill_1 FILLER_30_1197 ();
 sg13g2_fill_2 FILLER_30_1207 ();
 sg13g2_fill_8 FILLER_30_1235 ();
 sg13g2_fill_8 FILLER_30_1243 ();
 sg13g2_fill_8 FILLER_30_1251 ();
 sg13g2_fill_8 FILLER_30_1259 ();
 sg13g2_fill_8 FILLER_30_1267 ();
 sg13g2_fill_4 FILLER_30_1275 ();
 sg13g2_fill_2 FILLER_30_1279 ();
 sg13g2_fill_1 FILLER_30_1281 ();
 sg13g2_fill_8 FILLER_30_1307 ();
 sg13g2_fill_8 FILLER_30_1315 ();
 sg13g2_fill_8 FILLER_30_1323 ();
 sg13g2_fill_8 FILLER_30_1331 ();
 sg13g2_fill_8 FILLER_30_1339 ();
 sg13g2_fill_8 FILLER_30_1347 ();
 sg13g2_fill_8 FILLER_30_1355 ();
 sg13g2_fill_8 FILLER_30_1363 ();
 sg13g2_fill_8 FILLER_30_1371 ();
 sg13g2_fill_8 FILLER_30_1379 ();
 sg13g2_fill_8 FILLER_30_1387 ();
 sg13g2_fill_8 FILLER_30_1395 ();
 sg13g2_fill_8 FILLER_30_1403 ();
 sg13g2_fill_8 FILLER_30_1411 ();
 sg13g2_fill_8 FILLER_30_1419 ();
 sg13g2_fill_8 FILLER_30_1427 ();
 sg13g2_fill_8 FILLER_30_1435 ();
 sg13g2_fill_8 FILLER_30_1443 ();
 sg13g2_fill_8 FILLER_30_1451 ();
 sg13g2_fill_8 FILLER_30_1459 ();
 sg13g2_fill_8 FILLER_30_1467 ();
 sg13g2_fill_8 FILLER_30_1475 ();
 sg13g2_fill_8 FILLER_30_1483 ();
 sg13g2_fill_8 FILLER_30_1491 ();
 sg13g2_fill_8 FILLER_30_1499 ();
 sg13g2_fill_8 FILLER_30_1507 ();
 sg13g2_fill_8 FILLER_30_1515 ();
 sg13g2_fill_8 FILLER_30_1523 ();
 sg13g2_fill_8 FILLER_30_1531 ();
 sg13g2_fill_8 FILLER_30_1539 ();
 sg13g2_fill_8 FILLER_30_1547 ();
 sg13g2_fill_8 FILLER_30_1555 ();
 sg13g2_fill_8 FILLER_30_1563 ();
 sg13g2_fill_8 FILLER_30_1571 ();
 sg13g2_fill_8 FILLER_30_1579 ();
 sg13g2_fill_4 FILLER_30_1587 ();
 sg13g2_fill_1 FILLER_30_1591 ();
 sg13g2_fill_8 FILLER_31_0 ();
 sg13g2_fill_8 FILLER_31_8 ();
 sg13g2_fill_8 FILLER_31_16 ();
 sg13g2_fill_8 FILLER_31_24 ();
 sg13g2_fill_8 FILLER_31_32 ();
 sg13g2_fill_8 FILLER_31_40 ();
 sg13g2_fill_8 FILLER_31_48 ();
 sg13g2_fill_8 FILLER_31_56 ();
 sg13g2_fill_8 FILLER_31_64 ();
 sg13g2_fill_8 FILLER_31_72 ();
 sg13g2_fill_8 FILLER_31_80 ();
 sg13g2_fill_8 FILLER_31_88 ();
 sg13g2_fill_8 FILLER_31_96 ();
 sg13g2_fill_8 FILLER_31_104 ();
 sg13g2_fill_8 FILLER_31_112 ();
 sg13g2_fill_8 FILLER_31_120 ();
 sg13g2_fill_8 FILLER_31_128 ();
 sg13g2_fill_8 FILLER_31_136 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_fill_8 FILLER_31_183 ();
 sg13g2_fill_8 FILLER_31_191 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_4 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_fill_2 FILLER_31_242 ();
 sg13g2_fill_8 FILLER_31_254 ();
 sg13g2_fill_8 FILLER_31_262 ();
 sg13g2_fill_4 FILLER_31_270 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_8 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_303 ();
 sg13g2_fill_8 FILLER_31_329 ();
 sg13g2_fill_8 FILLER_31_337 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_8 FILLER_31_356 ();
 sg13g2_fill_8 FILLER_31_364 ();
 sg13g2_fill_4 FILLER_31_372 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_8 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_407 ();
 sg13g2_fill_4 FILLER_31_418 ();
 sg13g2_fill_2 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_424 ();
 sg13g2_fill_2 FILLER_31_454 ();
 sg13g2_fill_1 FILLER_31_462 ();
 sg13g2_fill_8 FILLER_31_539 ();
 sg13g2_fill_4 FILLER_31_547 ();
 sg13g2_fill_1 FILLER_31_551 ();
 sg13g2_fill_4 FILLER_31_568 ();
 sg13g2_fill_2 FILLER_31_572 ();
 sg13g2_fill_2 FILLER_31_604 ();
 sg13g2_fill_1 FILLER_31_606 ();
 sg13g2_fill_4 FILLER_31_724 ();
 sg13g2_fill_2 FILLER_31_728 ();
 sg13g2_fill_1 FILLER_31_730 ();
 sg13g2_fill_2 FILLER_31_781 ();
 sg13g2_fill_4 FILLER_31_809 ();
 sg13g2_fill_2 FILLER_31_813 ();
 sg13g2_fill_1 FILLER_31_815 ();
 sg13g2_fill_4 FILLER_31_860 ();
 sg13g2_fill_2 FILLER_31_864 ();
 sg13g2_fill_1 FILLER_31_866 ();
 sg13g2_fill_8 FILLER_31_893 ();
 sg13g2_fill_2 FILLER_31_905 ();
 sg13g2_fill_1 FILLER_31_913 ();
 sg13g2_fill_2 FILLER_31_932 ();
 sg13g2_fill_8 FILLER_31_940 ();
 sg13g2_fill_4 FILLER_31_948 ();
 sg13g2_fill_2 FILLER_31_952 ();
 sg13g2_fill_1 FILLER_31_954 ();
 sg13g2_fill_4 FILLER_31_980 ();
 sg13g2_fill_2 FILLER_31_984 ();
 sg13g2_fill_1 FILLER_31_986 ();
 sg13g2_fill_1 FILLER_31_1003 ();
 sg13g2_fill_8 FILLER_31_1020 ();
 sg13g2_fill_4 FILLER_31_1028 ();
 sg13g2_fill_2 FILLER_31_1032 ();
 sg13g2_fill_1 FILLER_31_1034 ();
 sg13g2_fill_8 FILLER_31_1040 ();
 sg13g2_fill_8 FILLER_31_1053 ();
 sg13g2_fill_8 FILLER_31_1061 ();
 sg13g2_fill_8 FILLER_31_1069 ();
 sg13g2_fill_4 FILLER_31_1077 ();
 sg13g2_fill_2 FILLER_31_1119 ();
 sg13g2_fill_8 FILLER_31_1126 ();
 sg13g2_fill_2 FILLER_31_1134 ();
 sg13g2_fill_8 FILLER_31_1146 ();
 sg13g2_fill_4 FILLER_31_1154 ();
 sg13g2_fill_1 FILLER_31_1158 ();
 sg13g2_fill_2 FILLER_31_1172 ();
 sg13g2_fill_2 FILLER_31_1200 ();
 sg13g2_fill_1 FILLER_31_1202 ();
 sg13g2_fill_8 FILLER_31_1213 ();
 sg13g2_fill_4 FILLER_31_1221 ();
 sg13g2_fill_2 FILLER_31_1225 ();
 sg13g2_fill_1 FILLER_31_1227 ();
 sg13g2_fill_8 FILLER_31_1319 ();
 sg13g2_fill_8 FILLER_31_1327 ();
 sg13g2_fill_8 FILLER_31_1335 ();
 sg13g2_fill_8 FILLER_31_1343 ();
 sg13g2_fill_8 FILLER_31_1351 ();
 sg13g2_fill_8 FILLER_31_1359 ();
 sg13g2_fill_8 FILLER_31_1367 ();
 sg13g2_fill_8 FILLER_31_1375 ();
 sg13g2_fill_8 FILLER_31_1383 ();
 sg13g2_fill_8 FILLER_31_1391 ();
 sg13g2_fill_8 FILLER_31_1399 ();
 sg13g2_fill_8 FILLER_31_1407 ();
 sg13g2_fill_8 FILLER_31_1415 ();
 sg13g2_fill_8 FILLER_31_1423 ();
 sg13g2_fill_8 FILLER_31_1431 ();
 sg13g2_fill_8 FILLER_31_1439 ();
 sg13g2_fill_8 FILLER_31_1447 ();
 sg13g2_fill_8 FILLER_31_1455 ();
 sg13g2_fill_8 FILLER_31_1463 ();
 sg13g2_fill_8 FILLER_31_1471 ();
 sg13g2_fill_8 FILLER_31_1479 ();
 sg13g2_fill_8 FILLER_31_1487 ();
 sg13g2_fill_8 FILLER_31_1495 ();
 sg13g2_fill_8 FILLER_31_1503 ();
 sg13g2_fill_8 FILLER_31_1511 ();
 sg13g2_fill_8 FILLER_31_1519 ();
 sg13g2_fill_8 FILLER_31_1527 ();
 sg13g2_fill_8 FILLER_31_1535 ();
 sg13g2_fill_8 FILLER_31_1543 ();
 sg13g2_fill_8 FILLER_31_1551 ();
 sg13g2_fill_8 FILLER_31_1559 ();
 sg13g2_fill_8 FILLER_31_1567 ();
 sg13g2_fill_8 FILLER_31_1575 ();
 sg13g2_fill_8 FILLER_31_1583 ();
 sg13g2_fill_1 FILLER_31_1591 ();
 sg13g2_fill_8 FILLER_32_0 ();
 sg13g2_fill_8 FILLER_32_8 ();
 sg13g2_fill_8 FILLER_32_16 ();
 sg13g2_fill_8 FILLER_32_24 ();
 sg13g2_fill_8 FILLER_32_32 ();
 sg13g2_fill_8 FILLER_32_40 ();
 sg13g2_fill_8 FILLER_32_48 ();
 sg13g2_fill_8 FILLER_32_56 ();
 sg13g2_fill_8 FILLER_32_64 ();
 sg13g2_fill_8 FILLER_32_72 ();
 sg13g2_fill_8 FILLER_32_80 ();
 sg13g2_fill_8 FILLER_32_88 ();
 sg13g2_fill_8 FILLER_32_96 ();
 sg13g2_fill_8 FILLER_32_104 ();
 sg13g2_fill_8 FILLER_32_112 ();
 sg13g2_fill_8 FILLER_32_120 ();
 sg13g2_fill_8 FILLER_32_128 ();
 sg13g2_fill_8 FILLER_32_136 ();
 sg13g2_fill_2 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_146 ();
 sg13g2_fill_8 FILLER_32_173 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_209 ();
 sg13g2_fill_8 FILLER_32_262 ();
 sg13g2_fill_8 FILLER_32_270 ();
 sg13g2_fill_8 FILLER_32_278 ();
 sg13g2_fill_8 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_294 ();
 sg13g2_fill_4 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_325 ();
 sg13g2_fill_1 FILLER_32_327 ();
 sg13g2_fill_8 FILLER_32_364 ();
 sg13g2_fill_4 FILLER_32_372 ();
 sg13g2_fill_1 FILLER_32_376 ();
 sg13g2_fill_8 FILLER_32_387 ();
 sg13g2_fill_4 FILLER_32_395 ();
 sg13g2_fill_2 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_419 ();
 sg13g2_fill_2 FILLER_32_452 ();
 sg13g2_fill_8 FILLER_32_483 ();
 sg13g2_fill_4 FILLER_32_491 ();
 sg13g2_fill_2 FILLER_32_495 ();
 sg13g2_fill_2 FILLER_32_514 ();
 sg13g2_fill_1 FILLER_32_523 ();
 sg13g2_fill_8 FILLER_32_531 ();
 sg13g2_fill_8 FILLER_32_539 ();
 sg13g2_fill_8 FILLER_32_554 ();
 sg13g2_fill_4 FILLER_32_562 ();
 sg13g2_fill_1 FILLER_32_566 ();
 sg13g2_fill_2 FILLER_32_572 ();
 sg13g2_fill_1 FILLER_32_574 ();
 sg13g2_fill_4 FILLER_32_605 ();
 sg13g2_fill_1 FILLER_32_609 ();
 sg13g2_fill_8 FILLER_32_666 ();
 sg13g2_fill_2 FILLER_32_674 ();
 sg13g2_fill_1 FILLER_32_690 ();
 sg13g2_fill_4 FILLER_32_717 ();
 sg13g2_fill_2 FILLER_32_721 ();
 sg13g2_fill_4 FILLER_32_730 ();
 sg13g2_fill_2 FILLER_32_734 ();
 sg13g2_fill_1 FILLER_32_736 ();
 sg13g2_fill_2 FILLER_32_747 ();
 sg13g2_fill_8 FILLER_32_754 ();
 sg13g2_fill_8 FILLER_32_762 ();
 sg13g2_fill_2 FILLER_32_770 ();
 sg13g2_fill_8 FILLER_32_830 ();
 sg13g2_fill_8 FILLER_32_838 ();
 sg13g2_fill_8 FILLER_32_846 ();
 sg13g2_fill_4 FILLER_32_854 ();
 sg13g2_fill_2 FILLER_32_858 ();
 sg13g2_fill_8 FILLER_32_871 ();
 sg13g2_fill_4 FILLER_32_879 ();
 sg13g2_fill_8 FILLER_32_893 ();
 sg13g2_fill_1 FILLER_32_901 ();
 sg13g2_fill_8 FILLER_32_906 ();
 sg13g2_fill_4 FILLER_32_914 ();
 sg13g2_fill_8 FILLER_32_923 ();
 sg13g2_fill_1 FILLER_32_931 ();
 sg13g2_fill_1 FILLER_32_963 ();
 sg13g2_fill_8 FILLER_32_1003 ();
 sg13g2_fill_8 FILLER_32_1011 ();
 sg13g2_fill_2 FILLER_32_1019 ();
 sg13g2_fill_1 FILLER_32_1021 ();
 sg13g2_fill_4 FILLER_32_1057 ();
 sg13g2_fill_1 FILLER_32_1061 ();
 sg13g2_fill_2 FILLER_32_1078 ();
 sg13g2_fill_1 FILLER_32_1080 ();
 sg13g2_fill_2 FILLER_32_1114 ();
 sg13g2_fill_8 FILLER_32_1146 ();
 sg13g2_fill_1 FILLER_32_1154 ();
 sg13g2_fill_2 FILLER_32_1161 ();
 sg13g2_fill_1 FILLER_32_1163 ();
 sg13g2_fill_2 FILLER_32_1190 ();
 sg13g2_fill_8 FILLER_32_1219 ();
 sg13g2_fill_4 FILLER_32_1227 ();
 sg13g2_fill_1 FILLER_32_1236 ();
 sg13g2_fill_4 FILLER_32_1263 ();
 sg13g2_fill_4 FILLER_32_1278 ();
 sg13g2_fill_8 FILLER_32_1312 ();
 sg13g2_fill_8 FILLER_32_1324 ();
 sg13g2_fill_8 FILLER_32_1332 ();
 sg13g2_fill_8 FILLER_32_1340 ();
 sg13g2_fill_8 FILLER_32_1348 ();
 sg13g2_fill_8 FILLER_32_1356 ();
 sg13g2_fill_8 FILLER_32_1364 ();
 sg13g2_fill_8 FILLER_32_1372 ();
 sg13g2_fill_8 FILLER_32_1380 ();
 sg13g2_fill_8 FILLER_32_1388 ();
 sg13g2_fill_8 FILLER_32_1396 ();
 sg13g2_fill_8 FILLER_32_1404 ();
 sg13g2_fill_8 FILLER_32_1412 ();
 sg13g2_fill_8 FILLER_32_1420 ();
 sg13g2_fill_8 FILLER_32_1428 ();
 sg13g2_fill_8 FILLER_32_1436 ();
 sg13g2_fill_8 FILLER_32_1444 ();
 sg13g2_fill_8 FILLER_32_1452 ();
 sg13g2_fill_8 FILLER_32_1460 ();
 sg13g2_fill_8 FILLER_32_1468 ();
 sg13g2_fill_8 FILLER_32_1476 ();
 sg13g2_fill_8 FILLER_32_1484 ();
 sg13g2_fill_8 FILLER_32_1492 ();
 sg13g2_fill_8 FILLER_32_1500 ();
 sg13g2_fill_8 FILLER_32_1508 ();
 sg13g2_fill_8 FILLER_32_1516 ();
 sg13g2_fill_8 FILLER_32_1524 ();
 sg13g2_fill_8 FILLER_32_1532 ();
 sg13g2_fill_8 FILLER_32_1540 ();
 sg13g2_fill_8 FILLER_32_1548 ();
 sg13g2_fill_8 FILLER_32_1556 ();
 sg13g2_fill_8 FILLER_32_1564 ();
 sg13g2_fill_8 FILLER_32_1572 ();
 sg13g2_fill_8 FILLER_32_1580 ();
 sg13g2_fill_4 FILLER_32_1588 ();
 sg13g2_fill_8 FILLER_33_0 ();
 sg13g2_fill_8 FILLER_33_8 ();
 sg13g2_fill_8 FILLER_33_16 ();
 sg13g2_fill_8 FILLER_33_24 ();
 sg13g2_fill_8 FILLER_33_32 ();
 sg13g2_fill_8 FILLER_33_40 ();
 sg13g2_fill_8 FILLER_33_48 ();
 sg13g2_fill_8 FILLER_33_56 ();
 sg13g2_fill_8 FILLER_33_64 ();
 sg13g2_fill_8 FILLER_33_72 ();
 sg13g2_fill_8 FILLER_33_80 ();
 sg13g2_fill_8 FILLER_33_88 ();
 sg13g2_fill_8 FILLER_33_96 ();
 sg13g2_fill_8 FILLER_33_104 ();
 sg13g2_fill_8 FILLER_33_112 ();
 sg13g2_fill_8 FILLER_33_156 ();
 sg13g2_fill_2 FILLER_33_164 ();
 sg13g2_fill_8 FILLER_33_186 ();
 sg13g2_fill_4 FILLER_33_194 ();
 sg13g2_fill_4 FILLER_33_208 ();
 sg13g2_fill_4 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_fill_4 FILLER_33_280 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_fill_8 FILLER_33_296 ();
 sg13g2_fill_4 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_318 ();
 sg13g2_fill_8 FILLER_33_345 ();
 sg13g2_fill_2 FILLER_33_353 ();
 sg13g2_fill_1 FILLER_33_355 ();
 sg13g2_fill_4 FILLER_33_382 ();
 sg13g2_fill_2 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_33_404 ();
 sg13g2_fill_8 FILLER_33_413 ();
 sg13g2_fill_1 FILLER_33_435 ();
 sg13g2_fill_2 FILLER_33_449 ();
 sg13g2_fill_1 FILLER_33_451 ();
 sg13g2_fill_8 FILLER_33_508 ();
 sg13g2_fill_8 FILLER_33_516 ();
 sg13g2_fill_4 FILLER_33_524 ();
 sg13g2_fill_2 FILLER_33_528 ();
 sg13g2_fill_1 FILLER_33_546 ();
 sg13g2_fill_4 FILLER_33_563 ();
 sg13g2_fill_8 FILLER_33_592 ();
 sg13g2_fill_4 FILLER_33_600 ();
 sg13g2_fill_2 FILLER_33_604 ();
 sg13g2_fill_1 FILLER_33_606 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_fill_8 FILLER_33_652 ();
 sg13g2_fill_2 FILLER_33_660 ();
 sg13g2_fill_1 FILLER_33_662 ();
 sg13g2_fill_2 FILLER_33_675 ();
 sg13g2_fill_1 FILLER_33_677 ();
 sg13g2_fill_4 FILLER_33_684 ();
 sg13g2_fill_1 FILLER_33_688 ();
 sg13g2_fill_4 FILLER_33_704 ();
 sg13g2_fill_2 FILLER_33_708 ();
 sg13g2_fill_2 FILLER_33_749 ();
 sg13g2_fill_2 FILLER_33_756 ();
 sg13g2_fill_8 FILLER_33_763 ();
 sg13g2_fill_8 FILLER_33_771 ();
 sg13g2_fill_8 FILLER_33_779 ();
 sg13g2_fill_8 FILLER_33_787 ();
 sg13g2_fill_8 FILLER_33_795 ();
 sg13g2_fill_8 FILLER_33_803 ();
 sg13g2_fill_8 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_819 ();
 sg13g2_fill_8 FILLER_33_828 ();
 sg13g2_fill_2 FILLER_33_836 ();
 sg13g2_fill_8 FILLER_33_849 ();
 sg13g2_fill_8 FILLER_33_857 ();
 sg13g2_fill_8 FILLER_33_865 ();
 sg13g2_fill_4 FILLER_33_873 ();
 sg13g2_fill_1 FILLER_33_877 ();
 sg13g2_fill_2 FILLER_33_903 ();
 sg13g2_fill_8 FILLER_33_911 ();
 sg13g2_fill_4 FILLER_33_919 ();
 sg13g2_fill_2 FILLER_33_923 ();
 sg13g2_fill_1 FILLER_33_925 ();
 sg13g2_fill_8 FILLER_33_930 ();
 sg13g2_fill_8 FILLER_33_938 ();
 sg13g2_fill_2 FILLER_33_946 ();
 sg13g2_fill_1 FILLER_33_948 ();
 sg13g2_fill_2 FILLER_33_955 ();
 sg13g2_fill_8 FILLER_33_992 ();
 sg13g2_fill_8 FILLER_33_1000 ();
 sg13g2_fill_2 FILLER_33_1008 ();
 sg13g2_fill_2 FILLER_33_1016 ();
 sg13g2_fill_1 FILLER_33_1018 ();
 sg13g2_fill_1 FILLER_33_1071 ();
 sg13g2_fill_2 FILLER_33_1080 ();
 sg13g2_fill_1 FILLER_33_1082 ();
 sg13g2_fill_2 FILLER_33_1109 ();
 sg13g2_fill_1 FILLER_33_1111 ();
 sg13g2_fill_1 FILLER_33_1118 ();
 sg13g2_fill_8 FILLER_33_1127 ();
 sg13g2_fill_8 FILLER_33_1135 ();
 sg13g2_fill_2 FILLER_33_1143 ();
 sg13g2_fill_8 FILLER_33_1177 ();
 sg13g2_fill_8 FILLER_33_1185 ();
 sg13g2_fill_2 FILLER_33_1193 ();
 sg13g2_fill_1 FILLER_33_1195 ();
 sg13g2_fill_1 FILLER_33_1226 ();
 sg13g2_fill_4 FILLER_33_1233 ();
 sg13g2_fill_8 FILLER_33_1247 ();
 sg13g2_fill_8 FILLER_33_1255 ();
 sg13g2_fill_4 FILLER_33_1263 ();
 sg13g2_fill_2 FILLER_33_1267 ();
 sg13g2_fill_1 FILLER_33_1269 ();
 sg13g2_fill_8 FILLER_33_1284 ();
 sg13g2_fill_8 FILLER_33_1292 ();
 sg13g2_fill_8 FILLER_33_1300 ();
 sg13g2_fill_8 FILLER_33_1308 ();
 sg13g2_fill_1 FILLER_33_1316 ();
 sg13g2_fill_8 FILLER_33_1323 ();
 sg13g2_fill_8 FILLER_33_1331 ();
 sg13g2_fill_8 FILLER_33_1339 ();
 sg13g2_fill_8 FILLER_33_1347 ();
 sg13g2_fill_8 FILLER_33_1355 ();
 sg13g2_fill_8 FILLER_33_1363 ();
 sg13g2_fill_8 FILLER_33_1371 ();
 sg13g2_fill_8 FILLER_33_1379 ();
 sg13g2_fill_8 FILLER_33_1387 ();
 sg13g2_fill_8 FILLER_33_1395 ();
 sg13g2_fill_8 FILLER_33_1403 ();
 sg13g2_fill_8 FILLER_33_1411 ();
 sg13g2_fill_8 FILLER_33_1419 ();
 sg13g2_fill_8 FILLER_33_1427 ();
 sg13g2_fill_8 FILLER_33_1435 ();
 sg13g2_fill_8 FILLER_33_1443 ();
 sg13g2_fill_8 FILLER_33_1451 ();
 sg13g2_fill_8 FILLER_33_1459 ();
 sg13g2_fill_8 FILLER_33_1467 ();
 sg13g2_fill_8 FILLER_33_1475 ();
 sg13g2_fill_8 FILLER_33_1483 ();
 sg13g2_fill_8 FILLER_33_1491 ();
 sg13g2_fill_8 FILLER_33_1499 ();
 sg13g2_fill_8 FILLER_33_1507 ();
 sg13g2_fill_8 FILLER_33_1515 ();
 sg13g2_fill_8 FILLER_33_1523 ();
 sg13g2_fill_8 FILLER_33_1531 ();
 sg13g2_fill_8 FILLER_33_1539 ();
 sg13g2_fill_8 FILLER_33_1547 ();
 sg13g2_fill_8 FILLER_33_1555 ();
 sg13g2_fill_8 FILLER_33_1563 ();
 sg13g2_fill_8 FILLER_33_1571 ();
 sg13g2_fill_8 FILLER_33_1579 ();
 sg13g2_fill_4 FILLER_33_1587 ();
 sg13g2_fill_1 FILLER_33_1591 ();
 sg13g2_fill_8 FILLER_34_0 ();
 sg13g2_fill_8 FILLER_34_8 ();
 sg13g2_fill_8 FILLER_34_16 ();
 sg13g2_fill_8 FILLER_34_24 ();
 sg13g2_fill_8 FILLER_34_32 ();
 sg13g2_fill_8 FILLER_34_40 ();
 sg13g2_fill_8 FILLER_34_48 ();
 sg13g2_fill_8 FILLER_34_56 ();
 sg13g2_fill_8 FILLER_34_64 ();
 sg13g2_fill_8 FILLER_34_72 ();
 sg13g2_fill_8 FILLER_34_80 ();
 sg13g2_fill_8 FILLER_34_88 ();
 sg13g2_fill_4 FILLER_34_96 ();
 sg13g2_fill_2 FILLER_34_100 ();
 sg13g2_fill_8 FILLER_34_128 ();
 sg13g2_fill_8 FILLER_34_136 ();
 sg13g2_fill_4 FILLER_34_144 ();
 sg13g2_fill_8 FILLER_34_173 ();
 sg13g2_fill_8 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_189 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_8 FILLER_34_202 ();
 sg13g2_fill_8 FILLER_34_210 ();
 sg13g2_fill_4 FILLER_34_218 ();
 sg13g2_fill_4 FILLER_34_225 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_8 FILLER_34_256 ();
 sg13g2_fill_4 FILLER_34_264 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_297 ();
 sg13g2_fill_4 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_4 FILLER_34_339 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_8 FILLER_34_369 ();
 sg13g2_fill_8 FILLER_34_395 ();
 sg13g2_fill_8 FILLER_34_403 ();
 sg13g2_fill_8 FILLER_34_411 ();
 sg13g2_fill_8 FILLER_34_419 ();
 sg13g2_fill_8 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_441 ();
 sg13g2_fill_2 FILLER_34_490 ();
 sg13g2_fill_4 FILLER_34_502 ();
 sg13g2_fill_2 FILLER_34_506 ();
 sg13g2_fill_8 FILLER_34_544 ();
 sg13g2_fill_8 FILLER_34_552 ();
 sg13g2_fill_8 FILLER_34_560 ();
 sg13g2_fill_2 FILLER_34_611 ();
 sg13g2_fill_1 FILLER_34_622 ();
 sg13g2_fill_8 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_637 ();
 sg13g2_fill_4 FILLER_34_644 ();
 sg13g2_fill_8 FILLER_34_653 ();
 sg13g2_fill_8 FILLER_34_661 ();
 sg13g2_fill_8 FILLER_34_669 ();
 sg13g2_fill_1 FILLER_34_677 ();
 sg13g2_fill_8 FILLER_34_701 ();
 sg13g2_fill_4 FILLER_34_709 ();
 sg13g2_fill_2 FILLER_34_713 ();
 sg13g2_fill_8 FILLER_34_785 ();
 sg13g2_fill_4 FILLER_34_793 ();
 sg13g2_fill_2 FILLER_34_803 ();
 sg13g2_fill_4 FILLER_34_816 ();
 sg13g2_fill_2 FILLER_34_820 ();
 sg13g2_fill_1 FILLER_34_822 ();
 sg13g2_fill_4 FILLER_34_847 ();
 sg13g2_fill_1 FILLER_34_851 ();
 sg13g2_fill_4 FILLER_34_888 ();
 sg13g2_fill_2 FILLER_34_912 ();
 sg13g2_fill_1 FILLER_34_914 ();
 sg13g2_fill_4 FILLER_34_939 ();
 sg13g2_fill_1 FILLER_34_957 ();
 sg13g2_fill_2 FILLER_34_971 ();
 sg13g2_fill_8 FILLER_34_981 ();
 sg13g2_fill_1 FILLER_34_989 ();
 sg13g2_fill_4 FILLER_34_1016 ();
 sg13g2_fill_2 FILLER_34_1020 ();
 sg13g2_fill_8 FILLER_34_1027 ();
 sg13g2_fill_2 FILLER_34_1035 ();
 sg13g2_fill_1 FILLER_34_1037 ();
 sg13g2_fill_1 FILLER_34_1048 ();
 sg13g2_fill_1 FILLER_34_1068 ();
 sg13g2_fill_8 FILLER_34_1085 ();
 sg13g2_fill_2 FILLER_34_1093 ();
 sg13g2_fill_4 FILLER_34_1120 ();
 sg13g2_fill_2 FILLER_34_1124 ();
 sg13g2_fill_8 FILLER_34_1184 ();
 sg13g2_fill_4 FILLER_34_1192 ();
 sg13g2_fill_2 FILLER_34_1196 ();
 sg13g2_fill_1 FILLER_34_1198 ();
 sg13g2_fill_2 FILLER_34_1209 ();
 sg13g2_fill_1 FILLER_34_1211 ();
 sg13g2_fill_1 FILLER_34_1238 ();
 sg13g2_fill_2 FILLER_34_1275 ();
 sg13g2_fill_1 FILLER_34_1277 ();
 sg13g2_fill_8 FILLER_34_1330 ();
 sg13g2_fill_8 FILLER_34_1338 ();
 sg13g2_fill_8 FILLER_34_1346 ();
 sg13g2_fill_8 FILLER_34_1354 ();
 sg13g2_fill_8 FILLER_34_1362 ();
 sg13g2_fill_8 FILLER_34_1370 ();
 sg13g2_fill_8 FILLER_34_1378 ();
 sg13g2_fill_8 FILLER_34_1386 ();
 sg13g2_fill_8 FILLER_34_1394 ();
 sg13g2_fill_8 FILLER_34_1402 ();
 sg13g2_fill_8 FILLER_34_1410 ();
 sg13g2_fill_8 FILLER_34_1418 ();
 sg13g2_fill_8 FILLER_34_1426 ();
 sg13g2_fill_8 FILLER_34_1434 ();
 sg13g2_fill_8 FILLER_34_1442 ();
 sg13g2_fill_8 FILLER_34_1450 ();
 sg13g2_fill_8 FILLER_34_1458 ();
 sg13g2_fill_8 FILLER_34_1466 ();
 sg13g2_fill_8 FILLER_34_1474 ();
 sg13g2_fill_8 FILLER_34_1482 ();
 sg13g2_fill_8 FILLER_34_1490 ();
 sg13g2_fill_8 FILLER_34_1498 ();
 sg13g2_fill_8 FILLER_34_1506 ();
 sg13g2_fill_8 FILLER_34_1514 ();
 sg13g2_fill_8 FILLER_34_1522 ();
 sg13g2_fill_8 FILLER_34_1530 ();
 sg13g2_fill_8 FILLER_34_1538 ();
 sg13g2_fill_8 FILLER_34_1546 ();
 sg13g2_fill_8 FILLER_34_1554 ();
 sg13g2_fill_8 FILLER_34_1562 ();
 sg13g2_fill_8 FILLER_34_1570 ();
 sg13g2_fill_8 FILLER_34_1578 ();
 sg13g2_fill_4 FILLER_34_1586 ();
 sg13g2_fill_2 FILLER_34_1590 ();
 sg13g2_fill_8 FILLER_35_0 ();
 sg13g2_fill_8 FILLER_35_8 ();
 sg13g2_fill_8 FILLER_35_16 ();
 sg13g2_fill_8 FILLER_35_24 ();
 sg13g2_fill_8 FILLER_35_32 ();
 sg13g2_fill_8 FILLER_35_40 ();
 sg13g2_fill_8 FILLER_35_48 ();
 sg13g2_fill_8 FILLER_35_56 ();
 sg13g2_fill_8 FILLER_35_64 ();
 sg13g2_fill_8 FILLER_35_72 ();
 sg13g2_fill_8 FILLER_35_80 ();
 sg13g2_fill_8 FILLER_35_88 ();
 sg13g2_fill_8 FILLER_35_96 ();
 sg13g2_fill_8 FILLER_35_104 ();
 sg13g2_fill_4 FILLER_35_112 ();
 sg13g2_fill_8 FILLER_35_136 ();
 sg13g2_fill_4 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_4 FILLER_35_187 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_1 FILLER_35_193 ();
 sg13g2_fill_8 FILLER_35_220 ();
 sg13g2_fill_8 FILLER_35_228 ();
 sg13g2_fill_8 FILLER_35_236 ();
 sg13g2_fill_8 FILLER_35_244 ();
 sg13g2_fill_4 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_8 FILLER_35_297 ();
 sg13g2_fill_8 FILLER_35_305 ();
 sg13g2_fill_8 FILLER_35_313 ();
 sg13g2_fill_8 FILLER_35_321 ();
 sg13g2_fill_8 FILLER_35_383 ();
 sg13g2_fill_8 FILLER_35_391 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_8 FILLER_35_514 ();
 sg13g2_fill_8 FILLER_35_522 ();
 sg13g2_fill_2 FILLER_35_530 ();
 sg13g2_fill_4 FILLER_35_542 ();
 sg13g2_fill_1 FILLER_35_546 ();
 sg13g2_fill_8 FILLER_35_573 ();
 sg13g2_fill_8 FILLER_35_581 ();
 sg13g2_fill_8 FILLER_35_589 ();
 sg13g2_fill_2 FILLER_35_603 ();
 sg13g2_fill_1 FILLER_35_609 ();
 sg13g2_fill_8 FILLER_35_701 ();
 sg13g2_fill_8 FILLER_35_709 ();
 sg13g2_fill_2 FILLER_35_717 ();
 sg13g2_fill_1 FILLER_35_719 ();
 sg13g2_fill_8 FILLER_35_733 ();
 sg13g2_fill_2 FILLER_35_766 ();
 sg13g2_fill_1 FILLER_35_768 ();
 sg13g2_fill_4 FILLER_35_805 ();
 sg13g2_fill_1 FILLER_35_814 ();
 sg13g2_fill_4 FILLER_35_837 ();
 sg13g2_fill_8 FILLER_35_852 ();
 sg13g2_fill_4 FILLER_35_860 ();
 sg13g2_fill_1 FILLER_35_864 ();
 sg13g2_fill_2 FILLER_35_871 ();
 sg13g2_fill_1 FILLER_35_873 ();
 sg13g2_fill_1 FILLER_35_880 ();
 sg13g2_fill_2 FILLER_35_891 ();
 sg13g2_fill_4 FILLER_35_898 ();
 sg13g2_fill_8 FILLER_35_911 ();
 sg13g2_fill_2 FILLER_35_919 ();
 sg13g2_fill_4 FILLER_35_979 ();
 sg13g2_fill_1 FILLER_35_1009 ();
 sg13g2_fill_4 FILLER_35_1020 ();
 sg13g2_fill_2 FILLER_35_1047 ();
 sg13g2_fill_1 FILLER_35_1077 ();
 sg13g2_fill_4 FILLER_35_1082 ();
 sg13g2_fill_2 FILLER_35_1117 ();
 sg13g2_fill_1 FILLER_35_1119 ();
 sg13g2_fill_8 FILLER_35_1186 ();
 sg13g2_fill_8 FILLER_35_1194 ();
 sg13g2_fill_8 FILLER_35_1202 ();
 sg13g2_fill_4 FILLER_35_1210 ();
 sg13g2_fill_2 FILLER_35_1214 ();
 sg13g2_fill_8 FILLER_35_1221 ();
 sg13g2_fill_8 FILLER_35_1229 ();
 sg13g2_fill_8 FILLER_35_1237 ();
 sg13g2_fill_4 FILLER_35_1249 ();
 sg13g2_fill_8 FILLER_35_1258 ();
 sg13g2_fill_4 FILLER_35_1266 ();
 sg13g2_fill_1 FILLER_35_1270 ();
 sg13g2_fill_8 FILLER_35_1276 ();
 sg13g2_fill_8 FILLER_35_1284 ();
 sg13g2_fill_2 FILLER_35_1292 ();
 sg13g2_fill_8 FILLER_35_1302 ();
 sg13g2_fill_4 FILLER_35_1310 ();
 sg13g2_fill_2 FILLER_35_1314 ();
 sg13g2_fill_1 FILLER_35_1316 ();
 sg13g2_fill_1 FILLER_35_1323 ();
 sg13g2_fill_8 FILLER_35_1329 ();
 sg13g2_fill_4 FILLER_35_1337 ();
 sg13g2_fill_8 FILLER_35_1353 ();
 sg13g2_fill_8 FILLER_35_1361 ();
 sg13g2_fill_8 FILLER_35_1373 ();
 sg13g2_fill_8 FILLER_35_1381 ();
 sg13g2_fill_8 FILLER_35_1389 ();
 sg13g2_fill_8 FILLER_35_1397 ();
 sg13g2_fill_8 FILLER_35_1405 ();
 sg13g2_fill_8 FILLER_35_1413 ();
 sg13g2_fill_8 FILLER_35_1421 ();
 sg13g2_fill_8 FILLER_35_1429 ();
 sg13g2_fill_8 FILLER_35_1437 ();
 sg13g2_fill_8 FILLER_35_1445 ();
 sg13g2_fill_8 FILLER_35_1453 ();
 sg13g2_fill_8 FILLER_35_1461 ();
 sg13g2_fill_8 FILLER_35_1469 ();
 sg13g2_fill_8 FILLER_35_1477 ();
 sg13g2_fill_8 FILLER_35_1485 ();
 sg13g2_fill_8 FILLER_35_1493 ();
 sg13g2_fill_8 FILLER_35_1501 ();
 sg13g2_fill_8 FILLER_35_1509 ();
 sg13g2_fill_8 FILLER_35_1517 ();
 sg13g2_fill_8 FILLER_35_1525 ();
 sg13g2_fill_8 FILLER_35_1533 ();
 sg13g2_fill_8 FILLER_35_1541 ();
 sg13g2_fill_8 FILLER_35_1549 ();
 sg13g2_fill_8 FILLER_35_1557 ();
 sg13g2_fill_8 FILLER_35_1565 ();
 sg13g2_fill_8 FILLER_35_1573 ();
 sg13g2_fill_8 FILLER_35_1581 ();
 sg13g2_fill_2 FILLER_35_1589 ();
 sg13g2_fill_1 FILLER_35_1591 ();
 sg13g2_fill_8 FILLER_36_0 ();
 sg13g2_fill_8 FILLER_36_8 ();
 sg13g2_fill_8 FILLER_36_16 ();
 sg13g2_fill_8 FILLER_36_24 ();
 sg13g2_fill_8 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_40 ();
 sg13g2_fill_1 FILLER_36_42 ();
 sg13g2_fill_8 FILLER_36_69 ();
 sg13g2_fill_1 FILLER_36_77 ();
 sg13g2_fill_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_92 ();
 sg13g2_fill_8 FILLER_36_128 ();
 sg13g2_fill_2 FILLER_36_136 ();
 sg13g2_fill_8 FILLER_36_158 ();
 sg13g2_fill_4 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_170 ();
 sg13g2_fill_1 FILLER_36_172 ();
 sg13g2_fill_8 FILLER_36_183 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_fill_4 FILLER_36_229 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_4 FILLER_36_294 ();
 sg13g2_fill_2 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_395 ();
 sg13g2_fill_8 FILLER_36_411 ();
 sg13g2_fill_4 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_423 ();
 sg13g2_fill_8 FILLER_36_434 ();
 sg13g2_fill_1 FILLER_36_503 ();
 sg13g2_fill_8 FILLER_36_514 ();
 sg13g2_fill_8 FILLER_36_522 ();
 sg13g2_fill_2 FILLER_36_530 ();
 sg13g2_fill_1 FILLER_36_532 ();
 sg13g2_fill_4 FILLER_36_543 ();
 sg13g2_fill_8 FILLER_36_573 ();
 sg13g2_fill_8 FILLER_36_581 ();
 sg13g2_fill_2 FILLER_36_589 ();
 sg13g2_fill_4 FILLER_36_603 ();
 sg13g2_fill_2 FILLER_36_607 ();
 sg13g2_fill_1 FILLER_36_609 ();
 sg13g2_fill_8 FILLER_36_629 ();
 sg13g2_fill_8 FILLER_36_637 ();
 sg13g2_fill_8 FILLER_36_645 ();
 sg13g2_fill_8 FILLER_36_653 ();
 sg13g2_fill_2 FILLER_36_661 ();
 sg13g2_fill_2 FILLER_36_668 ();
 sg13g2_fill_2 FILLER_36_675 ();
 sg13g2_fill_1 FILLER_36_677 ();
 sg13g2_fill_2 FILLER_36_683 ();
 sg13g2_fill_2 FILLER_36_693 ();
 sg13g2_fill_1 FILLER_36_695 ();
 sg13g2_fill_8 FILLER_36_726 ();
 sg13g2_fill_2 FILLER_36_734 ();
 sg13g2_fill_8 FILLER_36_764 ();
 sg13g2_fill_8 FILLER_36_772 ();
 sg13g2_fill_2 FILLER_36_780 ();
 sg13g2_fill_8 FILLER_36_786 ();
 sg13g2_fill_2 FILLER_36_794 ();
 sg13g2_fill_1 FILLER_36_796 ();
 sg13g2_fill_4 FILLER_36_802 ();
 sg13g2_fill_2 FILLER_36_819 ();
 sg13g2_fill_8 FILLER_36_832 ();
 sg13g2_fill_1 FILLER_36_840 ();
 sg13g2_fill_2 FILLER_36_846 ();
 sg13g2_fill_1 FILLER_36_848 ();
 sg13g2_fill_2 FILLER_36_892 ();
 sg13g2_fill_8 FILLER_36_900 ();
 sg13g2_fill_8 FILLER_36_908 ();
 sg13g2_fill_4 FILLER_36_916 ();
 sg13g2_fill_8 FILLER_36_924 ();
 sg13g2_fill_1 FILLER_36_932 ();
 sg13g2_fill_1 FILLER_36_938 ();
 sg13g2_fill_1 FILLER_36_969 ();
 sg13g2_fill_8 FILLER_36_996 ();
 sg13g2_fill_1 FILLER_36_1019 ();
 sg13g2_fill_2 FILLER_36_1050 ();
 sg13g2_fill_2 FILLER_36_1116 ();
 sg13g2_fill_2 FILLER_36_1152 ();
 sg13g2_fill_8 FILLER_36_1158 ();
 sg13g2_fill_8 FILLER_36_1166 ();
 sg13g2_fill_2 FILLER_36_1174 ();
 sg13g2_fill_4 FILLER_36_1212 ();
 sg13g2_fill_1 FILLER_36_1216 ();
 sg13g2_fill_2 FILLER_36_1225 ();
 sg13g2_fill_1 FILLER_36_1227 ();
 sg13g2_fill_1 FILLER_36_1252 ();
 sg13g2_fill_8 FILLER_36_1283 ();
 sg13g2_fill_8 FILLER_36_1291 ();
 sg13g2_fill_4 FILLER_36_1299 ();
 sg13g2_fill_2 FILLER_36_1303 ();
 sg13g2_fill_1 FILLER_36_1305 ();
 sg13g2_fill_4 FILLER_36_1310 ();
 sg13g2_fill_1 FILLER_36_1324 ();
 sg13g2_fill_2 FILLER_36_1335 ();
 sg13g2_fill_1 FILLER_36_1337 ();
 sg13g2_fill_2 FILLER_36_1346 ();
 sg13g2_fill_4 FILLER_36_1356 ();
 sg13g2_fill_8 FILLER_36_1381 ();
 sg13g2_fill_8 FILLER_36_1389 ();
 sg13g2_fill_8 FILLER_36_1397 ();
 sg13g2_fill_8 FILLER_36_1405 ();
 sg13g2_fill_8 FILLER_36_1413 ();
 sg13g2_fill_8 FILLER_36_1421 ();
 sg13g2_fill_8 FILLER_36_1429 ();
 sg13g2_fill_8 FILLER_36_1437 ();
 sg13g2_fill_8 FILLER_36_1445 ();
 sg13g2_fill_8 FILLER_36_1453 ();
 sg13g2_fill_8 FILLER_36_1461 ();
 sg13g2_fill_8 FILLER_36_1469 ();
 sg13g2_fill_8 FILLER_36_1477 ();
 sg13g2_fill_8 FILLER_36_1485 ();
 sg13g2_fill_8 FILLER_36_1493 ();
 sg13g2_fill_8 FILLER_36_1501 ();
 sg13g2_fill_8 FILLER_36_1509 ();
 sg13g2_fill_8 FILLER_36_1517 ();
 sg13g2_fill_8 FILLER_36_1525 ();
 sg13g2_fill_8 FILLER_36_1533 ();
 sg13g2_fill_8 FILLER_36_1541 ();
 sg13g2_fill_8 FILLER_36_1549 ();
 sg13g2_fill_8 FILLER_36_1557 ();
 sg13g2_fill_8 FILLER_36_1565 ();
 sg13g2_fill_8 FILLER_36_1573 ();
 sg13g2_fill_8 FILLER_36_1581 ();
 sg13g2_fill_2 FILLER_36_1589 ();
 sg13g2_fill_1 FILLER_36_1591 ();
 sg13g2_fill_8 FILLER_37_0 ();
 sg13g2_fill_8 FILLER_37_8 ();
 sg13g2_fill_8 FILLER_37_16 ();
 sg13g2_fill_4 FILLER_37_24 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_8 FILLER_37_117 ();
 sg13g2_fill_8 FILLER_37_125 ();
 sg13g2_fill_4 FILLER_37_133 ();
 sg13g2_fill_1 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_fill_4 FILLER_37_203 ();
 sg13g2_fill_2 FILLER_37_207 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_1 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_257 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_fill_8 FILLER_37_270 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_8 FILLER_37_290 ();
 sg13g2_fill_4 FILLER_37_298 ();
 sg13g2_fill_8 FILLER_37_312 ();
 sg13g2_fill_8 FILLER_37_320 ();
 sg13g2_fill_8 FILLER_37_328 ();
 sg13g2_fill_4 FILLER_37_336 ();
 sg13g2_fill_1 FILLER_37_379 ();
 sg13g2_fill_4 FILLER_37_390 ();
 sg13g2_fill_2 FILLER_37_394 ();
 sg13g2_fill_1 FILLER_37_396 ();
 sg13g2_fill_4 FILLER_37_438 ();
 sg13g2_fill_1 FILLER_37_442 ();
 sg13g2_fill_8 FILLER_37_459 ();
 sg13g2_fill_4 FILLER_37_467 ();
 sg13g2_fill_2 FILLER_37_471 ();
 sg13g2_fill_2 FILLER_37_508 ();
 sg13g2_fill_1 FILLER_37_510 ();
 sg13g2_fill_4 FILLER_37_517 ();
 sg13g2_fill_1 FILLER_37_521 ();
 sg13g2_fill_8 FILLER_37_537 ();
 sg13g2_fill_2 FILLER_37_545 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_8 FILLER_37_561 ();
 sg13g2_fill_4 FILLER_37_607 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_8 FILLER_37_618 ();
 sg13g2_fill_8 FILLER_37_626 ();
 sg13g2_fill_2 FILLER_37_634 ();
 sg13g2_fill_2 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_685 ();
 sg13g2_fill_1 FILLER_37_697 ();
 sg13g2_fill_8 FILLER_37_702 ();
 sg13g2_fill_2 FILLER_37_710 ();
 sg13g2_fill_1 FILLER_37_712 ();
 sg13g2_fill_8 FILLER_37_759 ();
 sg13g2_fill_4 FILLER_37_767 ();
 sg13g2_fill_2 FILLER_37_771 ();
 sg13g2_fill_2 FILLER_37_786 ();
 sg13g2_fill_8 FILLER_37_795 ();
 sg13g2_fill_8 FILLER_37_803 ();
 sg13g2_fill_2 FILLER_37_811 ();
 sg13g2_fill_1 FILLER_37_813 ();
 sg13g2_fill_2 FILLER_37_826 ();
 sg13g2_fill_1 FILLER_37_828 ();
 sg13g2_fill_4 FILLER_37_833 ();
 sg13g2_fill_1 FILLER_37_837 ();
 sg13g2_fill_8 FILLER_37_853 ();
 sg13g2_fill_8 FILLER_37_861 ();
 sg13g2_fill_4 FILLER_37_873 ();
 sg13g2_fill_2 FILLER_37_877 ();
 sg13g2_fill_1 FILLER_37_879 ();
 sg13g2_fill_1 FILLER_37_886 ();
 sg13g2_fill_8 FILLER_37_931 ();
 sg13g2_fill_4 FILLER_37_939 ();
 sg13g2_fill_1 FILLER_37_943 ();
 sg13g2_fill_2 FILLER_37_947 ();
 sg13g2_fill_1 FILLER_37_949 ();
 sg13g2_fill_2 FILLER_37_967 ();
 sg13g2_fill_4 FILLER_37_1010 ();
 sg13g2_fill_2 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1026 ();
 sg13g2_fill_4 FILLER_37_1059 ();
 sg13g2_fill_4 FILLER_37_1069 ();
 sg13g2_fill_4 FILLER_37_1137 ();
 sg13g2_fill_1 FILLER_37_1141 ();
 sg13g2_fill_8 FILLER_37_1151 ();
 sg13g2_fill_1 FILLER_37_1159 ();
 sg13g2_fill_8 FILLER_37_1168 ();
 sg13g2_fill_2 FILLER_37_1176 ();
 sg13g2_fill_4 FILLER_37_1184 ();
 sg13g2_fill_2 FILLER_37_1218 ();
 sg13g2_fill_1 FILLER_37_1228 ();
 sg13g2_fill_2 FILLER_37_1259 ();
 sg13g2_fill_4 FILLER_37_1269 ();
 sg13g2_fill_2 FILLER_37_1273 ();
 sg13g2_fill_4 FILLER_37_1311 ();
 sg13g2_fill_2 FILLER_37_1315 ();
 sg13g2_fill_1 FILLER_37_1317 ();
 sg13g2_fill_2 FILLER_37_1324 ();
 sg13g2_fill_8 FILLER_37_1331 ();
 sg13g2_fill_4 FILLER_37_1339 ();
 sg13g2_fill_4 FILLER_37_1347 ();
 sg13g2_fill_2 FILLER_37_1351 ();
 sg13g2_fill_8 FILLER_37_1357 ();
 sg13g2_fill_8 FILLER_37_1365 ();
 sg13g2_fill_8 FILLER_37_1373 ();
 sg13g2_fill_8 FILLER_37_1381 ();
 sg13g2_fill_8 FILLER_37_1389 ();
 sg13g2_fill_8 FILLER_37_1397 ();
 sg13g2_fill_8 FILLER_37_1405 ();
 sg13g2_fill_8 FILLER_37_1413 ();
 sg13g2_fill_8 FILLER_37_1421 ();
 sg13g2_fill_8 FILLER_37_1429 ();
 sg13g2_fill_8 FILLER_37_1437 ();
 sg13g2_fill_8 FILLER_37_1445 ();
 sg13g2_fill_8 FILLER_37_1453 ();
 sg13g2_fill_8 FILLER_37_1461 ();
 sg13g2_fill_8 FILLER_37_1469 ();
 sg13g2_fill_8 FILLER_37_1477 ();
 sg13g2_fill_8 FILLER_37_1485 ();
 sg13g2_fill_8 FILLER_37_1493 ();
 sg13g2_fill_8 FILLER_37_1501 ();
 sg13g2_fill_8 FILLER_37_1509 ();
 sg13g2_fill_8 FILLER_37_1517 ();
 sg13g2_fill_8 FILLER_37_1525 ();
 sg13g2_fill_8 FILLER_37_1533 ();
 sg13g2_fill_8 FILLER_37_1541 ();
 sg13g2_fill_8 FILLER_37_1549 ();
 sg13g2_fill_8 FILLER_37_1557 ();
 sg13g2_fill_8 FILLER_37_1565 ();
 sg13g2_fill_8 FILLER_37_1573 ();
 sg13g2_fill_8 FILLER_37_1581 ();
 sg13g2_fill_2 FILLER_37_1589 ();
 sg13g2_fill_1 FILLER_37_1591 ();
 sg13g2_fill_8 FILLER_38_0 ();
 sg13g2_fill_8 FILLER_38_8 ();
 sg13g2_fill_8 FILLER_38_16 ();
 sg13g2_fill_1 FILLER_38_24 ();
 sg13g2_fill_8 FILLER_38_45 ();
 sg13g2_fill_1 FILLER_38_53 ();
 sg13g2_fill_8 FILLER_38_74 ();
 sg13g2_fill_8 FILLER_38_144 ();
 sg13g2_fill_8 FILLER_38_152 ();
 sg13g2_fill_8 FILLER_38_160 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_fill_8 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_fill_4 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_208 ();
 sg13g2_fill_1 FILLER_38_210 ();
 sg13g2_fill_4 FILLER_38_221 ();
 sg13g2_fill_8 FILLER_38_231 ();
 sg13g2_fill_8 FILLER_38_239 ();
 sg13g2_fill_2 FILLER_38_247 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_8 FILLER_38_296 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_306 ();
 sg13g2_fill_4 FILLER_38_327 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_fill_8 FILLER_38_342 ();
 sg13g2_fill_8 FILLER_38_350 ();
 sg13g2_fill_4 FILLER_38_358 ();
 sg13g2_fill_2 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_8 FILLER_38_391 ();
 sg13g2_fill_4 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_403 ();
 sg13g2_fill_1 FILLER_38_405 ();
 sg13g2_fill_4 FILLER_38_414 ();
 sg13g2_fill_2 FILLER_38_418 ();
 sg13g2_fill_8 FILLER_38_462 ();
 sg13g2_fill_2 FILLER_38_470 ();
 sg13g2_fill_1 FILLER_38_472 ();
 sg13g2_fill_2 FILLER_38_499 ();
 sg13g2_fill_1 FILLER_38_501 ();
 sg13g2_fill_8 FILLER_38_518 ();
 sg13g2_fill_4 FILLER_38_526 ();
 sg13g2_fill_4 FILLER_38_540 ();
 sg13g2_fill_4 FILLER_38_551 ();
 sg13g2_fill_1 FILLER_38_555 ();
 sg13g2_fill_8 FILLER_38_566 ();
 sg13g2_fill_8 FILLER_38_574 ();
 sg13g2_fill_8 FILLER_38_582 ();
 sg13g2_fill_4 FILLER_38_590 ();
 sg13g2_fill_2 FILLER_38_594 ();
 sg13g2_fill_2 FILLER_38_601 ();
 sg13g2_fill_1 FILLER_38_603 ();
 sg13g2_fill_8 FILLER_38_622 ();
 sg13g2_fill_2 FILLER_38_630 ();
 sg13g2_fill_8 FILLER_38_640 ();
 sg13g2_fill_8 FILLER_38_703 ();
 sg13g2_fill_8 FILLER_38_711 ();
 sg13g2_fill_8 FILLER_38_719 ();
 sg13g2_fill_4 FILLER_38_727 ();
 sg13g2_fill_1 FILLER_38_731 ();
 sg13g2_fill_1 FILLER_38_774 ();
 sg13g2_fill_2 FILLER_38_804 ();
 sg13g2_fill_1 FILLER_38_806 ();
 sg13g2_fill_1 FILLER_38_822 ();
 sg13g2_fill_4 FILLER_38_828 ();
 sg13g2_fill_2 FILLER_38_832 ();
 sg13g2_fill_1 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_38_853 ();
 sg13g2_fill_8 FILLER_38_895 ();
 sg13g2_fill_2 FILLER_38_903 ();
 sg13g2_fill_8 FILLER_38_923 ();
 sg13g2_fill_8 FILLER_38_931 ();
 sg13g2_fill_8 FILLER_38_939 ();
 sg13g2_fill_8 FILLER_38_947 ();
 sg13g2_fill_8 FILLER_38_955 ();
 sg13g2_fill_1 FILLER_38_963 ();
 sg13g2_fill_8 FILLER_38_970 ();
 sg13g2_fill_8 FILLER_38_978 ();
 sg13g2_fill_8 FILLER_38_986 ();
 sg13g2_fill_8 FILLER_38_994 ();
 sg13g2_fill_1 FILLER_38_1002 ();
 sg13g2_fill_2 FILLER_38_1045 ();
 sg13g2_fill_1 FILLER_38_1047 ();
 sg13g2_fill_2 FILLER_38_1088 ();
 sg13g2_fill_8 FILLER_38_1095 ();
 sg13g2_fill_8 FILLER_38_1103 ();
 sg13g2_fill_8 FILLER_38_1111 ();
 sg13g2_fill_8 FILLER_38_1119 ();
 sg13g2_fill_8 FILLER_38_1127 ();
 sg13g2_fill_8 FILLER_38_1135 ();
 sg13g2_fill_2 FILLER_38_1143 ();
 sg13g2_fill_1 FILLER_38_1145 ();
 sg13g2_fill_8 FILLER_38_1160 ();
 sg13g2_fill_4 FILLER_38_1168 ();
 sg13g2_fill_2 FILLER_38_1172 ();
 sg13g2_fill_1 FILLER_38_1174 ();
 sg13g2_fill_8 FILLER_38_1211 ();
 sg13g2_fill_2 FILLER_38_1219 ();
 sg13g2_fill_1 FILLER_38_1226 ();
 sg13g2_fill_1 FILLER_38_1258 ();
 sg13g2_fill_8 FILLER_38_1265 ();
 sg13g2_fill_2 FILLER_38_1273 ();
 sg13g2_fill_1 FILLER_38_1311 ();
 sg13g2_fill_8 FILLER_38_1324 ();
 sg13g2_fill_4 FILLER_38_1332 ();
 sg13g2_fill_2 FILLER_38_1336 ();
 sg13g2_fill_1 FILLER_38_1338 ();
 sg13g2_fill_4 FILLER_38_1351 ();
 sg13g2_fill_1 FILLER_38_1373 ();
 sg13g2_fill_8 FILLER_38_1383 ();
 sg13g2_fill_8 FILLER_38_1391 ();
 sg13g2_fill_8 FILLER_38_1399 ();
 sg13g2_fill_8 FILLER_38_1407 ();
 sg13g2_fill_8 FILLER_38_1415 ();
 sg13g2_fill_8 FILLER_38_1423 ();
 sg13g2_fill_8 FILLER_38_1431 ();
 sg13g2_fill_8 FILLER_38_1439 ();
 sg13g2_fill_8 FILLER_38_1447 ();
 sg13g2_fill_8 FILLER_38_1455 ();
 sg13g2_fill_8 FILLER_38_1463 ();
 sg13g2_fill_8 FILLER_38_1471 ();
 sg13g2_fill_8 FILLER_38_1479 ();
 sg13g2_fill_8 FILLER_38_1487 ();
 sg13g2_fill_8 FILLER_38_1495 ();
 sg13g2_fill_8 FILLER_38_1503 ();
 sg13g2_fill_8 FILLER_38_1511 ();
 sg13g2_fill_8 FILLER_38_1519 ();
 sg13g2_fill_8 FILLER_38_1527 ();
 sg13g2_fill_8 FILLER_38_1535 ();
 sg13g2_fill_8 FILLER_38_1543 ();
 sg13g2_fill_8 FILLER_38_1551 ();
 sg13g2_fill_8 FILLER_38_1559 ();
 sg13g2_fill_8 FILLER_38_1567 ();
 sg13g2_fill_8 FILLER_38_1575 ();
 sg13g2_fill_8 FILLER_38_1583 ();
 sg13g2_fill_1 FILLER_38_1591 ();
 sg13g2_fill_8 FILLER_39_0 ();
 sg13g2_fill_8 FILLER_39_8 ();
 sg13g2_fill_8 FILLER_39_16 ();
 sg13g2_fill_8 FILLER_39_24 ();
 sg13g2_fill_8 FILLER_39_57 ();
 sg13g2_fill_2 FILLER_39_65 ();
 sg13g2_fill_1 FILLER_39_67 ();
 sg13g2_fill_4 FILLER_39_78 ();
 sg13g2_fill_2 FILLER_39_82 ();
 sg13g2_fill_1 FILLER_39_84 ();
 sg13g2_fill_8 FILLER_39_95 ();
 sg13g2_fill_8 FILLER_39_103 ();
 sg13g2_fill_8 FILLER_39_111 ();
 sg13g2_fill_8 FILLER_39_119 ();
 sg13g2_fill_4 FILLER_39_163 ();
 sg13g2_fill_2 FILLER_39_167 ();
 sg13g2_fill_2 FILLER_39_179 ();
 sg13g2_fill_1 FILLER_39_201 ();
 sg13g2_fill_8 FILLER_39_212 ();
 sg13g2_fill_4 FILLER_39_220 ();
 sg13g2_fill_8 FILLER_39_230 ();
 sg13g2_fill_8 FILLER_39_238 ();
 sg13g2_fill_2 FILLER_39_246 ();
 sg13g2_fill_1 FILLER_39_248 ();
 sg13g2_fill_4 FILLER_39_259 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_8 FILLER_39_270 ();
 sg13g2_fill_8 FILLER_39_278 ();
 sg13g2_fill_1 FILLER_39_286 ();
 sg13g2_fill_4 FILLER_39_303 ();
 sg13g2_fill_2 FILLER_39_307 ();
 sg13g2_fill_2 FILLER_39_329 ();
 sg13g2_fill_8 FILLER_39_357 ();
 sg13g2_fill_8 FILLER_39_365 ();
 sg13g2_fill_8 FILLER_39_373 ();
 sg13g2_fill_4 FILLER_39_381 ();
 sg13g2_fill_2 FILLER_39_385 ();
 sg13g2_fill_8 FILLER_39_395 ();
 sg13g2_fill_8 FILLER_39_413 ();
 sg13g2_fill_8 FILLER_39_421 ();
 sg13g2_fill_8 FILLER_39_465 ();
 sg13g2_fill_4 FILLER_39_473 ();
 sg13g2_fill_1 FILLER_39_477 ();
 sg13g2_fill_4 FILLER_39_488 ();
 sg13g2_fill_2 FILLER_39_492 ();
 sg13g2_fill_4 FILLER_39_499 ();
 sg13g2_fill_1 FILLER_39_503 ();
 sg13g2_fill_4 FILLER_39_512 ();
 sg13g2_fill_2 FILLER_39_516 ();
 sg13g2_fill_1 FILLER_39_518 ();
 sg13g2_fill_8 FILLER_39_560 ();
 sg13g2_fill_8 FILLER_39_568 ();
 sg13g2_fill_2 FILLER_39_602 ();
 sg13g2_fill_1 FILLER_39_604 ();
 sg13g2_fill_4 FILLER_39_631 ();
 sg13g2_fill_2 FILLER_39_635 ();
 sg13g2_fill_1 FILLER_39_637 ();
 sg13g2_fill_1 FILLER_39_661 ();
 sg13g2_fill_4 FILLER_39_716 ();
 sg13g2_fill_2 FILLER_39_720 ();
 sg13g2_fill_1 FILLER_39_722 ();
 sg13g2_fill_1 FILLER_39_734 ();
 sg13g2_fill_2 FILLER_39_783 ();
 sg13g2_fill_1 FILLER_39_807 ();
 sg13g2_fill_2 FILLER_39_814 ();
 sg13g2_fill_4 FILLER_39_834 ();
 sg13g2_fill_4 FILLER_39_849 ();
 sg13g2_fill_1 FILLER_39_884 ();
 sg13g2_fill_8 FILLER_39_895 ();
 sg13g2_fill_4 FILLER_39_903 ();
 sg13g2_fill_1 FILLER_39_907 ();
 sg13g2_fill_1 FILLER_39_913 ();
 sg13g2_fill_8 FILLER_39_920 ();
 sg13g2_fill_2 FILLER_39_928 ();
 sg13g2_fill_1 FILLER_39_930 ();
 sg13g2_fill_8 FILLER_39_974 ();
 sg13g2_fill_4 FILLER_39_1008 ();
 sg13g2_fill_4 FILLER_39_1067 ();
 sg13g2_fill_1 FILLER_39_1071 ();
 sg13g2_fill_4 FILLER_39_1084 ();
 sg13g2_fill_4 FILLER_39_1093 ();
 sg13g2_fill_2 FILLER_39_1097 ();
 sg13g2_fill_1 FILLER_39_1099 ();
 sg13g2_fill_8 FILLER_39_1126 ();
 sg13g2_fill_4 FILLER_39_1134 ();
 sg13g2_fill_1 FILLER_39_1138 ();
 sg13g2_fill_8 FILLER_39_1179 ();
 sg13g2_fill_8 FILLER_39_1187 ();
 sg13g2_fill_8 FILLER_39_1195 ();
 sg13g2_fill_1 FILLER_39_1203 ();
 sg13g2_fill_8 FILLER_39_1210 ();
 sg13g2_fill_2 FILLER_39_1218 ();
 sg13g2_fill_1 FILLER_39_1220 ();
 sg13g2_fill_8 FILLER_39_1284 ();
 sg13g2_fill_8 FILLER_39_1292 ();
 sg13g2_fill_8 FILLER_39_1300 ();
 sg13g2_fill_8 FILLER_39_1308 ();
 sg13g2_fill_4 FILLER_39_1321 ();
 sg13g2_fill_1 FILLER_39_1325 ();
 sg13g2_fill_1 FILLER_39_1334 ();
 sg13g2_fill_4 FILLER_39_1356 ();
 sg13g2_fill_2 FILLER_39_1360 ();
 sg13g2_fill_1 FILLER_39_1362 ();
 sg13g2_fill_8 FILLER_39_1387 ();
 sg13g2_fill_8 FILLER_39_1395 ();
 sg13g2_fill_8 FILLER_39_1403 ();
 sg13g2_fill_8 FILLER_39_1411 ();
 sg13g2_fill_8 FILLER_39_1419 ();
 sg13g2_fill_8 FILLER_39_1427 ();
 sg13g2_fill_8 FILLER_39_1435 ();
 sg13g2_fill_8 FILLER_39_1443 ();
 sg13g2_fill_8 FILLER_39_1451 ();
 sg13g2_fill_8 FILLER_39_1459 ();
 sg13g2_fill_8 FILLER_39_1467 ();
 sg13g2_fill_8 FILLER_39_1475 ();
 sg13g2_fill_8 FILLER_39_1483 ();
 sg13g2_fill_8 FILLER_39_1491 ();
 sg13g2_fill_8 FILLER_39_1499 ();
 sg13g2_fill_8 FILLER_39_1507 ();
 sg13g2_fill_8 FILLER_39_1515 ();
 sg13g2_fill_8 FILLER_39_1523 ();
 sg13g2_fill_8 FILLER_39_1531 ();
 sg13g2_fill_8 FILLER_39_1539 ();
 sg13g2_fill_8 FILLER_39_1547 ();
 sg13g2_fill_8 FILLER_39_1555 ();
 sg13g2_fill_8 FILLER_39_1563 ();
 sg13g2_fill_8 FILLER_39_1571 ();
 sg13g2_fill_8 FILLER_39_1579 ();
 sg13g2_fill_4 FILLER_39_1587 ();
 sg13g2_fill_1 FILLER_39_1591 ();
 sg13g2_fill_8 FILLER_40_0 ();
 sg13g2_fill_8 FILLER_40_68 ();
 sg13g2_fill_8 FILLER_40_76 ();
 sg13g2_fill_8 FILLER_40_84 ();
 sg13g2_fill_4 FILLER_40_92 ();
 sg13g2_fill_2 FILLER_40_96 ();
 sg13g2_fill_8 FILLER_40_142 ();
 sg13g2_fill_8 FILLER_40_150 ();
 sg13g2_fill_4 FILLER_40_158 ();
 sg13g2_fill_2 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_164 ();
 sg13g2_fill_8 FILLER_40_173 ();
 sg13g2_fill_4 FILLER_40_181 ();
 sg13g2_fill_4 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_201 ();
 sg13g2_fill_4 FILLER_40_229 ();
 sg13g2_fill_1 FILLER_40_251 ();
 sg13g2_fill_4 FILLER_40_262 ();
 sg13g2_fill_8 FILLER_40_274 ();
 sg13g2_fill_8 FILLER_40_282 ();
 sg13g2_fill_2 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_8 FILLER_40_309 ();
 sg13g2_fill_4 FILLER_40_317 ();
 sg13g2_fill_8 FILLER_40_333 ();
 sg13g2_fill_1 FILLER_40_341 ();
 sg13g2_fill_8 FILLER_40_362 ();
 sg13g2_fill_8 FILLER_40_370 ();
 sg13g2_fill_2 FILLER_40_378 ();
 sg13g2_fill_4 FILLER_40_396 ();
 sg13g2_fill_2 FILLER_40_400 ();
 sg13g2_fill_8 FILLER_40_442 ();
 sg13g2_fill_8 FILLER_40_450 ();
 sg13g2_fill_4 FILLER_40_458 ();
 sg13g2_fill_1 FILLER_40_462 ();
 sg13g2_fill_8 FILLER_40_489 ();
 sg13g2_fill_8 FILLER_40_497 ();
 sg13g2_fill_8 FILLER_40_505 ();
 sg13g2_fill_8 FILLER_40_513 ();
 sg13g2_fill_4 FILLER_40_521 ();
 sg13g2_fill_8 FILLER_40_533 ();
 sg13g2_fill_2 FILLER_40_541 ();
 sg13g2_fill_1 FILLER_40_543 ();
 sg13g2_fill_4 FILLER_40_580 ();
 sg13g2_fill_8 FILLER_40_592 ();
 sg13g2_fill_8 FILLER_40_600 ();
 sg13g2_fill_1 FILLER_40_625 ();
 sg13g2_fill_1 FILLER_40_681 ();
 sg13g2_fill_2 FILLER_40_695 ();
 sg13g2_fill_8 FILLER_40_730 ();
 sg13g2_fill_4 FILLER_40_738 ();
 sg13g2_fill_1 FILLER_40_742 ();
 sg13g2_fill_2 FILLER_40_750 ();
 sg13g2_fill_1 FILLER_40_752 ();
 sg13g2_fill_4 FILLER_40_759 ();
 sg13g2_fill_1 FILLER_40_763 ();
 sg13g2_fill_2 FILLER_40_793 ();
 sg13g2_fill_1 FILLER_40_819 ();
 sg13g2_fill_2 FILLER_40_826 ();
 sg13g2_fill_8 FILLER_40_849 ();
 sg13g2_fill_2 FILLER_40_862 ();
 sg13g2_fill_1 FILLER_40_864 ();
 sg13g2_fill_4 FILLER_40_890 ();
 sg13g2_fill_2 FILLER_40_905 ();
 sg13g2_fill_1 FILLER_40_907 ();
 sg13g2_fill_8 FILLER_40_919 ();
 sg13g2_fill_1 FILLER_40_927 ();
 sg13g2_fill_2 FILLER_40_954 ();
 sg13g2_fill_1 FILLER_40_968 ();
 sg13g2_fill_4 FILLER_40_995 ();
 sg13g2_fill_4 FILLER_40_1022 ();
 sg13g2_fill_1 FILLER_40_1026 ();
 sg13g2_fill_8 FILLER_40_1032 ();
 sg13g2_fill_2 FILLER_40_1040 ();
 sg13g2_fill_1 FILLER_40_1042 ();
 sg13g2_fill_2 FILLER_40_1074 ();
 sg13g2_fill_1 FILLER_40_1081 ();
 sg13g2_fill_2 FILLER_40_1097 ();
 sg13g2_fill_1 FILLER_40_1099 ();
 sg13g2_fill_8 FILLER_40_1161 ();
 sg13g2_fill_8 FILLER_40_1169 ();
 sg13g2_fill_8 FILLER_40_1182 ();
 sg13g2_fill_8 FILLER_40_1190 ();
 sg13g2_fill_2 FILLER_40_1220 ();
 sg13g2_fill_4 FILLER_40_1291 ();
 sg13g2_fill_8 FILLER_40_1306 ();
 sg13g2_fill_1 FILLER_40_1314 ();
 sg13g2_fill_4 FILLER_40_1337 ();
 sg13g2_fill_1 FILLER_40_1341 ();
 sg13g2_fill_8 FILLER_40_1354 ();
 sg13g2_fill_4 FILLER_40_1362 ();
 sg13g2_fill_4 FILLER_40_1374 ();
 sg13g2_fill_2 FILLER_40_1378 ();
 sg13g2_fill_4 FILLER_40_1398 ();
 sg13g2_fill_2 FILLER_40_1402 ();
 sg13g2_fill_8 FILLER_40_1412 ();
 sg13g2_fill_8 FILLER_40_1420 ();
 sg13g2_fill_8 FILLER_40_1428 ();
 sg13g2_fill_8 FILLER_40_1436 ();
 sg13g2_fill_8 FILLER_40_1444 ();
 sg13g2_fill_8 FILLER_40_1452 ();
 sg13g2_fill_8 FILLER_40_1460 ();
 sg13g2_fill_8 FILLER_40_1468 ();
 sg13g2_fill_8 FILLER_40_1476 ();
 sg13g2_fill_4 FILLER_40_1484 ();
 sg13g2_fill_8 FILLER_40_1528 ();
 sg13g2_fill_8 FILLER_40_1536 ();
 sg13g2_fill_8 FILLER_40_1544 ();
 sg13g2_fill_8 FILLER_40_1552 ();
 sg13g2_fill_8 FILLER_40_1560 ();
 sg13g2_fill_8 FILLER_40_1568 ();
 sg13g2_fill_8 FILLER_40_1576 ();
 sg13g2_fill_8 FILLER_40_1584 ();
 sg13g2_fill_8 FILLER_41_0 ();
 sg13g2_fill_8 FILLER_41_8 ();
 sg13g2_fill_8 FILLER_41_16 ();
 sg13g2_fill_4 FILLER_41_24 ();
 sg13g2_fill_1 FILLER_41_28 ();
 sg13g2_fill_4 FILLER_41_45 ();
 sg13g2_fill_1 FILLER_41_49 ();
 sg13g2_fill_4 FILLER_41_60 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_4 FILLER_41_110 ();
 sg13g2_fill_8 FILLER_41_134 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_fill_8 FILLER_41_169 ();
 sg13g2_fill_8 FILLER_41_177 ();
 sg13g2_fill_8 FILLER_41_185 ();
 sg13g2_fill_8 FILLER_41_203 ();
 sg13g2_fill_4 FILLER_41_211 ();
 sg13g2_fill_4 FILLER_41_225 ();
 sg13g2_fill_4 FILLER_41_286 ();
 sg13g2_fill_1 FILLER_41_290 ();
 sg13g2_fill_8 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_325 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_4 FILLER_41_361 ();
 sg13g2_fill_2 FILLER_41_373 ();
 sg13g2_fill_1 FILLER_41_375 ();
 sg13g2_fill_2 FILLER_41_386 ();
 sg13g2_fill_2 FILLER_41_394 ();
 sg13g2_fill_1 FILLER_41_396 ();
 sg13g2_fill_8 FILLER_41_404 ();
 sg13g2_fill_4 FILLER_41_412 ();
 sg13g2_fill_1 FILLER_41_416 ();
 sg13g2_fill_1 FILLER_41_433 ();
 sg13g2_fill_8 FILLER_41_450 ();
 sg13g2_fill_8 FILLER_41_458 ();
 sg13g2_fill_1 FILLER_41_466 ();
 sg13g2_fill_8 FILLER_41_475 ();
 sg13g2_fill_8 FILLER_41_483 ();
 sg13g2_fill_2 FILLER_41_491 ();
 sg13g2_fill_1 FILLER_41_493 ();
 sg13g2_fill_8 FILLER_41_538 ();
 sg13g2_fill_8 FILLER_41_546 ();
 sg13g2_fill_8 FILLER_41_554 ();
 sg13g2_fill_8 FILLER_41_562 ();
 sg13g2_fill_4 FILLER_41_570 ();
 sg13g2_fill_2 FILLER_41_574 ();
 sg13g2_fill_1 FILLER_41_576 ();
 sg13g2_fill_4 FILLER_41_603 ();
 sg13g2_fill_2 FILLER_41_607 ();
 sg13g2_fill_4 FILLER_41_620 ();
 sg13g2_fill_2 FILLER_41_624 ();
 sg13g2_fill_8 FILLER_41_630 ();
 sg13g2_fill_2 FILLER_41_638 ();
 sg13g2_fill_1 FILLER_41_640 ();
 sg13g2_fill_2 FILLER_41_648 ();
 sg13g2_fill_1 FILLER_41_650 ();
 sg13g2_fill_2 FILLER_41_661 ();
 sg13g2_fill_1 FILLER_41_671 ();
 sg13g2_fill_4 FILLER_41_691 ();
 sg13g2_fill_2 FILLER_41_695 ();
 sg13g2_fill_8 FILLER_41_701 ();
 sg13g2_fill_8 FILLER_41_709 ();
 sg13g2_fill_8 FILLER_41_723 ();
 sg13g2_fill_2 FILLER_41_750 ();
 sg13g2_fill_2 FILLER_41_783 ();
 sg13g2_fill_1 FILLER_41_805 ();
 sg13g2_fill_1 FILLER_41_814 ();
 sg13g2_fill_1 FILLER_41_833 ();
 sg13g2_fill_2 FILLER_41_850 ();
 sg13g2_fill_1 FILLER_41_852 ();
 sg13g2_fill_4 FILLER_41_889 ();
 sg13g2_fill_8 FILLER_41_902 ();
 sg13g2_fill_8 FILLER_41_910 ();
 sg13g2_fill_8 FILLER_41_918 ();
 sg13g2_fill_2 FILLER_41_926 ();
 sg13g2_fill_1 FILLER_41_928 ();
 sg13g2_fill_1 FILLER_41_949 ();
 sg13g2_fill_2 FILLER_41_956 ();
 sg13g2_fill_1 FILLER_41_964 ();
 sg13g2_fill_8 FILLER_41_975 ();
 sg13g2_fill_8 FILLER_41_983 ();
 sg13g2_fill_4 FILLER_41_991 ();
 sg13g2_fill_2 FILLER_41_995 ();
 sg13g2_fill_1 FILLER_41_997 ();
 sg13g2_fill_4 FILLER_41_1047 ();
 sg13g2_fill_2 FILLER_41_1051 ();
 sg13g2_fill_4 FILLER_41_1064 ();
 sg13g2_fill_2 FILLER_41_1068 ();
 sg13g2_fill_1 FILLER_41_1070 ();
 sg13g2_fill_8 FILLER_41_1076 ();
 sg13g2_fill_2 FILLER_41_1084 ();
 sg13g2_fill_2 FILLER_41_1090 ();
 sg13g2_fill_8 FILLER_41_1107 ();
 sg13g2_fill_2 FILLER_41_1115 ();
 sg13g2_fill_8 FILLER_41_1121 ();
 sg13g2_fill_8 FILLER_41_1129 ();
 sg13g2_fill_4 FILLER_41_1137 ();
 sg13g2_fill_2 FILLER_41_1141 ();
 sg13g2_fill_1 FILLER_41_1143 ();
 sg13g2_fill_1 FILLER_41_1150 ();
 sg13g2_fill_8 FILLER_41_1181 ();
 sg13g2_fill_8 FILLER_41_1189 ();
 sg13g2_fill_4 FILLER_41_1197 ();
 sg13g2_fill_2 FILLER_41_1201 ();
 sg13g2_fill_1 FILLER_41_1203 ();
 sg13g2_fill_1 FILLER_41_1215 ();
 sg13g2_fill_4 FILLER_41_1271 ();
 sg13g2_fill_2 FILLER_41_1275 ();
 sg13g2_fill_1 FILLER_41_1277 ();
 sg13g2_fill_2 FILLER_41_1320 ();
 sg13g2_fill_2 FILLER_41_1326 ();
 sg13g2_fill_1 FILLER_41_1328 ();
 sg13g2_fill_8 FILLER_41_1334 ();
 sg13g2_fill_4 FILLER_41_1342 ();
 sg13g2_fill_2 FILLER_41_1346 ();
 sg13g2_fill_1 FILLER_41_1348 ();
 sg13g2_fill_1 FILLER_41_1361 ();
 sg13g2_fill_8 FILLER_41_1366 ();
 sg13g2_fill_4 FILLER_41_1374 ();
 sg13g2_fill_2 FILLER_41_1378 ();
 sg13g2_fill_1 FILLER_41_1380 ();
 sg13g2_fill_1 FILLER_41_1401 ();
 sg13g2_fill_4 FILLER_41_1413 ();
 sg13g2_fill_2 FILLER_41_1417 ();
 sg13g2_fill_1 FILLER_41_1419 ();
 sg13g2_fill_4 FILLER_41_1442 ();
 sg13g2_fill_2 FILLER_41_1446 ();
 sg13g2_fill_1 FILLER_41_1448 ();
 sg13g2_fill_8 FILLER_41_1457 ();
 sg13g2_fill_8 FILLER_41_1465 ();
 sg13g2_fill_8 FILLER_41_1473 ();
 sg13g2_fill_4 FILLER_41_1481 ();
 sg13g2_fill_1 FILLER_41_1485 ();
 sg13g2_fill_8 FILLER_41_1526 ();
 sg13g2_fill_8 FILLER_41_1534 ();
 sg13g2_fill_8 FILLER_41_1542 ();
 sg13g2_fill_8 FILLER_41_1550 ();
 sg13g2_fill_8 FILLER_41_1558 ();
 sg13g2_fill_8 FILLER_41_1566 ();
 sg13g2_fill_8 FILLER_41_1574 ();
 sg13g2_fill_8 FILLER_41_1582 ();
 sg13g2_fill_2 FILLER_41_1590 ();
 sg13g2_fill_8 FILLER_42_0 ();
 sg13g2_fill_8 FILLER_42_8 ();
 sg13g2_fill_8 FILLER_42_16 ();
 sg13g2_fill_8 FILLER_42_24 ();
 sg13g2_fill_8 FILLER_42_32 ();
 sg13g2_fill_8 FILLER_42_40 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_8 FILLER_42_60 ();
 sg13g2_fill_8 FILLER_42_94 ();
 sg13g2_fill_4 FILLER_42_107 ();
 sg13g2_fill_2 FILLER_42_111 ();
 sg13g2_fill_2 FILLER_42_138 ();
 sg13g2_fill_4 FILLER_42_186 ();
 sg13g2_fill_2 FILLER_42_190 ();
 sg13g2_fill_1 FILLER_42_192 ();
 sg13g2_fill_4 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_8 FILLER_42_249 ();
 sg13g2_fill_8 FILLER_42_257 ();
 sg13g2_fill_2 FILLER_42_265 ();
 sg13g2_fill_8 FILLER_42_287 ();
 sg13g2_fill_8 FILLER_42_295 ();
 sg13g2_fill_2 FILLER_42_303 ();
 sg13g2_fill_1 FILLER_42_305 ();
 sg13g2_fill_1 FILLER_42_334 ();
 sg13g2_fill_2 FILLER_42_341 ();
 sg13g2_fill_1 FILLER_42_343 ();
 sg13g2_fill_4 FILLER_42_352 ();
 sg13g2_fill_8 FILLER_42_410 ();
 sg13g2_fill_8 FILLER_42_418 ();
 sg13g2_fill_4 FILLER_42_426 ();
 sg13g2_fill_1 FILLER_42_430 ();
 sg13g2_fill_1 FILLER_42_519 ();
 sg13g2_fill_4 FILLER_42_556 ();
 sg13g2_fill_1 FILLER_42_560 ();
 sg13g2_fill_2 FILLER_42_569 ();
 sg13g2_fill_2 FILLER_42_621 ();
 sg13g2_fill_1 FILLER_42_623 ();
 sg13g2_fill_4 FILLER_42_664 ();
 sg13g2_fill_2 FILLER_42_668 ();
 sg13g2_fill_1 FILLER_42_670 ();
 sg13g2_fill_1 FILLER_42_749 ();
 sg13g2_fill_8 FILLER_42_760 ();
 sg13g2_fill_8 FILLER_42_768 ();
 sg13g2_fill_8 FILLER_42_776 ();
 sg13g2_fill_2 FILLER_42_784 ();
 sg13g2_fill_4 FILLER_42_791 ();
 sg13g2_fill_1 FILLER_42_795 ();
 sg13g2_fill_8 FILLER_42_804 ();
 sg13g2_fill_8 FILLER_42_812 ();
 sg13g2_fill_2 FILLER_42_820 ();
 sg13g2_fill_1 FILLER_42_822 ();
 sg13g2_fill_2 FILLER_42_826 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_fill_1 FILLER_42_839 ();
 sg13g2_fill_8 FILLER_42_845 ();
 sg13g2_fill_2 FILLER_42_853 ();
 sg13g2_fill_1 FILLER_42_855 ();
 sg13g2_fill_4 FILLER_42_877 ();
 sg13g2_fill_2 FILLER_42_881 ();
 sg13g2_fill_1 FILLER_42_883 ();
 sg13g2_fill_2 FILLER_42_907 ();
 sg13g2_fill_4 FILLER_42_917 ();
 sg13g2_fill_8 FILLER_42_989 ();
 sg13g2_fill_8 FILLER_42_997 ();
 sg13g2_fill_8 FILLER_42_1005 ();
 sg13g2_fill_8 FILLER_42_1013 ();
 sg13g2_fill_4 FILLER_42_1021 ();
 sg13g2_fill_2 FILLER_42_1025 ();
 sg13g2_fill_8 FILLER_42_1057 ();
 sg13g2_fill_1 FILLER_42_1065 ();
 sg13g2_fill_2 FILLER_42_1081 ();
 sg13g2_fill_8 FILLER_42_1089 ();
 sg13g2_fill_1 FILLER_42_1101 ();
 sg13g2_fill_8 FILLER_42_1131 ();
 sg13g2_fill_8 FILLER_42_1139 ();
 sg13g2_fill_2 FILLER_42_1147 ();
 sg13g2_fill_8 FILLER_42_1161 ();
 sg13g2_fill_2 FILLER_42_1173 ();
 sg13g2_fill_1 FILLER_42_1175 ();
 sg13g2_fill_1 FILLER_42_1206 ();
 sg13g2_fill_8 FILLER_42_1229 ();
 sg13g2_fill_2 FILLER_42_1237 ();
 sg13g2_fill_4 FILLER_42_1249 ();
 sg13g2_fill_1 FILLER_42_1253 ();
 sg13g2_fill_4 FILLER_42_1284 ();
 sg13g2_fill_1 FILLER_42_1288 ();
 sg13g2_fill_4 FILLER_42_1323 ();
 sg13g2_fill_8 FILLER_42_1332 ();
 sg13g2_fill_2 FILLER_42_1340 ();
 sg13g2_fill_1 FILLER_42_1342 ();
 sg13g2_fill_4 FILLER_42_1351 ();
 sg13g2_fill_4 FILLER_42_1372 ();
 sg13g2_fill_8 FILLER_42_1380 ();
 sg13g2_fill_8 FILLER_42_1388 ();
 sg13g2_fill_8 FILLER_42_1396 ();
 sg13g2_fill_4 FILLER_42_1404 ();
 sg13g2_fill_2 FILLER_42_1408 ();
 sg13g2_fill_4 FILLER_42_1418 ();
 sg13g2_fill_1 FILLER_42_1422 ();
 sg13g2_fill_4 FILLER_42_1434 ();
 sg13g2_fill_8 FILLER_42_1460 ();
 sg13g2_fill_4 FILLER_42_1468 ();
 sg13g2_fill_2 FILLER_42_1472 ();
 sg13g2_fill_8 FILLER_42_1485 ();
 sg13g2_fill_8 FILLER_42_1493 ();
 sg13g2_fill_8 FILLER_42_1501 ();
 sg13g2_fill_8 FILLER_42_1509 ();
 sg13g2_fill_8 FILLER_42_1517 ();
 sg13g2_fill_8 FILLER_42_1525 ();
 sg13g2_fill_8 FILLER_42_1533 ();
 sg13g2_fill_1 FILLER_42_1541 ();
 sg13g2_fill_8 FILLER_42_1552 ();
 sg13g2_fill_2 FILLER_42_1560 ();
 sg13g2_fill_8 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_8 ();
 sg13g2_fill_1 FILLER_43_10 ();
 sg13g2_fill_2 FILLER_43_47 ();
 sg13g2_fill_4 FILLER_43_59 ();
 sg13g2_fill_2 FILLER_43_63 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_fill_8 FILLER_43_76 ();
 sg13g2_fill_4 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_98 ();
 sg13g2_fill_1 FILLER_43_100 ();
 sg13g2_fill_8 FILLER_43_159 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_fill_8 FILLER_43_209 ();
 sg13g2_fill_8 FILLER_43_217 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_fill_8 FILLER_43_262 ();
 sg13g2_fill_4 FILLER_43_270 ();
 sg13g2_fill_1 FILLER_43_274 ();
 sg13g2_fill_1 FILLER_43_285 ();
 sg13g2_fill_8 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_307 ();
 sg13g2_fill_1 FILLER_43_325 ();
 sg13g2_fill_8 FILLER_43_351 ();
 sg13g2_fill_8 FILLER_43_359 ();
 sg13g2_fill_8 FILLER_43_367 ();
 sg13g2_fill_4 FILLER_43_375 ();
 sg13g2_fill_1 FILLER_43_379 ();
 sg13g2_fill_8 FILLER_43_421 ();
 sg13g2_fill_8 FILLER_43_429 ();
 sg13g2_fill_2 FILLER_43_437 ();
 sg13g2_fill_1 FILLER_43_439 ();
 sg13g2_fill_8 FILLER_43_447 ();
 sg13g2_fill_2 FILLER_43_455 ();
 sg13g2_fill_1 FILLER_43_457 ();
 sg13g2_fill_4 FILLER_43_462 ();
 sg13g2_fill_4 FILLER_43_481 ();
 sg13g2_fill_2 FILLER_43_485 ();
 sg13g2_fill_1 FILLER_43_487 ();
 sg13g2_fill_8 FILLER_43_498 ();
 sg13g2_fill_4 FILLER_43_506 ();
 sg13g2_fill_1 FILLER_43_510 ();
 sg13g2_fill_1 FILLER_43_541 ();
 sg13g2_fill_4 FILLER_43_604 ();
 sg13g2_fill_2 FILLER_43_608 ();
 sg13g2_fill_1 FILLER_43_610 ();
 sg13g2_fill_1 FILLER_43_618 ();
 sg13g2_fill_4 FILLER_43_628 ();
 sg13g2_fill_1 FILLER_43_632 ();
 sg13g2_fill_8 FILLER_43_636 ();
 sg13g2_fill_1 FILLER_43_644 ();
 sg13g2_fill_8 FILLER_43_648 ();
 sg13g2_fill_1 FILLER_43_656 ();
 sg13g2_fill_8 FILLER_43_660 ();
 sg13g2_fill_4 FILLER_43_668 ();
 sg13g2_fill_2 FILLER_43_672 ();
 sg13g2_fill_1 FILLER_43_674 ();
 sg13g2_fill_8 FILLER_43_680 ();
 sg13g2_fill_4 FILLER_43_688 ();
 sg13g2_fill_2 FILLER_43_692 ();
 sg13g2_fill_1 FILLER_43_694 ();
 sg13g2_fill_8 FILLER_43_700 ();
 sg13g2_fill_8 FILLER_43_708 ();
 sg13g2_fill_8 FILLER_43_716 ();
 sg13g2_fill_1 FILLER_43_724 ();
 sg13g2_fill_4 FILLER_43_735 ();
 sg13g2_fill_2 FILLER_43_739 ();
 sg13g2_fill_1 FILLER_43_741 ();
 sg13g2_fill_8 FILLER_43_752 ();
 sg13g2_fill_8 FILLER_43_777 ();
 sg13g2_fill_2 FILLER_43_804 ();
 sg13g2_fill_1 FILLER_43_806 ();
 sg13g2_fill_2 FILLER_43_817 ();
 sg13g2_fill_1 FILLER_43_819 ();
 sg13g2_fill_4 FILLER_43_829 ();
 sg13g2_fill_1 FILLER_43_833 ();
 sg13g2_fill_1 FILLER_43_837 ();
 sg13g2_fill_8 FILLER_43_848 ();
 sg13g2_fill_2 FILLER_43_856 ();
 sg13g2_fill_1 FILLER_43_858 ();
 sg13g2_fill_8 FILLER_43_865 ();
 sg13g2_fill_1 FILLER_43_873 ();
 sg13g2_fill_4 FILLER_43_878 ();
 sg13g2_fill_2 FILLER_43_882 ();
 sg13g2_fill_2 FILLER_43_895 ();
 sg13g2_fill_1 FILLER_43_905 ();
 sg13g2_fill_1 FILLER_43_916 ();
 sg13g2_fill_4 FILLER_43_934 ();
 sg13g2_fill_1 FILLER_43_938 ();
 sg13g2_fill_1 FILLER_43_953 ();
 sg13g2_fill_2 FILLER_43_958 ();
 sg13g2_fill_1 FILLER_43_960 ();
 sg13g2_fill_1 FILLER_43_976 ();
 sg13g2_fill_8 FILLER_43_1003 ();
 sg13g2_fill_8 FILLER_43_1011 ();
 sg13g2_fill_4 FILLER_43_1019 ();
 sg13g2_fill_1 FILLER_43_1023 ();
 sg13g2_fill_1 FILLER_43_1034 ();
 sg13g2_fill_4 FILLER_43_1066 ();
 sg13g2_fill_4 FILLER_43_1099 ();
 sg13g2_fill_8 FILLER_43_1205 ();
 sg13g2_fill_2 FILLER_43_1213 ();
 sg13g2_fill_1 FILLER_43_1215 ();
 sg13g2_fill_8 FILLER_43_1230 ();
 sg13g2_fill_4 FILLER_43_1238 ();
 sg13g2_fill_1 FILLER_43_1248 ();
 sg13g2_fill_4 FILLER_43_1294 ();
 sg13g2_fill_1 FILLER_43_1298 ();
 sg13g2_fill_4 FILLER_43_1311 ();
 sg13g2_fill_2 FILLER_43_1315 ();
 sg13g2_fill_1 FILLER_43_1317 ();
 sg13g2_fill_2 FILLER_43_1333 ();
 sg13g2_fill_1 FILLER_43_1343 ();
 sg13g2_fill_2 FILLER_43_1353 ();
 sg13g2_fill_1 FILLER_43_1355 ();
 sg13g2_fill_2 FILLER_43_1360 ();
 sg13g2_fill_1 FILLER_43_1362 ();
 sg13g2_fill_2 FILLER_43_1384 ();
 sg13g2_fill_1 FILLER_43_1386 ();
 sg13g2_fill_1 FILLER_43_1395 ();
 sg13g2_fill_8 FILLER_43_1400 ();
 sg13g2_fill_8 FILLER_43_1449 ();
 sg13g2_fill_4 FILLER_43_1457 ();
 sg13g2_fill_2 FILLER_43_1461 ();
 sg13g2_fill_1 FILLER_43_1463 ();
 sg13g2_fill_2 FILLER_43_1483 ();
 sg13g2_fill_1 FILLER_43_1485 ();
 sg13g2_fill_4 FILLER_43_1497 ();
 sg13g2_fill_2 FILLER_43_1501 ();
 sg13g2_fill_1 FILLER_43_1503 ();
 sg13g2_fill_8 FILLER_43_1544 ();
 sg13g2_fill_8 FILLER_43_1582 ();
 sg13g2_fill_2 FILLER_43_1590 ();
 sg13g2_fill_8 FILLER_44_0 ();
 sg13g2_fill_8 FILLER_44_8 ();
 sg13g2_fill_4 FILLER_44_16 ();
 sg13g2_fill_2 FILLER_44_46 ();
 sg13g2_fill_4 FILLER_44_58 ();
 sg13g2_fill_1 FILLER_44_62 ();
 sg13g2_fill_1 FILLER_44_89 ();
 sg13g2_fill_8 FILLER_44_126 ();
 sg13g2_fill_8 FILLER_44_134 ();
 sg13g2_fill_4 FILLER_44_142 ();
 sg13g2_fill_2 FILLER_44_146 ();
 sg13g2_fill_8 FILLER_44_154 ();
 sg13g2_fill_4 FILLER_44_162 ();
 sg13g2_fill_8 FILLER_44_205 ();
 sg13g2_fill_8 FILLER_44_213 ();
 sg13g2_fill_1 FILLER_44_221 ();
 sg13g2_fill_4 FILLER_44_232 ();
 sg13g2_fill_2 FILLER_44_236 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_8 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_273 ();
 sg13g2_fill_1 FILLER_44_275 ();
 sg13g2_fill_2 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_313 ();
 sg13g2_fill_1 FILLER_44_315 ();
 sg13g2_fill_8 FILLER_44_361 ();
 sg13g2_fill_2 FILLER_44_379 ();
 sg13g2_fill_1 FILLER_44_402 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_fill_4 FILLER_44_435 ();
 sg13g2_fill_2 FILLER_44_439 ();
 sg13g2_fill_1 FILLER_44_441 ();
 sg13g2_fill_2 FILLER_44_483 ();
 sg13g2_fill_8 FILLER_44_506 ();
 sg13g2_fill_4 FILLER_44_514 ();
 sg13g2_fill_1 FILLER_44_518 ();
 sg13g2_fill_4 FILLER_44_532 ();
 sg13g2_fill_8 FILLER_44_546 ();
 sg13g2_fill_8 FILLER_44_554 ();
 sg13g2_fill_2 FILLER_44_562 ();
 sg13g2_fill_8 FILLER_44_569 ();
 sg13g2_fill_8 FILLER_44_577 ();
 sg13g2_fill_8 FILLER_44_585 ();
 sg13g2_fill_8 FILLER_44_593 ();
 sg13g2_fill_4 FILLER_44_601 ();
 sg13g2_fill_1 FILLER_44_605 ();
 sg13g2_fill_2 FILLER_44_707 ();
 sg13g2_fill_1 FILLER_44_709 ();
 sg13g2_fill_4 FILLER_44_743 ();
 sg13g2_fill_2 FILLER_44_747 ();
 sg13g2_fill_1 FILLER_44_818 ();
 sg13g2_fill_2 FILLER_44_836 ();
 sg13g2_fill_1 FILLER_44_838 ();
 sg13g2_fill_2 FILLER_44_860 ();
 sg13g2_fill_1 FILLER_44_862 ();
 sg13g2_fill_4 FILLER_44_868 ();
 sg13g2_fill_1 FILLER_44_872 ();
 sg13g2_fill_2 FILLER_44_882 ();
 sg13g2_fill_1 FILLER_44_884 ();
 sg13g2_fill_1 FILLER_44_913 ();
 sg13g2_fill_8 FILLER_44_922 ();
 sg13g2_fill_8 FILLER_44_930 ();
 sg13g2_fill_4 FILLER_44_938 ();
 sg13g2_fill_2 FILLER_44_942 ();
 sg13g2_fill_2 FILLER_44_980 ();
 sg13g2_fill_8 FILLER_44_1082 ();
 sg13g2_fill_4 FILLER_44_1090 ();
 sg13g2_fill_2 FILLER_44_1094 ();
 sg13g2_fill_4 FILLER_44_1102 ();
 sg13g2_fill_4 FILLER_44_1119 ();
 sg13g2_fill_2 FILLER_44_1123 ();
 sg13g2_fill_4 FILLER_44_1134 ();
 sg13g2_fill_8 FILLER_44_1142 ();
 sg13g2_fill_8 FILLER_44_1150 ();
 sg13g2_fill_4 FILLER_44_1158 ();
 sg13g2_fill_2 FILLER_44_1162 ();
 sg13g2_fill_2 FILLER_44_1182 ();
 sg13g2_fill_1 FILLER_44_1184 ();
 sg13g2_fill_4 FILLER_44_1245 ();
 sg13g2_fill_2 FILLER_44_1284 ();
 sg13g2_fill_8 FILLER_44_1322 ();
 sg13g2_fill_4 FILLER_44_1330 ();
 sg13g2_fill_2 FILLER_44_1334 ();
 sg13g2_fill_1 FILLER_44_1336 ();
 sg13g2_fill_4 FILLER_44_1350 ();
 sg13g2_fill_2 FILLER_44_1354 ();
 sg13g2_fill_1 FILLER_44_1356 ();
 sg13g2_fill_4 FILLER_44_1360 ();
 sg13g2_fill_2 FILLER_44_1364 ();
 sg13g2_fill_1 FILLER_44_1366 ();
 sg13g2_fill_8 FILLER_44_1371 ();
 sg13g2_fill_8 FILLER_44_1379 ();
 sg13g2_fill_4 FILLER_44_1387 ();
 sg13g2_fill_2 FILLER_44_1391 ();
 sg13g2_fill_1 FILLER_44_1404 ();
 sg13g2_fill_8 FILLER_44_1422 ();
 sg13g2_fill_8 FILLER_44_1430 ();
 sg13g2_fill_1 FILLER_44_1438 ();
 sg13g2_fill_4 FILLER_44_1479 ();
 sg13g2_fill_2 FILLER_44_1483 ();
 sg13g2_fill_8 FILLER_44_1496 ();
 sg13g2_fill_8 FILLER_44_1504 ();
 sg13g2_fill_8 FILLER_44_1512 ();
 sg13g2_fill_2 FILLER_44_1520 ();
 sg13g2_fill_2 FILLER_44_1547 ();
 sg13g2_fill_8 FILLER_44_1559 ();
 sg13g2_fill_8 FILLER_45_0 ();
 sg13g2_fill_8 FILLER_45_8 ();
 sg13g2_fill_8 FILLER_45_16 ();
 sg13g2_fill_8 FILLER_45_24 ();
 sg13g2_fill_4 FILLER_45_32 ();
 sg13g2_fill_8 FILLER_45_46 ();
 sg13g2_fill_4 FILLER_45_54 ();
 sg13g2_fill_1 FILLER_45_58 ();
 sg13g2_fill_8 FILLER_45_79 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_fill_8 FILLER_45_127 ();
 sg13g2_fill_8 FILLER_45_135 ();
 sg13g2_fill_1 FILLER_45_143 ();
 sg13g2_fill_4 FILLER_45_164 ();
 sg13g2_fill_1 FILLER_45_168 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_8 FILLER_45_243 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_4 FILLER_45_280 ();
 sg13g2_fill_4 FILLER_45_289 ();
 sg13g2_fill_1 FILLER_45_314 ();
 sg13g2_fill_4 FILLER_45_368 ();
 sg13g2_fill_2 FILLER_45_385 ();
 sg13g2_fill_1 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_414 ();
 sg13g2_fill_2 FILLER_45_452 ();
 sg13g2_fill_4 FILLER_45_515 ();
 sg13g2_fill_2 FILLER_45_544 ();
 sg13g2_fill_8 FILLER_45_582 ();
 sg13g2_fill_8 FILLER_45_590 ();
 sg13g2_fill_8 FILLER_45_598 ();
 sg13g2_fill_2 FILLER_45_606 ();
 sg13g2_fill_4 FILLER_45_618 ();
 sg13g2_fill_1 FILLER_45_622 ();
 sg13g2_fill_4 FILLER_45_632 ();
 sg13g2_fill_1 FILLER_45_673 ();
 sg13g2_fill_1 FILLER_45_689 ();
 sg13g2_fill_8 FILLER_45_694 ();
 sg13g2_fill_8 FILLER_45_718 ();
 sg13g2_fill_1 FILLER_45_726 ();
 sg13g2_fill_1 FILLER_45_761 ();
 sg13g2_fill_2 FILLER_45_801 ();
 sg13g2_fill_1 FILLER_45_803 ();
 sg13g2_fill_2 FILLER_45_810 ();
 sg13g2_fill_2 FILLER_45_817 ();
 sg13g2_fill_1 FILLER_45_819 ();
 sg13g2_fill_2 FILLER_45_838 ();
 sg13g2_fill_8 FILLER_45_844 ();
 sg13g2_fill_1 FILLER_45_852 ();
 sg13g2_fill_4 FILLER_45_863 ();
 sg13g2_fill_8 FILLER_45_906 ();
 sg13g2_fill_1 FILLER_45_914 ();
 sg13g2_fill_4 FILLER_45_931 ();
 sg13g2_fill_4 FILLER_45_938 ();
 sg13g2_fill_2 FILLER_45_942 ();
 sg13g2_fill_8 FILLER_45_947 ();
 sg13g2_fill_8 FILLER_45_955 ();
 sg13g2_fill_8 FILLER_45_963 ();
 sg13g2_fill_8 FILLER_45_971 ();
 sg13g2_fill_4 FILLER_45_979 ();
 sg13g2_fill_1 FILLER_45_983 ();
 sg13g2_fill_8 FILLER_45_997 ();
 sg13g2_fill_1 FILLER_45_1005 ();
 sg13g2_fill_8 FILLER_45_1011 ();
 sg13g2_fill_8 FILLER_45_1019 ();
 sg13g2_fill_4 FILLER_45_1027 ();
 sg13g2_fill_2 FILLER_45_1031 ();
 sg13g2_fill_1 FILLER_45_1033 ();
 sg13g2_fill_2 FILLER_45_1046 ();
 sg13g2_fill_8 FILLER_45_1076 ();
 sg13g2_fill_2 FILLER_45_1084 ();
 sg13g2_fill_4 FILLER_45_1120 ();
 sg13g2_fill_2 FILLER_45_1124 ();
 sg13g2_fill_2 FILLER_45_1136 ();
 sg13g2_fill_8 FILLER_45_1144 ();
 sg13g2_fill_8 FILLER_45_1152 ();
 sg13g2_fill_8 FILLER_45_1160 ();
 sg13g2_fill_2 FILLER_45_1178 ();
 sg13g2_fill_8 FILLER_45_1210 ();
 sg13g2_fill_2 FILLER_45_1218 ();
 sg13g2_fill_4 FILLER_45_1229 ();
 sg13g2_fill_2 FILLER_45_1273 ();
 sg13g2_fill_1 FILLER_45_1275 ();
 sg13g2_fill_4 FILLER_45_1289 ();
 sg13g2_fill_2 FILLER_45_1293 ();
 sg13g2_fill_4 FILLER_45_1301 ();
 sg13g2_fill_1 FILLER_45_1305 ();
 sg13g2_fill_8 FILLER_45_1315 ();
 sg13g2_fill_1 FILLER_45_1350 ();
 sg13g2_fill_2 FILLER_45_1358 ();
 sg13g2_fill_4 FILLER_45_1372 ();
 sg13g2_fill_1 FILLER_45_1376 ();
 sg13g2_fill_4 FILLER_45_1393 ();
 sg13g2_fill_1 FILLER_45_1397 ();
 sg13g2_fill_8 FILLER_45_1409 ();
 sg13g2_fill_8 FILLER_45_1417 ();
 sg13g2_fill_8 FILLER_45_1468 ();
 sg13g2_fill_8 FILLER_45_1476 ();
 sg13g2_fill_2 FILLER_45_1484 ();
 sg13g2_fill_1 FILLER_45_1486 ();
 sg13g2_fill_2 FILLER_45_1498 ();
 sg13g2_fill_8 FILLER_45_1543 ();
 sg13g2_fill_1 FILLER_45_1551 ();
 sg13g2_fill_8 FILLER_46_0 ();
 sg13g2_fill_8 FILLER_46_8 ();
 sg13g2_fill_8 FILLER_46_16 ();
 sg13g2_fill_8 FILLER_46_24 ();
 sg13g2_fill_2 FILLER_46_32 ();
 sg13g2_fill_8 FILLER_46_44 ();
 sg13g2_fill_8 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_60 ();
 sg13g2_fill_4 FILLER_46_87 ();
 sg13g2_fill_2 FILLER_46_91 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_8 FILLER_46_160 ();
 sg13g2_fill_8 FILLER_46_168 ();
 sg13g2_fill_8 FILLER_46_176 ();
 sg13g2_fill_4 FILLER_46_184 ();
 sg13g2_fill_2 FILLER_46_188 ();
 sg13g2_fill_1 FILLER_46_190 ();
 sg13g2_fill_8 FILLER_46_196 ();
 sg13g2_fill_8 FILLER_46_240 ();
 sg13g2_fill_4 FILLER_46_248 ();
 sg13g2_fill_8 FILLER_46_262 ();
 sg13g2_fill_8 FILLER_46_270 ();
 sg13g2_fill_8 FILLER_46_278 ();
 sg13g2_fill_8 FILLER_46_286 ();
 sg13g2_fill_8 FILLER_46_294 ();
 sg13g2_fill_8 FILLER_46_302 ();
 sg13g2_fill_8 FILLER_46_335 ();
 sg13g2_fill_8 FILLER_46_343 ();
 sg13g2_fill_4 FILLER_46_351 ();
 sg13g2_fill_1 FILLER_46_355 ();
 sg13g2_fill_8 FILLER_46_362 ();
 sg13g2_fill_1 FILLER_46_370 ();
 sg13g2_fill_8 FILLER_46_381 ();
 sg13g2_fill_8 FILLER_46_389 ();
 sg13g2_fill_8 FILLER_46_397 ();
 sg13g2_fill_4 FILLER_46_405 ();
 sg13g2_fill_2 FILLER_46_409 ();
 sg13g2_fill_8 FILLER_46_434 ();
 sg13g2_fill_8 FILLER_46_442 ();
 sg13g2_fill_8 FILLER_46_450 ();
 sg13g2_fill_8 FILLER_46_458 ();
 sg13g2_fill_8 FILLER_46_466 ();
 sg13g2_fill_2 FILLER_46_474 ();
 sg13g2_fill_8 FILLER_46_486 ();
 sg13g2_fill_4 FILLER_46_494 ();
 sg13g2_fill_2 FILLER_46_498 ();
 sg13g2_fill_2 FILLER_46_526 ();
 sg13g2_fill_4 FILLER_46_534 ();
 sg13g2_fill_2 FILLER_46_538 ();
 sg13g2_fill_4 FILLER_46_565 ();
 sg13g2_fill_1 FILLER_46_569 ();
 sg13g2_fill_4 FILLER_46_578 ();
 sg13g2_fill_2 FILLER_46_612 ();
 sg13g2_fill_1 FILLER_46_614 ();
 sg13g2_fill_8 FILLER_46_672 ();
 sg13g2_fill_8 FILLER_46_680 ();
 sg13g2_fill_2 FILLER_46_688 ();
 sg13g2_fill_8 FILLER_46_695 ();
 sg13g2_fill_2 FILLER_46_703 ();
 sg13g2_fill_1 FILLER_46_705 ();
 sg13g2_fill_1 FILLER_46_716 ();
 sg13g2_fill_8 FILLER_46_722 ();
 sg13g2_fill_8 FILLER_46_730 ();
 sg13g2_fill_8 FILLER_46_738 ();
 sg13g2_fill_4 FILLER_46_746 ();
 sg13g2_fill_2 FILLER_46_750 ();
 sg13g2_fill_1 FILLER_46_752 ();
 sg13g2_fill_1 FILLER_46_758 ();
 sg13g2_fill_2 FILLER_46_774 ();
 sg13g2_fill_1 FILLER_46_801 ();
 sg13g2_fill_8 FILLER_46_810 ();
 sg13g2_fill_4 FILLER_46_818 ();
 sg13g2_fill_2 FILLER_46_822 ();
 sg13g2_fill_1 FILLER_46_824 ();
 sg13g2_fill_8 FILLER_46_828 ();
 sg13g2_fill_8 FILLER_46_836 ();
 sg13g2_fill_4 FILLER_46_844 ();
 sg13g2_fill_1 FILLER_46_848 ();
 sg13g2_fill_4 FILLER_46_854 ();
 sg13g2_fill_4 FILLER_46_866 ();
 sg13g2_fill_2 FILLER_46_870 ();
 sg13g2_fill_1 FILLER_46_872 ();
 sg13g2_fill_2 FILLER_46_878 ();
 sg13g2_fill_2 FILLER_46_896 ();
 sg13g2_fill_4 FILLER_46_916 ();
 sg13g2_fill_2 FILLER_46_973 ();
 sg13g2_fill_1 FILLER_46_975 ();
 sg13g2_fill_8 FILLER_46_980 ();
 sg13g2_fill_8 FILLER_46_988 ();
 sg13g2_fill_8 FILLER_46_996 ();
 sg13g2_fill_4 FILLER_46_1004 ();
 sg13g2_fill_8 FILLER_46_1034 ();
 sg13g2_fill_2 FILLER_46_1059 ();
 sg13g2_fill_1 FILLER_46_1064 ();
 sg13g2_fill_8 FILLER_46_1099 ();
 sg13g2_fill_4 FILLER_46_1107 ();
 sg13g2_fill_2 FILLER_46_1111 ();
 sg13g2_fill_1 FILLER_46_1113 ();
 sg13g2_fill_1 FILLER_46_1132 ();
 sg13g2_fill_4 FILLER_46_1163 ();
 sg13g2_fill_4 FILLER_46_1207 ();
 sg13g2_fill_2 FILLER_46_1221 ();
 sg13g2_fill_1 FILLER_46_1223 ();
 sg13g2_fill_4 FILLER_46_1232 ();
 sg13g2_fill_1 FILLER_46_1236 ();
 sg13g2_fill_1 FILLER_46_1243 ();
 sg13g2_fill_4 FILLER_46_1250 ();
 sg13g2_fill_2 FILLER_46_1254 ();
 sg13g2_fill_1 FILLER_46_1256 ();
 sg13g2_fill_8 FILLER_46_1298 ();
 sg13g2_fill_4 FILLER_46_1306 ();
 sg13g2_fill_1 FILLER_46_1310 ();
 sg13g2_fill_2 FILLER_46_1316 ();
 sg13g2_fill_1 FILLER_46_1331 ();
 sg13g2_fill_1 FILLER_46_1352 ();
 sg13g2_fill_2 FILLER_46_1367 ();
 sg13g2_fill_1 FILLER_46_1369 ();
 sg13g2_fill_1 FILLER_46_1392 ();
 sg13g2_fill_4 FILLER_46_1445 ();
 sg13g2_fill_2 FILLER_46_1479 ();
 sg13g2_fill_1 FILLER_46_1481 ();
 sg13g2_fill_1 FILLER_46_1493 ();
 sg13g2_fill_8 FILLER_46_1504 ();
 sg13g2_fill_8 FILLER_46_1512 ();
 sg13g2_fill_8 FILLER_46_1560 ();
 sg13g2_fill_4 FILLER_46_1568 ();
 sg13g2_fill_2 FILLER_46_1572 ();
 sg13g2_fill_8 FILLER_46_1580 ();
 sg13g2_fill_4 FILLER_46_1588 ();
 sg13g2_fill_8 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_8 ();
 sg13g2_fill_1 FILLER_47_10 ();
 sg13g2_fill_8 FILLER_47_115 ();
 sg13g2_fill_1 FILLER_47_123 ();
 sg13g2_fill_8 FILLER_47_130 ();
 sg13g2_fill_2 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_140 ();
 sg13g2_fill_4 FILLER_47_177 ();
 sg13g2_fill_8 FILLER_47_186 ();
 sg13g2_fill_8 FILLER_47_194 ();
 sg13g2_fill_8 FILLER_47_202 ();
 sg13g2_fill_8 FILLER_47_210 ();
 sg13g2_fill_8 FILLER_47_218 ();
 sg13g2_fill_8 FILLER_47_226 ();
 sg13g2_fill_8 FILLER_47_234 ();
 sg13g2_fill_8 FILLER_47_242 ();
 sg13g2_fill_8 FILLER_47_258 ();
 sg13g2_fill_4 FILLER_47_266 ();
 sg13g2_fill_2 FILLER_47_270 ();
 sg13g2_fill_8 FILLER_47_297 ();
 sg13g2_fill_4 FILLER_47_305 ();
 sg13g2_fill_1 FILLER_47_309 ();
 sg13g2_fill_2 FILLER_47_381 ();
 sg13g2_fill_1 FILLER_47_383 ();
 sg13g2_fill_4 FILLER_47_397 ();
 sg13g2_fill_2 FILLER_47_401 ();
 sg13g2_fill_8 FILLER_47_416 ();
 sg13g2_fill_8 FILLER_47_454 ();
 sg13g2_fill_8 FILLER_47_462 ();
 sg13g2_fill_4 FILLER_47_470 ();
 sg13g2_fill_4 FILLER_47_484 ();
 sg13g2_fill_2 FILLER_47_488 ();
 sg13g2_fill_1 FILLER_47_490 ();
 sg13g2_fill_1 FILLER_47_527 ();
 sg13g2_fill_8 FILLER_47_544 ();
 sg13g2_fill_8 FILLER_47_552 ();
 sg13g2_fill_8 FILLER_47_560 ();
 sg13g2_fill_8 FILLER_47_568 ();
 sg13g2_fill_8 FILLER_47_576 ();
 sg13g2_fill_2 FILLER_47_584 ();
 sg13g2_fill_4 FILLER_47_612 ();
 sg13g2_fill_1 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_625 ();
 sg13g2_fill_8 FILLER_47_664 ();
 sg13g2_fill_4 FILLER_47_672 ();
 sg13g2_fill_4 FILLER_47_683 ();
 sg13g2_fill_2 FILLER_47_687 ();
 sg13g2_fill_8 FILLER_47_695 ();
 sg13g2_fill_4 FILLER_47_703 ();
 sg13g2_fill_1 FILLER_47_707 ();
 sg13g2_fill_8 FILLER_47_742 ();
 sg13g2_fill_2 FILLER_47_750 ();
 sg13g2_fill_4 FILLER_47_804 ();
 sg13g2_fill_2 FILLER_47_808 ();
 sg13g2_fill_4 FILLER_47_814 ();
 sg13g2_fill_2 FILLER_47_818 ();
 sg13g2_fill_1 FILLER_47_820 ();
 sg13g2_fill_1 FILLER_47_844 ();
 sg13g2_fill_8 FILLER_47_856 ();
 sg13g2_fill_8 FILLER_47_869 ();
 sg13g2_fill_4 FILLER_47_877 ();
 sg13g2_fill_1 FILLER_47_881 ();
 sg13g2_fill_4 FILLER_47_893 ();
 sg13g2_fill_1 FILLER_47_897 ();
 sg13g2_fill_2 FILLER_47_910 ();
 sg13g2_fill_2 FILLER_47_945 ();
 sg13g2_fill_4 FILLER_47_987 ();
 sg13g2_fill_2 FILLER_47_991 ();
 sg13g2_fill_1 FILLER_47_993 ();
 sg13g2_fill_4 FILLER_47_1015 ();
 sg13g2_fill_1 FILLER_47_1067 ();
 sg13g2_fill_1 FILLER_47_1078 ();
 sg13g2_fill_4 FILLER_47_1085 ();
 sg13g2_fill_2 FILLER_47_1089 ();
 sg13g2_fill_1 FILLER_47_1091 ();
 sg13g2_fill_2 FILLER_47_1128 ();
 sg13g2_fill_1 FILLER_47_1130 ();
 sg13g2_fill_2 FILLER_47_1169 ();
 sg13g2_fill_8 FILLER_47_1179 ();
 sg13g2_fill_8 FILLER_47_1187 ();
 sg13g2_fill_8 FILLER_47_1195 ();
 sg13g2_fill_1 FILLER_47_1203 ();
 sg13g2_fill_2 FILLER_47_1235 ();
 sg13g2_fill_1 FILLER_47_1237 ();
 sg13g2_fill_1 FILLER_47_1286 ();
 sg13g2_fill_1 FILLER_47_1313 ();
 sg13g2_fill_1 FILLER_47_1328 ();
 sg13g2_fill_2 FILLER_47_1346 ();
 sg13g2_fill_1 FILLER_47_1363 ();
 sg13g2_fill_2 FILLER_47_1372 ();
 sg13g2_fill_4 FILLER_47_1390 ();
 sg13g2_fill_2 FILLER_47_1394 ();
 sg13g2_fill_8 FILLER_47_1407 ();
 sg13g2_fill_8 FILLER_47_1415 ();
 sg13g2_fill_4 FILLER_47_1423 ();
 sg13g2_fill_1 FILLER_47_1427 ();
 sg13g2_fill_8 FILLER_47_1439 ();
 sg13g2_fill_2 FILLER_47_1447 ();
 sg13g2_fill_8 FILLER_47_1460 ();
 sg13g2_fill_4 FILLER_47_1490 ();
 sg13g2_fill_1 FILLER_47_1494 ();
 sg13g2_fill_2 FILLER_47_1520 ();
 sg13g2_fill_1 FILLER_47_1522 ();
 sg13g2_fill_2 FILLER_47_1548 ();
 sg13g2_fill_1 FILLER_47_1550 ();
 sg13g2_fill_1 FILLER_47_1561 ();
 sg13g2_fill_8 FILLER_48_0 ();
 sg13g2_fill_8 FILLER_48_8 ();
 sg13g2_fill_8 FILLER_48_16 ();
 sg13g2_fill_1 FILLER_48_24 ();
 sg13g2_fill_4 FILLER_48_71 ();
 sg13g2_fill_1 FILLER_48_75 ();
 sg13g2_fill_8 FILLER_48_86 ();
 sg13g2_fill_8 FILLER_48_94 ();
 sg13g2_fill_8 FILLER_48_102 ();
 sg13g2_fill_8 FILLER_48_110 ();
 sg13g2_fill_8 FILLER_48_118 ();
 sg13g2_fill_8 FILLER_48_126 ();
 sg13g2_fill_8 FILLER_48_134 ();
 sg13g2_fill_8 FILLER_48_142 ();
 sg13g2_fill_8 FILLER_48_150 ();
 sg13g2_fill_8 FILLER_48_158 ();
 sg13g2_fill_8 FILLER_48_166 ();
 sg13g2_fill_8 FILLER_48_174 ();
 sg13g2_fill_8 FILLER_48_182 ();
 sg13g2_fill_8 FILLER_48_190 ();
 sg13g2_fill_8 FILLER_48_198 ();
 sg13g2_fill_8 FILLER_48_206 ();
 sg13g2_fill_8 FILLER_48_214 ();
 sg13g2_fill_1 FILLER_48_222 ();
 sg13g2_fill_2 FILLER_48_228 ();
 sg13g2_fill_4 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_338 ();
 sg13g2_fill_2 FILLER_48_342 ();
 sg13g2_fill_1 FILLER_48_344 ();
 sg13g2_fill_1 FILLER_48_381 ();
 sg13g2_fill_4 FILLER_48_403 ();
 sg13g2_fill_8 FILLER_48_420 ();
 sg13g2_fill_8 FILLER_48_428 ();
 sg13g2_fill_1 FILLER_48_436 ();
 sg13g2_fill_8 FILLER_48_481 ();
 sg13g2_fill_4 FILLER_48_489 ();
 sg13g2_fill_8 FILLER_48_503 ();
 sg13g2_fill_8 FILLER_48_511 ();
 sg13g2_fill_4 FILLER_48_519 ();
 sg13g2_fill_2 FILLER_48_523 ();
 sg13g2_fill_2 FILLER_48_535 ();
 sg13g2_fill_1 FILLER_48_537 ();
 sg13g2_fill_8 FILLER_48_582 ();
 sg13g2_fill_8 FILLER_48_590 ();
 sg13g2_fill_8 FILLER_48_598 ();
 sg13g2_fill_1 FILLER_48_606 ();
 sg13g2_fill_2 FILLER_48_623 ();
 sg13g2_fill_2 FILLER_48_636 ();
 sg13g2_fill_1 FILLER_48_638 ();
 sg13g2_fill_2 FILLER_48_675 ();
 sg13g2_fill_4 FILLER_48_682 ();
 sg13g2_fill_1 FILLER_48_686 ();
 sg13g2_fill_2 FILLER_48_714 ();
 sg13g2_fill_4 FILLER_48_722 ();
 sg13g2_fill_2 FILLER_48_726 ();
 sg13g2_fill_1 FILLER_48_728 ();
 sg13g2_fill_8 FILLER_48_755 ();
 sg13g2_fill_8 FILLER_48_763 ();
 sg13g2_fill_8 FILLER_48_774 ();
 sg13g2_fill_8 FILLER_48_782 ();
 sg13g2_fill_2 FILLER_48_790 ();
 sg13g2_fill_8 FILLER_48_798 ();
 sg13g2_fill_2 FILLER_48_811 ();
 sg13g2_fill_2 FILLER_48_833 ();
 sg13g2_fill_1 FILLER_48_841 ();
 sg13g2_fill_2 FILLER_48_846 ();
 sg13g2_fill_1 FILLER_48_856 ();
 sg13g2_fill_2 FILLER_48_878 ();
 sg13g2_fill_1 FILLER_48_880 ();
 sg13g2_fill_2 FILLER_48_886 ();
 sg13g2_fill_1 FILLER_48_888 ();
 sg13g2_fill_1 FILLER_48_913 ();
 sg13g2_fill_1 FILLER_48_946 ();
 sg13g2_fill_1 FILLER_48_968 ();
 sg13g2_fill_4 FILLER_48_1005 ();
 sg13g2_fill_2 FILLER_48_1009 ();
 sg13g2_fill_2 FILLER_48_1036 ();
 sg13g2_fill_1 FILLER_48_1038 ();
 sg13g2_fill_4 FILLER_48_1045 ();
 sg13g2_fill_2 FILLER_48_1049 ();
 sg13g2_fill_1 FILLER_48_1051 ();
 sg13g2_fill_8 FILLER_48_1072 ();
 sg13g2_fill_4 FILLER_48_1080 ();
 sg13g2_fill_8 FILLER_48_1088 ();
 sg13g2_fill_8 FILLER_48_1096 ();
 sg13g2_fill_4 FILLER_48_1104 ();
 sg13g2_fill_2 FILLER_48_1108 ();
 sg13g2_fill_8 FILLER_48_1141 ();
 sg13g2_fill_4 FILLER_48_1149 ();
 sg13g2_fill_1 FILLER_48_1153 ();
 sg13g2_fill_8 FILLER_48_1157 ();
 sg13g2_fill_8 FILLER_48_1165 ();
 sg13g2_fill_8 FILLER_48_1173 ();
 sg13g2_fill_8 FILLER_48_1181 ();
 sg13g2_fill_8 FILLER_48_1189 ();
 sg13g2_fill_8 FILLER_48_1197 ();
 sg13g2_fill_8 FILLER_48_1205 ();
 sg13g2_fill_8 FILLER_48_1213 ();
 sg13g2_fill_1 FILLER_48_1221 ();
 sg13g2_fill_8 FILLER_48_1228 ();
 sg13g2_fill_2 FILLER_48_1236 ();
 sg13g2_fill_4 FILLER_48_1244 ();
 sg13g2_fill_1 FILLER_48_1248 ();
 sg13g2_fill_8 FILLER_48_1255 ();
 sg13g2_fill_8 FILLER_48_1263 ();
 sg13g2_fill_4 FILLER_48_1271 ();
 sg13g2_fill_1 FILLER_48_1275 ();
 sg13g2_fill_1 FILLER_48_1320 ();
 sg13g2_fill_2 FILLER_48_1337 ();
 sg13g2_fill_1 FILLER_48_1358 ();
 sg13g2_fill_8 FILLER_48_1379 ();
 sg13g2_fill_2 FILLER_48_1387 ();
 sg13g2_fill_1 FILLER_48_1389 ();
 sg13g2_fill_4 FILLER_48_1394 ();
 sg13g2_fill_8 FILLER_48_1403 ();
 sg13g2_fill_8 FILLER_48_1411 ();
 sg13g2_fill_8 FILLER_48_1419 ();
 sg13g2_fill_2 FILLER_48_1427 ();
 sg13g2_fill_1 FILLER_48_1429 ();
 sg13g2_fill_2 FILLER_48_1441 ();
 sg13g2_fill_1 FILLER_48_1443 ();
 sg13g2_fill_2 FILLER_48_1454 ();
 sg13g2_fill_1 FILLER_48_1456 ();
 sg13g2_fill_8 FILLER_48_1462 ();
 sg13g2_fill_8 FILLER_48_1470 ();
 sg13g2_fill_4 FILLER_48_1478 ();
 sg13g2_fill_8 FILLER_48_1504 ();
 sg13g2_fill_8 FILLER_48_1512 ();
 sg13g2_fill_8 FILLER_48_1520 ();
 sg13g2_fill_8 FILLER_48_1528 ();
 sg13g2_fill_8 FILLER_48_1536 ();
 sg13g2_fill_4 FILLER_48_1544 ();
 sg13g2_fill_1 FILLER_48_1548 ();
 sg13g2_fill_2 FILLER_48_1589 ();
 sg13g2_fill_1 FILLER_48_1591 ();
 sg13g2_fill_8 FILLER_49_0 ();
 sg13g2_fill_8 FILLER_49_8 ();
 sg13g2_fill_8 FILLER_49_16 ();
 sg13g2_fill_4 FILLER_49_24 ();
 sg13g2_fill_8 FILLER_49_38 ();
 sg13g2_fill_8 FILLER_49_46 ();
 sg13g2_fill_4 FILLER_49_54 ();
 sg13g2_fill_2 FILLER_49_58 ();
 sg13g2_fill_8 FILLER_49_70 ();
 sg13g2_fill_4 FILLER_49_78 ();
 sg13g2_fill_8 FILLER_49_92 ();
 sg13g2_fill_8 FILLER_49_100 ();
 sg13g2_fill_2 FILLER_49_108 ();
 sg13g2_fill_1 FILLER_49_110 ();
 sg13g2_fill_1 FILLER_49_121 ();
 sg13g2_fill_8 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_167 ();
 sg13g2_fill_8 FILLER_49_220 ();
 sg13g2_fill_4 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_232 ();
 sg13g2_fill_8 FILLER_49_244 ();
 sg13g2_fill_8 FILLER_49_252 ();
 sg13g2_fill_8 FILLER_49_260 ();
 sg13g2_fill_8 FILLER_49_268 ();
 sg13g2_fill_8 FILLER_49_276 ();
 sg13g2_fill_1 FILLER_49_284 ();
 sg13g2_fill_8 FILLER_49_311 ();
 sg13g2_fill_4 FILLER_49_319 ();
 sg13g2_fill_2 FILLER_49_323 ();
 sg13g2_fill_1 FILLER_49_325 ();
 sg13g2_fill_2 FILLER_49_344 ();
 sg13g2_fill_1 FILLER_49_346 ();
 sg13g2_fill_8 FILLER_49_365 ();
 sg13g2_fill_8 FILLER_49_373 ();
 sg13g2_fill_8 FILLER_49_381 ();
 sg13g2_fill_8 FILLER_49_389 ();
 sg13g2_fill_8 FILLER_49_407 ();
 sg13g2_fill_8 FILLER_49_415 ();
 sg13g2_fill_8 FILLER_49_433 ();
 sg13g2_fill_4 FILLER_49_441 ();
 sg13g2_fill_2 FILLER_49_445 ();
 sg13g2_fill_2 FILLER_49_483 ();
 sg13g2_fill_1 FILLER_49_491 ();
 sg13g2_fill_8 FILLER_49_502 ();
 sg13g2_fill_1 FILLER_49_510 ();
 sg13g2_fill_4 FILLER_49_521 ();
 sg13g2_fill_2 FILLER_49_525 ();
 sg13g2_fill_4 FILLER_49_537 ();
 sg13g2_fill_1 FILLER_49_547 ();
 sg13g2_fill_1 FILLER_49_584 ();
 sg13g2_fill_1 FILLER_49_621 ();
 sg13g2_fill_4 FILLER_49_627 ();
 sg13g2_fill_2 FILLER_49_631 ();
 sg13g2_fill_1 FILLER_49_633 ();
 sg13g2_fill_2 FILLER_49_639 ();
 sg13g2_fill_4 FILLER_49_648 ();
 sg13g2_fill_4 FILLER_49_655 ();
 sg13g2_fill_1 FILLER_49_659 ();
 sg13g2_fill_4 FILLER_49_701 ();
 sg13g2_fill_1 FILLER_49_705 ();
 sg13g2_fill_4 FILLER_49_721 ();
 sg13g2_fill_2 FILLER_49_725 ();
 sg13g2_fill_1 FILLER_49_727 ();
 sg13g2_fill_2 FILLER_49_746 ();
 sg13g2_fill_1 FILLER_49_748 ();
 sg13g2_fill_2 FILLER_49_757 ();
 sg13g2_fill_2 FILLER_49_778 ();
 sg13g2_fill_1 FILLER_49_780 ();
 sg13g2_fill_2 FILLER_49_786 ();
 sg13g2_fill_1 FILLER_49_788 ();
 sg13g2_fill_4 FILLER_49_793 ();
 sg13g2_fill_8 FILLER_49_802 ();
 sg13g2_fill_2 FILLER_49_810 ();
 sg13g2_fill_1 FILLER_49_812 ();
 sg13g2_fill_4 FILLER_49_818 ();
 sg13g2_fill_4 FILLER_49_830 ();
 sg13g2_fill_1 FILLER_49_834 ();
 sg13g2_fill_2 FILLER_49_857 ();
 sg13g2_fill_4 FILLER_49_891 ();
 sg13g2_fill_1 FILLER_49_895 ();
 sg13g2_fill_2 FILLER_49_902 ();
 sg13g2_fill_2 FILLER_49_907 ();
 sg13g2_fill_1 FILLER_49_941 ();
 sg13g2_fill_2 FILLER_49_948 ();
 sg13g2_fill_1 FILLER_49_960 ();
 sg13g2_fill_1 FILLER_49_969 ();
 sg13g2_fill_1 FILLER_49_978 ();
 sg13g2_fill_8 FILLER_49_990 ();
 sg13g2_fill_2 FILLER_49_998 ();
 sg13g2_fill_1 FILLER_49_1000 ();
 sg13g2_fill_4 FILLER_49_1041 ();
 sg13g2_fill_1 FILLER_49_1045 ();
 sg13g2_fill_2 FILLER_49_1072 ();
 sg13g2_fill_8 FILLER_49_1108 ();
 sg13g2_fill_2 FILLER_49_1129 ();
 sg13g2_fill_2 FILLER_49_1136 ();
 sg13g2_fill_1 FILLER_49_1138 ();
 sg13g2_fill_1 FILLER_49_1145 ();
 sg13g2_fill_4 FILLER_49_1160 ();
 sg13g2_fill_2 FILLER_49_1223 ();
 sg13g2_fill_1 FILLER_49_1225 ();
 sg13g2_fill_4 FILLER_49_1229 ();
 sg13g2_fill_2 FILLER_49_1233 ();
 sg13g2_fill_2 FILLER_49_1271 ();
 sg13g2_fill_8 FILLER_49_1276 ();
 sg13g2_fill_4 FILLER_49_1284 ();
 sg13g2_fill_2 FILLER_49_1288 ();
 sg13g2_fill_1 FILLER_49_1290 ();
 sg13g2_fill_2 FILLER_49_1321 ();
 sg13g2_fill_2 FILLER_49_1335 ();
 sg13g2_fill_2 FILLER_49_1349 ();
 sg13g2_fill_1 FILLER_49_1359 ();
 sg13g2_fill_1 FILLER_49_1371 ();
 sg13g2_fill_4 FILLER_49_1443 ();
 sg13g2_fill_2 FILLER_49_1447 ();
 sg13g2_fill_4 FILLER_49_1490 ();
 sg13g2_fill_2 FILLER_49_1494 ();
 sg13g2_fill_1 FILLER_49_1496 ();
 sg13g2_fill_4 FILLER_49_1505 ();
 sg13g2_fill_2 FILLER_49_1519 ();
 sg13g2_fill_1 FILLER_49_1521 ();
 sg13g2_fill_1 FILLER_49_1530 ();
 sg13g2_fill_8 FILLER_49_1536 ();
 sg13g2_fill_4 FILLER_49_1544 ();
 sg13g2_fill_1 FILLER_49_1548 ();
 sg13g2_fill_2 FILLER_49_1589 ();
 sg13g2_fill_1 FILLER_49_1591 ();
 sg13g2_fill_8 FILLER_50_0 ();
 sg13g2_fill_4 FILLER_50_8 ();
 sg13g2_fill_8 FILLER_50_38 ();
 sg13g2_fill_4 FILLER_50_56 ();
 sg13g2_fill_4 FILLER_50_76 ();
 sg13g2_fill_2 FILLER_50_85 ();
 sg13g2_fill_1 FILLER_50_97 ();
 sg13g2_fill_8 FILLER_50_124 ();
 sg13g2_fill_1 FILLER_50_132 ();
 sg13g2_fill_4 FILLER_50_153 ();
 sg13g2_fill_1 FILLER_50_157 ();
 sg13g2_fill_4 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_50_234 ();
 sg13g2_fill_8 FILLER_50_266 ();
 sg13g2_fill_8 FILLER_50_274 ();
 sg13g2_fill_2 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_2 FILLER_50_326 ();
 sg13g2_fill_1 FILLER_50_328 ();
 sg13g2_fill_2 FILLER_50_354 ();
 sg13g2_fill_1 FILLER_50_356 ();
 sg13g2_fill_8 FILLER_50_365 ();
 sg13g2_fill_8 FILLER_50_373 ();
 sg13g2_fill_8 FILLER_50_389 ();
 sg13g2_fill_2 FILLER_50_397 ();
 sg13g2_fill_8 FILLER_50_451 ();
 sg13g2_fill_1 FILLER_50_459 ();
 sg13g2_fill_4 FILLER_50_470 ();
 sg13g2_fill_2 FILLER_50_474 ();
 sg13g2_fill_2 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_488 ();
 sg13g2_fill_2 FILLER_50_547 ();
 sg13g2_fill_1 FILLER_50_549 ();
 sg13g2_fill_4 FILLER_50_566 ();
 sg13g2_fill_8 FILLER_50_580 ();
 sg13g2_fill_8 FILLER_50_588 ();
 sg13g2_fill_8 FILLER_50_596 ();
 sg13g2_fill_4 FILLER_50_604 ();
 sg13g2_fill_2 FILLER_50_608 ();
 sg13g2_fill_1 FILLER_50_610 ();
 sg13g2_fill_4 FILLER_50_623 ();
 sg13g2_fill_1 FILLER_50_641 ();
 sg13g2_fill_2 FILLER_50_664 ();
 sg13g2_fill_1 FILLER_50_666 ();
 sg13g2_fill_8 FILLER_50_672 ();
 sg13g2_fill_2 FILLER_50_685 ();
 sg13g2_fill_8 FILLER_50_692 ();
 sg13g2_fill_2 FILLER_50_700 ();
 sg13g2_fill_8 FILLER_50_705 ();
 sg13g2_fill_8 FILLER_50_713 ();
 sg13g2_fill_8 FILLER_50_721 ();
 sg13g2_fill_4 FILLER_50_729 ();
 sg13g2_fill_2 FILLER_50_733 ();
 sg13g2_fill_1 FILLER_50_735 ();
 sg13g2_fill_4 FILLER_50_741 ();
 sg13g2_fill_2 FILLER_50_745 ();
 sg13g2_fill_1 FILLER_50_747 ();
 sg13g2_fill_8 FILLER_50_788 ();
 sg13g2_fill_1 FILLER_50_796 ();
 sg13g2_fill_2 FILLER_50_808 ();
 sg13g2_fill_2 FILLER_50_819 ();
 sg13g2_fill_2 FILLER_50_837 ();
 sg13g2_fill_8 FILLER_50_843 ();
 sg13g2_fill_8 FILLER_50_851 ();
 sg13g2_fill_8 FILLER_50_859 ();
 sg13g2_fill_8 FILLER_50_867 ();
 sg13g2_fill_1 FILLER_50_875 ();
 sg13g2_fill_4 FILLER_50_888 ();
 sg13g2_fill_1 FILLER_50_901 ();
 sg13g2_fill_1 FILLER_50_905 ();
 sg13g2_fill_2 FILLER_50_912 ();
 sg13g2_fill_1 FILLER_50_965 ();
 sg13g2_fill_1 FILLER_50_984 ();
 sg13g2_fill_4 FILLER_50_1032 ();
 sg13g2_fill_4 FILLER_50_1047 ();
 sg13g2_fill_1 FILLER_50_1051 ();
 sg13g2_fill_2 FILLER_50_1058 ();
 sg13g2_fill_8 FILLER_50_1064 ();
 sg13g2_fill_1 FILLER_50_1072 ();
 sg13g2_fill_4 FILLER_50_1078 ();
 sg13g2_fill_4 FILLER_50_1096 ();
 sg13g2_fill_2 FILLER_50_1100 ();
 sg13g2_fill_1 FILLER_50_1102 ();
 sg13g2_fill_4 FILLER_50_1123 ();
 sg13g2_fill_1 FILLER_50_1127 ();
 sg13g2_fill_4 FILLER_50_1152 ();
 sg13g2_fill_1 FILLER_50_1168 ();
 sg13g2_fill_8 FILLER_50_1175 ();
 sg13g2_fill_2 FILLER_50_1183 ();
 sg13g2_fill_1 FILLER_50_1195 ();
 sg13g2_fill_2 FILLER_50_1220 ();
 sg13g2_fill_8 FILLER_50_1242 ();
 sg13g2_fill_8 FILLER_50_1250 ();
 sg13g2_fill_8 FILLER_50_1258 ();
 sg13g2_fill_8 FILLER_50_1266 ();
 sg13g2_fill_2 FILLER_50_1274 ();
 sg13g2_fill_1 FILLER_50_1276 ();
 sg13g2_fill_2 FILLER_50_1307 ();
 sg13g2_fill_2 FILLER_50_1332 ();
 sg13g2_fill_1 FILLER_50_1343 ();
 sg13g2_fill_2 FILLER_50_1350 ();
 sg13g2_fill_1 FILLER_50_1363 ();
 sg13g2_fill_8 FILLER_50_1385 ();
 sg13g2_fill_2 FILLER_50_1393 ();
 sg13g2_fill_1 FILLER_50_1395 ();
 sg13g2_fill_2 FILLER_50_1399 ();
 sg13g2_fill_8 FILLER_50_1407 ();
 sg13g2_fill_8 FILLER_50_1415 ();
 sg13g2_fill_4 FILLER_50_1423 ();
 sg13g2_fill_4 FILLER_50_1449 ();
 sg13g2_fill_1 FILLER_50_1453 ();
 sg13g2_fill_8 FILLER_50_1458 ();
 sg13g2_fill_8 FILLER_50_1466 ();
 sg13g2_fill_8 FILLER_50_1474 ();
 sg13g2_fill_8 FILLER_50_1482 ();
 sg13g2_fill_8 FILLER_50_1490 ();
 sg13g2_fill_4 FILLER_50_1498 ();
 sg13g2_fill_1 FILLER_50_1502 ();
 sg13g2_fill_8 FILLER_50_1563 ();
 sg13g2_fill_8 FILLER_50_1571 ();
 sg13g2_fill_8 FILLER_50_1579 ();
 sg13g2_fill_4 FILLER_50_1587 ();
 sg13g2_fill_1 FILLER_50_1591 ();
 sg13g2_fill_8 FILLER_51_0 ();
 sg13g2_fill_8 FILLER_51_8 ();
 sg13g2_fill_8 FILLER_51_16 ();
 sg13g2_fill_4 FILLER_51_24 ();
 sg13g2_fill_1 FILLER_51_69 ();
 sg13g2_fill_1 FILLER_51_76 ();
 sg13g2_fill_2 FILLER_51_87 ();
 sg13g2_fill_1 FILLER_51_89 ();
 sg13g2_fill_8 FILLER_51_101 ();
 sg13g2_fill_4 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_113 ();
 sg13g2_fill_8 FILLER_51_129 ();
 sg13g2_fill_8 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_145 ();
 sg13g2_fill_1 FILLER_51_147 ();
 sg13g2_fill_4 FILLER_51_174 ();
 sg13g2_fill_2 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_211 ();
 sg13g2_fill_1 FILLER_51_213 ();
 sg13g2_fill_4 FILLER_51_219 ();
 sg13g2_fill_2 FILLER_51_223 ();
 sg13g2_fill_1 FILLER_51_225 ();
 sg13g2_fill_8 FILLER_51_302 ();
 sg13g2_fill_8 FILLER_51_310 ();
 sg13g2_fill_8 FILLER_51_318 ();
 sg13g2_fill_8 FILLER_51_326 ();
 sg13g2_fill_8 FILLER_51_334 ();
 sg13g2_fill_4 FILLER_51_342 ();
 sg13g2_fill_8 FILLER_51_393 ();
 sg13g2_fill_8 FILLER_51_401 ();
 sg13g2_fill_8 FILLER_51_409 ();
 sg13g2_fill_8 FILLER_51_417 ();
 sg13g2_fill_4 FILLER_51_425 ();
 sg13g2_fill_2 FILLER_51_429 ();
 sg13g2_fill_1 FILLER_51_431 ();
 sg13g2_fill_8 FILLER_51_452 ();
 sg13g2_fill_8 FILLER_51_460 ();
 sg13g2_fill_4 FILLER_51_468 ();
 sg13g2_fill_1 FILLER_51_472 ();
 sg13g2_fill_8 FILLER_51_498 ();
 sg13g2_fill_8 FILLER_51_506 ();
 sg13g2_fill_8 FILLER_51_514 ();
 sg13g2_fill_2 FILLER_51_522 ();
 sg13g2_fill_4 FILLER_51_534 ();
 sg13g2_fill_4 FILLER_51_579 ();
 sg13g2_fill_1 FILLER_51_583 ();
 sg13g2_fill_2 FILLER_51_622 ();
 sg13g2_fill_2 FILLER_51_637 ();
 sg13g2_fill_1 FILLER_51_667 ();
 sg13g2_fill_1 FILLER_51_693 ();
 sg13g2_fill_8 FILLER_51_731 ();
 sg13g2_fill_1 FILLER_51_739 ();
 sg13g2_fill_8 FILLER_51_762 ();
 sg13g2_fill_4 FILLER_51_770 ();
 sg13g2_fill_2 FILLER_51_774 ();
 sg13g2_fill_2 FILLER_51_784 ();
 sg13g2_fill_4 FILLER_51_791 ();
 sg13g2_fill_1 FILLER_51_795 ();
 sg13g2_fill_1 FILLER_51_812 ();
 sg13g2_fill_2 FILLER_51_829 ();
 sg13g2_fill_1 FILLER_51_836 ();
 sg13g2_fill_1 FILLER_51_842 ();
 sg13g2_fill_1 FILLER_51_854 ();
 sg13g2_fill_2 FILLER_51_866 ();
 sg13g2_fill_4 FILLER_51_873 ();
 sg13g2_fill_4 FILLER_51_882 ();
 sg13g2_fill_2 FILLER_51_886 ();
 sg13g2_fill_1 FILLER_51_888 ();
 sg13g2_fill_1 FILLER_51_908 ();
 sg13g2_fill_1 FILLER_51_912 ();
 sg13g2_fill_2 FILLER_51_931 ();
 sg13g2_fill_2 FILLER_51_936 ();
 sg13g2_fill_2 FILLER_51_960 ();
 sg13g2_fill_2 FILLER_51_988 ();
 sg13g2_fill_8 FILLER_51_1005 ();
 sg13g2_fill_8 FILLER_51_1013 ();
 sg13g2_fill_2 FILLER_51_1021 ();
 sg13g2_fill_1 FILLER_51_1023 ();
 sg13g2_fill_8 FILLER_51_1041 ();
 sg13g2_fill_1 FILLER_51_1049 ();
 sg13g2_fill_8 FILLER_51_1056 ();
 sg13g2_fill_4 FILLER_51_1064 ();
 sg13g2_fill_2 FILLER_51_1073 ();
 sg13g2_fill_8 FILLER_51_1080 ();
 sg13g2_fill_1 FILLER_51_1088 ();
 sg13g2_fill_8 FILLER_51_1094 ();
 sg13g2_fill_8 FILLER_51_1102 ();
 sg13g2_fill_1 FILLER_51_1126 ();
 sg13g2_fill_2 FILLER_51_1135 ();
 sg13g2_fill_8 FILLER_51_1145 ();
 sg13g2_fill_1 FILLER_51_1153 ();
 sg13g2_fill_1 FILLER_51_1158 ();
 sg13g2_fill_1 FILLER_51_1170 ();
 sg13g2_fill_2 FILLER_51_1179 ();
 sg13g2_fill_4 FILLER_51_1197 ();
 sg13g2_fill_2 FILLER_51_1201 ();
 sg13g2_fill_4 FILLER_51_1240 ();
 sg13g2_fill_4 FILLER_51_1252 ();
 sg13g2_fill_2 FILLER_51_1256 ();
 sg13g2_fill_1 FILLER_51_1258 ();
 sg13g2_fill_4 FILLER_51_1262 ();
 sg13g2_fill_2 FILLER_51_1266 ();
 sg13g2_fill_1 FILLER_51_1268 ();
 sg13g2_fill_8 FILLER_51_1283 ();
 sg13g2_fill_2 FILLER_51_1297 ();
 sg13g2_fill_1 FILLER_51_1299 ();
 sg13g2_fill_2 FILLER_51_1316 ();
 sg13g2_fill_2 FILLER_51_1321 ();
 sg13g2_fill_2 FILLER_51_1357 ();
 sg13g2_fill_1 FILLER_51_1370 ();
 sg13g2_fill_8 FILLER_51_1418 ();
 sg13g2_fill_8 FILLER_51_1426 ();
 sg13g2_fill_8 FILLER_51_1434 ();
 sg13g2_fill_8 FILLER_51_1442 ();
 sg13g2_fill_8 FILLER_51_1450 ();
 sg13g2_fill_8 FILLER_51_1458 ();
 sg13g2_fill_8 FILLER_51_1466 ();
 sg13g2_fill_8 FILLER_51_1474 ();
 sg13g2_fill_2 FILLER_51_1482 ();
 sg13g2_fill_1 FILLER_51_1484 ();
 sg13g2_fill_8 FILLER_51_1495 ();
 sg13g2_fill_8 FILLER_51_1503 ();
 sg13g2_fill_8 FILLER_51_1511 ();
 sg13g2_fill_8 FILLER_51_1519 ();
 sg13g2_fill_2 FILLER_51_1527 ();
 sg13g2_fill_1 FILLER_51_1529 ();
 sg13g2_fill_8 FILLER_51_1565 ();
 sg13g2_fill_8 FILLER_51_1573 ();
 sg13g2_fill_8 FILLER_51_1581 ();
 sg13g2_fill_2 FILLER_51_1589 ();
 sg13g2_fill_1 FILLER_51_1591 ();
 sg13g2_fill_8 FILLER_52_0 ();
 sg13g2_fill_4 FILLER_52_8 ();
 sg13g2_fill_1 FILLER_52_12 ();
 sg13g2_fill_1 FILLER_52_57 ();
 sg13g2_fill_8 FILLER_52_64 ();
 sg13g2_fill_8 FILLER_52_72 ();
 sg13g2_fill_1 FILLER_52_80 ();
 sg13g2_fill_8 FILLER_52_92 ();
 sg13g2_fill_8 FILLER_52_100 ();
 sg13g2_fill_2 FILLER_52_108 ();
 sg13g2_fill_2 FILLER_52_120 ();
 sg13g2_fill_1 FILLER_52_122 ();
 sg13g2_fill_2 FILLER_52_133 ();
 sg13g2_fill_4 FILLER_52_160 ();
 sg13g2_fill_2 FILLER_52_164 ();
 sg13g2_fill_2 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_189 ();
 sg13g2_fill_8 FILLER_52_211 ();
 sg13g2_fill_4 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_223 ();
 sg13g2_fill_4 FILLER_52_234 ();
 sg13g2_fill_2 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_240 ();
 sg13g2_fill_8 FILLER_52_267 ();
 sg13g2_fill_2 FILLER_52_275 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_fill_8 FILLER_52_288 ();
 sg13g2_fill_2 FILLER_52_332 ();
 sg13g2_fill_8 FILLER_52_354 ();
 sg13g2_fill_8 FILLER_52_362 ();
 sg13g2_fill_2 FILLER_52_370 ();
 sg13g2_fill_2 FILLER_52_385 ();
 sg13g2_fill_8 FILLER_52_423 ();
 sg13g2_fill_8 FILLER_52_431 ();
 sg13g2_fill_2 FILLER_52_439 ();
 sg13g2_fill_8 FILLER_52_447 ();
 sg13g2_fill_8 FILLER_52_455 ();
 sg13g2_fill_1 FILLER_52_463 ();
 sg13g2_fill_4 FILLER_52_469 ();
 sg13g2_fill_1 FILLER_52_473 ();
 sg13g2_fill_1 FILLER_52_479 ();
 sg13g2_fill_2 FILLER_52_486 ();
 sg13g2_fill_1 FILLER_52_488 ();
 sg13g2_fill_8 FILLER_52_515 ();
 sg13g2_fill_4 FILLER_52_523 ();
 sg13g2_fill_1 FILLER_52_527 ();
 sg13g2_fill_8 FILLER_52_588 ();
 sg13g2_fill_4 FILLER_52_596 ();
 sg13g2_fill_2 FILLER_52_600 ();
 sg13g2_fill_1 FILLER_52_602 ();
 sg13g2_fill_1 FILLER_52_648 ();
 sg13g2_fill_8 FILLER_52_699 ();
 sg13g2_fill_1 FILLER_52_772 ();
 sg13g2_fill_2 FILLER_52_777 ();
 sg13g2_fill_1 FILLER_52_798 ();
 sg13g2_fill_1 FILLER_52_807 ();
 sg13g2_fill_2 FILLER_52_834 ();
 sg13g2_fill_1 FILLER_52_864 ();
 sg13g2_fill_2 FILLER_52_889 ();
 sg13g2_fill_1 FILLER_52_908 ();
 sg13g2_fill_2 FILLER_52_928 ();
 sg13g2_fill_2 FILLER_52_942 ();
 sg13g2_fill_1 FILLER_52_984 ();
 sg13g2_fill_2 FILLER_52_990 ();
 sg13g2_fill_2 FILLER_52_1018 ();
 sg13g2_fill_2 FILLER_52_1045 ();
 sg13g2_fill_8 FILLER_52_1060 ();
 sg13g2_fill_1 FILLER_52_1068 ();
 sg13g2_fill_8 FILLER_52_1088 ();
 sg13g2_fill_8 FILLER_52_1096 ();
 sg13g2_fill_8 FILLER_52_1120 ();
 sg13g2_fill_8 FILLER_52_1137 ();
 sg13g2_fill_4 FILLER_52_1145 ();
 sg13g2_fill_2 FILLER_52_1149 ();
 sg13g2_fill_1 FILLER_52_1151 ();
 sg13g2_fill_4 FILLER_52_1169 ();
 sg13g2_fill_1 FILLER_52_1173 ();
 sg13g2_fill_1 FILLER_52_1182 ();
 sg13g2_fill_1 FILLER_52_1186 ();
 sg13g2_fill_1 FILLER_52_1222 ();
 sg13g2_fill_1 FILLER_52_1231 ();
 sg13g2_fill_4 FILLER_52_1253 ();
 sg13g2_fill_1 FILLER_52_1265 ();
 sg13g2_fill_2 FILLER_52_1277 ();
 sg13g2_fill_2 FILLER_52_1290 ();
 sg13g2_fill_4 FILLER_52_1300 ();
 sg13g2_fill_2 FILLER_52_1304 ();
 sg13g2_fill_1 FILLER_52_1351 ();
 sg13g2_fill_1 FILLER_52_1374 ();
 sg13g2_fill_2 FILLER_52_1415 ();
 sg13g2_fill_2 FILLER_52_1447 ();
 sg13g2_fill_1 FILLER_52_1449 ();
 sg13g2_fill_1 FILLER_52_1490 ();
 sg13g2_fill_4 FILLER_52_1524 ();
 sg13g2_fill_2 FILLER_52_1528 ();
 sg13g2_fill_8 FILLER_52_1553 ();
 sg13g2_fill_1 FILLER_52_1561 ();
 sg13g2_fill_8 FILLER_53_0 ();
 sg13g2_fill_8 FILLER_53_8 ();
 sg13g2_fill_8 FILLER_53_16 ();
 sg13g2_fill_4 FILLER_53_24 ();
 sg13g2_fill_4 FILLER_53_51 ();
 sg13g2_fill_1 FILLER_53_55 ();
 sg13g2_fill_8 FILLER_53_62 ();
 sg13g2_fill_8 FILLER_53_70 ();
 sg13g2_fill_1 FILLER_53_78 ();
 sg13g2_fill_8 FILLER_53_85 ();
 sg13g2_fill_4 FILLER_53_93 ();
 sg13g2_fill_2 FILLER_53_97 ();
 sg13g2_fill_2 FILLER_53_172 ();
 sg13g2_fill_4 FILLER_53_207 ();
 sg13g2_fill_2 FILLER_53_211 ();
 sg13g2_fill_2 FILLER_53_239 ();
 sg13g2_fill_8 FILLER_53_262 ();
 sg13g2_fill_8 FILLER_53_270 ();
 sg13g2_fill_4 FILLER_53_278 ();
 sg13g2_fill_1 FILLER_53_282 ();
 sg13g2_fill_4 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_307 ();
 sg13g2_fill_8 FILLER_53_335 ();
 sg13g2_fill_1 FILLER_53_343 ();
 sg13g2_fill_8 FILLER_53_380 ();
 sg13g2_fill_4 FILLER_53_388 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_fill_2 FILLER_53_429 ();
 sg13g2_fill_1 FILLER_53_431 ();
 sg13g2_fill_8 FILLER_53_452 ();
 sg13g2_fill_1 FILLER_53_460 ();
 sg13g2_fill_8 FILLER_53_474 ();
 sg13g2_fill_1 FILLER_53_482 ();
 sg13g2_fill_1 FILLER_53_493 ();
 sg13g2_fill_8 FILLER_53_499 ();
 sg13g2_fill_2 FILLER_53_507 ();
 sg13g2_fill_1 FILLER_53_509 ();
 sg13g2_fill_4 FILLER_53_520 ();
 sg13g2_fill_2 FILLER_53_524 ();
 sg13g2_fill_1 FILLER_53_526 ();
 sg13g2_fill_8 FILLER_53_537 ();
 sg13g2_fill_8 FILLER_53_545 ();
 sg13g2_fill_8 FILLER_53_553 ();
 sg13g2_fill_8 FILLER_53_561 ();
 sg13g2_fill_8 FILLER_53_569 ();
 sg13g2_fill_8 FILLER_53_577 ();
 sg13g2_fill_8 FILLER_53_585 ();
 sg13g2_fill_1 FILLER_53_593 ();
 sg13g2_fill_1 FILLER_53_632 ();
 sg13g2_fill_2 FILLER_53_666 ();
 sg13g2_fill_2 FILLER_53_691 ();
 sg13g2_fill_1 FILLER_53_698 ();
 sg13g2_fill_8 FILLER_53_708 ();
 sg13g2_fill_4 FILLER_53_716 ();
 sg13g2_fill_2 FILLER_53_720 ();
 sg13g2_fill_1 FILLER_53_722 ();
 sg13g2_fill_4 FILLER_53_731 ();
 sg13g2_fill_2 FILLER_53_735 ();
 sg13g2_fill_1 FILLER_53_737 ();
 sg13g2_fill_1 FILLER_53_762 ();
 sg13g2_fill_4 FILLER_53_799 ();
 sg13g2_fill_2 FILLER_53_803 ();
 sg13g2_fill_1 FILLER_53_805 ();
 sg13g2_fill_2 FILLER_53_812 ();
 sg13g2_fill_2 FILLER_53_836 ();
 sg13g2_fill_4 FILLER_53_847 ();
 sg13g2_fill_1 FILLER_53_851 ();
 sg13g2_fill_8 FILLER_53_861 ();
 sg13g2_fill_4 FILLER_53_869 ();
 sg13g2_fill_2 FILLER_53_873 ();
 sg13g2_fill_2 FILLER_53_889 ();
 sg13g2_fill_2 FILLER_53_897 ();
 sg13g2_fill_1 FILLER_53_908 ();
 sg13g2_fill_2 FILLER_53_934 ();
 sg13g2_fill_1 FILLER_53_973 ();
 sg13g2_fill_2 FILLER_53_1011 ();
 sg13g2_fill_1 FILLER_53_1013 ();
 sg13g2_fill_1 FILLER_53_1039 ();
 sg13g2_fill_1 FILLER_53_1072 ();
 sg13g2_fill_4 FILLER_53_1077 ();
 sg13g2_fill_8 FILLER_53_1090 ();
 sg13g2_fill_8 FILLER_53_1098 ();
 sg13g2_fill_1 FILLER_53_1106 ();
 sg13g2_fill_8 FILLER_53_1117 ();
 sg13g2_fill_1 FILLER_53_1125 ();
 sg13g2_fill_8 FILLER_53_1134 ();
 sg13g2_fill_8 FILLER_53_1142 ();
 sg13g2_fill_1 FILLER_53_1163 ();
 sg13g2_fill_2 FILLER_53_1175 ();
 sg13g2_fill_1 FILLER_53_1191 ();
 sg13g2_fill_2 FILLER_53_1207 ();
 sg13g2_fill_2 FILLER_53_1219 ();
 sg13g2_fill_1 FILLER_53_1226 ();
 sg13g2_fill_4 FILLER_53_1245 ();
 sg13g2_fill_8 FILLER_53_1260 ();
 sg13g2_fill_4 FILLER_53_1268 ();
 sg13g2_fill_1 FILLER_53_1272 ();
 sg13g2_fill_2 FILLER_53_1284 ();
 sg13g2_fill_1 FILLER_53_1286 ();
 sg13g2_fill_1 FILLER_53_1317 ();
 sg13g2_fill_2 FILLER_53_1340 ();
 sg13g2_fill_2 FILLER_53_1356 ();
 sg13g2_fill_2 FILLER_53_1407 ();
 sg13g2_fill_2 FILLER_53_1419 ();
 sg13g2_fill_1 FILLER_53_1421 ();
 sg13g2_fill_4 FILLER_53_1452 ();
 sg13g2_fill_2 FILLER_53_1456 ();
 sg13g2_fill_2 FILLER_53_1488 ();
 sg13g2_fill_1 FILLER_53_1490 ();
 sg13g2_fill_4 FILLER_53_1501 ();
 sg13g2_fill_2 FILLER_53_1505 ();
 sg13g2_fill_1 FILLER_53_1507 ();
 sg13g2_fill_8 FILLER_53_1563 ();
 sg13g2_fill_8 FILLER_53_1571 ();
 sg13g2_fill_8 FILLER_53_1579 ();
 sg13g2_fill_4 FILLER_53_1587 ();
 sg13g2_fill_1 FILLER_53_1591 ();
 sg13g2_fill_8 FILLER_54_0 ();
 sg13g2_fill_2 FILLER_54_8 ();
 sg13g2_fill_1 FILLER_54_10 ();
 sg13g2_fill_4 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_69 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_8 FILLER_54_194 ();
 sg13g2_fill_4 FILLER_54_202 ();
 sg13g2_fill_8 FILLER_54_214 ();
 sg13g2_fill_8 FILLER_54_222 ();
 sg13g2_fill_8 FILLER_54_230 ();
 sg13g2_fill_1 FILLER_54_248 ();
 sg13g2_fill_2 FILLER_54_270 ();
 sg13g2_fill_4 FILLER_54_282 ();
 sg13g2_fill_2 FILLER_54_286 ();
 sg13g2_fill_1 FILLER_54_288 ();
 sg13g2_fill_8 FILLER_54_315 ();
 sg13g2_fill_1 FILLER_54_323 ();
 sg13g2_fill_8 FILLER_54_344 ();
 sg13g2_fill_8 FILLER_54_352 ();
 sg13g2_fill_8 FILLER_54_360 ();
 sg13g2_fill_8 FILLER_54_368 ();
 sg13g2_fill_2 FILLER_54_376 ();
 sg13g2_fill_1 FILLER_54_378 ();
 sg13g2_fill_2 FILLER_54_466 ();
 sg13g2_fill_1 FILLER_54_504 ();
 sg13g2_fill_2 FILLER_54_531 ();
 sg13g2_fill_4 FILLER_54_576 ();
 sg13g2_fill_1 FILLER_54_580 ();
 sg13g2_fill_8 FILLER_54_598 ();
 sg13g2_fill_2 FILLER_54_606 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_fill_1 FILLER_54_626 ();
 sg13g2_fill_2 FILLER_54_645 ();
 sg13g2_fill_1 FILLER_54_676 ();
 sg13g2_fill_4 FILLER_54_690 ();
 sg13g2_fill_1 FILLER_54_716 ();
 sg13g2_fill_4 FILLER_54_722 ();
 sg13g2_fill_2 FILLER_54_726 ();
 sg13g2_fill_4 FILLER_54_734 ();
 sg13g2_fill_2 FILLER_54_738 ();
 sg13g2_fill_8 FILLER_54_776 ();
 sg13g2_fill_4 FILLER_54_784 ();
 sg13g2_fill_2 FILLER_54_788 ();
 sg13g2_fill_1 FILLER_54_790 ();
 sg13g2_fill_1 FILLER_54_805 ();
 sg13g2_fill_1 FILLER_54_815 ();
 sg13g2_fill_8 FILLER_54_829 ();
 sg13g2_fill_8 FILLER_54_837 ();
 sg13g2_fill_8 FILLER_54_845 ();
 sg13g2_fill_4 FILLER_54_853 ();
 sg13g2_fill_1 FILLER_54_857 ();
 sg13g2_fill_8 FILLER_54_863 ();
 sg13g2_fill_8 FILLER_54_871 ();
 sg13g2_fill_2 FILLER_54_879 ();
 sg13g2_fill_1 FILLER_54_881 ();
 sg13g2_fill_1 FILLER_54_916 ();
 sg13g2_fill_1 FILLER_54_927 ();
 sg13g2_fill_2 FILLER_54_940 ();
 sg13g2_fill_1 FILLER_54_948 ();
 sg13g2_fill_2 FILLER_54_980 ();
 sg13g2_fill_1 FILLER_54_1008 ();
 sg13g2_fill_1 FILLER_54_1039 ();
 sg13g2_fill_2 FILLER_54_1082 ();
 sg13g2_fill_4 FILLER_54_1096 ();
 sg13g2_fill_2 FILLER_54_1116 ();
 sg13g2_fill_4 FILLER_54_1139 ();
 sg13g2_fill_1 FILLER_54_1143 ();
 sg13g2_fill_8 FILLER_54_1149 ();
 sg13g2_fill_4 FILLER_54_1157 ();
 sg13g2_fill_2 FILLER_54_1172 ();
 sg13g2_fill_2 FILLER_54_1183 ();
 sg13g2_fill_2 FILLER_54_1198 ();
 sg13g2_fill_2 FILLER_54_1243 ();
 sg13g2_fill_4 FILLER_54_1261 ();
 sg13g2_fill_2 FILLER_54_1265 ();
 sg13g2_fill_8 FILLER_54_1291 ();
 sg13g2_fill_8 FILLER_54_1299 ();
 sg13g2_fill_8 FILLER_54_1307 ();
 sg13g2_fill_2 FILLER_54_1315 ();
 sg13g2_fill_1 FILLER_54_1317 ();
 sg13g2_fill_2 FILLER_54_1330 ();
 sg13g2_fill_2 FILLER_54_1353 ();
 sg13g2_fill_1 FILLER_54_1365 ();
 sg13g2_fill_1 FILLER_54_1375 ();
 sg13g2_fill_1 FILLER_54_1389 ();
 sg13g2_fill_1 FILLER_54_1406 ();
 sg13g2_fill_2 FILLER_54_1415 ();
 sg13g2_fill_4 FILLER_54_1445 ();
 sg13g2_fill_2 FILLER_54_1449 ();
 sg13g2_fill_2 FILLER_54_1489 ();
 sg13g2_fill_8 FILLER_54_1521 ();
 sg13g2_fill_8 FILLER_54_1529 ();
 sg13g2_fill_8 FILLER_54_1537 ();
 sg13g2_fill_4 FILLER_54_1545 ();
 sg13g2_fill_2 FILLER_54_1549 ();
 sg13g2_fill_1 FILLER_54_1561 ();
 sg13g2_fill_8 FILLER_55_0 ();
 sg13g2_fill_8 FILLER_55_8 ();
 sg13g2_fill_8 FILLER_55_16 ();
 sg13g2_fill_8 FILLER_55_24 ();
 sg13g2_fill_8 FILLER_55_32 ();
 sg13g2_fill_4 FILLER_55_50 ();
 sg13g2_fill_2 FILLER_55_54 ();
 sg13g2_fill_1 FILLER_55_56 ();
 sg13g2_fill_1 FILLER_55_67 ();
 sg13g2_fill_4 FILLER_55_83 ();
 sg13g2_fill_1 FILLER_55_87 ();
 sg13g2_fill_8 FILLER_55_113 ();
 sg13g2_fill_8 FILLER_55_121 ();
 sg13g2_fill_8 FILLER_55_129 ();
 sg13g2_fill_4 FILLER_55_137 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_fill_4 FILLER_55_153 ();
 sg13g2_fill_2 FILLER_55_165 ();
 sg13g2_fill_1 FILLER_55_195 ();
 sg13g2_fill_8 FILLER_55_232 ();
 sg13g2_fill_8 FILLER_55_240 ();
 sg13g2_fill_8 FILLER_55_248 ();
 sg13g2_fill_4 FILLER_55_256 ();
 sg13g2_fill_2 FILLER_55_260 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_4 FILLER_55_297 ();
 sg13g2_fill_2 FILLER_55_326 ();
 sg13g2_fill_4 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_342 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_fill_4 FILLER_55_381 ();
 sg13g2_fill_2 FILLER_55_395 ();
 sg13g2_fill_1 FILLER_55_397 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_fill_1 FILLER_55_409 ();
 sg13g2_fill_2 FILLER_55_420 ();
 sg13g2_fill_8 FILLER_55_439 ();
 sg13g2_fill_1 FILLER_55_447 ();
 sg13g2_fill_8 FILLER_55_454 ();
 sg13g2_fill_8 FILLER_55_462 ();
 sg13g2_fill_8 FILLER_55_470 ();
 sg13g2_fill_8 FILLER_55_478 ();
 sg13g2_fill_4 FILLER_55_486 ();
 sg13g2_fill_2 FILLER_55_490 ();
 sg13g2_fill_1 FILLER_55_497 ();
 sg13g2_fill_8 FILLER_55_502 ();
 sg13g2_fill_8 FILLER_55_516 ();
 sg13g2_fill_8 FILLER_55_524 ();
 sg13g2_fill_2 FILLER_55_537 ();
 sg13g2_fill_1 FILLER_55_539 ();
 sg13g2_fill_4 FILLER_55_549 ();
 sg13g2_fill_2 FILLER_55_553 ();
 sg13g2_fill_1 FILLER_55_555 ();
 sg13g2_fill_2 FILLER_55_673 ();
 sg13g2_fill_1 FILLER_55_675 ();
 sg13g2_fill_1 FILLER_55_707 ();
 sg13g2_fill_1 FILLER_55_714 ();
 sg13g2_fill_1 FILLER_55_748 ();
 sg13g2_fill_4 FILLER_55_755 ();
 sg13g2_fill_2 FILLER_55_759 ();
 sg13g2_fill_1 FILLER_55_788 ();
 sg13g2_fill_1 FILLER_55_843 ();
 sg13g2_fill_4 FILLER_55_848 ();
 sg13g2_fill_1 FILLER_55_852 ();
 sg13g2_fill_4 FILLER_55_869 ();
 sg13g2_fill_2 FILLER_55_873 ();
 sg13g2_fill_1 FILLER_55_929 ();
 sg13g2_fill_1 FILLER_55_941 ();
 sg13g2_fill_1 FILLER_55_956 ();
 sg13g2_fill_1 FILLER_55_965 ();
 sg13g2_fill_1 FILLER_55_1033 ();
 sg13g2_fill_1 FILLER_55_1045 ();
 sg13g2_fill_4 FILLER_55_1059 ();
 sg13g2_fill_2 FILLER_55_1063 ();
 sg13g2_fill_1 FILLER_55_1065 ();
 sg13g2_fill_8 FILLER_55_1071 ();
 sg13g2_fill_4 FILLER_55_1100 ();
 sg13g2_fill_1 FILLER_55_1104 ();
 sg13g2_fill_1 FILLER_55_1110 ();
 sg13g2_fill_8 FILLER_55_1115 ();
 sg13g2_fill_1 FILLER_55_1123 ();
 sg13g2_fill_2 FILLER_55_1132 ();
 sg13g2_fill_4 FILLER_55_1162 ();
 sg13g2_fill_1 FILLER_55_1166 ();
 sg13g2_fill_1 FILLER_55_1191 ();
 sg13g2_fill_2 FILLER_55_1214 ();
 sg13g2_fill_4 FILLER_55_1235 ();
 sg13g2_fill_1 FILLER_55_1239 ();
 sg13g2_fill_4 FILLER_55_1245 ();
 sg13g2_fill_2 FILLER_55_1249 ();
 sg13g2_fill_8 FILLER_55_1276 ();
 sg13g2_fill_2 FILLER_55_1292 ();
 sg13g2_fill_1 FILLER_55_1294 ();
 sg13g2_fill_4 FILLER_55_1303 ();
 sg13g2_fill_1 FILLER_55_1307 ();
 sg13g2_fill_1 FILLER_55_1323 ();
 sg13g2_fill_2 FILLER_55_1340 ();
 sg13g2_fill_2 FILLER_55_1358 ();
 sg13g2_fill_1 FILLER_55_1372 ();
 sg13g2_fill_1 FILLER_55_1380 ();
 sg13g2_fill_4 FILLER_55_1413 ();
 sg13g2_fill_2 FILLER_55_1417 ();
 sg13g2_fill_2 FILLER_55_1449 ();
 sg13g2_fill_1 FILLER_55_1451 ();
 sg13g2_fill_8 FILLER_55_1505 ();
 sg13g2_fill_8 FILLER_55_1513 ();
 sg13g2_fill_8 FILLER_55_1521 ();
 sg13g2_fill_8 FILLER_55_1539 ();
 sg13g2_fill_8 FILLER_55_1547 ();
 sg13g2_fill_4 FILLER_55_1555 ();
 sg13g2_fill_2 FILLER_55_1559 ();
 sg13g2_fill_1 FILLER_55_1561 ();
 sg13g2_fill_8 FILLER_56_0 ();
 sg13g2_fill_8 FILLER_56_8 ();
 sg13g2_fill_2 FILLER_56_16 ();
 sg13g2_fill_2 FILLER_56_80 ();
 sg13g2_fill_4 FILLER_56_103 ();
 sg13g2_fill_2 FILLER_56_107 ();
 sg13g2_fill_4 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_175 ();
 sg13g2_fill_8 FILLER_56_185 ();
 sg13g2_fill_8 FILLER_56_193 ();
 sg13g2_fill_8 FILLER_56_201 ();
 sg13g2_fill_8 FILLER_56_209 ();
 sg13g2_fill_4 FILLER_56_217 ();
 sg13g2_fill_8 FILLER_56_250 ();
 sg13g2_fill_8 FILLER_56_273 ();
 sg13g2_fill_4 FILLER_56_281 ();
 sg13g2_fill_2 FILLER_56_285 ();
 sg13g2_fill_1 FILLER_56_287 ();
 sg13g2_fill_2 FILLER_56_340 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_fill_8 FILLER_56_385 ();
 sg13g2_fill_8 FILLER_56_393 ();
 sg13g2_fill_8 FILLER_56_401 ();
 sg13g2_fill_4 FILLER_56_409 ();
 sg13g2_fill_2 FILLER_56_413 ();
 sg13g2_fill_4 FILLER_56_419 ();
 sg13g2_fill_8 FILLER_56_428 ();
 sg13g2_fill_1 FILLER_56_436 ();
 sg13g2_fill_1 FILLER_56_441 ();
 sg13g2_fill_8 FILLER_56_447 ();
 sg13g2_fill_8 FILLER_56_455 ();
 sg13g2_fill_2 FILLER_56_463 ();
 sg13g2_fill_1 FILLER_56_465 ();
 sg13g2_fill_2 FILLER_56_502 ();
 sg13g2_fill_1 FILLER_56_504 ();
 sg13g2_fill_4 FILLER_56_515 ();
 sg13g2_fill_1 FILLER_56_519 ();
 sg13g2_fill_2 FILLER_56_530 ();
 sg13g2_fill_1 FILLER_56_532 ();
 sg13g2_fill_1 FILLER_56_544 ();
 sg13g2_fill_1 FILLER_56_554 ();
 sg13g2_fill_4 FILLER_56_565 ();
 sg13g2_fill_8 FILLER_56_574 ();
 sg13g2_fill_8 FILLER_56_582 ();
 sg13g2_fill_8 FILLER_56_590 ();
 sg13g2_fill_4 FILLER_56_598 ();
 sg13g2_fill_2 FILLER_56_627 ();
 sg13g2_fill_1 FILLER_56_639 ();
 sg13g2_fill_2 FILLER_56_674 ();
 sg13g2_fill_2 FILLER_56_702 ();
 sg13g2_fill_1 FILLER_56_704 ();
 sg13g2_fill_2 FILLER_56_711 ();
 sg13g2_fill_1 FILLER_56_713 ();
 sg13g2_fill_8 FILLER_56_724 ();
 sg13g2_fill_4 FILLER_56_732 ();
 sg13g2_fill_2 FILLER_56_736 ();
 sg13g2_fill_1 FILLER_56_738 ();
 sg13g2_fill_4 FILLER_56_760 ();
 sg13g2_fill_2 FILLER_56_796 ();
 sg13g2_fill_2 FILLER_56_857 ();
 sg13g2_fill_2 FILLER_56_872 ();
 sg13g2_fill_1 FILLER_56_874 ();
 sg13g2_fill_1 FILLER_56_896 ();
 sg13g2_fill_1 FILLER_56_923 ();
 sg13g2_fill_2 FILLER_56_984 ();
 sg13g2_fill_1 FILLER_56_986 ();
 sg13g2_fill_8 FILLER_56_990 ();
 sg13g2_fill_8 FILLER_56_998 ();
 sg13g2_fill_8 FILLER_56_1006 ();
 sg13g2_fill_8 FILLER_56_1014 ();
 sg13g2_fill_4 FILLER_56_1022 ();
 sg13g2_fill_8 FILLER_56_1061 ();
 sg13g2_fill_8 FILLER_56_1069 ();
 sg13g2_fill_1 FILLER_56_1082 ();
 sg13g2_fill_8 FILLER_56_1088 ();
 sg13g2_fill_2 FILLER_56_1096 ();
 sg13g2_fill_1 FILLER_56_1098 ();
 sg13g2_fill_1 FILLER_56_1113 ();
 sg13g2_fill_8 FILLER_56_1119 ();
 sg13g2_fill_8 FILLER_56_1127 ();
 sg13g2_fill_4 FILLER_56_1135 ();
 sg13g2_fill_2 FILLER_56_1149 ();
 sg13g2_fill_4 FILLER_56_1158 ();
 sg13g2_fill_2 FILLER_56_1162 ();
 sg13g2_fill_8 FILLER_56_1169 ();
 sg13g2_fill_2 FILLER_56_1177 ();
 sg13g2_fill_2 FILLER_56_1192 ();
 sg13g2_fill_8 FILLER_56_1220 ();
 sg13g2_fill_1 FILLER_56_1228 ();
 sg13g2_fill_8 FILLER_56_1244 ();
 sg13g2_fill_8 FILLER_56_1252 ();
 sg13g2_fill_8 FILLER_56_1260 ();
 sg13g2_fill_2 FILLER_56_1268 ();
 sg13g2_fill_8 FILLER_56_1278 ();
 sg13g2_fill_4 FILLER_56_1286 ();
 sg13g2_fill_4 FILLER_56_1294 ();
 sg13g2_fill_2 FILLER_56_1298 ();
 sg13g2_fill_2 FILLER_56_1314 ();
 sg13g2_fill_1 FILLER_56_1325 ();
 sg13g2_fill_1 FILLER_56_1345 ();
 sg13g2_fill_2 FILLER_56_1373 ();
 sg13g2_fill_2 FILLER_56_1380 ();
 sg13g2_fill_1 FILLER_56_1392 ();
 sg13g2_fill_8 FILLER_56_1398 ();
 sg13g2_fill_2 FILLER_56_1406 ();
 sg13g2_fill_1 FILLER_56_1428 ();
 sg13g2_fill_4 FILLER_56_1476 ();
 sg13g2_fill_2 FILLER_56_1480 ();
 sg13g2_fill_1 FILLER_56_1492 ();
 sg13g2_fill_1 FILLER_56_1503 ();
 sg13g2_fill_2 FILLER_56_1564 ();
 sg13g2_fill_1 FILLER_56_1566 ();
 sg13g2_fill_8 FILLER_57_0 ();
 sg13g2_fill_8 FILLER_57_8 ();
 sg13g2_fill_8 FILLER_57_16 ();
 sg13g2_fill_8 FILLER_57_24 ();
 sg13g2_fill_8 FILLER_57_32 ();
 sg13g2_fill_8 FILLER_57_40 ();
 sg13g2_fill_8 FILLER_57_48 ();
 sg13g2_fill_8 FILLER_57_56 ();
 sg13g2_fill_4 FILLER_57_64 ();
 sg13g2_fill_2 FILLER_57_68 ();
 sg13g2_fill_8 FILLER_57_80 ();
 sg13g2_fill_1 FILLER_57_88 ();
 sg13g2_fill_8 FILLER_57_94 ();
 sg13g2_fill_1 FILLER_57_102 ();
 sg13g2_fill_8 FILLER_57_139 ();
 sg13g2_fill_8 FILLER_57_147 ();
 sg13g2_fill_8 FILLER_57_155 ();
 sg13g2_fill_2 FILLER_57_163 ();
 sg13g2_fill_1 FILLER_57_165 ();
 sg13g2_fill_1 FILLER_57_174 ();
 sg13g2_fill_1 FILLER_57_183 ();
 sg13g2_fill_1 FILLER_57_194 ();
 sg13g2_fill_1 FILLER_57_221 ();
 sg13g2_fill_4 FILLER_57_243 ();
 sg13g2_fill_2 FILLER_57_281 ();
 sg13g2_fill_8 FILLER_57_310 ();
 sg13g2_fill_8 FILLER_57_318 ();
 sg13g2_fill_8 FILLER_57_326 ();
 sg13g2_fill_2 FILLER_57_334 ();
 sg13g2_fill_2 FILLER_57_340 ();
 sg13g2_fill_1 FILLER_57_342 ();
 sg13g2_fill_8 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_370 ();
 sg13g2_fill_8 FILLER_57_391 ();
 sg13g2_fill_8 FILLER_57_399 ();
 sg13g2_fill_8 FILLER_57_407 ();
 sg13g2_fill_4 FILLER_57_415 ();
 sg13g2_fill_2 FILLER_57_419 ();
 sg13g2_fill_8 FILLER_57_429 ();
 sg13g2_fill_4 FILLER_57_437 ();
 sg13g2_fill_8 FILLER_57_467 ();
 sg13g2_fill_1 FILLER_57_475 ();
 sg13g2_fill_4 FILLER_57_502 ();
 sg13g2_fill_1 FILLER_57_506 ();
 sg13g2_fill_2 FILLER_57_517 ();
 sg13g2_fill_1 FILLER_57_519 ();
 sg13g2_fill_8 FILLER_57_536 ();
 sg13g2_fill_8 FILLER_57_544 ();
 sg13g2_fill_4 FILLER_57_552 ();
 sg13g2_fill_1 FILLER_57_556 ();
 sg13g2_fill_8 FILLER_57_600 ();
 sg13g2_fill_2 FILLER_57_608 ();
 sg13g2_fill_1 FILLER_57_610 ();
 sg13g2_fill_8 FILLER_57_619 ();
 sg13g2_fill_8 FILLER_57_627 ();
 sg13g2_fill_8 FILLER_57_638 ();
 sg13g2_fill_4 FILLER_57_646 ();
 sg13g2_fill_1 FILLER_57_650 ();
 sg13g2_fill_8 FILLER_57_654 ();
 sg13g2_fill_1 FILLER_57_674 ();
 sg13g2_fill_4 FILLER_57_678 ();
 sg13g2_fill_4 FILLER_57_717 ();
 sg13g2_fill_2 FILLER_57_721 ();
 sg13g2_fill_4 FILLER_57_735 ();
 sg13g2_fill_2 FILLER_57_764 ();
 sg13g2_fill_1 FILLER_57_784 ();
 sg13g2_fill_4 FILLER_57_799 ();
 sg13g2_fill_1 FILLER_57_808 ();
 sg13g2_fill_2 FILLER_57_827 ();
 sg13g2_fill_8 FILLER_57_834 ();
 sg13g2_fill_8 FILLER_57_848 ();
 sg13g2_fill_8 FILLER_57_856 ();
 sg13g2_fill_8 FILLER_57_876 ();
 sg13g2_fill_2 FILLER_57_884 ();
 sg13g2_fill_1 FILLER_57_907 ();
 sg13g2_fill_1 FILLER_57_913 ();
 sg13g2_fill_2 FILLER_57_930 ();
 sg13g2_fill_1 FILLER_57_946 ();
 sg13g2_fill_8 FILLER_57_1004 ();
 sg13g2_fill_4 FILLER_57_1012 ();
 sg13g2_fill_2 FILLER_57_1016 ();
 sg13g2_fill_1 FILLER_57_1018 ();
 sg13g2_fill_8 FILLER_57_1024 ();
 sg13g2_fill_4 FILLER_57_1032 ();
 sg13g2_fill_1 FILLER_57_1036 ();
 sg13g2_fill_1 FILLER_57_1053 ();
 sg13g2_fill_4 FILLER_57_1068 ();
 sg13g2_fill_2 FILLER_57_1072 ();
 sg13g2_fill_1 FILLER_57_1095 ();
 sg13g2_fill_4 FILLER_57_1111 ();
 sg13g2_fill_2 FILLER_57_1134 ();
 sg13g2_fill_1 FILLER_57_1136 ();
 sg13g2_fill_8 FILLER_57_1150 ();
 sg13g2_fill_2 FILLER_57_1166 ();
 sg13g2_fill_2 FILLER_57_1181 ();
 sg13g2_fill_1 FILLER_57_1183 ();
 sg13g2_fill_1 FILLER_57_1192 ();
 sg13g2_fill_4 FILLER_57_1201 ();
 sg13g2_fill_4 FILLER_57_1226 ();
 sg13g2_fill_2 FILLER_57_1251 ();
 sg13g2_fill_2 FILLER_57_1258 ();
 sg13g2_fill_1 FILLER_57_1260 ();
 sg13g2_fill_8 FILLER_57_1266 ();
 sg13g2_fill_2 FILLER_57_1274 ();
 sg13g2_fill_1 FILLER_57_1276 ();
 sg13g2_fill_2 FILLER_57_1298 ();
 sg13g2_fill_8 FILLER_57_1305 ();
 sg13g2_fill_1 FILLER_57_1319 ();
 sg13g2_fill_2 FILLER_57_1353 ();
 sg13g2_fill_1 FILLER_57_1363 ();
 sg13g2_fill_2 FILLER_57_1391 ();
 sg13g2_fill_8 FILLER_57_1423 ();
 sg13g2_fill_8 FILLER_57_1431 ();
 sg13g2_fill_8 FILLER_57_1439 ();
 sg13g2_fill_8 FILLER_57_1447 ();
 sg13g2_fill_1 FILLER_57_1455 ();
 sg13g2_fill_8 FILLER_57_1469 ();
 sg13g2_fill_2 FILLER_57_1537 ();
 sg13g2_fill_2 FILLER_57_1559 ();
 sg13g2_fill_1 FILLER_57_1591 ();
 sg13g2_fill_8 FILLER_58_0 ();
 sg13g2_fill_8 FILLER_58_8 ();
 sg13g2_fill_8 FILLER_58_16 ();
 sg13g2_fill_4 FILLER_58_24 ();
 sg13g2_fill_2 FILLER_58_28 ();
 sg13g2_fill_1 FILLER_58_30 ();
 sg13g2_fill_2 FILLER_58_41 ();
 sg13g2_fill_1 FILLER_58_43 ();
 sg13g2_fill_8 FILLER_58_54 ();
 sg13g2_fill_2 FILLER_58_62 ();
 sg13g2_fill_2 FILLER_58_116 ();
 sg13g2_fill_8 FILLER_58_128 ();
 sg13g2_fill_8 FILLER_58_136 ();
 sg13g2_fill_8 FILLER_58_154 ();
 sg13g2_fill_4 FILLER_58_162 ();
 sg13g2_fill_2 FILLER_58_166 ();
 sg13g2_fill_2 FILLER_58_176 ();
 sg13g2_fill_1 FILLER_58_178 ();
 sg13g2_fill_8 FILLER_58_205 ();
 sg13g2_fill_2 FILLER_58_213 ();
 sg13g2_fill_1 FILLER_58_215 ();
 sg13g2_fill_2 FILLER_58_226 ();
 sg13g2_fill_1 FILLER_58_228 ();
 sg13g2_fill_2 FILLER_58_282 ();
 sg13g2_fill_4 FILLER_58_305 ();
 sg13g2_fill_2 FILLER_58_309 ();
 sg13g2_fill_8 FILLER_58_321 ();
 sg13g2_fill_8 FILLER_58_374 ();
 sg13g2_fill_8 FILLER_58_418 ();
 sg13g2_fill_8 FILLER_58_426 ();
 sg13g2_fill_2 FILLER_58_434 ();
 sg13g2_fill_8 FILLER_58_451 ();
 sg13g2_fill_8 FILLER_58_459 ();
 sg13g2_fill_4 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_471 ();
 sg13g2_fill_8 FILLER_58_482 ();
 sg13g2_fill_8 FILLER_58_490 ();
 sg13g2_fill_2 FILLER_58_498 ();
 sg13g2_fill_8 FILLER_58_506 ();
 sg13g2_fill_4 FILLER_58_514 ();
 sg13g2_fill_4 FILLER_58_524 ();
 sg13g2_fill_4 FILLER_58_538 ();
 sg13g2_fill_2 FILLER_58_542 ();
 sg13g2_fill_1 FILLER_58_544 ();
 sg13g2_fill_1 FILLER_58_564 ();
 sg13g2_fill_8 FILLER_58_575 ();
 sg13g2_fill_1 FILLER_58_583 ();
 sg13g2_fill_8 FILLER_58_614 ();
 sg13g2_fill_2 FILLER_58_622 ();
 sg13g2_fill_1 FILLER_58_624 ();
 sg13g2_fill_8 FILLER_58_649 ();
 sg13g2_fill_2 FILLER_58_671 ();
 sg13g2_fill_2 FILLER_58_699 ();
 sg13g2_fill_1 FILLER_58_701 ();
 sg13g2_fill_2 FILLER_58_737 ();
 sg13g2_fill_2 FILLER_58_764 ();
 sg13g2_fill_2 FILLER_58_774 ();
 sg13g2_fill_2 FILLER_58_806 ();
 sg13g2_fill_1 FILLER_58_808 ();
 sg13g2_fill_1 FILLER_58_822 ();
 sg13g2_fill_4 FILLER_58_828 ();
 sg13g2_fill_1 FILLER_58_832 ();
 sg13g2_fill_8 FILLER_58_837 ();
 sg13g2_fill_4 FILLER_58_845 ();
 sg13g2_fill_2 FILLER_58_849 ();
 sg13g2_fill_8 FILLER_58_857 ();
 sg13g2_fill_4 FILLER_58_865 ();
 sg13g2_fill_2 FILLER_58_869 ();
 sg13g2_fill_2 FILLER_58_899 ();
 sg13g2_fill_4 FILLER_58_944 ();
 sg13g2_fill_1 FILLER_58_948 ();
 sg13g2_fill_1 FILLER_58_957 ();
 sg13g2_fill_4 FILLER_58_963 ();
 sg13g2_fill_1 FILLER_58_967 ();
 sg13g2_fill_2 FILLER_58_972 ();
 sg13g2_fill_1 FILLER_58_974 ();
 sg13g2_fill_8 FILLER_58_983 ();
 sg13g2_fill_1 FILLER_58_1001 ();
 sg13g2_fill_1 FILLER_58_1007 ();
 sg13g2_fill_2 FILLER_58_1021 ();
 sg13g2_fill_1 FILLER_58_1023 ();
 sg13g2_fill_8 FILLER_58_1032 ();
 sg13g2_fill_8 FILLER_58_1040 ();
 sg13g2_fill_8 FILLER_58_1048 ();
 sg13g2_fill_4 FILLER_58_1056 ();
 sg13g2_fill_2 FILLER_58_1060 ();
 sg13g2_fill_1 FILLER_58_1062 ();
 sg13g2_fill_2 FILLER_58_1080 ();
 sg13g2_fill_8 FILLER_58_1087 ();
 sg13g2_fill_2 FILLER_58_1095 ();
 sg13g2_fill_8 FILLER_58_1110 ();
 sg13g2_fill_8 FILLER_58_1118 ();
 sg13g2_fill_1 FILLER_58_1126 ();
 sg13g2_fill_4 FILLER_58_1135 ();
 sg13g2_fill_8 FILLER_58_1147 ();
 sg13g2_fill_8 FILLER_58_1155 ();
 sg13g2_fill_4 FILLER_58_1163 ();
 sg13g2_fill_8 FILLER_58_1171 ();
 sg13g2_fill_4 FILLER_58_1179 ();
 sg13g2_fill_1 FILLER_58_1183 ();
 sg13g2_fill_1 FILLER_58_1192 ();
 sg13g2_fill_8 FILLER_58_1214 ();
 sg13g2_fill_2 FILLER_58_1222 ();
 sg13g2_fill_4 FILLER_58_1253 ();
 sg13g2_fill_8 FILLER_58_1265 ();
 sg13g2_fill_1 FILLER_58_1273 ();
 sg13g2_fill_2 FILLER_58_1291 ();
 sg13g2_fill_1 FILLER_58_1293 ();
 sg13g2_fill_8 FILLER_58_1304 ();
 sg13g2_fill_2 FILLER_58_1312 ();
 sg13g2_fill_1 FILLER_58_1341 ();
 sg13g2_fill_2 FILLER_58_1374 ();
 sg13g2_fill_1 FILLER_58_1396 ();
 sg13g2_fill_8 FILLER_58_1403 ();
 sg13g2_fill_4 FILLER_58_1411 ();
 sg13g2_fill_1 FILLER_58_1415 ();
 sg13g2_fill_4 FILLER_58_1479 ();
 sg13g2_fill_2 FILLER_58_1483 ();
 sg13g2_fill_1 FILLER_58_1485 ();
 sg13g2_fill_8 FILLER_58_1489 ();
 sg13g2_fill_8 FILLER_58_1497 ();
 sg13g2_fill_8 FILLER_58_1505 ();
 sg13g2_fill_2 FILLER_58_1513 ();
 sg13g2_fill_1 FILLER_58_1515 ();
 sg13g2_fill_1 FILLER_58_1546 ();
 sg13g2_fill_8 FILLER_58_1557 ();
 sg13g2_fill_8 FILLER_58_1565 ();
 sg13g2_fill_8 FILLER_58_1573 ();
 sg13g2_fill_8 FILLER_58_1581 ();
 sg13g2_fill_2 FILLER_58_1589 ();
 sg13g2_fill_1 FILLER_58_1591 ();
 sg13g2_fill_8 FILLER_59_0 ();
 sg13g2_fill_4 FILLER_59_8 ();
 sg13g2_fill_8 FILLER_59_38 ();
 sg13g2_fill_1 FILLER_59_46 ();
 sg13g2_fill_4 FILLER_59_73 ();
 sg13g2_fill_2 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_102 ();
 sg13g2_fill_1 FILLER_59_104 ();
 sg13g2_fill_8 FILLER_59_110 ();
 sg13g2_fill_2 FILLER_59_118 ();
 sg13g2_fill_4 FILLER_59_141 ();
 sg13g2_fill_1 FILLER_59_145 ();
 sg13g2_fill_4 FILLER_59_172 ();
 sg13g2_fill_2 FILLER_59_176 ();
 sg13g2_fill_1 FILLER_59_178 ();
 sg13g2_fill_2 FILLER_59_197 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_fill_4 FILLER_59_216 ();
 sg13g2_fill_8 FILLER_59_225 ();
 sg13g2_fill_4 FILLER_59_233 ();
 sg13g2_fill_1 FILLER_59_237 ();
 sg13g2_fill_4 FILLER_59_264 ();
 sg13g2_fill_2 FILLER_59_268 ();
 sg13g2_fill_8 FILLER_59_296 ();
 sg13g2_fill_8 FILLER_59_304 ();
 sg13g2_fill_4 FILLER_59_348 ();
 sg13g2_fill_1 FILLER_59_352 ();
 sg13g2_fill_8 FILLER_59_369 ();
 sg13g2_fill_8 FILLER_59_384 ();
 sg13g2_fill_4 FILLER_59_392 ();
 sg13g2_fill_4 FILLER_59_432 ();
 sg13g2_fill_1 FILLER_59_436 ();
 sg13g2_fill_8 FILLER_59_473 ();
 sg13g2_fill_2 FILLER_59_481 ();
 sg13g2_fill_1 FILLER_59_483 ();
 sg13g2_fill_4 FILLER_59_510 ();
 sg13g2_fill_1 FILLER_59_514 ();
 sg13g2_fill_1 FILLER_59_524 ();
 sg13g2_fill_8 FILLER_59_544 ();
 sg13g2_fill_4 FILLER_59_552 ();
 sg13g2_fill_8 FILLER_59_592 ();
 sg13g2_fill_4 FILLER_59_600 ();
 sg13g2_fill_1 FILLER_59_604 ();
 sg13g2_fill_2 FILLER_59_615 ();
 sg13g2_fill_2 FILLER_59_634 ();
 sg13g2_fill_2 FILLER_59_682 ();
 sg13g2_fill_1 FILLER_59_684 ();
 sg13g2_fill_1 FILLER_59_727 ();
 sg13g2_fill_2 FILLER_59_736 ();
 sg13g2_fill_1 FILLER_59_738 ();
 sg13g2_fill_1 FILLER_59_775 ();
 sg13g2_fill_4 FILLER_59_788 ();
 sg13g2_fill_1 FILLER_59_792 ();
 sg13g2_fill_8 FILLER_59_799 ();
 sg13g2_fill_1 FILLER_59_807 ();
 sg13g2_fill_8 FILLER_59_840 ();
 sg13g2_fill_4 FILLER_59_875 ();
 sg13g2_fill_2 FILLER_59_879 ();
 sg13g2_fill_1 FILLER_59_881 ();
 sg13g2_fill_8 FILLER_59_887 ();
 sg13g2_fill_1 FILLER_59_895 ();
 sg13g2_fill_8 FILLER_59_904 ();
 sg13g2_fill_2 FILLER_59_912 ();
 sg13g2_fill_4 FILLER_59_922 ();
 sg13g2_fill_2 FILLER_59_926 ();
 sg13g2_fill_8 FILLER_59_932 ();
 sg13g2_fill_8 FILLER_59_948 ();
 sg13g2_fill_8 FILLER_59_956 ();
 sg13g2_fill_4 FILLER_59_964 ();
 sg13g2_fill_2 FILLER_59_968 ();
 sg13g2_fill_1 FILLER_59_970 ();
 sg13g2_fill_4 FILLER_59_997 ();
 sg13g2_fill_2 FILLER_59_1001 ();
 sg13g2_fill_8 FILLER_59_1011 ();
 sg13g2_fill_4 FILLER_59_1019 ();
 sg13g2_fill_2 FILLER_59_1023 ();
 sg13g2_fill_1 FILLER_59_1025 ();
 sg13g2_fill_8 FILLER_59_1039 ();
 sg13g2_fill_4 FILLER_59_1047 ();
 sg13g2_fill_4 FILLER_59_1060 ();
 sg13g2_fill_4 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1075 ();
 sg13g2_fill_1 FILLER_59_1077 ();
 sg13g2_fill_8 FILLER_59_1086 ();
 sg13g2_fill_8 FILLER_59_1094 ();
 sg13g2_fill_4 FILLER_59_1102 ();
 sg13g2_fill_2 FILLER_59_1106 ();
 sg13g2_fill_4 FILLER_59_1138 ();
 sg13g2_fill_8 FILLER_59_1146 ();
 sg13g2_fill_8 FILLER_59_1154 ();
 sg13g2_fill_8 FILLER_59_1183 ();
 sg13g2_fill_8 FILLER_59_1191 ();
 sg13g2_fill_8 FILLER_59_1199 ();
 sg13g2_fill_8 FILLER_59_1207 ();
 sg13g2_fill_2 FILLER_59_1215 ();
 sg13g2_fill_1 FILLER_59_1217 ();
 sg13g2_fill_8 FILLER_59_1230 ();
 sg13g2_fill_8 FILLER_59_1238 ();
 sg13g2_fill_8 FILLER_59_1246 ();
 sg13g2_fill_4 FILLER_59_1254 ();
 sg13g2_fill_2 FILLER_59_1258 ();
 sg13g2_fill_4 FILLER_59_1266 ();
 sg13g2_fill_1 FILLER_59_1270 ();
 sg13g2_fill_8 FILLER_59_1287 ();
 sg13g2_fill_4 FILLER_59_1295 ();
 sg13g2_fill_4 FILLER_59_1303 ();
 sg13g2_fill_2 FILLER_59_1307 ();
 sg13g2_fill_4 FILLER_59_1313 ();
 sg13g2_fill_2 FILLER_59_1317 ();
 sg13g2_fill_1 FILLER_59_1319 ();
 sg13g2_fill_8 FILLER_59_1326 ();
 sg13g2_fill_2 FILLER_59_1334 ();
 sg13g2_fill_2 FILLER_59_1340 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_fill_2 FILLER_59_1383 ();
 sg13g2_fill_1 FILLER_59_1390 ();
 sg13g2_fill_8 FILLER_59_1397 ();
 sg13g2_fill_1 FILLER_59_1405 ();
 sg13g2_fill_8 FILLER_59_1424 ();
 sg13g2_fill_4 FILLER_59_1432 ();
 sg13g2_fill_2 FILLER_59_1436 ();
 sg13g2_fill_8 FILLER_59_1448 ();
 sg13g2_fill_8 FILLER_59_1456 ();
 sg13g2_fill_8 FILLER_59_1464 ();
 sg13g2_fill_8 FILLER_59_1472 ();
 sg13g2_fill_4 FILLER_59_1480 ();
 sg13g2_fill_2 FILLER_59_1484 ();
 sg13g2_fill_8 FILLER_59_1494 ();
 sg13g2_fill_2 FILLER_59_1502 ();
 sg13g2_fill_8 FILLER_59_1534 ();
 sg13g2_fill_4 FILLER_59_1542 ();
 sg13g2_fill_1 FILLER_59_1546 ();
 sg13g2_fill_2 FILLER_59_1557 ();
 sg13g2_fill_2 FILLER_59_1589 ();
 sg13g2_fill_1 FILLER_59_1591 ();
 sg13g2_fill_8 FILLER_60_0 ();
 sg13g2_fill_8 FILLER_60_8 ();
 sg13g2_fill_8 FILLER_60_42 ();
 sg13g2_fill_1 FILLER_60_50 ();
 sg13g2_fill_8 FILLER_60_76 ();
 sg13g2_fill_1 FILLER_60_120 ();
 sg13g2_fill_8 FILLER_60_142 ();
 sg13g2_fill_8 FILLER_60_150 ();
 sg13g2_fill_4 FILLER_60_158 ();
 sg13g2_fill_8 FILLER_60_170 ();
 sg13g2_fill_8 FILLER_60_178 ();
 sg13g2_fill_8 FILLER_60_186 ();
 sg13g2_fill_4 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_fill_1 FILLER_60_200 ();
 sg13g2_fill_8 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_245 ();
 sg13g2_fill_8 FILLER_60_253 ();
 sg13g2_fill_8 FILLER_60_261 ();
 sg13g2_fill_8 FILLER_60_269 ();
 sg13g2_fill_8 FILLER_60_277 ();
 sg13g2_fill_8 FILLER_60_285 ();
 sg13g2_fill_8 FILLER_60_293 ();
 sg13g2_fill_8 FILLER_60_309 ();
 sg13g2_fill_8 FILLER_60_317 ();
 sg13g2_fill_8 FILLER_60_325 ();
 sg13g2_fill_8 FILLER_60_333 ();
 sg13g2_fill_1 FILLER_60_341 ();
 sg13g2_fill_4 FILLER_60_348 ();
 sg13g2_fill_1 FILLER_60_352 ();
 sg13g2_fill_8 FILLER_60_360 ();
 sg13g2_fill_4 FILLER_60_368 ();
 sg13g2_fill_4 FILLER_60_377 ();
 sg13g2_fill_1 FILLER_60_381 ();
 sg13g2_fill_8 FILLER_60_387 ();
 sg13g2_fill_8 FILLER_60_395 ();
 sg13g2_fill_8 FILLER_60_408 ();
 sg13g2_fill_4 FILLER_60_416 ();
 sg13g2_fill_4 FILLER_60_434 ();
 sg13g2_fill_2 FILLER_60_438 ();
 sg13g2_fill_1 FILLER_60_440 ();
 sg13g2_fill_2 FILLER_60_451 ();
 sg13g2_fill_8 FILLER_60_494 ();
 sg13g2_fill_8 FILLER_60_502 ();
 sg13g2_fill_2 FILLER_60_510 ();
 sg13g2_fill_1 FILLER_60_512 ();
 sg13g2_fill_4 FILLER_60_528 ();
 sg13g2_fill_1 FILLER_60_532 ();
 sg13g2_fill_8 FILLER_60_538 ();
 sg13g2_fill_4 FILLER_60_546 ();
 sg13g2_fill_1 FILLER_60_550 ();
 sg13g2_fill_8 FILLER_60_587 ();
 sg13g2_fill_8 FILLER_60_595 ();
 sg13g2_fill_4 FILLER_60_603 ();
 sg13g2_fill_1 FILLER_60_607 ();
 sg13g2_fill_2 FILLER_60_619 ();
 sg13g2_fill_1 FILLER_60_621 ();
 sg13g2_fill_8 FILLER_60_696 ();
 sg13g2_fill_8 FILLER_60_704 ();
 sg13g2_fill_4 FILLER_60_712 ();
 sg13g2_fill_2 FILLER_60_716 ();
 sg13g2_fill_2 FILLER_60_742 ();
 sg13g2_fill_1 FILLER_60_750 ();
 sg13g2_fill_1 FILLER_60_756 ();
 sg13g2_fill_2 FILLER_60_792 ();
 sg13g2_fill_8 FILLER_60_799 ();
 sg13g2_fill_4 FILLER_60_820 ();
 sg13g2_fill_2 FILLER_60_824 ();
 sg13g2_fill_2 FILLER_60_829 ();
 sg13g2_fill_1 FILLER_60_831 ();
 sg13g2_fill_8 FILLER_60_868 ();
 sg13g2_fill_4 FILLER_60_876 ();
 sg13g2_fill_2 FILLER_60_880 ();
 sg13g2_fill_4 FILLER_60_903 ();
 sg13g2_fill_8 FILLER_60_911 ();
 sg13g2_fill_8 FILLER_60_919 ();
 sg13g2_fill_2 FILLER_60_927 ();
 sg13g2_fill_8 FILLER_60_934 ();
 sg13g2_fill_2 FILLER_60_942 ();
 sg13g2_fill_4 FILLER_60_972 ();
 sg13g2_fill_2 FILLER_60_976 ();
 sg13g2_fill_4 FILLER_60_982 ();
 sg13g2_fill_4 FILLER_60_995 ();
 sg13g2_fill_1 FILLER_60_1007 ();
 sg13g2_fill_4 FILLER_60_1019 ();
 sg13g2_fill_1 FILLER_60_1023 ();
 sg13g2_fill_1 FILLER_60_1047 ();
 sg13g2_fill_4 FILLER_60_1079 ();
 sg13g2_fill_1 FILLER_60_1083 ();
 sg13g2_fill_4 FILLER_60_1089 ();
 sg13g2_fill_8 FILLER_60_1114 ();
 sg13g2_fill_8 FILLER_60_1122 ();
 sg13g2_fill_8 FILLER_60_1172 ();
 sg13g2_fill_2 FILLER_60_1188 ();
 sg13g2_fill_1 FILLER_60_1190 ();
 sg13g2_fill_4 FILLER_60_1212 ();
 sg13g2_fill_1 FILLER_60_1216 ();
 sg13g2_fill_4 FILLER_60_1238 ();
 sg13g2_fill_2 FILLER_60_1242 ();
 sg13g2_fill_4 FILLER_60_1295 ();
 sg13g2_fill_2 FILLER_60_1307 ();
 sg13g2_fill_1 FILLER_60_1309 ();
 sg13g2_fill_1 FILLER_60_1321 ();
 sg13g2_fill_8 FILLER_60_1337 ();
 sg13g2_fill_4 FILLER_60_1345 ();
 sg13g2_fill_2 FILLER_60_1349 ();
 sg13g2_fill_1 FILLER_60_1351 ();
 sg13g2_fill_1 FILLER_60_1386 ();
 sg13g2_fill_8 FILLER_60_1397 ();
 sg13g2_fill_2 FILLER_60_1405 ();
 sg13g2_fill_1 FILLER_60_1407 ();
 sg13g2_fill_8 FILLER_60_1412 ();
 sg13g2_fill_8 FILLER_60_1420 ();
 sg13g2_fill_8 FILLER_60_1428 ();
 sg13g2_fill_8 FILLER_60_1436 ();
 sg13g2_fill_8 FILLER_60_1444 ();
 sg13g2_fill_4 FILLER_60_1462 ();
 sg13g2_fill_1 FILLER_60_1466 ();
 sg13g2_fill_8 FILLER_60_1517 ();
 sg13g2_fill_8 FILLER_60_1525 ();
 sg13g2_fill_1 FILLER_60_1533 ();
 sg13g2_fill_2 FILLER_60_1589 ();
 sg13g2_fill_1 FILLER_60_1591 ();
 sg13g2_fill_8 FILLER_61_0 ();
 sg13g2_fill_8 FILLER_61_8 ();
 sg13g2_fill_8 FILLER_61_16 ();
 sg13g2_fill_4 FILLER_61_24 ();
 sg13g2_fill_2 FILLER_61_28 ();
 sg13g2_fill_1 FILLER_61_30 ();
 sg13g2_fill_2 FILLER_61_41 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_fill_8 FILLER_61_80 ();
 sg13g2_fill_8 FILLER_61_88 ();
 sg13g2_fill_8 FILLER_61_96 ();
 sg13g2_fill_8 FILLER_61_104 ();
 sg13g2_fill_8 FILLER_61_112 ();
 sg13g2_fill_8 FILLER_61_120 ();
 sg13g2_fill_8 FILLER_61_128 ();
 sg13g2_fill_8 FILLER_61_136 ();
 sg13g2_fill_2 FILLER_61_144 ();
 sg13g2_fill_8 FILLER_61_188 ();
 sg13g2_fill_8 FILLER_61_196 ();
 sg13g2_fill_1 FILLER_61_204 ();
 sg13g2_fill_8 FILLER_61_213 ();
 sg13g2_fill_8 FILLER_61_221 ();
 sg13g2_fill_4 FILLER_61_229 ();
 sg13g2_fill_8 FILLER_61_243 ();
 sg13g2_fill_1 FILLER_61_251 ();
 sg13g2_fill_8 FILLER_61_273 ();
 sg13g2_fill_8 FILLER_61_289 ();
 sg13g2_fill_8 FILLER_61_297 ();
 sg13g2_fill_2 FILLER_61_346 ();
 sg13g2_fill_1 FILLER_61_348 ();
 sg13g2_fill_4 FILLER_61_357 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_fill_2 FILLER_61_379 ();
 sg13g2_fill_2 FILLER_61_438 ();
 sg13g2_fill_1 FILLER_61_450 ();
 sg13g2_fill_1 FILLER_61_456 ();
 sg13g2_fill_2 FILLER_61_473 ();
 sg13g2_fill_4 FILLER_61_485 ();
 sg13g2_fill_2 FILLER_61_489 ();
 sg13g2_fill_1 FILLER_61_491 ();
 sg13g2_fill_8 FILLER_61_512 ();
 sg13g2_fill_8 FILLER_61_520 ();
 sg13g2_fill_8 FILLER_61_528 ();
 sg13g2_fill_2 FILLER_61_536 ();
 sg13g2_fill_2 FILLER_61_547 ();
 sg13g2_fill_1 FILLER_61_549 ();
 sg13g2_fill_8 FILLER_61_556 ();
 sg13g2_fill_8 FILLER_61_564 ();
 sg13g2_fill_8 FILLER_61_572 ();
 sg13g2_fill_8 FILLER_61_580 ();
 sg13g2_fill_4 FILLER_61_588 ();
 sg13g2_fill_2 FILLER_61_617 ();
 sg13g2_fill_1 FILLER_61_656 ();
 sg13g2_fill_8 FILLER_61_697 ();
 sg13g2_fill_8 FILLER_61_705 ();
 sg13g2_fill_4 FILLER_61_713 ();
 sg13g2_fill_1 FILLER_61_732 ();
 sg13g2_fill_1 FILLER_61_759 ();
 sg13g2_fill_1 FILLER_61_772 ();
 sg13g2_fill_2 FILLER_61_783 ();
 sg13g2_fill_1 FILLER_61_795 ();
 sg13g2_fill_8 FILLER_61_799 ();
 sg13g2_fill_2 FILLER_61_807 ();
 sg13g2_fill_8 FILLER_61_841 ();
 sg13g2_fill_8 FILLER_61_849 ();
 sg13g2_fill_1 FILLER_61_857 ();
 sg13g2_fill_8 FILLER_61_868 ();
 sg13g2_fill_8 FILLER_61_876 ();
 sg13g2_fill_8 FILLER_61_888 ();
 sg13g2_fill_1 FILLER_61_896 ();
 sg13g2_fill_2 FILLER_61_901 ();
 sg13g2_fill_4 FILLER_61_923 ();
 sg13g2_fill_8 FILLER_61_961 ();
 sg13g2_fill_2 FILLER_61_969 ();
 sg13g2_fill_1 FILLER_61_971 ();
 sg13g2_fill_2 FILLER_61_977 ();
 sg13g2_fill_8 FILLER_61_988 ();
 sg13g2_fill_8 FILLER_61_996 ();
 sg13g2_fill_4 FILLER_61_1004 ();
 sg13g2_fill_4 FILLER_61_1015 ();
 sg13g2_fill_2 FILLER_61_1019 ();
 sg13g2_fill_1 FILLER_61_1021 ();
 sg13g2_fill_8 FILLER_61_1035 ();
 sg13g2_fill_8 FILLER_61_1043 ();
 sg13g2_fill_1 FILLER_61_1051 ();
 sg13g2_fill_2 FILLER_61_1098 ();
 sg13g2_fill_1 FILLER_61_1100 ();
 sg13g2_fill_8 FILLER_61_1122 ();
 sg13g2_fill_8 FILLER_61_1130 ();
 sg13g2_fill_8 FILLER_61_1138 ();
 sg13g2_fill_4 FILLER_61_1146 ();
 sg13g2_fill_2 FILLER_61_1150 ();
 sg13g2_fill_1 FILLER_61_1152 ();
 sg13g2_fill_8 FILLER_61_1174 ();
 sg13g2_fill_4 FILLER_61_1190 ();
 sg13g2_fill_1 FILLER_61_1194 ();
 sg13g2_fill_8 FILLER_61_1237 ();
 sg13g2_fill_2 FILLER_61_1245 ();
 sg13g2_fill_1 FILLER_61_1247 ();
 sg13g2_fill_2 FILLER_61_1269 ();
 sg13g2_fill_1 FILLER_61_1271 ();
 sg13g2_fill_4 FILLER_61_1277 ();
 sg13g2_fill_1 FILLER_61_1297 ();
 sg13g2_fill_4 FILLER_61_1303 ();
 sg13g2_fill_2 FILLER_61_1307 ();
 sg13g2_fill_1 FILLER_61_1309 ();
 sg13g2_fill_2 FILLER_61_1328 ();
 sg13g2_fill_1 FILLER_61_1336 ();
 sg13g2_fill_4 FILLER_61_1354 ();
 sg13g2_fill_2 FILLER_61_1358 ();
 sg13g2_fill_8 FILLER_61_1373 ();
 sg13g2_fill_2 FILLER_61_1381 ();
 sg13g2_fill_1 FILLER_61_1383 ();
 sg13g2_fill_8 FILLER_61_1389 ();
 sg13g2_fill_4 FILLER_61_1397 ();
 sg13g2_fill_1 FILLER_61_1401 ();
 sg13g2_fill_2 FILLER_61_1411 ();
 sg13g2_fill_1 FILLER_61_1413 ();
 sg13g2_fill_4 FILLER_61_1444 ();
 sg13g2_fill_2 FILLER_61_1448 ();
 sg13g2_fill_1 FILLER_61_1450 ();
 sg13g2_fill_8 FILLER_61_1491 ();
 sg13g2_fill_8 FILLER_61_1499 ();
 sg13g2_fill_8 FILLER_61_1507 ();
 sg13g2_fill_8 FILLER_61_1545 ();
 sg13g2_fill_2 FILLER_61_1553 ();
 sg13g2_fill_1 FILLER_61_1555 ();
 sg13g2_fill_8 FILLER_61_1564 ();
 sg13g2_fill_8 FILLER_61_1572 ();
 sg13g2_fill_8 FILLER_61_1580 ();
 sg13g2_fill_4 FILLER_61_1588 ();
 sg13g2_fill_8 FILLER_62_0 ();
 sg13g2_fill_8 FILLER_62_8 ();
 sg13g2_fill_8 FILLER_62_16 ();
 sg13g2_fill_4 FILLER_62_24 ();
 sg13g2_fill_1 FILLER_62_28 ();
 sg13g2_fill_4 FILLER_62_39 ();
 sg13g2_fill_8 FILLER_62_53 ();
 sg13g2_fill_8 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_69 ();
 sg13g2_fill_8 FILLER_62_80 ();
 sg13g2_fill_8 FILLER_62_88 ();
 sg13g2_fill_8 FILLER_62_96 ();
 sg13g2_fill_8 FILLER_62_104 ();
 sg13g2_fill_1 FILLER_62_112 ();
 sg13g2_fill_8 FILLER_62_149 ();
 sg13g2_fill_8 FILLER_62_157 ();
 sg13g2_fill_4 FILLER_62_165 ();
 sg13g2_fill_1 FILLER_62_190 ();
 sg13g2_fill_4 FILLER_62_199 ();
 sg13g2_fill_8 FILLER_62_260 ();
 sg13g2_fill_2 FILLER_62_268 ();
 sg13g2_fill_8 FILLER_62_313 ();
 sg13g2_fill_8 FILLER_62_321 ();
 sg13g2_fill_8 FILLER_62_329 ();
 sg13g2_fill_8 FILLER_62_337 ();
 sg13g2_fill_2 FILLER_62_350 ();
 sg13g2_fill_8 FILLER_62_360 ();
 sg13g2_fill_4 FILLER_62_368 ();
 sg13g2_fill_1 FILLER_62_372 ();
 sg13g2_fill_8 FILLER_62_378 ();
 sg13g2_fill_2 FILLER_62_386 ();
 sg13g2_fill_1 FILLER_62_388 ();
 sg13g2_fill_4 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_403 ();
 sg13g2_fill_8 FILLER_62_418 ();
 sg13g2_fill_4 FILLER_62_432 ();
 sg13g2_fill_4 FILLER_62_472 ();
 sg13g2_fill_2 FILLER_62_476 ();
 sg13g2_fill_1 FILLER_62_478 ();
 sg13g2_fill_8 FILLER_62_505 ();
 sg13g2_fill_2 FILLER_62_513 ();
 sg13g2_fill_1 FILLER_62_515 ();
 sg13g2_fill_8 FILLER_62_534 ();
 sg13g2_fill_4 FILLER_62_542 ();
 sg13g2_fill_8 FILLER_62_556 ();
 sg13g2_fill_8 FILLER_62_564 ();
 sg13g2_fill_8 FILLER_62_572 ();
 sg13g2_fill_1 FILLER_62_580 ();
 sg13g2_fill_4 FILLER_62_620 ();
 sg13g2_fill_2 FILLER_62_624 ();
 sg13g2_fill_1 FILLER_62_626 ();
 sg13g2_fill_8 FILLER_62_630 ();
 sg13g2_fill_4 FILLER_62_638 ();
 sg13g2_fill_1 FILLER_62_642 ();
 sg13g2_fill_8 FILLER_62_687 ();
 sg13g2_fill_2 FILLER_62_695 ();
 sg13g2_fill_1 FILLER_62_697 ();
 sg13g2_fill_2 FILLER_62_745 ();
 sg13g2_fill_2 FILLER_62_788 ();
 sg13g2_fill_2 FILLER_62_796 ();
 sg13g2_fill_1 FILLER_62_810 ();
 sg13g2_fill_1 FILLER_62_832 ();
 sg13g2_fill_1 FILLER_62_845 ();
 sg13g2_fill_8 FILLER_62_851 ();
 sg13g2_fill_4 FILLER_62_859 ();
 sg13g2_fill_1 FILLER_62_863 ();
 sg13g2_fill_2 FILLER_62_893 ();
 sg13g2_fill_1 FILLER_62_917 ();
 sg13g2_fill_1 FILLER_62_934 ();
 sg13g2_fill_8 FILLER_62_955 ();
 sg13g2_fill_8 FILLER_62_963 ();
 sg13g2_fill_4 FILLER_62_971 ();
 sg13g2_fill_1 FILLER_62_975 ();
 sg13g2_fill_2 FILLER_62_982 ();
 sg13g2_fill_8 FILLER_62_1044 ();
 sg13g2_fill_8 FILLER_62_1052 ();
 sg13g2_fill_8 FILLER_62_1060 ();
 sg13g2_fill_2 FILLER_62_1068 ();
 sg13g2_fill_1 FILLER_62_1070 ();
 sg13g2_fill_8 FILLER_62_1077 ();
 sg13g2_fill_4 FILLER_62_1085 ();
 sg13g2_fill_2 FILLER_62_1089 ();
 sg13g2_fill_8 FILLER_62_1095 ();
 sg13g2_fill_2 FILLER_62_1103 ();
 sg13g2_fill_8 FILLER_62_1110 ();
 sg13g2_fill_4 FILLER_62_1118 ();
 sg13g2_fill_4 FILLER_62_1142 ();
 sg13g2_fill_2 FILLER_62_1156 ();
 sg13g2_fill_1 FILLER_62_1158 ();
 sg13g2_fill_8 FILLER_62_1169 ();
 sg13g2_fill_8 FILLER_62_1177 ();
 sg13g2_fill_8 FILLER_62_1185 ();
 sg13g2_fill_8 FILLER_62_1193 ();
 sg13g2_fill_8 FILLER_62_1214 ();
 sg13g2_fill_4 FILLER_62_1222 ();
 sg13g2_fill_8 FILLER_62_1250 ();
 sg13g2_fill_8 FILLER_62_1258 ();
 sg13g2_fill_2 FILLER_62_1266 ();
 sg13g2_fill_4 FILLER_62_1289 ();
 sg13g2_fill_4 FILLER_62_1306 ();
 sg13g2_fill_2 FILLER_62_1310 ();
 sg13g2_fill_2 FILLER_62_1317 ();
 sg13g2_fill_2 FILLER_62_1322 ();
 sg13g2_fill_8 FILLER_62_1329 ();
 sg13g2_fill_1 FILLER_62_1346 ();
 sg13g2_fill_8 FILLER_62_1367 ();
 sg13g2_fill_1 FILLER_62_1375 ();
 sg13g2_fill_2 FILLER_62_1384 ();
 sg13g2_fill_8 FILLER_62_1400 ();
 sg13g2_fill_1 FILLER_62_1408 ();
 sg13g2_fill_8 FILLER_62_1477 ();
 sg13g2_fill_8 FILLER_62_1485 ();
 sg13g2_fill_8 FILLER_62_1493 ();
 sg13g2_fill_2 FILLER_62_1501 ();
 sg13g2_fill_8 FILLER_62_1543 ();
 sg13g2_fill_2 FILLER_62_1551 ();
 sg13g2_fill_1 FILLER_62_1553 ();
 sg13g2_fill_8 FILLER_63_0 ();
 sg13g2_fill_4 FILLER_63_8 ();
 sg13g2_fill_1 FILLER_63_12 ();
 sg13g2_fill_4 FILLER_63_39 ();
 sg13g2_fill_2 FILLER_63_43 ();
 sg13g2_fill_1 FILLER_63_45 ();
 sg13g2_fill_4 FILLER_63_68 ();
 sg13g2_fill_4 FILLER_63_82 ();
 sg13g2_fill_4 FILLER_63_127 ();
 sg13g2_fill_2 FILLER_63_131 ();
 sg13g2_fill_4 FILLER_63_143 ();
 sg13g2_fill_2 FILLER_63_147 ();
 sg13g2_fill_1 FILLER_63_149 ();
 sg13g2_fill_8 FILLER_63_171 ();
 sg13g2_fill_8 FILLER_63_179 ();
 sg13g2_fill_4 FILLER_63_187 ();
 sg13g2_fill_1 FILLER_63_191 ();
 sg13g2_fill_8 FILLER_63_218 ();
 sg13g2_fill_4 FILLER_63_226 ();
 sg13g2_fill_2 FILLER_63_230 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_4 FILLER_63_289 ();
 sg13g2_fill_1 FILLER_63_293 ();
 sg13g2_fill_8 FILLER_63_310 ();
 sg13g2_fill_2 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_346 ();
 sg13g2_fill_4 FILLER_63_357 ();
 sg13g2_fill_2 FILLER_63_361 ();
 sg13g2_fill_8 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_fill_1 FILLER_63_409 ();
 sg13g2_fill_8 FILLER_63_428 ();
 sg13g2_fill_8 FILLER_63_436 ();
 sg13g2_fill_8 FILLER_63_444 ();
 sg13g2_fill_8 FILLER_63_452 ();
 sg13g2_fill_8 FILLER_63_460 ();
 sg13g2_fill_2 FILLER_63_468 ();
 sg13g2_fill_8 FILLER_63_506 ();
 sg13g2_fill_4 FILLER_63_514 ();
 sg13g2_fill_4 FILLER_63_544 ();
 sg13g2_fill_1 FILLER_63_548 ();
 sg13g2_fill_8 FILLER_63_585 ();
 sg13g2_fill_1 FILLER_63_593 ();
 sg13g2_fill_8 FILLER_63_597 ();
 sg13g2_fill_8 FILLER_63_605 ();
 sg13g2_fill_8 FILLER_63_621 ();
 sg13g2_fill_8 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_637 ();
 sg13g2_fill_8 FILLER_63_646 ();
 sg13g2_fill_2 FILLER_63_654 ();
 sg13g2_fill_1 FILLER_63_656 ();
 sg13g2_fill_2 FILLER_63_665 ();
 sg13g2_fill_1 FILLER_63_667 ();
 sg13g2_fill_1 FILLER_63_674 ();
 sg13g2_fill_8 FILLER_63_678 ();
 sg13g2_fill_1 FILLER_63_686 ();
 sg13g2_fill_8 FILLER_63_713 ();
 sg13g2_fill_4 FILLER_63_733 ();
 sg13g2_fill_2 FILLER_63_737 ();
 sg13g2_fill_2 FILLER_63_756 ();
 sg13g2_fill_8 FILLER_63_772 ();
 sg13g2_fill_8 FILLER_63_780 ();
 sg13g2_fill_2 FILLER_63_788 ();
 sg13g2_fill_1 FILLER_63_790 ();
 sg13g2_fill_1 FILLER_63_797 ();
 sg13g2_fill_2 FILLER_63_857 ();
 sg13g2_fill_1 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_865 ();
 sg13g2_fill_8 FILLER_63_871 ();
 sg13g2_fill_4 FILLER_63_879 ();
 sg13g2_fill_2 FILLER_63_883 ();
 sg13g2_fill_2 FILLER_63_889 ();
 sg13g2_fill_1 FILLER_63_891 ();
 sg13g2_fill_2 FILLER_63_905 ();
 sg13g2_fill_4 FILLER_63_944 ();
 sg13g2_fill_4 FILLER_63_957 ();
 sg13g2_fill_2 FILLER_63_971 ();
 sg13g2_fill_1 FILLER_63_973 ();
 sg13g2_fill_8 FILLER_63_980 ();
 sg13g2_fill_2 FILLER_63_993 ();
 sg13g2_fill_8 FILLER_63_1010 ();
 sg13g2_fill_8 FILLER_63_1018 ();
 sg13g2_fill_1 FILLER_63_1026 ();
 sg13g2_fill_4 FILLER_63_1040 ();
 sg13g2_fill_2 FILLER_63_1065 ();
 sg13g2_fill_1 FILLER_63_1067 ();
 sg13g2_fill_2 FILLER_63_1073 ();
 sg13g2_fill_4 FILLER_63_1080 ();
 sg13g2_fill_2 FILLER_63_1084 ();
 sg13g2_fill_4 FILLER_63_1091 ();
 sg13g2_fill_2 FILLER_63_1095 ();
 sg13g2_fill_4 FILLER_63_1114 ();
 sg13g2_fill_2 FILLER_63_1128 ();
 sg13g2_fill_1 FILLER_63_1130 ();
 sg13g2_fill_2 FILLER_63_1152 ();
 sg13g2_fill_1 FILLER_63_1154 ();
 sg13g2_fill_8 FILLER_63_1197 ();
 sg13g2_fill_8 FILLER_63_1205 ();
 sg13g2_fill_8 FILLER_63_1213 ();
 sg13g2_fill_8 FILLER_63_1221 ();
 sg13g2_fill_8 FILLER_63_1229 ();
 sg13g2_fill_4 FILLER_63_1237 ();
 sg13g2_fill_2 FILLER_63_1241 ();
 sg13g2_fill_1 FILLER_63_1243 ();
 sg13g2_fill_8 FILLER_63_1265 ();
 sg13g2_fill_8 FILLER_63_1273 ();
 sg13g2_fill_2 FILLER_63_1281 ();
 sg13g2_fill_8 FILLER_63_1288 ();
 sg13g2_fill_8 FILLER_63_1296 ();
 sg13g2_fill_4 FILLER_63_1304 ();
 sg13g2_fill_1 FILLER_63_1308 ();
 sg13g2_fill_8 FILLER_63_1330 ();
 sg13g2_fill_2 FILLER_63_1338 ();
 sg13g2_fill_1 FILLER_63_1340 ();
 sg13g2_fill_8 FILLER_63_1351 ();
 sg13g2_fill_2 FILLER_63_1364 ();
 sg13g2_fill_1 FILLER_63_1375 ();
 sg13g2_fill_2 FILLER_63_1415 ();
 sg13g2_fill_1 FILLER_63_1417 ();
 sg13g2_fill_8 FILLER_63_1423 ();
 sg13g2_fill_8 FILLER_63_1431 ();
 sg13g2_fill_8 FILLER_63_1474 ();
 sg13g2_fill_2 FILLER_63_1500 ();
 sg13g2_fill_8 FILLER_63_1512 ();
 sg13g2_fill_8 FILLER_63_1520 ();
 sg13g2_fill_8 FILLER_63_1528 ();
 sg13g2_fill_8 FILLER_63_1536 ();
 sg13g2_fill_8 FILLER_63_1544 ();
 sg13g2_fill_4 FILLER_63_1587 ();
 sg13g2_fill_1 FILLER_63_1591 ();
 sg13g2_fill_8 FILLER_64_0 ();
 sg13g2_fill_8 FILLER_64_8 ();
 sg13g2_fill_8 FILLER_64_16 ();
 sg13g2_fill_4 FILLER_64_24 ();
 sg13g2_fill_2 FILLER_64_28 ();
 sg13g2_fill_4 FILLER_64_40 ();
 sg13g2_fill_2 FILLER_64_44 ();
 sg13g2_fill_1 FILLER_64_46 ();
 sg13g2_fill_8 FILLER_64_57 ();
 sg13g2_fill_4 FILLER_64_65 ();
 sg13g2_fill_2 FILLER_64_69 ();
 sg13g2_fill_1 FILLER_64_71 ();
 sg13g2_fill_8 FILLER_64_115 ();
 sg13g2_fill_8 FILLER_64_123 ();
 sg13g2_fill_4 FILLER_64_131 ();
 sg13g2_fill_8 FILLER_64_161 ();
 sg13g2_fill_8 FILLER_64_195 ();
 sg13g2_fill_1 FILLER_64_203 ();
 sg13g2_fill_4 FILLER_64_214 ();
 sg13g2_fill_2 FILLER_64_239 ();
 sg13g2_fill_8 FILLER_64_267 ();
 sg13g2_fill_8 FILLER_64_275 ();
 sg13g2_fill_1 FILLER_64_283 ();
 sg13g2_fill_8 FILLER_64_305 ();
 sg13g2_fill_2 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_315 ();
 sg13g2_fill_8 FILLER_64_326 ();
 sg13g2_fill_8 FILLER_64_334 ();
 sg13g2_fill_4 FILLER_64_342 ();
 sg13g2_fill_1 FILLER_64_346 ();
 sg13g2_fill_4 FILLER_64_357 ();
 sg13g2_fill_2 FILLER_64_361 ();
 sg13g2_fill_1 FILLER_64_389 ();
 sg13g2_fill_4 FILLER_64_400 ();
 sg13g2_fill_2 FILLER_64_404 ();
 sg13g2_fill_2 FILLER_64_426 ();
 sg13g2_fill_8 FILLER_64_454 ();
 sg13g2_fill_8 FILLER_64_467 ();
 sg13g2_fill_8 FILLER_64_475 ();
 sg13g2_fill_8 FILLER_64_483 ();
 sg13g2_fill_8 FILLER_64_491 ();
 sg13g2_fill_1 FILLER_64_499 ();
 sg13g2_fill_4 FILLER_64_518 ();
 sg13g2_fill_1 FILLER_64_522 ();
 sg13g2_fill_2 FILLER_64_539 ();
 sg13g2_fill_1 FILLER_64_541 ();
 sg13g2_fill_8 FILLER_64_652 ();
 sg13g2_fill_4 FILLER_64_660 ();
 sg13g2_fill_2 FILLER_64_664 ();
 sg13g2_fill_1 FILLER_64_666 ();
 sg13g2_fill_4 FILLER_64_686 ();
 sg13g2_fill_2 FILLER_64_690 ();
 sg13g2_fill_8 FILLER_64_739 ();
 sg13g2_fill_8 FILLER_64_747 ();
 sg13g2_fill_2 FILLER_64_755 ();
 sg13g2_fill_1 FILLER_64_757 ();
 sg13g2_fill_4 FILLER_64_767 ();
 sg13g2_fill_1 FILLER_64_771 ();
 sg13g2_fill_4 FILLER_64_775 ();
 sg13g2_fill_8 FILLER_64_785 ();
 sg13g2_fill_1 FILLER_64_793 ();
 sg13g2_fill_8 FILLER_64_799 ();
 sg13g2_fill_8 FILLER_64_829 ();
 sg13g2_fill_2 FILLER_64_844 ();
 sg13g2_fill_1 FILLER_64_846 ();
 sg13g2_fill_2 FILLER_64_864 ();
 sg13g2_fill_1 FILLER_64_866 ();
 sg13g2_fill_2 FILLER_64_884 ();
 sg13g2_fill_2 FILLER_64_901 ();
 sg13g2_fill_1 FILLER_64_942 ();
 sg13g2_fill_8 FILLER_64_974 ();
 sg13g2_fill_2 FILLER_64_982 ();
 sg13g2_fill_1 FILLER_64_984 ();
 sg13g2_fill_4 FILLER_64_990 ();
 sg13g2_fill_1 FILLER_64_1007 ();
 sg13g2_fill_4 FILLER_64_1033 ();
 sg13g2_fill_2 FILLER_64_1037 ();
 sg13g2_fill_1 FILLER_64_1039 ();
 sg13g2_fill_1 FILLER_64_1048 ();
 sg13g2_fill_8 FILLER_64_1053 ();
 sg13g2_fill_1 FILLER_64_1061 ();
 sg13g2_fill_2 FILLER_64_1099 ();
 sg13g2_fill_1 FILLER_64_1101 ();
 sg13g2_fill_8 FILLER_64_1110 ();
 sg13g2_fill_4 FILLER_64_1118 ();
 sg13g2_fill_2 FILLER_64_1122 ();
 sg13g2_fill_1 FILLER_64_1124 ();
 sg13g2_fill_4 FILLER_64_1146 ();
 sg13g2_fill_2 FILLER_64_1150 ();
 sg13g2_fill_8 FILLER_64_1162 ();
 sg13g2_fill_8 FILLER_64_1170 ();
 sg13g2_fill_1 FILLER_64_1178 ();
 sg13g2_fill_1 FILLER_64_1222 ();
 sg13g2_fill_2 FILLER_64_1248 ();
 sg13g2_fill_8 FILLER_64_1258 ();
 sg13g2_fill_2 FILLER_64_1287 ();
 sg13g2_fill_4 FILLER_64_1297 ();
 sg13g2_fill_1 FILLER_64_1301 ();
 sg13g2_fill_4 FILLER_64_1312 ();
 sg13g2_fill_1 FILLER_64_1316 ();
 sg13g2_fill_8 FILLER_64_1332 ();
 sg13g2_fill_4 FILLER_64_1340 ();
 sg13g2_fill_2 FILLER_64_1344 ();
 sg13g2_fill_1 FILLER_64_1346 ();
 sg13g2_fill_4 FILLER_64_1360 ();
 sg13g2_fill_2 FILLER_64_1364 ();
 sg13g2_fill_8 FILLER_64_1380 ();
 sg13g2_fill_4 FILLER_64_1388 ();
 sg13g2_fill_2 FILLER_64_1392 ();
 sg13g2_fill_4 FILLER_64_1454 ();
 sg13g2_fill_1 FILLER_64_1458 ();
 sg13g2_fill_4 FILLER_64_1492 ();
 sg13g2_fill_4 FILLER_64_1526 ();
 sg13g2_fill_1 FILLER_64_1530 ();
 sg13g2_fill_4 FILLER_64_1556 ();
 sg13g2_fill_2 FILLER_64_1560 ();
 sg13g2_fill_8 FILLER_64_1567 ();
 sg13g2_fill_8 FILLER_64_1575 ();
 sg13g2_fill_8 FILLER_64_1583 ();
 sg13g2_fill_1 FILLER_64_1591 ();
 sg13g2_fill_8 FILLER_65_0 ();
 sg13g2_fill_8 FILLER_65_8 ();
 sg13g2_fill_1 FILLER_65_16 ();
 sg13g2_fill_8 FILLER_65_43 ();
 sg13g2_fill_8 FILLER_65_51 ();
 sg13g2_fill_8 FILLER_65_59 ();
 sg13g2_fill_8 FILLER_65_87 ();
 sg13g2_fill_4 FILLER_65_95 ();
 sg13g2_fill_2 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_112 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_fill_8 FILLER_65_146 ();
 sg13g2_fill_2 FILLER_65_154 ();
 sg13g2_fill_1 FILLER_65_164 ();
 sg13g2_fill_2 FILLER_65_188 ();
 sg13g2_fill_1 FILLER_65_190 ();
 sg13g2_fill_8 FILLER_65_217 ();
 sg13g2_fill_8 FILLER_65_225 ();
 sg13g2_fill_4 FILLER_65_236 ();
 sg13g2_fill_1 FILLER_65_240 ();
 sg13g2_fill_8 FILLER_65_251 ();
 sg13g2_fill_2 FILLER_65_306 ();
 sg13g2_fill_1 FILLER_65_308 ();
 sg13g2_fill_2 FILLER_65_361 ();
 sg13g2_fill_1 FILLER_65_363 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_fill_1 FILLER_65_404 ();
 sg13g2_fill_1 FILLER_65_431 ();
 sg13g2_fill_2 FILLER_65_438 ();
 sg13g2_fill_4 FILLER_65_451 ();
 sg13g2_fill_8 FILLER_65_475 ();
 sg13g2_fill_8 FILLER_65_483 ();
 sg13g2_fill_2 FILLER_65_491 ();
 sg13g2_fill_2 FILLER_65_498 ();
 sg13g2_fill_4 FILLER_65_525 ();
 sg13g2_fill_1 FILLER_65_529 ();
 sg13g2_fill_2 FILLER_65_546 ();
 sg13g2_fill_8 FILLER_65_559 ();
 sg13g2_fill_8 FILLER_65_567 ();
 sg13g2_fill_8 FILLER_65_575 ();
 sg13g2_fill_8 FILLER_65_583 ();
 sg13g2_fill_8 FILLER_65_591 ();
 sg13g2_fill_8 FILLER_65_599 ();
 sg13g2_fill_8 FILLER_65_607 ();
 sg13g2_fill_1 FILLER_65_615 ();
 sg13g2_fill_8 FILLER_65_619 ();
 sg13g2_fill_8 FILLER_65_627 ();
 sg13g2_fill_2 FILLER_65_635 ();
 sg13g2_fill_1 FILLER_65_637 ();
 sg13g2_fill_2 FILLER_65_659 ();
 sg13g2_fill_8 FILLER_65_674 ();
 sg13g2_fill_4 FILLER_65_682 ();
 sg13g2_fill_1 FILLER_65_686 ();
 sg13g2_fill_4 FILLER_65_703 ();
 sg13g2_fill_1 FILLER_65_728 ();
 sg13g2_fill_4 FILLER_65_734 ();
 sg13g2_fill_2 FILLER_65_738 ();
 sg13g2_fill_1 FILLER_65_745 ();
 sg13g2_fill_2 FILLER_65_759 ();
 sg13g2_fill_1 FILLER_65_761 ();
 sg13g2_fill_2 FILLER_65_807 ();
 sg13g2_fill_2 FILLER_65_838 ();
 sg13g2_fill_4 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_858 ();
 sg13g2_fill_2 FILLER_65_867 ();
 sg13g2_fill_1 FILLER_65_869 ();
 sg13g2_fill_8 FILLER_65_876 ();
 sg13g2_fill_2 FILLER_65_923 ();
 sg13g2_fill_4 FILLER_65_975 ();
 sg13g2_fill_2 FILLER_65_979 ();
 sg13g2_fill_1 FILLER_65_981 ();
 sg13g2_fill_1 FILLER_65_1005 ();
 sg13g2_fill_8 FILLER_65_1036 ();
 sg13g2_fill_8 FILLER_65_1044 ();
 sg13g2_fill_8 FILLER_65_1052 ();
 sg13g2_fill_8 FILLER_65_1060 ();
 sg13g2_fill_8 FILLER_65_1085 ();
 sg13g2_fill_8 FILLER_65_1093 ();
 sg13g2_fill_8 FILLER_65_1101 ();
 sg13g2_fill_4 FILLER_65_1109 ();
 sg13g2_fill_1 FILLER_65_1113 ();
 sg13g2_fill_8 FILLER_65_1124 ();
 sg13g2_fill_8 FILLER_65_1132 ();
 sg13g2_fill_8 FILLER_65_1140 ();
 sg13g2_fill_4 FILLER_65_1148 ();
 sg13g2_fill_1 FILLER_65_1152 ();
 sg13g2_fill_4 FILLER_65_1161 ();
 sg13g2_fill_1 FILLER_65_1165 ();
 sg13g2_fill_1 FILLER_65_1181 ();
 sg13g2_fill_8 FILLER_65_1190 ();
 sg13g2_fill_2 FILLER_65_1198 ();
 sg13g2_fill_4 FILLER_65_1225 ();
 sg13g2_fill_2 FILLER_65_1239 ();
 sg13g2_fill_1 FILLER_65_1251 ();
 sg13g2_fill_8 FILLER_65_1262 ();
 sg13g2_fill_4 FILLER_65_1291 ();
 sg13g2_fill_2 FILLER_65_1295 ();
 sg13g2_fill_2 FILLER_65_1326 ();
 sg13g2_fill_1 FILLER_65_1328 ();
 sg13g2_fill_8 FILLER_65_1334 ();
 sg13g2_fill_1 FILLER_65_1342 ();
 sg13g2_fill_2 FILLER_65_1357 ();
 sg13g2_fill_1 FILLER_65_1359 ();
 sg13g2_fill_1 FILLER_65_1375 ();
 sg13g2_fill_2 FILLER_65_1379 ();
 sg13g2_fill_8 FILLER_65_1390 ();
 sg13g2_fill_8 FILLER_65_1401 ();
 sg13g2_fill_8 FILLER_65_1409 ();
 sg13g2_fill_8 FILLER_65_1417 ();
 sg13g2_fill_8 FILLER_65_1425 ();
 sg13g2_fill_8 FILLER_65_1433 ();
 sg13g2_fill_1 FILLER_65_1441 ();
 sg13g2_fill_8 FILLER_65_1450 ();
 sg13g2_fill_8 FILLER_65_1458 ();
 sg13g2_fill_2 FILLER_65_1466 ();
 sg13g2_fill_8 FILLER_65_1476 ();
 sg13g2_fill_2 FILLER_65_1484 ();
 sg13g2_fill_8 FILLER_65_1524 ();
 sg13g2_fill_8 FILLER_65_1532 ();
 sg13g2_fill_2 FILLER_65_1540 ();
 sg13g2_fill_8 FILLER_65_1547 ();
 sg13g2_fill_8 FILLER_65_1555 ();
 sg13g2_fill_8 FILLER_65_1571 ();
 sg13g2_fill_8 FILLER_65_1579 ();
 sg13g2_fill_4 FILLER_65_1587 ();
 sg13g2_fill_1 FILLER_65_1591 ();
 sg13g2_fill_8 FILLER_66_0 ();
 sg13g2_fill_8 FILLER_66_8 ();
 sg13g2_fill_8 FILLER_66_16 ();
 sg13g2_fill_8 FILLER_66_24 ();
 sg13g2_fill_4 FILLER_66_32 ();
 sg13g2_fill_1 FILLER_66_36 ();
 sg13g2_fill_8 FILLER_66_83 ();
 sg13g2_fill_8 FILLER_66_91 ();
 sg13g2_fill_1 FILLER_66_99 ();
 sg13g2_fill_4 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_124 ();
 sg13g2_fill_1 FILLER_66_126 ();
 sg13g2_fill_8 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_160 ();
 sg13g2_fill_4 FILLER_66_170 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_8 FILLER_66_200 ();
 sg13g2_fill_8 FILLER_66_208 ();
 sg13g2_fill_4 FILLER_66_216 ();
 sg13g2_fill_1 FILLER_66_220 ();
 sg13g2_fill_8 FILLER_66_231 ();
 sg13g2_fill_8 FILLER_66_239 ();
 sg13g2_fill_8 FILLER_66_247 ();
 sg13g2_fill_8 FILLER_66_255 ();
 sg13g2_fill_4 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_8 FILLER_66_278 ();
 sg13g2_fill_8 FILLER_66_286 ();
 sg13g2_fill_8 FILLER_66_294 ();
 sg13g2_fill_8 FILLER_66_302 ();
 sg13g2_fill_4 FILLER_66_310 ();
 sg13g2_fill_2 FILLER_66_314 ();
 sg13g2_fill_8 FILLER_66_326 ();
 sg13g2_fill_8 FILLER_66_334 ();
 sg13g2_fill_2 FILLER_66_342 ();
 sg13g2_fill_8 FILLER_66_360 ();
 sg13g2_fill_4 FILLER_66_368 ();
 sg13g2_fill_2 FILLER_66_372 ();
 sg13g2_fill_1 FILLER_66_374 ();
 sg13g2_fill_4 FILLER_66_436 ();
 sg13g2_fill_1 FILLER_66_502 ();
 sg13g2_fill_4 FILLER_66_529 ();
 sg13g2_fill_4 FILLER_66_541 ();
 sg13g2_fill_4 FILLER_66_565 ();
 sg13g2_fill_2 FILLER_66_569 ();
 sg13g2_fill_8 FILLER_66_579 ();
 sg13g2_fill_2 FILLER_66_587 ();
 sg13g2_fill_8 FILLER_66_622 ();
 sg13g2_fill_8 FILLER_66_630 ();
 sg13g2_fill_8 FILLER_66_638 ();
 sg13g2_fill_1 FILLER_66_651 ();
 sg13g2_fill_8 FILLER_66_668 ();
 sg13g2_fill_8 FILLER_66_676 ();
 sg13g2_fill_1 FILLER_66_684 ();
 sg13g2_fill_8 FILLER_66_703 ();
 sg13g2_fill_2 FILLER_66_711 ();
 sg13g2_fill_1 FILLER_66_713 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_fill_1 FILLER_66_811 ();
 sg13g2_fill_2 FILLER_66_844 ();
 sg13g2_fill_4 FILLER_66_872 ();
 sg13g2_fill_2 FILLER_66_876 ();
 sg13g2_fill_1 FILLER_66_878 ();
 sg13g2_fill_2 FILLER_66_905 ();
 sg13g2_fill_1 FILLER_66_950 ();
 sg13g2_fill_8 FILLER_66_1035 ();
 sg13g2_fill_1 FILLER_66_1043 ();
 sg13g2_fill_2 FILLER_66_1049 ();
 sg13g2_fill_1 FILLER_66_1051 ();
 sg13g2_fill_8 FILLER_66_1073 ();
 sg13g2_fill_8 FILLER_66_1089 ();
 sg13g2_fill_2 FILLER_66_1097 ();
 sg13g2_fill_2 FILLER_66_1120 ();
 sg13g2_fill_1 FILLER_66_1122 ();
 sg13g2_fill_4 FILLER_66_1136 ();
 sg13g2_fill_2 FILLER_66_1145 ();
 sg13g2_fill_1 FILLER_66_1147 ();
 sg13g2_fill_8 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1176 ();
 sg13g2_fill_1 FILLER_66_1178 ();
 sg13g2_fill_8 FILLER_66_1188 ();
 sg13g2_fill_8 FILLER_66_1206 ();
 sg13g2_fill_2 FILLER_66_1214 ();
 sg13g2_fill_1 FILLER_66_1216 ();
 sg13g2_fill_2 FILLER_66_1233 ();
 sg13g2_fill_1 FILLER_66_1235 ();
 sg13g2_fill_4 FILLER_66_1246 ();
 sg13g2_fill_1 FILLER_66_1250 ();
 sg13g2_fill_8 FILLER_66_1261 ();
 sg13g2_fill_4 FILLER_66_1290 ();
 sg13g2_fill_2 FILLER_66_1294 ();
 sg13g2_fill_1 FILLER_66_1296 ();
 sg13g2_fill_4 FILLER_66_1328 ();
 sg13g2_fill_1 FILLER_66_1340 ();
 sg13g2_fill_2 FILLER_66_1370 ();
 sg13g2_fill_4 FILLER_66_1410 ();
 sg13g2_fill_1 FILLER_66_1414 ();
 sg13g2_fill_2 FILLER_66_1425 ();
 sg13g2_fill_8 FILLER_66_1457 ();
 sg13g2_fill_8 FILLER_66_1465 ();
 sg13g2_fill_1 FILLER_66_1473 ();
 sg13g2_fill_4 FILLER_66_1504 ();
 sg13g2_fill_2 FILLER_66_1560 ();
 sg13g2_fill_8 FILLER_67_0 ();
 sg13g2_fill_8 FILLER_67_8 ();
 sg13g2_fill_8 FILLER_67_16 ();
 sg13g2_fill_2 FILLER_67_24 ();
 sg13g2_fill_8 FILLER_67_34 ();
 sg13g2_fill_8 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_50 ();
 sg13g2_fill_8 FILLER_67_108 ();
 sg13g2_fill_4 FILLER_67_137 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_fill_4 FILLER_67_194 ();
 sg13g2_fill_1 FILLER_67_198 ();
 sg13g2_fill_8 FILLER_67_251 ();
 sg13g2_fill_8 FILLER_67_259 ();
 sg13g2_fill_2 FILLER_67_267 ();
 sg13g2_fill_1 FILLER_67_269 ();
 sg13g2_fill_2 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_318 ();
 sg13g2_fill_2 FILLER_67_355 ();
 sg13g2_fill_1 FILLER_67_357 ();
 sg13g2_fill_4 FILLER_67_409 ();
 sg13g2_fill_1 FILLER_67_413 ();
 sg13g2_fill_1 FILLER_67_427 ();
 sg13g2_fill_1 FILLER_67_441 ();
 sg13g2_fill_8 FILLER_67_465 ();
 sg13g2_fill_8 FILLER_67_473 ();
 sg13g2_fill_8 FILLER_67_481 ();
 sg13g2_fill_8 FILLER_67_489 ();
 sg13g2_fill_8 FILLER_67_497 ();
 sg13g2_fill_2 FILLER_67_505 ();
 sg13g2_fill_1 FILLER_67_507 ();
 sg13g2_fill_1 FILLER_67_549 ();
 sg13g2_fill_4 FILLER_67_560 ();
 sg13g2_fill_1 FILLER_67_564 ();
 sg13g2_fill_4 FILLER_67_591 ();
 sg13g2_fill_4 FILLER_67_603 ();
 sg13g2_fill_2 FILLER_67_637 ();
 sg13g2_fill_8 FILLER_67_659 ();
 sg13g2_fill_2 FILLER_67_667 ();
 sg13g2_fill_1 FILLER_67_669 ();
 sg13g2_fill_1 FILLER_67_722 ();
 sg13g2_fill_2 FILLER_67_734 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_1 FILLER_67_778 ();
 sg13g2_fill_1 FILLER_67_834 ();
 sg13g2_fill_2 FILLER_67_890 ();
 sg13g2_fill_2 FILLER_67_898 ();
 sg13g2_fill_2 FILLER_67_906 ();
 sg13g2_fill_1 FILLER_67_922 ();
 sg13g2_fill_1 FILLER_67_958 ();
 sg13g2_fill_1 FILLER_67_988 ();
 sg13g2_fill_2 FILLER_67_1027 ();
 sg13g2_fill_1 FILLER_67_1029 ();
 sg13g2_fill_8 FILLER_67_1059 ();
 sg13g2_fill_4 FILLER_67_1067 ();
 sg13g2_fill_1 FILLER_67_1071 ();
 sg13g2_fill_2 FILLER_67_1097 ();
 sg13g2_fill_1 FILLER_67_1099 ();
 sg13g2_fill_4 FILLER_67_1105 ();
 sg13g2_fill_2 FILLER_67_1109 ();
 sg13g2_fill_2 FILLER_67_1116 ();
 sg13g2_fill_1 FILLER_67_1118 ();
 sg13g2_fill_2 FILLER_67_1133 ();
 sg13g2_fill_2 FILLER_67_1145 ();
 sg13g2_fill_1 FILLER_67_1147 ();
 sg13g2_fill_2 FILLER_67_1158 ();
 sg13g2_fill_8 FILLER_67_1200 ();
 sg13g2_fill_4 FILLER_67_1208 ();
 sg13g2_fill_1 FILLER_67_1212 ();
 sg13g2_fill_8 FILLER_67_1218 ();
 sg13g2_fill_8 FILLER_67_1226 ();
 sg13g2_fill_8 FILLER_67_1234 ();
 sg13g2_fill_8 FILLER_67_1242 ();
 sg13g2_fill_8 FILLER_67_1250 ();
 sg13g2_fill_8 FILLER_67_1258 ();
 sg13g2_fill_8 FILLER_67_1266 ();
 sg13g2_fill_8 FILLER_67_1274 ();
 sg13g2_fill_2 FILLER_67_1282 ();
 sg13g2_fill_8 FILLER_67_1294 ();
 sg13g2_fill_1 FILLER_67_1302 ();
 sg13g2_fill_8 FILLER_67_1306 ();
 sg13g2_fill_2 FILLER_67_1314 ();
 sg13g2_fill_1 FILLER_67_1316 ();
 sg13g2_fill_4 FILLER_67_1339 ();
 sg13g2_fill_2 FILLER_67_1353 ();
 sg13g2_fill_1 FILLER_67_1365 ();
 sg13g2_fill_1 FILLER_67_1405 ();
 sg13g2_fill_8 FILLER_67_1436 ();
 sg13g2_fill_1 FILLER_67_1444 ();
 sg13g2_fill_8 FILLER_67_1485 ();
 sg13g2_fill_4 FILLER_67_1493 ();
 sg13g2_fill_2 FILLER_67_1497 ();
 sg13g2_fill_8 FILLER_67_1505 ();
 sg13g2_fill_8 FILLER_67_1513 ();
 sg13g2_fill_4 FILLER_67_1521 ();
 sg13g2_fill_8 FILLER_67_1541 ();
 sg13g2_fill_4 FILLER_67_1556 ();
 sg13g2_fill_2 FILLER_67_1560 ();
 sg13g2_fill_8 FILLER_68_0 ();
 sg13g2_fill_4 FILLER_68_8 ();
 sg13g2_fill_2 FILLER_68_12 ();
 sg13g2_fill_8 FILLER_68_40 ();
 sg13g2_fill_8 FILLER_68_48 ();
 sg13g2_fill_4 FILLER_68_56 ();
 sg13g2_fill_2 FILLER_68_60 ();
 sg13g2_fill_1 FILLER_68_62 ();
 sg13g2_fill_8 FILLER_68_97 ();
 sg13g2_fill_4 FILLER_68_105 ();
 sg13g2_fill_2 FILLER_68_109 ();
 sg13g2_fill_1 FILLER_68_111 ();
 sg13g2_fill_4 FILLER_68_138 ();
 sg13g2_fill_2 FILLER_68_142 ();
 sg13g2_fill_2 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_fill_4 FILLER_68_209 ();
 sg13g2_fill_2 FILLER_68_213 ();
 sg13g2_fill_8 FILLER_68_225 ();
 sg13g2_fill_2 FILLER_68_233 ();
 sg13g2_fill_8 FILLER_68_297 ();
 sg13g2_fill_8 FILLER_68_305 ();
 sg13g2_fill_8 FILLER_68_313 ();
 sg13g2_fill_8 FILLER_68_321 ();
 sg13g2_fill_4 FILLER_68_329 ();
 sg13g2_fill_8 FILLER_68_363 ();
 sg13g2_fill_8 FILLER_68_371 ();
 sg13g2_fill_2 FILLER_68_379 ();
 sg13g2_fill_1 FILLER_68_381 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_68_422 ();
 sg13g2_fill_4 FILLER_68_453 ();
 sg13g2_fill_1 FILLER_68_457 ();
 sg13g2_fill_8 FILLER_68_468 ();
 sg13g2_fill_8 FILLER_68_512 ();
 sg13g2_fill_8 FILLER_68_520 ();
 sg13g2_fill_8 FILLER_68_528 ();
 sg13g2_fill_8 FILLER_68_536 ();
 sg13g2_fill_4 FILLER_68_544 ();
 sg13g2_fill_2 FILLER_68_548 ();
 sg13g2_fill_2 FILLER_68_560 ();
 sg13g2_fill_1 FILLER_68_588 ();
 sg13g2_fill_4 FILLER_68_597 ();
 sg13g2_fill_8 FILLER_68_630 ();
 sg13g2_fill_2 FILLER_68_638 ();
 sg13g2_fill_1 FILLER_68_640 ();
 sg13g2_fill_1 FILLER_68_646 ();
 sg13g2_fill_8 FILLER_68_659 ();
 sg13g2_fill_4 FILLER_68_667 ();
 sg13g2_fill_1 FILLER_68_671 ();
 sg13g2_fill_8 FILLER_68_684 ();
 sg13g2_fill_2 FILLER_68_692 ();
 sg13g2_fill_2 FILLER_68_703 ();
 sg13g2_fill_4 FILLER_68_735 ();
 sg13g2_fill_2 FILLER_68_739 ();
 sg13g2_fill_1 FILLER_68_741 ();
 sg13g2_fill_1 FILLER_68_789 ();
 sg13g2_fill_1 FILLER_68_821 ();
 sg13g2_fill_1 FILLER_68_847 ();
 sg13g2_fill_1 FILLER_68_863 ();
 sg13g2_fill_4 FILLER_68_869 ();
 sg13g2_fill_2 FILLER_68_873 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_fill_1 FILLER_68_911 ();
 sg13g2_fill_1 FILLER_68_934 ();
 sg13g2_fill_1 FILLER_68_951 ();
 sg13g2_fill_8 FILLER_68_1035 ();
 sg13g2_fill_1 FILLER_68_1043 ();
 sg13g2_fill_4 FILLER_68_1049 ();
 sg13g2_fill_8 FILLER_68_1071 ();
 sg13g2_fill_1 FILLER_68_1079 ();
 sg13g2_fill_2 FILLER_68_1098 ();
 sg13g2_fill_1 FILLER_68_1100 ();
 sg13g2_fill_4 FILLER_68_1111 ();
 sg13g2_fill_4 FILLER_68_1133 ();
 sg13g2_fill_2 FILLER_68_1137 ();
 sg13g2_fill_8 FILLER_68_1144 ();
 sg13g2_fill_4 FILLER_68_1152 ();
 sg13g2_fill_2 FILLER_68_1156 ();
 sg13g2_fill_2 FILLER_68_1163 ();
 sg13g2_fill_8 FILLER_68_1170 ();
 sg13g2_fill_2 FILLER_68_1178 ();
 sg13g2_fill_8 FILLER_68_1185 ();
 sg13g2_fill_2 FILLER_68_1193 ();
 sg13g2_fill_1 FILLER_68_1204 ();
 sg13g2_fill_4 FILLER_68_1210 ();
 sg13g2_fill_1 FILLER_68_1229 ();
 sg13g2_fill_8 FILLER_68_1270 ();
 sg13g2_fill_2 FILLER_68_1278 ();
 sg13g2_fill_1 FILLER_68_1280 ();
 sg13g2_fill_8 FILLER_68_1291 ();
 sg13g2_fill_1 FILLER_68_1299 ();
 sg13g2_fill_2 FILLER_68_1312 ();
 sg13g2_fill_1 FILLER_68_1322 ();
 sg13g2_fill_8 FILLER_68_1334 ();
 sg13g2_fill_8 FILLER_68_1342 ();
 sg13g2_fill_2 FILLER_68_1350 ();
 sg13g2_fill_2 FILLER_68_1364 ();
 sg13g2_fill_2 FILLER_68_1371 ();
 sg13g2_fill_1 FILLER_68_1384 ();
 sg13g2_fill_2 FILLER_68_1426 ();
 sg13g2_fill_1 FILLER_68_1449 ();
 sg13g2_fill_8 FILLER_68_1454 ();
 sg13g2_fill_4 FILLER_68_1462 ();
 sg13g2_fill_1 FILLER_68_1550 ();
 sg13g2_fill_1 FILLER_68_1591 ();
 sg13g2_fill_8 FILLER_69_0 ();
 sg13g2_fill_8 FILLER_69_8 ();
 sg13g2_fill_4 FILLER_69_16 ();
 sg13g2_fill_2 FILLER_69_20 ();
 sg13g2_fill_1 FILLER_69_22 ();
 sg13g2_fill_4 FILLER_69_59 ();
 sg13g2_fill_2 FILLER_69_63 ();
 sg13g2_fill_8 FILLER_69_126 ();
 sg13g2_fill_4 FILLER_69_134 ();
 sg13g2_fill_1 FILLER_69_138 ();
 sg13g2_fill_8 FILLER_69_149 ();
 sg13g2_fill_8 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_165 ();
 sg13g2_fill_8 FILLER_69_177 ();
 sg13g2_fill_4 FILLER_69_185 ();
 sg13g2_fill_8 FILLER_69_224 ();
 sg13g2_fill_4 FILLER_69_232 ();
 sg13g2_fill_2 FILLER_69_236 ();
 sg13g2_fill_8 FILLER_69_248 ();
 sg13g2_fill_2 FILLER_69_256 ();
 sg13g2_fill_1 FILLER_69_258 ();
 sg13g2_fill_4 FILLER_69_287 ();
 sg13g2_fill_2 FILLER_69_291 ();
 sg13g2_fill_1 FILLER_69_293 ();
 sg13g2_fill_8 FILLER_69_320 ();
 sg13g2_fill_8 FILLER_69_328 ();
 sg13g2_fill_2 FILLER_69_336 ();
 sg13g2_fill_1 FILLER_69_338 ();
 sg13g2_fill_8 FILLER_69_365 ();
 sg13g2_fill_8 FILLER_69_373 ();
 sg13g2_fill_4 FILLER_69_381 ();
 sg13g2_fill_1 FILLER_69_385 ();
 sg13g2_fill_4 FILLER_69_396 ();
 sg13g2_fill_2 FILLER_69_400 ();
 sg13g2_fill_8 FILLER_69_405 ();
 sg13g2_fill_2 FILLER_69_413 ();
 sg13g2_fill_4 FILLER_69_441 ();
 sg13g2_fill_2 FILLER_69_491 ();
 sg13g2_fill_8 FILLER_69_501 ();
 sg13g2_fill_8 FILLER_69_509 ();
 sg13g2_fill_8 FILLER_69_517 ();
 sg13g2_fill_8 FILLER_69_525 ();
 sg13g2_fill_8 FILLER_69_533 ();
 sg13g2_fill_8 FILLER_69_541 ();
 sg13g2_fill_8 FILLER_69_549 ();
 sg13g2_fill_8 FILLER_69_557 ();
 sg13g2_fill_8 FILLER_69_565 ();
 sg13g2_fill_8 FILLER_69_573 ();
 sg13g2_fill_2 FILLER_69_581 ();
 sg13g2_fill_1 FILLER_69_583 ();
 sg13g2_fill_2 FILLER_69_609 ();
 sg13g2_fill_1 FILLER_69_611 ();
 sg13g2_fill_8 FILLER_69_642 ();
 sg13g2_fill_2 FILLER_69_650 ();
 sg13g2_fill_1 FILLER_69_652 ();
 sg13g2_fill_2 FILLER_69_689 ();
 sg13g2_fill_1 FILLER_69_764 ();
 sg13g2_fill_1 FILLER_69_868 ();
 sg13g2_fill_2 FILLER_69_881 ();
 sg13g2_fill_1 FILLER_69_895 ();
 sg13g2_fill_2 FILLER_69_927 ();
 sg13g2_fill_1 FILLER_69_942 ();
 sg13g2_fill_2 FILLER_69_957 ();
 sg13g2_fill_1 FILLER_69_969 ();
 sg13g2_fill_2 FILLER_69_980 ();
 sg13g2_fill_8 FILLER_69_1036 ();
 sg13g2_fill_8 FILLER_69_1044 ();
 sg13g2_fill_4 FILLER_69_1052 ();
 sg13g2_fill_2 FILLER_69_1068 ();
 sg13g2_fill_2 FILLER_69_1076 ();
 sg13g2_fill_8 FILLER_69_1083 ();
 sg13g2_fill_8 FILLER_69_1091 ();
 sg13g2_fill_8 FILLER_69_1099 ();
 sg13g2_fill_8 FILLER_69_1129 ();
 sg13g2_fill_1 FILLER_69_1137 ();
 sg13g2_fill_8 FILLER_69_1142 ();
 sg13g2_fill_4 FILLER_69_1150 ();
 sg13g2_fill_8 FILLER_69_1159 ();
 sg13g2_fill_8 FILLER_69_1167 ();
 sg13g2_fill_4 FILLER_69_1180 ();
 sg13g2_fill_2 FILLER_69_1184 ();
 sg13g2_fill_1 FILLER_69_1186 ();
 sg13g2_fill_4 FILLER_69_1191 ();
 sg13g2_fill_4 FILLER_69_1204 ();
 sg13g2_fill_2 FILLER_69_1208 ();
 sg13g2_fill_4 FILLER_69_1257 ();
 sg13g2_fill_1 FILLER_69_1261 ();
 sg13g2_fill_8 FILLER_69_1319 ();
 sg13g2_fill_8 FILLER_69_1327 ();
 sg13g2_fill_8 FILLER_69_1335 ();
 sg13g2_fill_2 FILLER_69_1343 ();
 sg13g2_fill_1 FILLER_69_1345 ();
 sg13g2_fill_1 FILLER_69_1372 ();
 sg13g2_fill_1 FILLER_69_1406 ();
 sg13g2_fill_4 FILLER_69_1459 ();
 sg13g2_fill_2 FILLER_69_1463 ();
 sg13g2_fill_1 FILLER_69_1465 ();
 sg13g2_fill_2 FILLER_69_1476 ();
 sg13g2_fill_1 FILLER_69_1478 ();
 sg13g2_fill_8 FILLER_69_1487 ();
 sg13g2_fill_8 FILLER_69_1495 ();
 sg13g2_fill_8 FILLER_69_1503 ();
 sg13g2_fill_8 FILLER_69_1511 ();
 sg13g2_fill_8 FILLER_69_1519 ();
 sg13g2_fill_8 FILLER_69_1527 ();
 sg13g2_fill_4 FILLER_69_1535 ();
 sg13g2_fill_1 FILLER_69_1539 ();
 sg13g2_fill_4 FILLER_69_1553 ();
 sg13g2_fill_2 FILLER_69_1557 ();
 sg13g2_fill_2 FILLER_69_1589 ();
 sg13g2_fill_1 FILLER_69_1591 ();
 sg13g2_fill_8 FILLER_70_0 ();
 sg13g2_fill_8 FILLER_70_8 ();
 sg13g2_fill_8 FILLER_70_16 ();
 sg13g2_fill_2 FILLER_70_24 ();
 sg13g2_fill_1 FILLER_70_26 ();
 sg13g2_fill_8 FILLER_70_37 ();
 sg13g2_fill_4 FILLER_70_45 ();
 sg13g2_fill_4 FILLER_70_102 ();
 sg13g2_fill_8 FILLER_70_117 ();
 sg13g2_fill_4 FILLER_70_125 ();
 sg13g2_fill_8 FILLER_70_155 ();
 sg13g2_fill_4 FILLER_70_163 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_fill_4 FILLER_70_195 ();
 sg13g2_fill_8 FILLER_70_224 ();
 sg13g2_fill_4 FILLER_70_232 ();
 sg13g2_fill_2 FILLER_70_236 ();
 sg13g2_fill_8 FILLER_70_264 ();
 sg13g2_fill_4 FILLER_70_272 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_fill_1 FILLER_70_298 ();
 sg13g2_fill_2 FILLER_70_335 ();
 sg13g2_fill_1 FILLER_70_347 ();
 sg13g2_fill_2 FILLER_70_368 ();
 sg13g2_fill_1 FILLER_70_370 ();
 sg13g2_fill_8 FILLER_70_387 ();
 sg13g2_fill_4 FILLER_70_395 ();
 sg13g2_fill_2 FILLER_70_399 ();
 sg13g2_fill_8 FILLER_70_406 ();
 sg13g2_fill_8 FILLER_70_414 ();
 sg13g2_fill_8 FILLER_70_422 ();
 sg13g2_fill_8 FILLER_70_430 ();
 sg13g2_fill_8 FILLER_70_438 ();
 sg13g2_fill_1 FILLER_70_446 ();
 sg13g2_fill_8 FILLER_70_473 ();
 sg13g2_fill_2 FILLER_70_481 ();
 sg13g2_fill_8 FILLER_70_491 ();
 sg13g2_fill_4 FILLER_70_499 ();
 sg13g2_fill_2 FILLER_70_503 ();
 sg13g2_fill_8 FILLER_70_557 ();
 sg13g2_fill_2 FILLER_70_565 ();
 sg13g2_fill_1 FILLER_70_567 ();
 sg13g2_fill_2 FILLER_70_594 ();
 sg13g2_fill_1 FILLER_70_596 ();
 sg13g2_fill_1 FILLER_70_627 ();
 sg13g2_fill_4 FILLER_70_636 ();
 sg13g2_fill_8 FILLER_70_646 ();
 sg13g2_fill_1 FILLER_70_654 ();
 sg13g2_fill_8 FILLER_70_688 ();
 sg13g2_fill_4 FILLER_70_696 ();
 sg13g2_fill_1 FILLER_70_700 ();
 sg13g2_fill_2 FILLER_70_769 ();
 sg13g2_fill_1 FILLER_70_771 ();
 sg13g2_fill_1 FILLER_70_786 ();
 sg13g2_fill_1 FILLER_70_862 ();
 sg13g2_fill_2 FILLER_70_900 ();
 sg13g2_fill_2 FILLER_70_945 ();
 sg13g2_fill_2 FILLER_70_1002 ();
 sg13g2_fill_4 FILLER_70_1034 ();
 sg13g2_fill_2 FILLER_70_1038 ();
 sg13g2_fill_2 FILLER_70_1048 ();
 sg13g2_fill_1 FILLER_70_1050 ();
 sg13g2_fill_1 FILLER_70_1057 ();
 sg13g2_fill_2 FILLER_70_1062 ();
 sg13g2_fill_1 FILLER_70_1078 ();
 sg13g2_fill_1 FILLER_70_1092 ();
 sg13g2_fill_8 FILLER_70_1101 ();
 sg13g2_fill_8 FILLER_70_1109 ();
 sg13g2_fill_2 FILLER_70_1117 ();
 sg13g2_fill_2 FILLER_70_1123 ();
 sg13g2_fill_4 FILLER_70_1135 ();
 sg13g2_fill_1 FILLER_70_1139 ();
 sg13g2_fill_4 FILLER_70_1145 ();
 sg13g2_fill_1 FILLER_70_1149 ();
 sg13g2_fill_8 FILLER_70_1160 ();
 sg13g2_fill_1 FILLER_70_1168 ();
 sg13g2_fill_2 FILLER_70_1181 ();
 sg13g2_fill_4 FILLER_70_1187 ();
 sg13g2_fill_1 FILLER_70_1191 ();
 sg13g2_fill_8 FILLER_70_1195 ();
 sg13g2_fill_1 FILLER_70_1203 ();
 sg13g2_fill_8 FILLER_70_1213 ();
 sg13g2_fill_8 FILLER_70_1221 ();
 sg13g2_fill_2 FILLER_70_1229 ();
 sg13g2_fill_1 FILLER_70_1231 ();
 sg13g2_fill_2 FILLER_70_1237 ();
 sg13g2_fill_1 FILLER_70_1239 ();
 sg13g2_fill_8 FILLER_70_1245 ();
 sg13g2_fill_2 FILLER_70_1253 ();
 sg13g2_fill_1 FILLER_70_1255 ();
 sg13g2_fill_2 FILLER_70_1277 ();
 sg13g2_fill_8 FILLER_70_1289 ();
 sg13g2_fill_4 FILLER_70_1297 ();
 sg13g2_fill_1 FILLER_70_1301 ();
 sg13g2_fill_1 FILLER_70_1310 ();
 sg13g2_fill_4 FILLER_70_1322 ();
 sg13g2_fill_1 FILLER_70_1326 ();
 sg13g2_fill_4 FILLER_70_1335 ();
 sg13g2_fill_1 FILLER_70_1339 ();
 sg13g2_fill_1 FILLER_70_1354 ();
 sg13g2_fill_1 FILLER_70_1368 ();
 sg13g2_fill_1 FILLER_70_1374 ();
 sg13g2_fill_2 FILLER_70_1407 ();
 sg13g2_fill_2 FILLER_70_1414 ();
 sg13g2_fill_1 FILLER_70_1426 ();
 sg13g2_fill_8 FILLER_70_1436 ();
 sg13g2_fill_4 FILLER_70_1444 ();
 sg13g2_fill_8 FILLER_70_1456 ();
 sg13g2_fill_4 FILLER_70_1464 ();
 sg13g2_fill_1 FILLER_70_1468 ();
 sg13g2_fill_4 FILLER_70_1499 ();
 sg13g2_fill_2 FILLER_70_1503 ();
 sg13g2_fill_1 FILLER_70_1505 ();
 sg13g2_fill_2 FILLER_70_1536 ();
 sg13g2_fill_1 FILLER_70_1538 ();
 sg13g2_fill_2 FILLER_70_1545 ();
 sg13g2_fill_1 FILLER_70_1547 ();
 sg13g2_fill_8 FILLER_70_1556 ();
 sg13g2_fill_2 FILLER_70_1564 ();
 sg13g2_fill_8 FILLER_70_1570 ();
 sg13g2_fill_8 FILLER_70_1578 ();
 sg13g2_fill_4 FILLER_70_1586 ();
 sg13g2_fill_2 FILLER_70_1590 ();
 sg13g2_fill_8 FILLER_71_0 ();
 sg13g2_fill_8 FILLER_71_8 ();
 sg13g2_fill_8 FILLER_71_16 ();
 sg13g2_fill_8 FILLER_71_24 ();
 sg13g2_fill_8 FILLER_71_32 ();
 sg13g2_fill_8 FILLER_71_40 ();
 sg13g2_fill_1 FILLER_71_48 ();
 sg13g2_fill_2 FILLER_71_59 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_4 FILLER_71_93 ();
 sg13g2_fill_2 FILLER_71_97 ();
 sg13g2_fill_1 FILLER_71_99 ();
 sg13g2_fill_1 FILLER_71_105 ();
 sg13g2_fill_8 FILLER_71_111 ();
 sg13g2_fill_4 FILLER_71_119 ();
 sg13g2_fill_1 FILLER_71_123 ();
 sg13g2_fill_4 FILLER_71_160 ();
 sg13g2_fill_1 FILLER_71_164 ();
 sg13g2_fill_8 FILLER_71_173 ();
 sg13g2_fill_8 FILLER_71_181 ();
 sg13g2_fill_2 FILLER_71_197 ();
 sg13g2_fill_8 FILLER_71_246 ();
 sg13g2_fill_4 FILLER_71_254 ();
 sg13g2_fill_2 FILLER_71_258 ();
 sg13g2_fill_1 FILLER_71_260 ();
 sg13g2_fill_8 FILLER_71_287 ();
 sg13g2_fill_8 FILLER_71_295 ();
 sg13g2_fill_8 FILLER_71_303 ();
 sg13g2_fill_8 FILLER_71_311 ();
 sg13g2_fill_8 FILLER_71_319 ();
 sg13g2_fill_8 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_335 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_407 ();
 sg13g2_fill_2 FILLER_71_418 ();
 sg13g2_fill_8 FILLER_71_446 ();
 sg13g2_fill_8 FILLER_71_454 ();
 sg13g2_fill_8 FILLER_71_462 ();
 sg13g2_fill_8 FILLER_71_470 ();
 sg13g2_fill_8 FILLER_71_478 ();
 sg13g2_fill_4 FILLER_71_486 ();
 sg13g2_fill_8 FILLER_71_516 ();
 sg13g2_fill_1 FILLER_71_524 ();
 sg13g2_fill_2 FILLER_71_570 ();
 sg13g2_fill_1 FILLER_71_572 ();
 sg13g2_fill_4 FILLER_71_634 ();
 sg13g2_fill_2 FILLER_71_638 ();
 sg13g2_fill_2 FILLER_71_674 ();
 sg13g2_fill_4 FILLER_71_721 ();
 sg13g2_fill_4 FILLER_71_730 ();
 sg13g2_fill_2 FILLER_71_734 ();
 sg13g2_fill_1 FILLER_71_736 ();
 sg13g2_fill_8 FILLER_71_750 ();
 sg13g2_fill_1 FILLER_71_758 ();
 sg13g2_fill_4 FILLER_71_789 ();
 sg13g2_fill_2 FILLER_71_793 ();
 sg13g2_fill_1 FILLER_71_795 ();
 sg13g2_fill_2 FILLER_71_832 ();
 sg13g2_fill_8 FILLER_71_866 ();
 sg13g2_fill_2 FILLER_71_880 ();
 sg13g2_fill_2 FILLER_71_897 ();
 sg13g2_fill_2 FILLER_71_915 ();
 sg13g2_fill_1 FILLER_71_955 ();
 sg13g2_fill_2 FILLER_71_969 ();
 sg13g2_fill_1 FILLER_71_1066 ();
 sg13g2_fill_8 FILLER_71_1077 ();
 sg13g2_fill_8 FILLER_71_1085 ();
 sg13g2_fill_8 FILLER_71_1093 ();
 sg13g2_fill_4 FILLER_71_1101 ();
 sg13g2_fill_4 FILLER_71_1112 ();
 sg13g2_fill_1 FILLER_71_1116 ();
 sg13g2_fill_2 FILLER_71_1121 ();
 sg13g2_fill_1 FILLER_71_1123 ();
 sg13g2_fill_2 FILLER_71_1149 ();
 sg13g2_fill_1 FILLER_71_1151 ();
 sg13g2_fill_2 FILLER_71_1161 ();
 sg13g2_fill_4 FILLER_71_1172 ();
 sg13g2_fill_2 FILLER_71_1185 ();
 sg13g2_fill_2 FILLER_71_1218 ();
 sg13g2_fill_8 FILLER_71_1230 ();
 sg13g2_fill_8 FILLER_71_1238 ();
 sg13g2_fill_4 FILLER_71_1246 ();
 sg13g2_fill_2 FILLER_71_1250 ();
 sg13g2_fill_1 FILLER_71_1252 ();
 sg13g2_fill_8 FILLER_71_1257 ();
 sg13g2_fill_4 FILLER_71_1265 ();
 sg13g2_fill_8 FILLER_71_1273 ();
 sg13g2_fill_8 FILLER_71_1281 ();
 sg13g2_fill_8 FILLER_71_1289 ();
 sg13g2_fill_2 FILLER_71_1297 ();
 sg13g2_fill_2 FILLER_71_1308 ();
 sg13g2_fill_2 FILLER_71_1329 ();
 sg13g2_fill_2 FILLER_71_1356 ();
 sg13g2_fill_2 FILLER_71_1390 ();
 sg13g2_fill_2 FILLER_71_1409 ();
 sg13g2_fill_8 FILLER_71_1430 ();
 sg13g2_fill_4 FILLER_71_1438 ();
 sg13g2_fill_8 FILLER_71_1446 ();
 sg13g2_fill_8 FILLER_71_1454 ();
 sg13g2_fill_8 FILLER_71_1462 ();
 sg13g2_fill_4 FILLER_71_1497 ();
 sg13g2_fill_4 FILLER_71_1519 ();
 sg13g2_fill_1 FILLER_71_1523 ();
 sg13g2_fill_2 FILLER_71_1532 ();
 sg13g2_fill_2 FILLER_71_1560 ();
 sg13g2_fill_8 FILLER_72_0 ();
 sg13g2_fill_8 FILLER_72_8 ();
 sg13g2_fill_8 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_24 ();
 sg13g2_fill_8 FILLER_72_61 ();
 sg13g2_fill_8 FILLER_72_69 ();
 sg13g2_fill_8 FILLER_72_77 ();
 sg13g2_fill_2 FILLER_72_85 ();
 sg13g2_fill_1 FILLER_72_87 ();
 sg13g2_fill_8 FILLER_72_93 ();
 sg13g2_fill_8 FILLER_72_134 ();
 sg13g2_fill_4 FILLER_72_142 ();
 sg13g2_fill_1 FILLER_72_146 ();
 sg13g2_fill_2 FILLER_72_168 ();
 sg13g2_fill_1 FILLER_72_170 ();
 sg13g2_fill_2 FILLER_72_197 ();
 sg13g2_fill_8 FILLER_72_230 ();
 sg13g2_fill_8 FILLER_72_238 ();
 sg13g2_fill_4 FILLER_72_246 ();
 sg13g2_fill_1 FILLER_72_250 ();
 sg13g2_fill_8 FILLER_72_259 ();
 sg13g2_fill_8 FILLER_72_267 ();
 sg13g2_fill_8 FILLER_72_275 ();
 sg13g2_fill_2 FILLER_72_283 ();
 sg13g2_fill_2 FILLER_72_314 ();
 sg13g2_fill_1 FILLER_72_316 ();
 sg13g2_fill_8 FILLER_72_330 ();
 sg13g2_fill_8 FILLER_72_338 ();
 sg13g2_fill_8 FILLER_72_346 ();
 sg13g2_fill_8 FILLER_72_354 ();
 sg13g2_fill_2 FILLER_72_362 ();
 sg13g2_fill_4 FILLER_72_377 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_fill_8 FILLER_72_395 ();
 sg13g2_fill_4 FILLER_72_403 ();
 sg13g2_fill_2 FILLER_72_407 ();
 sg13g2_fill_1 FILLER_72_409 ();
 sg13g2_fill_8 FILLER_72_446 ();
 sg13g2_fill_4 FILLER_72_454 ();
 sg13g2_fill_2 FILLER_72_458 ();
 sg13g2_fill_2 FILLER_72_486 ();
 sg13g2_fill_1 FILLER_72_488 ();
 sg13g2_fill_4 FILLER_72_507 ();
 sg13g2_fill_2 FILLER_72_511 ();
 sg13g2_fill_1 FILLER_72_513 ();
 sg13g2_fill_8 FILLER_72_534 ();
 sg13g2_fill_1 FILLER_72_542 ();
 sg13g2_fill_2 FILLER_72_561 ();
 sg13g2_fill_8 FILLER_72_629 ();
 sg13g2_fill_8 FILLER_72_637 ();
 sg13g2_fill_8 FILLER_72_645 ();
 sg13g2_fill_8 FILLER_72_653 ();
 sg13g2_fill_1 FILLER_72_697 ();
 sg13g2_fill_2 FILLER_72_707 ();
 sg13g2_fill_2 FILLER_72_714 ();
 sg13g2_fill_1 FILLER_72_716 ();
 sg13g2_fill_2 FILLER_72_727 ();
 sg13g2_fill_1 FILLER_72_729 ();
 sg13g2_fill_4 FILLER_72_798 ();
 sg13g2_fill_1 FILLER_72_802 ();
 sg13g2_fill_2 FILLER_72_827 ();
 sg13g2_fill_2 FILLER_72_832 ();
 sg13g2_fill_4 FILLER_72_866 ();
 sg13g2_fill_2 FILLER_72_870 ();
 sg13g2_fill_1 FILLER_72_872 ();
 sg13g2_fill_1 FILLER_72_901 ();
 sg13g2_fill_2 FILLER_72_913 ();
 sg13g2_fill_1 FILLER_72_920 ();
 sg13g2_fill_2 FILLER_72_931 ();
 sg13g2_fill_2 FILLER_72_944 ();
 sg13g2_fill_1 FILLER_72_990 ();
 sg13g2_fill_8 FILLER_72_1010 ();
 sg13g2_fill_2 FILLER_72_1018 ();
 sg13g2_fill_8 FILLER_72_1024 ();
 sg13g2_fill_1 FILLER_72_1032 ();
 sg13g2_fill_8 FILLER_72_1037 ();
 sg13g2_fill_1 FILLER_72_1045 ();
 sg13g2_fill_4 FILLER_72_1050 ();
 sg13g2_fill_2 FILLER_72_1077 ();
 sg13g2_fill_1 FILLER_72_1079 ();
 sg13g2_fill_2 FILLER_72_1125 ();
 sg13g2_fill_1 FILLER_72_1127 ();
 sg13g2_fill_1 FILLER_72_1133 ();
 sg13g2_fill_4 FILLER_72_1138 ();
 sg13g2_fill_2 FILLER_72_1142 ();
 sg13g2_fill_8 FILLER_72_1172 ();
 sg13g2_fill_2 FILLER_72_1180 ();
 sg13g2_fill_8 FILLER_72_1186 ();
 sg13g2_fill_8 FILLER_72_1194 ();
 sg13g2_fill_8 FILLER_72_1202 ();
 sg13g2_fill_2 FILLER_72_1210 ();
 sg13g2_fill_1 FILLER_72_1212 ();
 sg13g2_fill_4 FILLER_72_1218 ();
 sg13g2_fill_2 FILLER_72_1222 ();
 sg13g2_fill_2 FILLER_72_1233 ();
 sg13g2_fill_1 FILLER_72_1248 ();
 sg13g2_fill_8 FILLER_72_1289 ();
 sg13g2_fill_4 FILLER_72_1297 ();
 sg13g2_fill_2 FILLER_72_1301 ();
 sg13g2_fill_2 FILLER_72_1343 ();
 sg13g2_fill_1 FILLER_72_1360 ();
 sg13g2_fill_2 FILLER_72_1364 ();
 sg13g2_fill_2 FILLER_72_1378 ();
 sg13g2_fill_4 FILLER_72_1431 ();
 sg13g2_fill_1 FILLER_72_1466 ();
 sg13g2_fill_4 FILLER_72_1485 ();
 sg13g2_fill_2 FILLER_72_1489 ();
 sg13g2_fill_8 FILLER_72_1503 ();
 sg13g2_fill_2 FILLER_72_1511 ();
 sg13g2_fill_1 FILLER_72_1513 ();
 sg13g2_fill_8 FILLER_72_1519 ();
 sg13g2_fill_8 FILLER_72_1527 ();
 sg13g2_fill_8 FILLER_72_1535 ();
 sg13g2_fill_2 FILLER_72_1543 ();
 sg13g2_fill_8 FILLER_72_1550 ();
 sg13g2_fill_1 FILLER_72_1558 ();
 sg13g2_fill_2 FILLER_72_1589 ();
 sg13g2_fill_1 FILLER_72_1591 ();
 sg13g2_fill_8 FILLER_73_0 ();
 sg13g2_fill_4 FILLER_73_8 ();
 sg13g2_fill_2 FILLER_73_12 ();
 sg13g2_fill_1 FILLER_73_14 ();
 sg13g2_fill_8 FILLER_73_73 ();
 sg13g2_fill_1 FILLER_73_81 ();
 sg13g2_fill_4 FILLER_73_88 ();
 sg13g2_fill_2 FILLER_73_126 ();
 sg13g2_fill_4 FILLER_73_138 ();
 sg13g2_fill_1 FILLER_73_173 ();
 sg13g2_fill_8 FILLER_73_184 ();
 sg13g2_fill_2 FILLER_73_192 ();
 sg13g2_fill_1 FILLER_73_212 ();
 sg13g2_fill_4 FILLER_73_249 ();
 sg13g2_fill_2 FILLER_73_253 ();
 sg13g2_fill_4 FILLER_73_312 ();
 sg13g2_fill_2 FILLER_73_316 ();
 sg13g2_fill_1 FILLER_73_318 ();
 sg13g2_fill_4 FILLER_73_332 ();
 sg13g2_fill_1 FILLER_73_336 ();
 sg13g2_fill_4 FILLER_73_345 ();
 sg13g2_fill_8 FILLER_73_362 ();
 sg13g2_fill_4 FILLER_73_370 ();
 sg13g2_fill_1 FILLER_73_374 ();
 sg13g2_fill_8 FILLER_73_380 ();
 sg13g2_fill_4 FILLER_73_388 ();
 sg13g2_fill_8 FILLER_73_397 ();
 sg13g2_fill_8 FILLER_73_405 ();
 sg13g2_fill_1 FILLER_73_428 ();
 sg13g2_fill_8 FILLER_73_469 ();
 sg13g2_fill_4 FILLER_73_477 ();
 sg13g2_fill_1 FILLER_73_481 ();
 sg13g2_fill_8 FILLER_73_534 ();
 sg13g2_fill_2 FILLER_73_542 ();
 sg13g2_fill_1 FILLER_73_544 ();
 sg13g2_fill_8 FILLER_73_587 ();
 sg13g2_fill_8 FILLER_73_595 ();
 sg13g2_fill_4 FILLER_73_603 ();
 sg13g2_fill_2 FILLER_73_607 ();
 sg13g2_fill_1 FILLER_73_609 ();
 sg13g2_fill_2 FILLER_73_646 ();
 sg13g2_fill_1 FILLER_73_648 ();
 sg13g2_fill_2 FILLER_73_675 ();
 sg13g2_fill_1 FILLER_73_677 ();
 sg13g2_fill_4 FILLER_73_734 ();
 sg13g2_fill_4 FILLER_73_768 ();
 sg13g2_fill_2 FILLER_73_772 ();
 sg13g2_fill_8 FILLER_73_837 ();
 sg13g2_fill_1 FILLER_73_845 ();
 sg13g2_fill_2 FILLER_73_898 ();
 sg13g2_fill_2 FILLER_73_905 ();
 sg13g2_fill_2 FILLER_73_944 ();
 sg13g2_fill_2 FILLER_73_992 ();
 sg13g2_fill_8 FILLER_73_1000 ();
 sg13g2_fill_8 FILLER_73_1008 ();
 sg13g2_fill_4 FILLER_73_1016 ();
 sg13g2_fill_2 FILLER_73_1020 ();
 sg13g2_fill_1 FILLER_73_1022 ();
 sg13g2_fill_1 FILLER_73_1028 ();
 sg13g2_fill_1 FILLER_73_1044 ();
 sg13g2_fill_8 FILLER_73_1068 ();
 sg13g2_fill_8 FILLER_73_1076 ();
 sg13g2_fill_8 FILLER_73_1084 ();
 sg13g2_fill_8 FILLER_73_1092 ();
 sg13g2_fill_4 FILLER_73_1100 ();
 sg13g2_fill_1 FILLER_73_1104 ();
 sg13g2_fill_8 FILLER_73_1126 ();
 sg13g2_fill_1 FILLER_73_1134 ();
 sg13g2_fill_8 FILLER_73_1139 ();
 sg13g2_fill_1 FILLER_73_1147 ();
 sg13g2_fill_8 FILLER_73_1157 ();
 sg13g2_fill_8 FILLER_73_1165 ();
 sg13g2_fill_1 FILLER_73_1173 ();
 sg13g2_fill_1 FILLER_73_1178 ();
 sg13g2_fill_2 FILLER_73_1192 ();
 sg13g2_fill_1 FILLER_73_1194 ();
 sg13g2_fill_8 FILLER_73_1224 ();
 sg13g2_fill_8 FILLER_73_1232 ();
 sg13g2_fill_4 FILLER_73_1240 ();
 sg13g2_fill_1 FILLER_73_1244 ();
 sg13g2_fill_4 FILLER_73_1249 ();
 sg13g2_fill_1 FILLER_73_1253 ();
 sg13g2_fill_8 FILLER_73_1263 ();
 sg13g2_fill_2 FILLER_73_1271 ();
 sg13g2_fill_1 FILLER_73_1273 ();
 sg13g2_fill_8 FILLER_73_1279 ();
 sg13g2_fill_8 FILLER_73_1287 ();
 sg13g2_fill_2 FILLER_73_1300 ();
 sg13g2_fill_8 FILLER_73_1305 ();
 sg13g2_fill_8 FILLER_73_1318 ();
 sg13g2_fill_4 FILLER_73_1326 ();
 sg13g2_fill_1 FILLER_73_1330 ();
 sg13g2_fill_2 FILLER_73_1337 ();
 sg13g2_fill_2 FILLER_73_1347 ();
 sg13g2_fill_2 FILLER_73_1356 ();
 sg13g2_fill_4 FILLER_73_1449 ();
 sg13g2_fill_4 FILLER_73_1461 ();
 sg13g2_fill_2 FILLER_73_1465 ();
 sg13g2_fill_1 FILLER_73_1467 ();
 sg13g2_fill_8 FILLER_73_1583 ();
 sg13g2_fill_1 FILLER_73_1591 ();
 sg13g2_fill_8 FILLER_74_0 ();
 sg13g2_fill_8 FILLER_74_8 ();
 sg13g2_fill_8 FILLER_74_16 ();
 sg13g2_fill_2 FILLER_74_24 ();
 sg13g2_fill_8 FILLER_74_36 ();
 sg13g2_fill_8 FILLER_74_44 ();
 sg13g2_fill_8 FILLER_74_52 ();
 sg13g2_fill_2 FILLER_74_60 ();
 sg13g2_fill_1 FILLER_74_62 ();
 sg13g2_fill_2 FILLER_74_98 ();
 sg13g2_fill_1 FILLER_74_100 ();
 sg13g2_fill_8 FILLER_74_111 ();
 sg13g2_fill_8 FILLER_74_119 ();
 sg13g2_fill_2 FILLER_74_127 ();
 sg13g2_fill_2 FILLER_74_155 ();
 sg13g2_fill_1 FILLER_74_157 ();
 sg13g2_fill_8 FILLER_74_166 ();
 sg13g2_fill_4 FILLER_74_174 ();
 sg13g2_fill_2 FILLER_74_178 ();
 sg13g2_fill_4 FILLER_74_201 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_8 FILLER_74_232 ();
 sg13g2_fill_1 FILLER_74_240 ();
 sg13g2_fill_8 FILLER_74_277 ();
 sg13g2_fill_8 FILLER_74_285 ();
 sg13g2_fill_8 FILLER_74_293 ();
 sg13g2_fill_1 FILLER_74_301 ();
 sg13g2_fill_2 FILLER_74_310 ();
 sg13g2_fill_1 FILLER_74_312 ();
 sg13g2_fill_4 FILLER_74_326 ();
 sg13g2_fill_2 FILLER_74_330 ();
 sg13g2_fill_1 FILLER_74_332 ();
 sg13g2_fill_8 FILLER_74_346 ();
 sg13g2_fill_1 FILLER_74_354 ();
 sg13g2_fill_8 FILLER_74_401 ();
 sg13g2_fill_8 FILLER_74_409 ();
 sg13g2_fill_8 FILLER_74_417 ();
 sg13g2_fill_8 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_433 ();
 sg13g2_fill_4 FILLER_74_452 ();
 sg13g2_fill_2 FILLER_74_456 ();
 sg13g2_fill_1 FILLER_74_458 ();
 sg13g2_fill_8 FILLER_74_485 ();
 sg13g2_fill_8 FILLER_74_493 ();
 sg13g2_fill_2 FILLER_74_501 ();
 sg13g2_fill_1 FILLER_74_503 ();
 sg13g2_fill_8 FILLER_74_510 ();
 sg13g2_fill_4 FILLER_74_518 ();
 sg13g2_fill_1 FILLER_74_522 ();
 sg13g2_fill_4 FILLER_74_531 ();
 sg13g2_fill_2 FILLER_74_535 ();
 sg13g2_fill_8 FILLER_74_547 ();
 sg13g2_fill_8 FILLER_74_555 ();
 sg13g2_fill_8 FILLER_74_563 ();
 sg13g2_fill_2 FILLER_74_571 ();
 sg13g2_fill_1 FILLER_74_573 ();
 sg13g2_fill_2 FILLER_74_590 ();
 sg13g2_fill_4 FILLER_74_602 ();
 sg13g2_fill_1 FILLER_74_606 ();
 sg13g2_fill_4 FILLER_74_633 ();
 sg13g2_fill_1 FILLER_74_637 ();
 sg13g2_fill_8 FILLER_74_646 ();
 sg13g2_fill_2 FILLER_74_654 ();
 sg13g2_fill_1 FILLER_74_656 ();
 sg13g2_fill_8 FILLER_74_665 ();
 sg13g2_fill_8 FILLER_74_673 ();
 sg13g2_fill_4 FILLER_74_681 ();
 sg13g2_fill_8 FILLER_74_693 ();
 sg13g2_fill_4 FILLER_74_701 ();
 sg13g2_fill_2 FILLER_74_705 ();
 sg13g2_fill_8 FILLER_74_746 ();
 sg13g2_fill_1 FILLER_74_754 ();
 sg13g2_fill_4 FILLER_74_798 ();
 sg13g2_fill_1 FILLER_74_802 ();
 sg13g2_fill_8 FILLER_74_813 ();
 sg13g2_fill_8 FILLER_74_821 ();
 sg13g2_fill_4 FILLER_74_829 ();
 sg13g2_fill_8 FILLER_74_863 ();
 sg13g2_fill_2 FILLER_74_871 ();
 sg13g2_fill_1 FILLER_74_897 ();
 sg13g2_fill_2 FILLER_74_908 ();
 sg13g2_fill_1 FILLER_74_922 ();
 sg13g2_fill_2 FILLER_74_962 ();
 sg13g2_fill_1 FILLER_74_985 ();
 sg13g2_fill_8 FILLER_74_1069 ();
 sg13g2_fill_4 FILLER_74_1077 ();
 sg13g2_fill_4 FILLER_74_1101 ();
 sg13g2_fill_1 FILLER_74_1105 ();
 sg13g2_fill_4 FILLER_74_1110 ();
 sg13g2_fill_1 FILLER_74_1114 ();
 sg13g2_fill_2 FILLER_74_1125 ();
 sg13g2_fill_4 FILLER_74_1132 ();
 sg13g2_fill_1 FILLER_74_1136 ();
 sg13g2_fill_1 FILLER_74_1142 ();
 sg13g2_fill_2 FILLER_74_1158 ();
 sg13g2_fill_1 FILLER_74_1160 ();
 sg13g2_fill_2 FILLER_74_1171 ();
 sg13g2_fill_1 FILLER_74_1173 ();
 sg13g2_fill_2 FILLER_74_1193 ();
 sg13g2_fill_8 FILLER_74_1203 ();
 sg13g2_fill_1 FILLER_74_1242 ();
 sg13g2_fill_4 FILLER_74_1257 ();
 sg13g2_fill_8 FILLER_74_1267 ();
 sg13g2_fill_2 FILLER_74_1275 ();
 sg13g2_fill_1 FILLER_74_1277 ();
 sg13g2_fill_4 FILLER_74_1282 ();
 sg13g2_fill_2 FILLER_74_1295 ();
 sg13g2_fill_8 FILLER_74_1306 ();
 sg13g2_fill_4 FILLER_74_1314 ();
 sg13g2_fill_2 FILLER_74_1318 ();
 sg13g2_fill_1 FILLER_74_1320 ();
 sg13g2_fill_4 FILLER_74_1331 ();
 sg13g2_fill_1 FILLER_74_1335 ();
 sg13g2_fill_4 FILLER_74_1341 ();
 sg13g2_fill_1 FILLER_74_1416 ();
 sg13g2_fill_2 FILLER_74_1422 ();
 sg13g2_fill_1 FILLER_74_1424 ();
 sg13g2_fill_4 FILLER_74_1429 ();
 sg13g2_fill_2 FILLER_74_1433 ();
 sg13g2_fill_1 FILLER_74_1435 ();
 sg13g2_fill_4 FILLER_74_1466 ();
 sg13g2_fill_2 FILLER_74_1470 ();
 sg13g2_fill_1 FILLER_74_1472 ();
 sg13g2_fill_8 FILLER_74_1480 ();
 sg13g2_fill_4 FILLER_74_1488 ();
 sg13g2_fill_2 FILLER_74_1492 ();
 sg13g2_fill_1 FILLER_74_1494 ();
 sg13g2_fill_2 FILLER_74_1500 ();
 sg13g2_fill_1 FILLER_74_1502 ();
 sg13g2_fill_1 FILLER_74_1510 ();
 sg13g2_fill_8 FILLER_74_1517 ();
 sg13g2_fill_8 FILLER_74_1525 ();
 sg13g2_fill_8 FILLER_74_1533 ();
 sg13g2_fill_8 FILLER_75_0 ();
 sg13g2_fill_8 FILLER_75_8 ();
 sg13g2_fill_8 FILLER_75_16 ();
 sg13g2_fill_8 FILLER_75_24 ();
 sg13g2_fill_8 FILLER_75_32 ();
 sg13g2_fill_8 FILLER_75_40 ();
 sg13g2_fill_4 FILLER_75_48 ();
 sg13g2_fill_8 FILLER_75_88 ();
 sg13g2_fill_4 FILLER_75_96 ();
 sg13g2_fill_2 FILLER_75_100 ();
 sg13g2_fill_1 FILLER_75_102 ();
 sg13g2_fill_8 FILLER_75_134 ();
 sg13g2_fill_8 FILLER_75_173 ();
 sg13g2_fill_1 FILLER_75_181 ();
 sg13g2_fill_8 FILLER_75_203 ();
 sg13g2_fill_8 FILLER_75_211 ();
 sg13g2_fill_8 FILLER_75_219 ();
 sg13g2_fill_4 FILLER_75_227 ();
 sg13g2_fill_1 FILLER_75_231 ();
 sg13g2_fill_8 FILLER_75_242 ();
 sg13g2_fill_8 FILLER_75_250 ();
 sg13g2_fill_8 FILLER_75_258 ();
 sg13g2_fill_2 FILLER_75_266 ();
 sg13g2_fill_1 FILLER_75_268 ();
 sg13g2_fill_8 FILLER_75_294 ();
 sg13g2_fill_4 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_306 ();
 sg13g2_fill_8 FILLER_75_317 ();
 sg13g2_fill_8 FILLER_75_325 ();
 sg13g2_fill_8 FILLER_75_333 ();
 sg13g2_fill_4 FILLER_75_341 ();
 sg13g2_fill_2 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_75_347 ();
 sg13g2_fill_8 FILLER_75_378 ();
 sg13g2_fill_4 FILLER_75_386 ();
 sg13g2_fill_2 FILLER_75_390 ();
 sg13g2_fill_8 FILLER_75_418 ();
 sg13g2_fill_1 FILLER_75_426 ();
 sg13g2_fill_2 FILLER_75_437 ();
 sg13g2_fill_8 FILLER_75_470 ();
 sg13g2_fill_1 FILLER_75_478 ();
 sg13g2_fill_8 FILLER_75_485 ();
 sg13g2_fill_4 FILLER_75_493 ();
 sg13g2_fill_1 FILLER_75_507 ();
 sg13g2_fill_8 FILLER_75_526 ();
 sg13g2_fill_1 FILLER_75_534 ();
 sg13g2_fill_4 FILLER_75_540 ();
 sg13g2_fill_4 FILLER_75_570 ();
 sg13g2_fill_2 FILLER_75_574 ();
 sg13g2_fill_1 FILLER_75_576 ();
 sg13g2_fill_8 FILLER_75_608 ();
 sg13g2_fill_8 FILLER_75_616 ();
 sg13g2_fill_8 FILLER_75_624 ();
 sg13g2_fill_8 FILLER_75_632 ();
 sg13g2_fill_4 FILLER_75_640 ();
 sg13g2_fill_4 FILLER_75_649 ();
 sg13g2_fill_1 FILLER_75_653 ();
 sg13g2_fill_8 FILLER_75_672 ();
 sg13g2_fill_2 FILLER_75_680 ();
 sg13g2_fill_4 FILLER_75_702 ();
 sg13g2_fill_1 FILLER_75_706 ();
 sg13g2_fill_8 FILLER_75_737 ();
 sg13g2_fill_4 FILLER_75_745 ();
 sg13g2_fill_2 FILLER_75_749 ();
 sg13g2_fill_1 FILLER_75_751 ();
 sg13g2_fill_1 FILLER_75_760 ();
 sg13g2_fill_8 FILLER_75_796 ();
 sg13g2_fill_2 FILLER_75_804 ();
 sg13g2_fill_8 FILLER_75_867 ();
 sg13g2_fill_1 FILLER_75_875 ();
 sg13g2_fill_1 FILLER_75_888 ();
 sg13g2_fill_1 FILLER_75_945 ();
 sg13g2_fill_2 FILLER_75_950 ();
 sg13g2_fill_4 FILLER_75_1011 ();
 sg13g2_fill_1 FILLER_75_1015 ();
 sg13g2_fill_4 FILLER_75_1019 ();
 sg13g2_fill_2 FILLER_75_1023 ();
 sg13g2_fill_1 FILLER_75_1028 ();
 sg13g2_fill_2 FILLER_75_1045 ();
 sg13g2_fill_1 FILLER_75_1066 ();
 sg13g2_fill_1 FILLER_75_1070 ();
 sg13g2_fill_2 FILLER_75_1087 ();
 sg13g2_fill_2 FILLER_75_1097 ();
 sg13g2_fill_8 FILLER_75_1113 ();
 sg13g2_fill_4 FILLER_75_1121 ();
 sg13g2_fill_1 FILLER_75_1125 ();
 sg13g2_fill_8 FILLER_75_1131 ();
 sg13g2_fill_8 FILLER_75_1139 ();
 sg13g2_fill_2 FILLER_75_1147 ();
 sg13g2_fill_2 FILLER_75_1154 ();
 sg13g2_fill_2 FILLER_75_1165 ();
 sg13g2_fill_2 FILLER_75_1186 ();
 sg13g2_fill_4 FILLER_75_1192 ();
 sg13g2_fill_2 FILLER_75_1196 ();
 sg13g2_fill_1 FILLER_75_1198 ();
 sg13g2_fill_4 FILLER_75_1204 ();
 sg13g2_fill_1 FILLER_75_1208 ();
 sg13g2_fill_2 FILLER_75_1219 ();
 sg13g2_fill_8 FILLER_75_1224 ();
 sg13g2_fill_8 FILLER_75_1232 ();
 sg13g2_fill_2 FILLER_75_1244 ();
 sg13g2_fill_1 FILLER_75_1246 ();
 sg13g2_fill_8 FILLER_75_1252 ();
 sg13g2_fill_2 FILLER_75_1260 ();
 sg13g2_fill_1 FILLER_75_1280 ();
 sg13g2_fill_2 FILLER_75_1313 ();
 sg13g2_fill_1 FILLER_75_1315 ();
 sg13g2_fill_1 FILLER_75_1321 ();
 sg13g2_fill_8 FILLER_75_1331 ();
 sg13g2_fill_8 FILLER_75_1339 ();
 sg13g2_fill_4 FILLER_75_1347 ();
 sg13g2_fill_1 FILLER_75_1363 ();
 sg13g2_fill_1 FILLER_75_1367 ();
 sg13g2_fill_2 FILLER_75_1374 ();
 sg13g2_fill_2 FILLER_75_1429 ();
 sg13g2_fill_1 FILLER_75_1431 ();
 sg13g2_fill_1 FILLER_75_1478 ();
 sg13g2_fill_2 FILLER_75_1487 ();
 sg13g2_fill_1 FILLER_75_1489 ();
 sg13g2_fill_1 FILLER_75_1498 ();
 sg13g2_fill_4 FILLER_75_1527 ();
 sg13g2_fill_2 FILLER_75_1531 ();
 sg13g2_fill_1 FILLER_75_1533 ();
 sg13g2_fill_1 FILLER_75_1548 ();
 sg13g2_fill_2 FILLER_75_1559 ();
 sg13g2_fill_1 FILLER_75_1561 ();
 sg13g2_fill_8 FILLER_76_0 ();
 sg13g2_fill_8 FILLER_76_8 ();
 sg13g2_fill_8 FILLER_76_16 ();
 sg13g2_fill_8 FILLER_76_24 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_fill_8 FILLER_76_59 ();
 sg13g2_fill_8 FILLER_76_67 ();
 sg13g2_fill_8 FILLER_76_75 ();
 sg13g2_fill_8 FILLER_76_104 ();
 sg13g2_fill_8 FILLER_76_112 ();
 sg13g2_fill_8 FILLER_76_120 ();
 sg13g2_fill_2 FILLER_76_128 ();
 sg13g2_fill_1 FILLER_76_130 ();
 sg13g2_fill_8 FILLER_76_152 ();
 sg13g2_fill_2 FILLER_76_160 ();
 sg13g2_fill_1 FILLER_76_162 ();
 sg13g2_fill_2 FILLER_76_199 ();
 sg13g2_fill_1 FILLER_76_201 ();
 sg13g2_fill_4 FILLER_76_228 ();
 sg13g2_fill_1 FILLER_76_232 ();
 sg13g2_fill_1 FILLER_76_259 ();
 sg13g2_fill_4 FILLER_76_333 ();
 sg13g2_fill_2 FILLER_76_376 ();
 sg13g2_fill_8 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_453 ();
 sg13g2_fill_4 FILLER_76_475 ();
 sg13g2_fill_4 FILLER_76_489 ();
 sg13g2_fill_2 FILLER_76_493 ();
 sg13g2_fill_1 FILLER_76_495 ();
 sg13g2_fill_4 FILLER_76_506 ();
 sg13g2_fill_2 FILLER_76_534 ();
 sg13g2_fill_2 FILLER_76_546 ();
 sg13g2_fill_1 FILLER_76_548 ();
 sg13g2_fill_8 FILLER_76_580 ();
 sg13g2_fill_2 FILLER_76_588 ();
 sg13g2_fill_8 FILLER_76_596 ();
 sg13g2_fill_8 FILLER_76_604 ();
 sg13g2_fill_8 FILLER_76_612 ();
 sg13g2_fill_8 FILLER_76_620 ();
 sg13g2_fill_8 FILLER_76_628 ();
 sg13g2_fill_2 FILLER_76_636 ();
 sg13g2_fill_4 FILLER_76_646 ();
 sg13g2_fill_2 FILLER_76_718 ();
 sg13g2_fill_4 FILLER_76_750 ();
 sg13g2_fill_2 FILLER_76_762 ();
 sg13g2_fill_2 FILLER_76_774 ();
 sg13g2_fill_8 FILLER_76_802 ();
 sg13g2_fill_2 FILLER_76_810 ();
 sg13g2_fill_1 FILLER_76_812 ();
 sg13g2_fill_2 FILLER_76_864 ();
 sg13g2_fill_1 FILLER_76_866 ();
 sg13g2_fill_1 FILLER_76_944 ();
 sg13g2_fill_2 FILLER_76_985 ();
 sg13g2_fill_1 FILLER_76_996 ();
 sg13g2_fill_2 FILLER_76_1087 ();
 sg13g2_fill_2 FILLER_76_1094 ();
 sg13g2_fill_8 FILLER_76_1105 ();
 sg13g2_fill_2 FILLER_76_1128 ();
 sg13g2_fill_1 FILLER_76_1130 ();
 sg13g2_fill_8 FILLER_76_1150 ();
 sg13g2_fill_4 FILLER_76_1158 ();
 sg13g2_fill_1 FILLER_76_1162 ();
 sg13g2_fill_4 FILLER_76_1167 ();
 sg13g2_fill_8 FILLER_76_1176 ();
 sg13g2_fill_4 FILLER_76_1241 ();
 sg13g2_fill_2 FILLER_76_1245 ();
 sg13g2_fill_4 FILLER_76_1252 ();
 sg13g2_fill_2 FILLER_76_1256 ();
 sg13g2_fill_8 FILLER_76_1263 ();
 sg13g2_fill_1 FILLER_76_1271 ();
 sg13g2_fill_4 FILLER_76_1280 ();
 sg13g2_fill_2 FILLER_76_1284 ();
 sg13g2_fill_1 FILLER_76_1286 ();
 sg13g2_fill_1 FILLER_76_1298 ();
 sg13g2_fill_2 FILLER_76_1312 ();
 sg13g2_fill_4 FILLER_76_1327 ();
 sg13g2_fill_1 FILLER_76_1331 ();
 sg13g2_fill_8 FILLER_76_1342 ();
 sg13g2_fill_2 FILLER_76_1371 ();
 sg13g2_fill_2 FILLER_76_1419 ();
 sg13g2_fill_2 FILLER_76_1452 ();
 sg13g2_fill_1 FILLER_76_1454 ();
 sg13g2_fill_1 FILLER_76_1497 ();
 sg13g2_fill_1 FILLER_76_1514 ();
 sg13g2_fill_8 FILLER_76_1561 ();
 sg13g2_fill_8 FILLER_76_1569 ();
 sg13g2_fill_8 FILLER_76_1577 ();
 sg13g2_fill_4 FILLER_76_1585 ();
 sg13g2_fill_2 FILLER_76_1589 ();
 sg13g2_fill_1 FILLER_76_1591 ();
 sg13g2_fill_8 FILLER_77_0 ();
 sg13g2_fill_8 FILLER_77_8 ();
 sg13g2_fill_8 FILLER_77_16 ();
 sg13g2_fill_4 FILLER_77_24 ();
 sg13g2_fill_1 FILLER_77_28 ();
 sg13g2_fill_8 FILLER_77_68 ();
 sg13g2_fill_1 FILLER_77_76 ();
 sg13g2_fill_8 FILLER_77_87 ();
 sg13g2_fill_4 FILLER_77_95 ();
 sg13g2_fill_1 FILLER_77_99 ();
 sg13g2_fill_8 FILLER_77_126 ();
 sg13g2_fill_4 FILLER_77_134 ();
 sg13g2_fill_8 FILLER_77_170 ();
 sg13g2_fill_4 FILLER_77_178 ();
 sg13g2_fill_8 FILLER_77_218 ();
 sg13g2_fill_4 FILLER_77_226 ();
 sg13g2_fill_1 FILLER_77_230 ();
 sg13g2_fill_2 FILLER_77_257 ();
 sg13g2_fill_8 FILLER_77_303 ();
 sg13g2_fill_8 FILLER_77_311 ();
 sg13g2_fill_4 FILLER_77_319 ();
 sg13g2_fill_4 FILLER_77_374 ();
 sg13g2_fill_8 FILLER_77_404 ();
 sg13g2_fill_8 FILLER_77_412 ();
 sg13g2_fill_8 FILLER_77_420 ();
 sg13g2_fill_4 FILLER_77_428 ();
 sg13g2_fill_8 FILLER_77_446 ();
 sg13g2_fill_8 FILLER_77_454 ();
 sg13g2_fill_2 FILLER_77_462 ();
 sg13g2_fill_8 FILLER_77_490 ();
 sg13g2_fill_2 FILLER_77_535 ();
 sg13g2_fill_1 FILLER_77_537 ();
 sg13g2_fill_8 FILLER_77_548 ();
 sg13g2_fill_8 FILLER_77_556 ();
 sg13g2_fill_2 FILLER_77_564 ();
 sg13g2_fill_1 FILLER_77_566 ();
 sg13g2_fill_8 FILLER_77_571 ();
 sg13g2_fill_4 FILLER_77_579 ();
 sg13g2_fill_2 FILLER_77_583 ();
 sg13g2_fill_1 FILLER_77_585 ();
 sg13g2_fill_8 FILLER_77_590 ();
 sg13g2_fill_1 FILLER_77_634 ();
 sg13g2_fill_8 FILLER_77_643 ();
 sg13g2_fill_8 FILLER_77_651 ();
 sg13g2_fill_8 FILLER_77_659 ();
 sg13g2_fill_8 FILLER_77_667 ();
 sg13g2_fill_8 FILLER_77_675 ();
 sg13g2_fill_8 FILLER_77_683 ();
 sg13g2_fill_4 FILLER_77_691 ();
 sg13g2_fill_2 FILLER_77_695 ();
 sg13g2_fill_2 FILLER_77_727 ();
 sg13g2_fill_1 FILLER_77_729 ();
 sg13g2_fill_8 FILLER_77_738 ();
 sg13g2_fill_8 FILLER_77_746 ();
 sg13g2_fill_8 FILLER_77_754 ();
 sg13g2_fill_1 FILLER_77_762 ();
 sg13g2_fill_2 FILLER_77_799 ();
 sg13g2_fill_8 FILLER_77_822 ();
 sg13g2_fill_2 FILLER_77_830 ();
 sg13g2_fill_4 FILLER_77_837 ();
 sg13g2_fill_4 FILLER_77_867 ();
 sg13g2_fill_2 FILLER_77_871 ();
 sg13g2_fill_2 FILLER_77_901 ();
 sg13g2_fill_1 FILLER_77_925 ();
 sg13g2_fill_1 FILLER_77_934 ();
 sg13g2_fill_2 FILLER_77_944 ();
 sg13g2_fill_1 FILLER_77_957 ();
 sg13g2_fill_2 FILLER_77_1043 ();
 sg13g2_fill_1 FILLER_77_1051 ();
 sg13g2_fill_2 FILLER_77_1068 ();
 sg13g2_fill_2 FILLER_77_1106 ();
 sg13g2_fill_1 FILLER_77_1108 ();
 sg13g2_fill_4 FILLER_77_1129 ();
 sg13g2_fill_2 FILLER_77_1133 ();
 sg13g2_fill_2 FILLER_77_1164 ();
 sg13g2_fill_8 FILLER_77_1177 ();
 sg13g2_fill_2 FILLER_77_1185 ();
 sg13g2_fill_1 FILLER_77_1187 ();
 sg13g2_fill_8 FILLER_77_1193 ();
 sg13g2_fill_8 FILLER_77_1201 ();
 sg13g2_fill_2 FILLER_77_1209 ();
 sg13g2_fill_8 FILLER_77_1221 ();
 sg13g2_fill_8 FILLER_77_1229 ();
 sg13g2_fill_4 FILLER_77_1237 ();
 sg13g2_fill_2 FILLER_77_1241 ();
 sg13g2_fill_8 FILLER_77_1267 ();
 sg13g2_fill_4 FILLER_77_1275 ();
 sg13g2_fill_8 FILLER_77_1293 ();
 sg13g2_fill_8 FILLER_77_1306 ();
 sg13g2_fill_8 FILLER_77_1314 ();
 sg13g2_fill_2 FILLER_77_1322 ();
 sg13g2_fill_2 FILLER_77_1329 ();
 sg13g2_fill_1 FILLER_77_1331 ();
 sg13g2_fill_2 FILLER_77_1344 ();
 sg13g2_fill_1 FILLER_77_1346 ();
 sg13g2_fill_2 FILLER_77_1355 ();
 sg13g2_fill_2 FILLER_77_1392 ();
 sg13g2_fill_1 FILLER_77_1419 ();
 sg13g2_fill_4 FILLER_77_1445 ();
 sg13g2_fill_1 FILLER_77_1449 ();
 sg13g2_fill_8 FILLER_77_1455 ();
 sg13g2_fill_1 FILLER_77_1463 ();
 sg13g2_fill_1 FILLER_77_1472 ();
 sg13g2_fill_8 FILLER_77_1477 ();
 sg13g2_fill_8 FILLER_77_1485 ();
 sg13g2_fill_8 FILLER_77_1493 ();
 sg13g2_fill_8 FILLER_77_1501 ();
 sg13g2_fill_2 FILLER_77_1509 ();
 sg13g2_fill_8 FILLER_77_1520 ();
 sg13g2_fill_8 FILLER_77_1528 ();
 sg13g2_fill_8 FILLER_77_1536 ();
 sg13g2_fill_1 FILLER_77_1544 ();
 sg13g2_fill_4 FILLER_77_1550 ();
 sg13g2_fill_2 FILLER_77_1554 ();
 sg13g2_fill_4 FILLER_77_1586 ();
 sg13g2_fill_2 FILLER_77_1590 ();
 sg13g2_fill_8 FILLER_78_0 ();
 sg13g2_fill_8 FILLER_78_8 ();
 sg13g2_fill_8 FILLER_78_16 ();
 sg13g2_fill_2 FILLER_78_24 ();
 sg13g2_fill_1 FILLER_78_26 ();
 sg13g2_fill_8 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_61 ();
 sg13g2_fill_2 FILLER_78_88 ();
 sg13g2_fill_4 FILLER_78_94 ();
 sg13g2_fill_1 FILLER_78_108 ();
 sg13g2_fill_2 FILLER_78_135 ();
 sg13g2_fill_1 FILLER_78_137 ();
 sg13g2_fill_8 FILLER_78_174 ();
 sg13g2_fill_8 FILLER_78_182 ();
 sg13g2_fill_8 FILLER_78_190 ();
 sg13g2_fill_8 FILLER_78_198 ();
 sg13g2_fill_4 FILLER_78_206 ();
 sg13g2_fill_2 FILLER_78_210 ();
 sg13g2_fill_1 FILLER_78_212 ();
 sg13g2_fill_8 FILLER_78_274 ();
 sg13g2_fill_8 FILLER_78_282 ();
 sg13g2_fill_1 FILLER_78_290 ();
 sg13g2_fill_2 FILLER_78_301 ();
 sg13g2_fill_1 FILLER_78_303 ();
 sg13g2_fill_1 FILLER_78_325 ();
 sg13g2_fill_1 FILLER_78_351 ();
 sg13g2_fill_8 FILLER_78_357 ();
 sg13g2_fill_4 FILLER_78_385 ();
 sg13g2_fill_2 FILLER_78_389 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_fill_8 FILLER_78_402 ();
 sg13g2_fill_8 FILLER_78_410 ();
 sg13g2_fill_2 FILLER_78_418 ();
 sg13g2_fill_1 FILLER_78_420 ();
 sg13g2_fill_8 FILLER_78_431 ();
 sg13g2_fill_8 FILLER_78_439 ();
 sg13g2_fill_2 FILLER_78_447 ();
 sg13g2_fill_8 FILLER_78_454 ();
 sg13g2_fill_8 FILLER_78_462 ();
 sg13g2_fill_8 FILLER_78_470 ();
 sg13g2_fill_4 FILLER_78_478 ();
 sg13g2_fill_4 FILLER_78_526 ();
 sg13g2_fill_2 FILLER_78_530 ();
 sg13g2_fill_1 FILLER_78_532 ();
 sg13g2_fill_8 FILLER_78_543 ();
 sg13g2_fill_8 FILLER_78_551 ();
 sg13g2_fill_8 FILLER_78_559 ();
 sg13g2_fill_8 FILLER_78_567 ();
 sg13g2_fill_1 FILLER_78_575 ();
 sg13g2_fill_8 FILLER_78_612 ();
 sg13g2_fill_4 FILLER_78_620 ();
 sg13g2_fill_4 FILLER_78_660 ();
 sg13g2_fill_1 FILLER_78_664 ();
 sg13g2_fill_8 FILLER_78_679 ();
 sg13g2_fill_4 FILLER_78_687 ();
 sg13g2_fill_1 FILLER_78_691 ();
 sg13g2_fill_8 FILLER_78_717 ();
 sg13g2_fill_4 FILLER_78_725 ();
 sg13g2_fill_8 FILLER_78_765 ();
 sg13g2_fill_2 FILLER_78_773 ();
 sg13g2_fill_8 FILLER_78_801 ();
 sg13g2_fill_8 FILLER_78_809 ();
 sg13g2_fill_4 FILLER_78_817 ();
 sg13g2_fill_2 FILLER_78_821 ();
 sg13g2_fill_1 FILLER_78_823 ();
 sg13g2_fill_4 FILLER_78_860 ();
 sg13g2_fill_2 FILLER_78_890 ();
 sg13g2_fill_2 FILLER_78_921 ();
 sg13g2_fill_2 FILLER_78_1021 ();
 sg13g2_fill_1 FILLER_78_1064 ();
 sg13g2_fill_2 FILLER_78_1080 ();
 sg13g2_fill_2 FILLER_78_1086 ();
 sg13g2_fill_1 FILLER_78_1095 ();
 sg13g2_fill_2 FILLER_78_1113 ();
 sg13g2_fill_8 FILLER_78_1120 ();
 sg13g2_fill_8 FILLER_78_1128 ();
 sg13g2_fill_8 FILLER_78_1136 ();
 sg13g2_fill_4 FILLER_78_1144 ();
 sg13g2_fill_1 FILLER_78_1148 ();
 sg13g2_fill_8 FILLER_78_1153 ();
 sg13g2_fill_8 FILLER_78_1161 ();
 sg13g2_fill_8 FILLER_78_1169 ();
 sg13g2_fill_2 FILLER_78_1177 ();
 sg13g2_fill_8 FILLER_78_1187 ();
 sg13g2_fill_8 FILLER_78_1195 ();
 sg13g2_fill_8 FILLER_78_1203 ();
 sg13g2_fill_8 FILLER_78_1215 ();
 sg13g2_fill_8 FILLER_78_1223 ();
 sg13g2_fill_2 FILLER_78_1231 ();
 sg13g2_fill_1 FILLER_78_1233 ();
 sg13g2_fill_8 FILLER_78_1238 ();
 sg13g2_fill_8 FILLER_78_1246 ();
 sg13g2_fill_1 FILLER_78_1254 ();
 sg13g2_fill_4 FILLER_78_1258 ();
 sg13g2_fill_2 FILLER_78_1262 ();
 sg13g2_fill_1 FILLER_78_1264 ();
 sg13g2_fill_8 FILLER_78_1270 ();
 sg13g2_fill_4 FILLER_78_1278 ();
 sg13g2_fill_1 FILLER_78_1282 ();
 sg13g2_fill_2 FILLER_78_1307 ();
 sg13g2_fill_4 FILLER_78_1336 ();
 sg13g2_fill_4 FILLER_78_1358 ();
 sg13g2_fill_2 FILLER_78_1362 ();
 sg13g2_fill_1 FILLER_78_1364 ();
 sg13g2_fill_2 FILLER_78_1374 ();
 sg13g2_fill_1 FILLER_78_1387 ();
 sg13g2_fill_4 FILLER_78_1414 ();
 sg13g2_fill_2 FILLER_78_1418 ();
 sg13g2_fill_8 FILLER_78_1445 ();
 sg13g2_fill_1 FILLER_78_1453 ();
 sg13g2_fill_8 FILLER_78_1462 ();
 sg13g2_fill_4 FILLER_78_1470 ();
 sg13g2_fill_1 FILLER_78_1474 ();
 sg13g2_fill_1 FILLER_78_1485 ();
 sg13g2_fill_1 FILLER_78_1490 ();
 sg13g2_fill_1 FILLER_78_1495 ();
 sg13g2_fill_1 FILLER_78_1510 ();
 sg13g2_fill_4 FILLER_78_1549 ();
 sg13g2_fill_2 FILLER_78_1553 ();
 sg13g2_fill_1 FILLER_78_1555 ();
 sg13g2_fill_4 FILLER_78_1586 ();
 sg13g2_fill_2 FILLER_78_1590 ();
 sg13g2_fill_8 FILLER_79_0 ();
 sg13g2_fill_8 FILLER_79_8 ();
 sg13g2_fill_4 FILLER_79_16 ();
 sg13g2_fill_2 FILLER_79_20 ();
 sg13g2_fill_1 FILLER_79_22 ();
 sg13g2_fill_8 FILLER_79_69 ();
 sg13g2_fill_8 FILLER_79_77 ();
 sg13g2_fill_4 FILLER_79_85 ();
 sg13g2_fill_1 FILLER_79_89 ();
 sg13g2_fill_8 FILLER_79_125 ();
 sg13g2_fill_8 FILLER_79_133 ();
 sg13g2_fill_8 FILLER_79_141 ();
 sg13g2_fill_8 FILLER_79_149 ();
 sg13g2_fill_8 FILLER_79_157 ();
 sg13g2_fill_8 FILLER_79_165 ();
 sg13g2_fill_8 FILLER_79_173 ();
 sg13g2_fill_2 FILLER_79_181 ();
 sg13g2_fill_1 FILLER_79_183 ();
 sg13g2_fill_8 FILLER_79_189 ();
 sg13g2_fill_8 FILLER_79_197 ();
 sg13g2_fill_2 FILLER_79_205 ();
 sg13g2_fill_1 FILLER_79_207 ();
 sg13g2_fill_2 FILLER_79_240 ();
 sg13g2_fill_8 FILLER_79_252 ();
 sg13g2_fill_8 FILLER_79_351 ();
 sg13g2_fill_4 FILLER_79_359 ();
 sg13g2_fill_2 FILLER_79_373 ();
 sg13g2_fill_8 FILLER_79_385 ();
 sg13g2_fill_8 FILLER_79_419 ();
 sg13g2_fill_1 FILLER_79_453 ();
 sg13g2_fill_8 FILLER_79_463 ();
 sg13g2_fill_4 FILLER_79_479 ();
 sg13g2_fill_1 FILLER_79_483 ();
 sg13g2_fill_8 FILLER_79_489 ();
 sg13g2_fill_2 FILLER_79_497 ();
 sg13g2_fill_8 FILLER_79_525 ();
 sg13g2_fill_4 FILLER_79_553 ();
 sg13g2_fill_2 FILLER_79_557 ();
 sg13g2_fill_8 FILLER_79_567 ();
 sg13g2_fill_8 FILLER_79_575 ();
 sg13g2_fill_8 FILLER_79_583 ();
 sg13g2_fill_8 FILLER_79_591 ();
 sg13g2_fill_8 FILLER_79_599 ();
 sg13g2_fill_1 FILLER_79_615 ();
 sg13g2_fill_8 FILLER_79_641 ();
 sg13g2_fill_8 FILLER_79_649 ();
 sg13g2_fill_1 FILLER_79_665 ();
 sg13g2_fill_2 FILLER_79_686 ();
 sg13g2_fill_8 FILLER_79_692 ();
 sg13g2_fill_4 FILLER_79_700 ();
 sg13g2_fill_4 FILLER_79_713 ();
 sg13g2_fill_2 FILLER_79_717 ();
 sg13g2_fill_1 FILLER_79_719 ();
 sg13g2_fill_8 FILLER_79_748 ();
 sg13g2_fill_8 FILLER_79_756 ();
 sg13g2_fill_8 FILLER_79_764 ();
 sg13g2_fill_8 FILLER_79_772 ();
 sg13g2_fill_8 FILLER_79_780 ();
 sg13g2_fill_8 FILLER_79_788 ();
 sg13g2_fill_2 FILLER_79_796 ();
 sg13g2_fill_8 FILLER_79_834 ();
 sg13g2_fill_4 FILLER_79_842 ();
 sg13g2_fill_2 FILLER_79_846 ();
 sg13g2_fill_1 FILLER_79_848 ();
 sg13g2_fill_8 FILLER_79_857 ();
 sg13g2_fill_8 FILLER_79_865 ();
 sg13g2_fill_2 FILLER_79_873 ();
 sg13g2_fill_1 FILLER_79_875 ();
 sg13g2_fill_2 FILLER_79_886 ();
 sg13g2_fill_1 FILLER_79_888 ();
 sg13g2_fill_1 FILLER_79_897 ();
 sg13g2_fill_2 FILLER_79_916 ();
 sg13g2_fill_2 FILLER_79_973 ();
 sg13g2_fill_1 FILLER_79_985 ();
 sg13g2_fill_1 FILLER_79_1038 ();
 sg13g2_fill_2 FILLER_79_1048 ();
 sg13g2_fill_1 FILLER_79_1085 ();
 sg13g2_fill_1 FILLER_79_1096 ();
 sg13g2_fill_1 FILLER_79_1101 ();
 sg13g2_fill_2 FILLER_79_1114 ();
 sg13g2_fill_4 FILLER_79_1136 ();
 sg13g2_fill_2 FILLER_79_1149 ();
 sg13g2_fill_1 FILLER_79_1169 ();
 sg13g2_fill_2 FILLER_79_1182 ();
 sg13g2_fill_1 FILLER_79_1184 ();
 sg13g2_fill_4 FILLER_79_1227 ();
 sg13g2_fill_1 FILLER_79_1231 ();
 sg13g2_fill_8 FILLER_79_1240 ();
 sg13g2_fill_1 FILLER_79_1248 ();
 sg13g2_fill_4 FILLER_79_1277 ();
 sg13g2_fill_2 FILLER_79_1281 ();
 sg13g2_fill_1 FILLER_79_1283 ();
 sg13g2_fill_1 FILLER_79_1290 ();
 sg13g2_fill_8 FILLER_79_1295 ();
 sg13g2_fill_8 FILLER_79_1303 ();
 sg13g2_fill_1 FILLER_79_1334 ();
 sg13g2_fill_2 FILLER_79_1340 ();
 sg13g2_fill_1 FILLER_79_1342 ();
 sg13g2_fill_8 FILLER_79_1353 ();
 sg13g2_fill_8 FILLER_79_1361 ();
 sg13g2_fill_1 FILLER_79_1369 ();
 sg13g2_fill_1 FILLER_79_1385 ();
 sg13g2_fill_2 FILLER_79_1407 ();
 sg13g2_fill_1 FILLER_79_1409 ();
 sg13g2_fill_8 FILLER_79_1436 ();
 sg13g2_fill_2 FILLER_79_1444 ();
 sg13g2_fill_4 FILLER_79_1454 ();
 sg13g2_fill_2 FILLER_79_1458 ();
 sg13g2_fill_1 FILLER_79_1460 ();
 sg13g2_fill_2 FILLER_79_1491 ();
 sg13g2_fill_1 FILLER_79_1493 ();
 sg13g2_fill_1 FILLER_79_1510 ();
 sg13g2_fill_2 FILLER_79_1516 ();
 sg13g2_fill_8 FILLER_79_1548 ();
 sg13g2_fill_4 FILLER_79_1556 ();
 sg13g2_fill_2 FILLER_79_1560 ();
 sg13g2_fill_8 FILLER_80_0 ();
 sg13g2_fill_8 FILLER_80_8 ();
 sg13g2_fill_8 FILLER_80_16 ();
 sg13g2_fill_2 FILLER_80_24 ();
 sg13g2_fill_8 FILLER_80_36 ();
 sg13g2_fill_8 FILLER_80_44 ();
 sg13g2_fill_1 FILLER_80_52 ();
 sg13g2_fill_4 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_103 ();
 sg13g2_fill_1 FILLER_80_105 ();
 sg13g2_fill_8 FILLER_80_116 ();
 sg13g2_fill_8 FILLER_80_134 ();
 sg13g2_fill_8 FILLER_80_142 ();
 sg13g2_fill_4 FILLER_80_171 ();
 sg13g2_fill_1 FILLER_80_175 ();
 sg13g2_fill_2 FILLER_80_184 ();
 sg13g2_fill_1 FILLER_80_186 ();
 sg13g2_fill_8 FILLER_80_200 ();
 sg13g2_fill_2 FILLER_80_208 ();
 sg13g2_fill_8 FILLER_80_218 ();
 sg13g2_fill_8 FILLER_80_226 ();
 sg13g2_fill_8 FILLER_80_234 ();
 sg13g2_fill_8 FILLER_80_242 ();
 sg13g2_fill_8 FILLER_80_250 ();
 sg13g2_fill_8 FILLER_80_258 ();
 sg13g2_fill_4 FILLER_80_266 ();
 sg13g2_fill_2 FILLER_80_270 ();
 sg13g2_fill_1 FILLER_80_272 ();
 sg13g2_fill_8 FILLER_80_283 ();
 sg13g2_fill_4 FILLER_80_291 ();
 sg13g2_fill_8 FILLER_80_300 ();
 sg13g2_fill_8 FILLER_80_308 ();
 sg13g2_fill_8 FILLER_80_316 ();
 sg13g2_fill_4 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_364 ();
 sg13g2_fill_4 FILLER_80_392 ();
 sg13g2_fill_2 FILLER_80_396 ();
 sg13g2_fill_8 FILLER_80_429 ();
 sg13g2_fill_4 FILLER_80_437 ();
 sg13g2_fill_2 FILLER_80_441 ();
 sg13g2_fill_1 FILLER_80_443 ();
 sg13g2_fill_4 FILLER_80_490 ();
 sg13g2_fill_8 FILLER_80_504 ();
 sg13g2_fill_8 FILLER_80_512 ();
 sg13g2_fill_2 FILLER_80_520 ();
 sg13g2_fill_1 FILLER_80_522 ();
 sg13g2_fill_4 FILLER_80_595 ();
 sg13g2_fill_1 FILLER_80_599 ();
 sg13g2_fill_4 FILLER_80_610 ();
 sg13g2_fill_2 FILLER_80_614 ();
 sg13g2_fill_1 FILLER_80_616 ();
 sg13g2_fill_4 FILLER_80_658 ();
 sg13g2_fill_1 FILLER_80_669 ();
 sg13g2_fill_1 FILLER_80_677 ();
 sg13g2_fill_4 FILLER_80_731 ();
 sg13g2_fill_2 FILLER_80_735 ();
 sg13g2_fill_4 FILLER_80_767 ();
 sg13g2_fill_2 FILLER_80_771 ();
 sg13g2_fill_1 FILLER_80_773 ();
 sg13g2_fill_8 FILLER_80_800 ();
 sg13g2_fill_1 FILLER_80_808 ();
 sg13g2_fill_8 FILLER_80_830 ();
 sg13g2_fill_4 FILLER_80_838 ();
 sg13g2_fill_2 FILLER_80_842 ();
 sg13g2_fill_2 FILLER_80_884 ();
 sg13g2_fill_1 FILLER_80_886 ();
 sg13g2_fill_2 FILLER_80_900 ();
 sg13g2_fill_1 FILLER_80_934 ();
 sg13g2_fill_2 FILLER_80_947 ();
 sg13g2_fill_2 FILLER_80_965 ();
 sg13g2_fill_1 FILLER_80_1046 ();
 sg13g2_fill_2 FILLER_80_1077 ();
 sg13g2_fill_2 FILLER_80_1104 ();
 sg13g2_fill_2 FILLER_80_1130 ();
 sg13g2_fill_1 FILLER_80_1132 ();
 sg13g2_fill_8 FILLER_80_1141 ();
 sg13g2_fill_1 FILLER_80_1149 ();
 sg13g2_fill_4 FILLER_80_1158 ();
 sg13g2_fill_2 FILLER_80_1162 ();
 sg13g2_fill_8 FILLER_80_1177 ();
 sg13g2_fill_4 FILLER_80_1185 ();
 sg13g2_fill_1 FILLER_80_1189 ();
 sg13g2_fill_2 FILLER_80_1194 ();
 sg13g2_fill_4 FILLER_80_1204 ();
 sg13g2_fill_1 FILLER_80_1208 ();
 sg13g2_fill_2 FILLER_80_1213 ();
 sg13g2_fill_4 FILLER_80_1228 ();
 sg13g2_fill_2 FILLER_80_1232 ();
 sg13g2_fill_1 FILLER_80_1258 ();
 sg13g2_fill_8 FILLER_80_1278 ();
 sg13g2_fill_1 FILLER_80_1286 ();
 sg13g2_fill_2 FILLER_80_1295 ();
 sg13g2_fill_8 FILLER_80_1302 ();
 sg13g2_fill_8 FILLER_80_1310 ();
 sg13g2_fill_1 FILLER_80_1318 ();
 sg13g2_fill_4 FILLER_80_1327 ();
 sg13g2_fill_8 FILLER_80_1349 ();
 sg13g2_fill_8 FILLER_80_1357 ();
 sg13g2_fill_1 FILLER_80_1369 ();
 sg13g2_fill_1 FILLER_80_1377 ();
 sg13g2_fill_2 FILLER_80_1407 ();
 sg13g2_fill_1 FILLER_80_1414 ();
 sg13g2_fill_8 FILLER_80_1461 ();
 sg13g2_fill_4 FILLER_80_1469 ();
 sg13g2_fill_1 FILLER_80_1473 ();
 sg13g2_fill_8 FILLER_80_1487 ();
 sg13g2_fill_4 FILLER_80_1495 ();
 sg13g2_fill_8 FILLER_80_1518 ();
 sg13g2_fill_8 FILLER_80_1526 ();
 sg13g2_fill_2 FILLER_80_1534 ();
 sg13g2_fill_1 FILLER_80_1536 ();
 sg13g2_fill_8 FILLER_80_1580 ();
 sg13g2_fill_4 FILLER_80_1588 ();
 sg13g2_fill_8 FILLER_81_0 ();
 sg13g2_fill_8 FILLER_81_8 ();
 sg13g2_fill_8 FILLER_81_16 ();
 sg13g2_fill_8 FILLER_81_24 ();
 sg13g2_fill_8 FILLER_81_32 ();
 sg13g2_fill_8 FILLER_81_40 ();
 sg13g2_fill_8 FILLER_81_48 ();
 sg13g2_fill_2 FILLER_81_56 ();
 sg13g2_fill_1 FILLER_81_58 ();
 sg13g2_fill_8 FILLER_81_81 ();
 sg13g2_fill_4 FILLER_81_89 ();
 sg13g2_fill_1 FILLER_81_93 ();
 sg13g2_fill_4 FILLER_81_120 ();
 sg13g2_fill_2 FILLER_81_124 ();
 sg13g2_fill_1 FILLER_81_126 ();
 sg13g2_fill_4 FILLER_81_174 ();
 sg13g2_fill_2 FILLER_81_178 ();
 sg13g2_fill_8 FILLER_81_216 ();
 sg13g2_fill_4 FILLER_81_224 ();
 sg13g2_fill_1 FILLER_81_228 ();
 sg13g2_fill_4 FILLER_81_263 ();
 sg13g2_fill_2 FILLER_81_267 ();
 sg13g2_fill_1 FILLER_81_269 ();
 sg13g2_fill_8 FILLER_81_280 ();
 sg13g2_fill_8 FILLER_81_288 ();
 sg13g2_fill_8 FILLER_81_296 ();
 sg13g2_fill_8 FILLER_81_304 ();
 sg13g2_fill_8 FILLER_81_312 ();
 sg13g2_fill_2 FILLER_81_320 ();
 sg13g2_fill_1 FILLER_81_322 ();
 sg13g2_fill_4 FILLER_81_331 ();
 sg13g2_fill_1 FILLER_81_335 ();
 sg13g2_fill_1 FILLER_81_362 ();
 sg13g2_fill_2 FILLER_81_404 ();
 sg13g2_fill_1 FILLER_81_406 ();
 sg13g2_fill_8 FILLER_81_410 ();
 sg13g2_fill_2 FILLER_81_418 ();
 sg13g2_fill_1 FILLER_81_420 ();
 sg13g2_fill_4 FILLER_81_441 ();
 sg13g2_fill_2 FILLER_81_445 ();
 sg13g2_fill_8 FILLER_81_461 ();
 sg13g2_fill_8 FILLER_81_479 ();
 sg13g2_fill_8 FILLER_81_487 ();
 sg13g2_fill_2 FILLER_81_495 ();
 sg13g2_fill_4 FILLER_81_507 ();
 sg13g2_fill_1 FILLER_81_511 ();
 sg13g2_fill_8 FILLER_81_519 ();
 sg13g2_fill_8 FILLER_81_527 ();
 sg13g2_fill_2 FILLER_81_535 ();
 sg13g2_fill_2 FILLER_81_549 ();
 sg13g2_fill_1 FILLER_81_551 ();
 sg13g2_fill_8 FILLER_81_638 ();
 sg13g2_fill_8 FILLER_81_646 ();
 sg13g2_fill_8 FILLER_81_654 ();
 sg13g2_fill_4 FILLER_81_662 ();
 sg13g2_fill_2 FILLER_81_666 ();
 sg13g2_fill_8 FILLER_81_681 ();
 sg13g2_fill_8 FILLER_81_689 ();
 sg13g2_fill_8 FILLER_81_697 ();
 sg13g2_fill_4 FILLER_81_705 ();
 sg13g2_fill_2 FILLER_81_709 ();
 sg13g2_fill_1 FILLER_81_711 ();
 sg13g2_fill_4 FILLER_81_718 ();
 sg13g2_fill_1 FILLER_81_722 ();
 sg13g2_fill_8 FILLER_81_736 ();
 sg13g2_fill_4 FILLER_81_744 ();
 sg13g2_fill_8 FILLER_81_763 ();
 sg13g2_fill_4 FILLER_81_781 ();
 sg13g2_fill_2 FILLER_81_785 ();
 sg13g2_fill_4 FILLER_81_818 ();
 sg13g2_fill_8 FILLER_81_858 ();
 sg13g2_fill_8 FILLER_81_866 ();
 sg13g2_fill_4 FILLER_81_874 ();
 sg13g2_fill_1 FILLER_81_878 ();
 sg13g2_fill_2 FILLER_81_889 ();
 sg13g2_fill_2 FILLER_81_954 ();
 sg13g2_fill_1 FILLER_81_973 ();
 sg13g2_fill_1 FILLER_81_982 ();
 sg13g2_fill_2 FILLER_81_1058 ();
 sg13g2_fill_1 FILLER_81_1086 ();
 sg13g2_fill_8 FILLER_81_1113 ();
 sg13g2_fill_2 FILLER_81_1121 ();
 sg13g2_fill_1 FILLER_81_1128 ();
 sg13g2_fill_8 FILLER_81_1164 ();
 sg13g2_fill_8 FILLER_81_1172 ();
 sg13g2_fill_1 FILLER_81_1180 ();
 sg13g2_fill_4 FILLER_81_1196 ();
 sg13g2_fill_2 FILLER_81_1204 ();
 sg13g2_fill_1 FILLER_81_1206 ();
 sg13g2_fill_2 FILLER_81_1225 ();
 sg13g2_fill_8 FILLER_81_1236 ();
 sg13g2_fill_8 FILLER_81_1244 ();
 sg13g2_fill_1 FILLER_81_1252 ();
 sg13g2_fill_8 FILLER_81_1258 ();
 sg13g2_fill_4 FILLER_81_1270 ();
 sg13g2_fill_1 FILLER_81_1274 ();
 sg13g2_fill_1 FILLER_81_1296 ();
 sg13g2_fill_4 FILLER_81_1305 ();
 sg13g2_fill_2 FILLER_81_1309 ();
 sg13g2_fill_1 FILLER_81_1311 ();
 sg13g2_fill_1 FILLER_81_1330 ();
 sg13g2_fill_4 FILLER_81_1334 ();
 sg13g2_fill_2 FILLER_81_1338 ();
 sg13g2_fill_1 FILLER_81_1340 ();
 sg13g2_fill_4 FILLER_81_1359 ();
 sg13g2_fill_8 FILLER_81_1378 ();
 sg13g2_fill_2 FILLER_81_1386 ();
 sg13g2_fill_1 FILLER_81_1388 ();
 sg13g2_fill_2 FILLER_81_1393 ();
 sg13g2_fill_1 FILLER_81_1395 ();
 sg13g2_fill_4 FILLER_81_1405 ();
 sg13g2_fill_1 FILLER_81_1409 ();
 sg13g2_fill_4 FILLER_81_1461 ();
 sg13g2_fill_1 FILLER_81_1465 ();
 sg13g2_fill_8 FILLER_81_1474 ();
 sg13g2_fill_4 FILLER_81_1482 ();
 sg13g2_fill_2 FILLER_81_1486 ();
 sg13g2_fill_8 FILLER_81_1499 ();
 sg13g2_fill_8 FILLER_81_1507 ();
 sg13g2_fill_4 FILLER_81_1515 ();
 sg13g2_fill_8 FILLER_81_1527 ();
 sg13g2_fill_8 FILLER_81_1541 ();
 sg13g2_fill_8 FILLER_81_1549 ();
 sg13g2_fill_2 FILLER_81_1557 ();
 sg13g2_fill_8 FILLER_81_1584 ();
 sg13g2_fill_8 FILLER_82_0 ();
 sg13g2_fill_8 FILLER_82_8 ();
 sg13g2_fill_8 FILLER_82_16 ();
 sg13g2_fill_2 FILLER_82_24 ();
 sg13g2_fill_4 FILLER_82_52 ();
 sg13g2_fill_8 FILLER_82_92 ();
 sg13g2_fill_8 FILLER_82_100 ();
 sg13g2_fill_8 FILLER_82_108 ();
 sg13g2_fill_4 FILLER_82_116 ();
 sg13g2_fill_1 FILLER_82_120 ();
 sg13g2_fill_8 FILLER_82_167 ();
 sg13g2_fill_4 FILLER_82_175 ();
 sg13g2_fill_8 FILLER_82_205 ();
 sg13g2_fill_8 FILLER_82_213 ();
 sg13g2_fill_4 FILLER_82_221 ();
 sg13g2_fill_8 FILLER_82_235 ();
 sg13g2_fill_2 FILLER_82_243 ();
 sg13g2_fill_1 FILLER_82_245 ();
 sg13g2_fill_1 FILLER_82_256 ();
 sg13g2_fill_2 FILLER_82_283 ();
 sg13g2_fill_8 FILLER_82_311 ();
 sg13g2_fill_8 FILLER_82_319 ();
 sg13g2_fill_2 FILLER_82_327 ();
 sg13g2_fill_1 FILLER_82_329 ();
 sg13g2_fill_8 FILLER_82_340 ();
 sg13g2_fill_8 FILLER_82_348 ();
 sg13g2_fill_1 FILLER_82_356 ();
 sg13g2_fill_8 FILLER_82_403 ();
 sg13g2_fill_4 FILLER_82_411 ();
 sg13g2_fill_4 FILLER_82_423 ();
 sg13g2_fill_2 FILLER_82_427 ();
 sg13g2_fill_1 FILLER_82_444 ();
 sg13g2_fill_8 FILLER_82_455 ();
 sg13g2_fill_4 FILLER_82_463 ();
 sg13g2_fill_2 FILLER_82_467 ();
 sg13g2_fill_8 FILLER_82_495 ();
 sg13g2_fill_8 FILLER_82_529 ();
 sg13g2_fill_4 FILLER_82_537 ();
 sg13g2_fill_2 FILLER_82_541 ();
 sg13g2_fill_2 FILLER_82_572 ();
 sg13g2_fill_1 FILLER_82_574 ();
 sg13g2_fill_8 FILLER_82_585 ();
 sg13g2_fill_2 FILLER_82_593 ();
 sg13g2_fill_8 FILLER_82_603 ();
 sg13g2_fill_1 FILLER_82_611 ();
 sg13g2_fill_4 FILLER_82_632 ();
 sg13g2_fill_4 FILLER_82_662 ();
 sg13g2_fill_8 FILLER_82_696 ();
 sg13g2_fill_4 FILLER_82_704 ();
 sg13g2_fill_2 FILLER_82_708 ();
 sg13g2_fill_2 FILLER_82_718 ();
 sg13g2_fill_4 FILLER_82_724 ();
 sg13g2_fill_2 FILLER_82_728 ();
 sg13g2_fill_1 FILLER_82_730 ();
 sg13g2_fill_2 FILLER_82_739 ();
 sg13g2_fill_2 FILLER_82_749 ();
 sg13g2_fill_4 FILLER_82_776 ();
 sg13g2_fill_1 FILLER_82_780 ();
 sg13g2_fill_8 FILLER_82_799 ();
 sg13g2_fill_8 FILLER_82_807 ();
 sg13g2_fill_2 FILLER_82_815 ();
 sg13g2_fill_1 FILLER_82_817 ();
 sg13g2_fill_8 FILLER_82_834 ();
 sg13g2_fill_4 FILLER_82_842 ();
 sg13g2_fill_4 FILLER_82_851 ();
 sg13g2_fill_2 FILLER_82_868 ();
 sg13g2_fill_1 FILLER_82_870 ();
 sg13g2_fill_1 FILLER_82_909 ();
 sg13g2_fill_1 FILLER_82_931 ();
 sg13g2_fill_1 FILLER_82_1033 ();
 sg13g2_fill_4 FILLER_82_1105 ();
 sg13g2_fill_1 FILLER_82_1109 ();
 sg13g2_fill_8 FILLER_82_1114 ();
 sg13g2_fill_4 FILLER_82_1122 ();
 sg13g2_fill_2 FILLER_82_1126 ();
 sg13g2_fill_2 FILLER_82_1138 ();
 sg13g2_fill_8 FILLER_82_1144 ();
 sg13g2_fill_4 FILLER_82_1156 ();
 sg13g2_fill_2 FILLER_82_1160 ();
 sg13g2_fill_1 FILLER_82_1162 ();
 sg13g2_fill_8 FILLER_82_1169 ();
 sg13g2_fill_1 FILLER_82_1182 ();
 sg13g2_fill_4 FILLER_82_1188 ();
 sg13g2_fill_1 FILLER_82_1192 ();
 sg13g2_fill_2 FILLER_82_1198 ();
 sg13g2_fill_1 FILLER_82_1200 ();
 sg13g2_fill_2 FILLER_82_1220 ();
 sg13g2_fill_1 FILLER_82_1222 ();
 sg13g2_fill_4 FILLER_82_1240 ();
 sg13g2_fill_1 FILLER_82_1244 ();
 sg13g2_fill_8 FILLER_82_1268 ();
 sg13g2_fill_4 FILLER_82_1276 ();
 sg13g2_fill_2 FILLER_82_1280 ();
 sg13g2_fill_4 FILLER_82_1297 ();
 sg13g2_fill_1 FILLER_82_1301 ();
 sg13g2_fill_8 FILLER_82_1324 ();
 sg13g2_fill_1 FILLER_82_1332 ();
 sg13g2_fill_2 FILLER_82_1338 ();
 sg13g2_fill_1 FILLER_82_1340 ();
 sg13g2_fill_2 FILLER_82_1367 ();
 sg13g2_fill_1 FILLER_82_1369 ();
 sg13g2_fill_2 FILLER_82_1373 ();
 sg13g2_fill_1 FILLER_82_1375 ();
 sg13g2_fill_1 FILLER_82_1381 ();
 sg13g2_fill_1 FILLER_82_1387 ();
 sg13g2_fill_1 FILLER_82_1391 ();
 sg13g2_fill_1 FILLER_82_1423 ();
 sg13g2_fill_8 FILLER_82_1428 ();
 sg13g2_fill_8 FILLER_82_1436 ();
 sg13g2_fill_8 FILLER_82_1444 ();
 sg13g2_fill_4 FILLER_82_1452 ();
 sg13g2_fill_1 FILLER_82_1456 ();
 sg13g2_fill_8 FILLER_82_1514 ();
 sg13g2_fill_1 FILLER_82_1522 ();
 sg13g2_fill_8 FILLER_82_1528 ();
 sg13g2_fill_4 FILLER_82_1536 ();
 sg13g2_fill_1 FILLER_82_1540 ();
 sg13g2_fill_8 FILLER_82_1549 ();
 sg13g2_fill_4 FILLER_82_1557 ();
 sg13g2_fill_1 FILLER_82_1561 ();
 sg13g2_fill_8 FILLER_83_0 ();
 sg13g2_fill_8 FILLER_83_8 ();
 sg13g2_fill_4 FILLER_83_16 ();
 sg13g2_fill_4 FILLER_83_56 ();
 sg13g2_fill_1 FILLER_83_60 ();
 sg13g2_fill_2 FILLER_83_74 ();
 sg13g2_fill_4 FILLER_83_101 ();
 sg13g2_fill_8 FILLER_83_131 ();
 sg13g2_fill_8 FILLER_83_139 ();
 sg13g2_fill_1 FILLER_83_147 ();
 sg13g2_fill_2 FILLER_83_173 ();
 sg13g2_fill_4 FILLER_83_185 ();
 sg13g2_fill_2 FILLER_83_189 ();
 sg13g2_fill_2 FILLER_83_261 ();
 sg13g2_fill_1 FILLER_83_335 ();
 sg13g2_fill_4 FILLER_83_362 ();
 sg13g2_fill_1 FILLER_83_366 ();
 sg13g2_fill_2 FILLER_83_392 ();
 sg13g2_fill_1 FILLER_83_394 ();
 sg13g2_fill_8 FILLER_83_466 ();
 sg13g2_fill_4 FILLER_83_474 ();
 sg13g2_fill_8 FILLER_83_483 ();
 sg13g2_fill_4 FILLER_83_491 ();
 sg13g2_fill_2 FILLER_83_495 ();
 sg13g2_fill_1 FILLER_83_497 ();
 sg13g2_fill_8 FILLER_83_511 ();
 sg13g2_fill_4 FILLER_83_519 ();
 sg13g2_fill_4 FILLER_83_565 ();
 sg13g2_fill_2 FILLER_83_569 ();
 sg13g2_fill_2 FILLER_83_581 ();
 sg13g2_fill_8 FILLER_83_593 ();
 sg13g2_fill_8 FILLER_83_601 ();
 sg13g2_fill_8 FILLER_83_609 ();
 sg13g2_fill_4 FILLER_83_617 ();
 sg13g2_fill_1 FILLER_83_637 ();
 sg13g2_fill_8 FILLER_83_671 ();
 sg13g2_fill_4 FILLER_83_679 ();
 sg13g2_fill_2 FILLER_83_789 ();
 sg13g2_fill_1 FILLER_83_791 ();
 sg13g2_fill_8 FILLER_83_802 ();
 sg13g2_fill_4 FILLER_83_815 ();
 sg13g2_fill_4 FILLER_83_832 ();
 sg13g2_fill_1 FILLER_83_836 ();
 sg13g2_fill_8 FILLER_83_863 ();
 sg13g2_fill_8 FILLER_83_871 ();
 sg13g2_fill_8 FILLER_83_879 ();
 sg13g2_fill_4 FILLER_83_887 ();
 sg13g2_fill_2 FILLER_83_891 ();
 sg13g2_fill_1 FILLER_83_893 ();
 sg13g2_fill_4 FILLER_83_897 ();
 sg13g2_fill_1 FILLER_83_901 ();
 sg13g2_fill_1 FILLER_83_912 ();
 sg13g2_fill_8 FILLER_83_924 ();
 sg13g2_fill_2 FILLER_83_932 ();
 sg13g2_fill_1 FILLER_83_934 ();
 sg13g2_fill_2 FILLER_83_964 ();
 sg13g2_fill_1 FILLER_83_971 ();
 sg13g2_fill_1 FILLER_83_981 ();
 sg13g2_fill_2 FILLER_83_1030 ();
 sg13g2_fill_2 FILLER_83_1040 ();
 sg13g2_fill_1 FILLER_83_1058 ();
 sg13g2_fill_1 FILLER_83_1067 ();
 sg13g2_fill_1 FILLER_83_1073 ();
 sg13g2_fill_2 FILLER_83_1124 ();
 sg13g2_fill_1 FILLER_83_1126 ();
 sg13g2_fill_8 FILLER_83_1149 ();
 sg13g2_fill_8 FILLER_83_1157 ();
 sg13g2_fill_4 FILLER_83_1165 ();
 sg13g2_fill_1 FILLER_83_1169 ();
 sg13g2_fill_8 FILLER_83_1191 ();
 sg13g2_fill_8 FILLER_83_1199 ();
 sg13g2_fill_8 FILLER_83_1207 ();
 sg13g2_fill_4 FILLER_83_1220 ();
 sg13g2_fill_8 FILLER_83_1228 ();
 sg13g2_fill_4 FILLER_83_1236 ();
 sg13g2_fill_1 FILLER_83_1240 ();
 sg13g2_fill_4 FILLER_83_1274 ();
 sg13g2_fill_2 FILLER_83_1278 ();
 sg13g2_fill_1 FILLER_83_1280 ();
 sg13g2_fill_2 FILLER_83_1300 ();
 sg13g2_fill_1 FILLER_83_1302 ();
 sg13g2_fill_8 FILLER_83_1307 ();
 sg13g2_fill_2 FILLER_83_1315 ();
 sg13g2_fill_8 FILLER_83_1321 ();
 sg13g2_fill_4 FILLER_83_1329 ();
 sg13g2_fill_2 FILLER_83_1333 ();
 sg13g2_fill_8 FILLER_83_1357 ();
 sg13g2_fill_4 FILLER_83_1365 ();
 sg13g2_fill_2 FILLER_83_1369 ();
 sg13g2_fill_1 FILLER_83_1376 ();
 sg13g2_fill_2 FILLER_83_1382 ();
 sg13g2_fill_1 FILLER_83_1384 ();
 sg13g2_fill_8 FILLER_83_1396 ();
 sg13g2_fill_8 FILLER_83_1404 ();
 sg13g2_fill_4 FILLER_83_1412 ();
 sg13g2_fill_2 FILLER_83_1416 ();
 sg13g2_fill_2 FILLER_83_1427 ();
 sg13g2_fill_1 FILLER_83_1429 ();
 sg13g2_fill_4 FILLER_83_1456 ();
 sg13g2_fill_2 FILLER_83_1460 ();
 sg13g2_fill_1 FILLER_83_1462 ();
 sg13g2_fill_1 FILLER_83_1472 ();
 sg13g2_fill_2 FILLER_83_1508 ();
 sg13g2_fill_2 FILLER_83_1553 ();
 sg13g2_fill_1 FILLER_83_1555 ();
 sg13g2_fill_4 FILLER_83_1586 ();
 sg13g2_fill_2 FILLER_83_1590 ();
 sg13g2_fill_8 FILLER_84_0 ();
 sg13g2_fill_8 FILLER_84_8 ();
 sg13g2_fill_8 FILLER_84_16 ();
 sg13g2_fill_2 FILLER_84_24 ();
 sg13g2_fill_1 FILLER_84_26 ();
 sg13g2_fill_8 FILLER_84_37 ();
 sg13g2_fill_4 FILLER_84_45 ();
 sg13g2_fill_1 FILLER_84_49 ();
 sg13g2_fill_1 FILLER_84_60 ();
 sg13g2_fill_2 FILLER_84_96 ();
 sg13g2_fill_8 FILLER_84_104 ();
 sg13g2_fill_8 FILLER_84_112 ();
 sg13g2_fill_8 FILLER_84_120 ();
 sg13g2_fill_2 FILLER_84_128 ();
 sg13g2_fill_8 FILLER_84_140 ();
 sg13g2_fill_8 FILLER_84_148 ();
 sg13g2_fill_8 FILLER_84_156 ();
 sg13g2_fill_2 FILLER_84_164 ();
 sg13g2_fill_8 FILLER_84_174 ();
 sg13g2_fill_2 FILLER_84_182 ();
 sg13g2_fill_1 FILLER_84_184 ();
 sg13g2_fill_8 FILLER_84_195 ();
 sg13g2_fill_4 FILLER_84_203 ();
 sg13g2_fill_2 FILLER_84_207 ();
 sg13g2_fill_2 FILLER_84_217 ();
 sg13g2_fill_1 FILLER_84_219 ();
 sg13g2_fill_8 FILLER_84_230 ();
 sg13g2_fill_8 FILLER_84_238 ();
 sg13g2_fill_8 FILLER_84_246 ();
 sg13g2_fill_8 FILLER_84_254 ();
 sg13g2_fill_8 FILLER_84_262 ();
 sg13g2_fill_4 FILLER_84_270 ();
 sg13g2_fill_2 FILLER_84_274 ();
 sg13g2_fill_8 FILLER_84_296 ();
 sg13g2_fill_2 FILLER_84_304 ();
 sg13g2_fill_2 FILLER_84_327 ();
 sg13g2_fill_1 FILLER_84_329 ();
 sg13g2_fill_1 FILLER_84_366 ();
 sg13g2_fill_2 FILLER_84_399 ();
 sg13g2_fill_1 FILLER_84_401 ();
 sg13g2_fill_8 FILLER_84_418 ();
 sg13g2_fill_8 FILLER_84_426 ();
 sg13g2_fill_8 FILLER_84_434 ();
 sg13g2_fill_4 FILLER_84_442 ();
 sg13g2_fill_2 FILLER_84_460 ();
 sg13g2_fill_1 FILLER_84_462 ();
 sg13g2_fill_8 FILLER_84_499 ();
 sg13g2_fill_4 FILLER_84_507 ();
 sg13g2_fill_2 FILLER_84_511 ();
 sg13g2_fill_1 FILLER_84_513 ();
 sg13g2_fill_1 FILLER_84_550 ();
 sg13g2_fill_8 FILLER_84_574 ();
 sg13g2_fill_2 FILLER_84_582 ();
 sg13g2_fill_8 FILLER_84_592 ();
 sg13g2_fill_4 FILLER_84_608 ();
 sg13g2_fill_2 FILLER_84_612 ();
 sg13g2_fill_4 FILLER_84_622 ();
 sg13g2_fill_2 FILLER_84_631 ();
 sg13g2_fill_8 FILLER_84_682 ();
 sg13g2_fill_8 FILLER_84_690 ();
 sg13g2_fill_8 FILLER_84_698 ();
 sg13g2_fill_8 FILLER_84_706 ();
 sg13g2_fill_8 FILLER_84_714 ();
 sg13g2_fill_2 FILLER_84_722 ();
 sg13g2_fill_1 FILLER_84_724 ();
 sg13g2_fill_8 FILLER_84_738 ();
 sg13g2_fill_8 FILLER_84_746 ();
 sg13g2_fill_4 FILLER_84_754 ();
 sg13g2_fill_2 FILLER_84_758 ();
 sg13g2_fill_1 FILLER_84_760 ();
 sg13g2_fill_8 FILLER_84_787 ();
 sg13g2_fill_8 FILLER_84_821 ();
 sg13g2_fill_4 FILLER_84_829 ();
 sg13g2_fill_1 FILLER_84_833 ();
 sg13g2_fill_1 FILLER_84_844 ();
 sg13g2_fill_2 FILLER_84_902 ();
 sg13g2_fill_8 FILLER_84_940 ();
 sg13g2_fill_2 FILLER_84_948 ();
 sg13g2_fill_1 FILLER_84_975 ();
 sg13g2_fill_2 FILLER_84_1005 ();
 sg13g2_fill_1 FILLER_84_1038 ();
 sg13g2_fill_1 FILLER_84_1044 ();
 sg13g2_fill_1 FILLER_84_1060 ();
 sg13g2_fill_2 FILLER_84_1090 ();
 sg13g2_fill_2 FILLER_84_1113 ();
 sg13g2_fill_1 FILLER_84_1123 ();
 sg13g2_fill_8 FILLER_84_1132 ();
 sg13g2_fill_2 FILLER_84_1140 ();
 sg13g2_fill_1 FILLER_84_1142 ();
 sg13g2_fill_8 FILLER_84_1148 ();
 sg13g2_fill_8 FILLER_84_1156 ();
 sg13g2_fill_2 FILLER_84_1164 ();
 sg13g2_fill_4 FILLER_84_1176 ();
 sg13g2_fill_2 FILLER_84_1180 ();
 sg13g2_fill_1 FILLER_84_1182 ();
 sg13g2_fill_2 FILLER_84_1193 ();
 sg13g2_fill_1 FILLER_84_1195 ();
 sg13g2_fill_8 FILLER_84_1236 ();
 sg13g2_fill_2 FILLER_84_1248 ();
 sg13g2_fill_8 FILLER_84_1254 ();
 sg13g2_fill_1 FILLER_84_1262 ();
 sg13g2_fill_8 FILLER_84_1277 ();
 sg13g2_fill_2 FILLER_84_1285 ();
 sg13g2_fill_1 FILLER_84_1287 ();
 sg13g2_fill_8 FILLER_84_1296 ();
 sg13g2_fill_2 FILLER_84_1304 ();
 sg13g2_fill_1 FILLER_84_1306 ();
 sg13g2_fill_4 FILLER_84_1336 ();
 sg13g2_fill_2 FILLER_84_1340 ();
 sg13g2_fill_1 FILLER_84_1342 ();
 sg13g2_fill_4 FILLER_84_1352 ();
 sg13g2_fill_2 FILLER_84_1356 ();
 sg13g2_fill_1 FILLER_84_1358 ();
 sg13g2_fill_2 FILLER_84_1381 ();
 sg13g2_fill_8 FILLER_84_1395 ();
 sg13g2_fill_8 FILLER_84_1403 ();
 sg13g2_fill_1 FILLER_84_1411 ();
 sg13g2_fill_2 FILLER_84_1417 ();
 sg13g2_fill_1 FILLER_84_1419 ();
 sg13g2_fill_1 FILLER_84_1467 ();
 sg13g2_fill_2 FILLER_84_1514 ();
 sg13g2_fill_2 FILLER_84_1523 ();
 sg13g2_fill_8 FILLER_84_1533 ();
 sg13g2_fill_4 FILLER_84_1541 ();
 sg13g2_fill_1 FILLER_84_1545 ();
 sg13g2_fill_8 FILLER_84_1551 ();
 sg13g2_fill_2 FILLER_84_1559 ();
 sg13g2_fill_1 FILLER_84_1561 ();
 sg13g2_fill_8 FILLER_85_0 ();
 sg13g2_fill_8 FILLER_85_8 ();
 sg13g2_fill_8 FILLER_85_16 ();
 sg13g2_fill_8 FILLER_85_24 ();
 sg13g2_fill_8 FILLER_85_32 ();
 sg13g2_fill_8 FILLER_85_40 ();
 sg13g2_fill_2 FILLER_85_48 ();
 sg13g2_fill_1 FILLER_85_50 ();
 sg13g2_fill_4 FILLER_85_77 ();
 sg13g2_fill_2 FILLER_85_81 ();
 sg13g2_fill_1 FILLER_85_104 ();
 sg13g2_fill_8 FILLER_85_186 ();
 sg13g2_fill_8 FILLER_85_194 ();
 sg13g2_fill_8 FILLER_85_202 ();
 sg13g2_fill_8 FILLER_85_210 ();
 sg13g2_fill_4 FILLER_85_218 ();
 sg13g2_fill_8 FILLER_85_232 ();
 sg13g2_fill_8 FILLER_85_240 ();
 sg13g2_fill_8 FILLER_85_274 ();
 sg13g2_fill_4 FILLER_85_282 ();
 sg13g2_fill_2 FILLER_85_294 ();
 sg13g2_fill_8 FILLER_85_342 ();
 sg13g2_fill_8 FILLER_85_350 ();
 sg13g2_fill_8 FILLER_85_358 ();
 sg13g2_fill_2 FILLER_85_366 ();
 sg13g2_fill_1 FILLER_85_383 ();
 sg13g2_fill_2 FILLER_85_391 ();
 sg13g2_fill_1 FILLER_85_393 ();
 sg13g2_fill_4 FILLER_85_430 ();
 sg13g2_fill_8 FILLER_85_472 ();
 sg13g2_fill_8 FILLER_85_480 ();
 sg13g2_fill_8 FILLER_85_498 ();
 sg13g2_fill_4 FILLER_85_506 ();
 sg13g2_fill_1 FILLER_85_510 ();
 sg13g2_fill_4 FILLER_85_526 ();
 sg13g2_fill_8 FILLER_85_540 ();
 sg13g2_fill_4 FILLER_85_548 ();
 sg13g2_fill_2 FILLER_85_552 ();
 sg13g2_fill_1 FILLER_85_554 ();
 sg13g2_fill_8 FILLER_85_565 ();
 sg13g2_fill_2 FILLER_85_573 ();
 sg13g2_fill_1 FILLER_85_575 ();
 sg13g2_fill_2 FILLER_85_593 ();
 sg13g2_fill_8 FILLER_85_637 ();
 sg13g2_fill_1 FILLER_85_645 ();
 sg13g2_fill_8 FILLER_85_652 ();
 sg13g2_fill_4 FILLER_85_660 ();
 sg13g2_fill_1 FILLER_85_664 ();
 sg13g2_fill_4 FILLER_85_699 ();
 sg13g2_fill_2 FILLER_85_703 ();
 sg13g2_fill_1 FILLER_85_705 ();
 sg13g2_fill_8 FILLER_85_716 ();
 sg13g2_fill_4 FILLER_85_724 ();
 sg13g2_fill_1 FILLER_85_728 ();
 sg13g2_fill_8 FILLER_85_737 ();
 sg13g2_fill_8 FILLER_85_745 ();
 sg13g2_fill_8 FILLER_85_753 ();
 sg13g2_fill_8 FILLER_85_761 ();
 sg13g2_fill_4 FILLER_85_769 ();
 sg13g2_fill_2 FILLER_85_773 ();
 sg13g2_fill_8 FILLER_85_785 ();
 sg13g2_fill_8 FILLER_85_793 ();
 sg13g2_fill_8 FILLER_85_801 ();
 sg13g2_fill_2 FILLER_85_809 ();
 sg13g2_fill_4 FILLER_85_892 ();
 sg13g2_fill_2 FILLER_85_896 ();
 sg13g2_fill_4 FILLER_85_945 ();
 sg13g2_fill_1 FILLER_85_949 ();
 sg13g2_fill_1 FILLER_85_975 ();
 sg13g2_fill_2 FILLER_85_1015 ();
 sg13g2_fill_2 FILLER_85_1026 ();
 sg13g2_fill_1 FILLER_85_1050 ();
 sg13g2_fill_1 FILLER_85_1071 ();
 sg13g2_fill_2 FILLER_85_1080 ();
 sg13g2_fill_1 FILLER_85_1087 ();
 sg13g2_fill_4 FILLER_85_1126 ();
 sg13g2_fill_1 FILLER_85_1130 ();
 sg13g2_fill_8 FILLER_85_1136 ();
 sg13g2_fill_8 FILLER_85_1144 ();
 sg13g2_fill_1 FILLER_85_1157 ();
 sg13g2_fill_1 FILLER_85_1167 ();
 sg13g2_fill_2 FILLER_85_1179 ();
 sg13g2_fill_1 FILLER_85_1181 ();
 sg13g2_fill_2 FILLER_85_1188 ();
 sg13g2_fill_4 FILLER_85_1202 ();
 sg13g2_fill_1 FILLER_85_1226 ();
 sg13g2_fill_4 FILLER_85_1242 ();
 sg13g2_fill_1 FILLER_85_1246 ();
 sg13g2_fill_8 FILLER_85_1275 ();
 sg13g2_fill_1 FILLER_85_1283 ();
 sg13g2_fill_4 FILLER_85_1292 ();
 sg13g2_fill_2 FILLER_85_1296 ();
 sg13g2_fill_1 FILLER_85_1298 ();
 sg13g2_fill_8 FILLER_85_1305 ();
 sg13g2_fill_1 FILLER_85_1313 ();
 sg13g2_fill_1 FILLER_85_1326 ();
 sg13g2_fill_8 FILLER_85_1344 ();
 sg13g2_fill_8 FILLER_85_1352 ();
 sg13g2_fill_8 FILLER_85_1360 ();
 sg13g2_fill_2 FILLER_85_1368 ();
 sg13g2_fill_2 FILLER_85_1383 ();
 sg13g2_fill_8 FILLER_85_1390 ();
 sg13g2_fill_2 FILLER_85_1398 ();
 sg13g2_fill_2 FILLER_85_1405 ();
 sg13g2_fill_1 FILLER_85_1407 ();
 sg13g2_fill_8 FILLER_85_1412 ();
 sg13g2_fill_2 FILLER_85_1420 ();
 sg13g2_fill_1 FILLER_85_1422 ();
 sg13g2_fill_2 FILLER_85_1432 ();
 sg13g2_fill_4 FILLER_85_1459 ();
 sg13g2_fill_2 FILLER_85_1463 ();
 sg13g2_fill_1 FILLER_85_1465 ();
 sg13g2_fill_2 FILLER_85_1484 ();
 sg13g2_fill_1 FILLER_85_1497 ();
 sg13g2_fill_2 FILLER_85_1522 ();
 sg13g2_fill_4 FILLER_85_1569 ();
 sg13g2_fill_1 FILLER_85_1573 ();
 sg13g2_fill_8 FILLER_85_1582 ();
 sg13g2_fill_2 FILLER_85_1590 ();
 sg13g2_fill_8 FILLER_86_0 ();
 sg13g2_fill_8 FILLER_86_8 ();
 sg13g2_fill_8 FILLER_86_16 ();
 sg13g2_fill_8 FILLER_86_24 ();
 sg13g2_fill_8 FILLER_86_32 ();
 sg13g2_fill_2 FILLER_86_40 ();
 sg13g2_fill_1 FILLER_86_42 ();
 sg13g2_fill_8 FILLER_86_89 ();
 sg13g2_fill_8 FILLER_86_97 ();
 sg13g2_fill_2 FILLER_86_105 ();
 sg13g2_fill_1 FILLER_86_107 ();
 sg13g2_fill_8 FILLER_86_116 ();
 sg13g2_fill_1 FILLER_86_124 ();
 sg13g2_fill_8 FILLER_86_135 ();
 sg13g2_fill_8 FILLER_86_143 ();
 sg13g2_fill_1 FILLER_86_172 ();
 sg13g2_fill_4 FILLER_86_191 ();
 sg13g2_fill_2 FILLER_86_195 ();
 sg13g2_fill_4 FILLER_86_218 ();
 sg13g2_fill_2 FILLER_86_222 ();
 sg13g2_fill_8 FILLER_86_260 ();
 sg13g2_fill_1 FILLER_86_268 ();
 sg13g2_fill_2 FILLER_86_303 ();
 sg13g2_fill_1 FILLER_86_305 ();
 sg13g2_fill_8 FILLER_86_309 ();
 sg13g2_fill_8 FILLER_86_317 ();
 sg13g2_fill_4 FILLER_86_325 ();
 sg13g2_fill_2 FILLER_86_329 ();
 sg13g2_fill_1 FILLER_86_331 ();
 sg13g2_fill_8 FILLER_86_358 ();
 sg13g2_fill_4 FILLER_86_366 ();
 sg13g2_fill_2 FILLER_86_370 ();
 sg13g2_fill_1 FILLER_86_372 ();
 sg13g2_fill_8 FILLER_86_393 ();
 sg13g2_fill_4 FILLER_86_448 ();
 sg13g2_fill_8 FILLER_86_457 ();
 sg13g2_fill_4 FILLER_86_465 ();
 sg13g2_fill_8 FILLER_86_515 ();
 sg13g2_fill_4 FILLER_86_523 ();
 sg13g2_fill_2 FILLER_86_527 ();
 sg13g2_fill_1 FILLER_86_529 ();
 sg13g2_fill_8 FILLER_86_535 ();
 sg13g2_fill_8 FILLER_86_543 ();
 sg13g2_fill_2 FILLER_86_551 ();
 sg13g2_fill_1 FILLER_86_553 ();
 sg13g2_fill_4 FILLER_86_580 ();
 sg13g2_fill_2 FILLER_86_584 ();
 sg13g2_fill_4 FILLER_86_597 ();
 sg13g2_fill_2 FILLER_86_601 ();
 sg13g2_fill_1 FILLER_86_603 ();
 sg13g2_fill_8 FILLER_86_609 ();
 sg13g2_fill_4 FILLER_86_617 ();
 sg13g2_fill_2 FILLER_86_621 ();
 sg13g2_fill_1 FILLER_86_623 ();
 sg13g2_fill_8 FILLER_86_655 ();
 sg13g2_fill_8 FILLER_86_663 ();
 sg13g2_fill_8 FILLER_86_671 ();
 sg13g2_fill_2 FILLER_86_679 ();
 sg13g2_fill_1 FILLER_86_681 ();
 sg13g2_fill_4 FILLER_86_687 ();
 sg13g2_fill_1 FILLER_86_750 ();
 sg13g2_fill_8 FILLER_86_769 ();
 sg13g2_fill_4 FILLER_86_777 ();
 sg13g2_fill_2 FILLER_86_781 ();
 sg13g2_fill_2 FILLER_86_793 ();
 sg13g2_fill_4 FILLER_86_803 ();
 sg13g2_fill_1 FILLER_86_807 ();
 sg13g2_fill_4 FILLER_86_833 ();
 sg13g2_fill_1 FILLER_86_837 ();
 sg13g2_fill_4 FILLER_86_885 ();
 sg13g2_fill_8 FILLER_86_915 ();
 sg13g2_fill_4 FILLER_86_923 ();
 sg13g2_fill_2 FILLER_86_927 ();
 sg13g2_fill_4 FILLER_86_935 ();
 sg13g2_fill_2 FILLER_86_939 ();
 sg13g2_fill_2 FILLER_86_974 ();
 sg13g2_fill_2 FILLER_86_1006 ();
 sg13g2_fill_1 FILLER_86_1029 ();
 sg13g2_fill_2 FILLER_86_1058 ();
 sg13g2_fill_1 FILLER_86_1104 ();
 sg13g2_fill_4 FILLER_86_1121 ();
 sg13g2_fill_2 FILLER_86_1146 ();
 sg13g2_fill_1 FILLER_86_1148 ();
 sg13g2_fill_1 FILLER_86_1172 ();
 sg13g2_fill_8 FILLER_86_1201 ();
 sg13g2_fill_2 FILLER_86_1209 ();
 sg13g2_fill_4 FILLER_86_1216 ();
 sg13g2_fill_2 FILLER_86_1220 ();
 sg13g2_fill_1 FILLER_86_1222 ();
 sg13g2_fill_8 FILLER_86_1239 ();
 sg13g2_fill_2 FILLER_86_1253 ();
 sg13g2_fill_1 FILLER_86_1255 ();
 sg13g2_fill_8 FILLER_86_1261 ();
 sg13g2_fill_4 FILLER_86_1269 ();
 sg13g2_fill_2 FILLER_86_1273 ();
 sg13g2_fill_1 FILLER_86_1275 ();
 sg13g2_fill_2 FILLER_86_1280 ();
 sg13g2_fill_2 FILLER_86_1290 ();
 sg13g2_fill_8 FILLER_86_1317 ();
 sg13g2_fill_4 FILLER_86_1325 ();
 sg13g2_fill_2 FILLER_86_1329 ();
 sg13g2_fill_1 FILLER_86_1331 ();
 sg13g2_fill_8 FILLER_86_1338 ();
 sg13g2_fill_1 FILLER_86_1346 ();
 sg13g2_fill_8 FILLER_86_1374 ();
 sg13g2_fill_2 FILLER_86_1387 ();
 sg13g2_fill_4 FILLER_86_1394 ();
 sg13g2_fill_2 FILLER_86_1398 ();
 sg13g2_fill_4 FILLER_86_1430 ();
 sg13g2_fill_4 FILLER_86_1438 ();
 sg13g2_fill_2 FILLER_86_1442 ();
 sg13g2_fill_8 FILLER_86_1453 ();
 sg13g2_fill_8 FILLER_86_1461 ();
 sg13g2_fill_4 FILLER_86_1469 ();
 sg13g2_fill_2 FILLER_86_1473 ();
 sg13g2_fill_1 FILLER_86_1475 ();
 sg13g2_fill_1 FILLER_86_1492 ();
 sg13g2_fill_2 FILLER_86_1534 ();
 sg13g2_fill_1 FILLER_86_1536 ();
 sg13g2_fill_8 FILLER_87_0 ();
 sg13g2_fill_8 FILLER_87_8 ();
 sg13g2_fill_8 FILLER_87_16 ();
 sg13g2_fill_8 FILLER_87_24 ();
 sg13g2_fill_8 FILLER_87_32 ();
 sg13g2_fill_8 FILLER_87_40 ();
 sg13g2_fill_8 FILLER_87_48 ();
 sg13g2_fill_8 FILLER_87_56 ();
 sg13g2_fill_8 FILLER_87_64 ();
 sg13g2_fill_8 FILLER_87_72 ();
 sg13g2_fill_8 FILLER_87_80 ();
 sg13g2_fill_8 FILLER_87_88 ();
 sg13g2_fill_1 FILLER_87_96 ();
 sg13g2_fill_8 FILLER_87_115 ();
 sg13g2_fill_8 FILLER_87_123 ();
 sg13g2_fill_2 FILLER_87_131 ();
 sg13g2_fill_1 FILLER_87_133 ();
 sg13g2_fill_8 FILLER_87_160 ();
 sg13g2_fill_4 FILLER_87_168 ();
 sg13g2_fill_1 FILLER_87_172 ();
 sg13g2_fill_1 FILLER_87_181 ();
 sg13g2_fill_8 FILLER_87_229 ();
 sg13g2_fill_8 FILLER_87_237 ();
 sg13g2_fill_8 FILLER_87_245 ();
 sg13g2_fill_8 FILLER_87_253 ();
 sg13g2_fill_2 FILLER_87_261 ();
 sg13g2_fill_1 FILLER_87_263 ();
 sg13g2_fill_8 FILLER_87_274 ();
 sg13g2_fill_8 FILLER_87_282 ();
 sg13g2_fill_8 FILLER_87_290 ();
 sg13g2_fill_8 FILLER_87_298 ();
 sg13g2_fill_8 FILLER_87_311 ();
 sg13g2_fill_4 FILLER_87_319 ();
 sg13g2_fill_8 FILLER_87_395 ();
 sg13g2_fill_8 FILLER_87_403 ();
 sg13g2_fill_8 FILLER_87_411 ();
 sg13g2_fill_4 FILLER_87_419 ();
 sg13g2_fill_2 FILLER_87_423 ();
 sg13g2_fill_8 FILLER_87_435 ();
 sg13g2_fill_8 FILLER_87_443 ();
 sg13g2_fill_8 FILLER_87_451 ();
 sg13g2_fill_1 FILLER_87_459 ();
 sg13g2_fill_8 FILLER_87_473 ();
 sg13g2_fill_1 FILLER_87_481 ();
 sg13g2_fill_4 FILLER_87_488 ();
 sg13g2_fill_8 FILLER_87_517 ();
 sg13g2_fill_4 FILLER_87_525 ();
 sg13g2_fill_1 FILLER_87_529 ();
 sg13g2_fill_2 FILLER_87_538 ();
 sg13g2_fill_1 FILLER_87_540 ();
 sg13g2_fill_8 FILLER_87_561 ();
 sg13g2_fill_8 FILLER_87_569 ();
 sg13g2_fill_8 FILLER_87_577 ();
 sg13g2_fill_8 FILLER_87_585 ();
 sg13g2_fill_8 FILLER_87_593 ();
 sg13g2_fill_8 FILLER_87_601 ();
 sg13g2_fill_4 FILLER_87_609 ();
 sg13g2_fill_2 FILLER_87_613 ();
 sg13g2_fill_1 FILLER_87_615 ();
 sg13g2_fill_2 FILLER_87_620 ();
 sg13g2_fill_8 FILLER_87_678 ();
 sg13g2_fill_8 FILLER_87_686 ();
 sg13g2_fill_8 FILLER_87_708 ();
 sg13g2_fill_8 FILLER_87_716 ();
 sg13g2_fill_4 FILLER_87_782 ();
 sg13g2_fill_2 FILLER_87_786 ();
 sg13g2_fill_4 FILLER_87_835 ();
 sg13g2_fill_1 FILLER_87_839 ();
 sg13g2_fill_2 FILLER_87_881 ();
 sg13g2_fill_1 FILLER_87_886 ();
 sg13g2_fill_2 FILLER_87_890 ();
 sg13g2_fill_2 FILLER_87_1009 ();
 sg13g2_fill_2 FILLER_87_1022 ();
 sg13g2_fill_2 FILLER_87_1038 ();
 sg13g2_fill_2 FILLER_87_1054 ();
 sg13g2_fill_2 FILLER_87_1078 ();
 sg13g2_fill_8 FILLER_87_1122 ();
 sg13g2_fill_4 FILLER_87_1130 ();
 sg13g2_fill_2 FILLER_87_1154 ();
 sg13g2_fill_1 FILLER_87_1156 ();
 sg13g2_fill_8 FILLER_87_1166 ();
 sg13g2_fill_1 FILLER_87_1174 ();
 sg13g2_fill_8 FILLER_87_1190 ();
 sg13g2_fill_8 FILLER_87_1198 ();
 sg13g2_fill_2 FILLER_87_1206 ();
 sg13g2_fill_1 FILLER_87_1208 ();
 sg13g2_fill_4 FILLER_87_1214 ();
 sg13g2_fill_2 FILLER_87_1218 ();
 sg13g2_fill_1 FILLER_87_1226 ();
 sg13g2_fill_4 FILLER_87_1233 ();
 sg13g2_fill_2 FILLER_87_1249 ();
 sg13g2_fill_4 FILLER_87_1256 ();
 sg13g2_fill_2 FILLER_87_1265 ();
 sg13g2_fill_1 FILLER_87_1267 ();
 sg13g2_fill_8 FILLER_87_1272 ();
 sg13g2_fill_8 FILLER_87_1280 ();
 sg13g2_fill_4 FILLER_87_1288 ();
 sg13g2_fill_2 FILLER_87_1297 ();
 sg13g2_fill_1 FILLER_87_1299 ();
 sg13g2_fill_4 FILLER_87_1309 ();
 sg13g2_fill_2 FILLER_87_1313 ();
 sg13g2_fill_1 FILLER_87_1315 ();
 sg13g2_fill_1 FILLER_87_1328 ();
 sg13g2_fill_2 FILLER_87_1334 ();
 sg13g2_fill_1 FILLER_87_1336 ();
 sg13g2_fill_2 FILLER_87_1350 ();
 sg13g2_fill_1 FILLER_87_1352 ();
 sg13g2_fill_8 FILLER_87_1357 ();
 sg13g2_fill_4 FILLER_87_1365 ();
 sg13g2_fill_1 FILLER_87_1369 ();
 sg13g2_fill_2 FILLER_87_1398 ();
 sg13g2_fill_1 FILLER_87_1486 ();
 sg13g2_fill_8 FILLER_87_1493 ();
 sg13g2_fill_4 FILLER_87_1501 ();
 sg13g2_fill_1 FILLER_87_1505 ();
 sg13g2_fill_4 FILLER_87_1517 ();
 sg13g2_fill_2 FILLER_87_1521 ();
 sg13g2_fill_1 FILLER_87_1523 ();
 sg13g2_fill_4 FILLER_87_1532 ();
 sg13g2_fill_2 FILLER_87_1536 ();
 sg13g2_fill_8 FILLER_87_1543 ();
 sg13g2_fill_8 FILLER_87_1551 ();
 sg13g2_fill_2 FILLER_87_1559 ();
 sg13g2_fill_1 FILLER_87_1561 ();
 sg13g2_fill_8 FILLER_88_0 ();
 sg13g2_fill_8 FILLER_88_8 ();
 sg13g2_fill_8 FILLER_88_16 ();
 sg13g2_fill_8 FILLER_88_24 ();
 sg13g2_fill_8 FILLER_88_32 ();
 sg13g2_fill_8 FILLER_88_40 ();
 sg13g2_fill_8 FILLER_88_48 ();
 sg13g2_fill_4 FILLER_88_56 ();
 sg13g2_fill_2 FILLER_88_60 ();
 sg13g2_fill_2 FILLER_88_70 ();
 sg13g2_fill_1 FILLER_88_72 ();
 sg13g2_fill_8 FILLER_88_83 ();
 sg13g2_fill_4 FILLER_88_117 ();
 sg13g2_fill_1 FILLER_88_121 ();
 sg13g2_fill_8 FILLER_88_197 ();
 sg13g2_fill_8 FILLER_88_205 ();
 sg13g2_fill_8 FILLER_88_213 ();
 sg13g2_fill_2 FILLER_88_221 ();
 sg13g2_fill_4 FILLER_88_249 ();
 sg13g2_fill_4 FILLER_88_259 ();
 sg13g2_fill_8 FILLER_88_293 ();
 sg13g2_fill_4 FILLER_88_301 ();
 sg13g2_fill_1 FILLER_88_305 ();
 sg13g2_fill_8 FILLER_88_309 ();
 sg13g2_fill_8 FILLER_88_317 ();
 sg13g2_fill_8 FILLER_88_325 ();
 sg13g2_fill_8 FILLER_88_333 ();
 sg13g2_fill_8 FILLER_88_341 ();
 sg13g2_fill_8 FILLER_88_349 ();
 sg13g2_fill_4 FILLER_88_386 ();
 sg13g2_fill_8 FILLER_88_400 ();
 sg13g2_fill_8 FILLER_88_408 ();
 sg13g2_fill_8 FILLER_88_416 ();
 sg13g2_fill_8 FILLER_88_424 ();
 sg13g2_fill_8 FILLER_88_432 ();
 sg13g2_fill_2 FILLER_88_440 ();
 sg13g2_fill_1 FILLER_88_442 ();
 sg13g2_fill_8 FILLER_88_492 ();
 sg13g2_fill_8 FILLER_88_500 ();
 sg13g2_fill_4 FILLER_88_508 ();
 sg13g2_fill_1 FILLER_88_512 ();
 sg13g2_fill_4 FILLER_88_549 ();
 sg13g2_fill_2 FILLER_88_553 ();
 sg13g2_fill_1 FILLER_88_555 ();
 sg13g2_fill_4 FILLER_88_582 ();
 sg13g2_fill_2 FILLER_88_586 ();
 sg13g2_fill_8 FILLER_88_640 ();
 sg13g2_fill_8 FILLER_88_648 ();
 sg13g2_fill_2 FILLER_88_656 ();
 sg13g2_fill_8 FILLER_88_694 ();
 sg13g2_fill_2 FILLER_88_702 ();
 sg13g2_fill_1 FILLER_88_704 ();
 sg13g2_fill_8 FILLER_88_713 ();
 sg13g2_fill_8 FILLER_88_721 ();
 sg13g2_fill_8 FILLER_88_729 ();
 sg13g2_fill_8 FILLER_88_737 ();
 sg13g2_fill_8 FILLER_88_745 ();
 sg13g2_fill_8 FILLER_88_753 ();
 sg13g2_fill_8 FILLER_88_761 ();
 sg13g2_fill_4 FILLER_88_769 ();
 sg13g2_fill_2 FILLER_88_773 ();
 sg13g2_fill_1 FILLER_88_775 ();
 sg13g2_fill_8 FILLER_88_814 ();
 sg13g2_fill_8 FILLER_88_822 ();
 sg13g2_fill_8 FILLER_88_830 ();
 sg13g2_fill_8 FILLER_88_838 ();
 sg13g2_fill_8 FILLER_88_846 ();
 sg13g2_fill_8 FILLER_88_854 ();
 sg13g2_fill_8 FILLER_88_862 ();
 sg13g2_fill_4 FILLER_88_870 ();
 sg13g2_fill_2 FILLER_88_874 ();
 sg13g2_fill_1 FILLER_88_876 ();
 sg13g2_fill_1 FILLER_88_883 ();
 sg13g2_fill_1 FILLER_88_896 ();
 sg13g2_fill_1 FILLER_88_928 ();
 sg13g2_fill_8 FILLER_88_939 ();
 sg13g2_fill_1 FILLER_88_947 ();
 sg13g2_fill_1 FILLER_88_1027 ();
 sg13g2_fill_2 FILLER_88_1051 ();
 sg13g2_fill_1 FILLER_88_1071 ();
 sg13g2_fill_1 FILLER_88_1114 ();
 sg13g2_fill_1 FILLER_88_1129 ();
 sg13g2_fill_1 FILLER_88_1154 ();
 sg13g2_fill_8 FILLER_88_1168 ();
 sg13g2_fill_8 FILLER_88_1176 ();
 sg13g2_fill_2 FILLER_88_1184 ();
 sg13g2_fill_8 FILLER_88_1194 ();
 sg13g2_fill_2 FILLER_88_1202 ();
 sg13g2_fill_1 FILLER_88_1223 ();
 sg13g2_fill_8 FILLER_88_1232 ();
 sg13g2_fill_8 FILLER_88_1240 ();
 sg13g2_fill_8 FILLER_88_1248 ();
 sg13g2_fill_1 FILLER_88_1261 ();
 sg13g2_fill_8 FILLER_88_1272 ();
 sg13g2_fill_4 FILLER_88_1280 ();
 sg13g2_fill_2 FILLER_88_1284 ();
 sg13g2_fill_1 FILLER_88_1286 ();
 sg13g2_fill_4 FILLER_88_1299 ();
 sg13g2_fill_8 FILLER_88_1308 ();
 sg13g2_fill_8 FILLER_88_1316 ();
 sg13g2_fill_8 FILLER_88_1324 ();
 sg13g2_fill_4 FILLER_88_1332 ();
 sg13g2_fill_2 FILLER_88_1342 ();
 sg13g2_fill_8 FILLER_88_1365 ();
 sg13g2_fill_1 FILLER_88_1373 ();
 sg13g2_fill_2 FILLER_88_1378 ();
 sg13g2_fill_8 FILLER_88_1384 ();
 sg13g2_fill_2 FILLER_88_1392 ();
 sg13g2_fill_2 FILLER_88_1397 ();
 sg13g2_fill_1 FILLER_88_1399 ();
 sg13g2_fill_2 FILLER_88_1405 ();
 sg13g2_fill_1 FILLER_88_1407 ();
 sg13g2_fill_8 FILLER_88_1417 ();
 sg13g2_fill_4 FILLER_88_1430 ();
 sg13g2_fill_2 FILLER_88_1434 ();
 sg13g2_fill_1 FILLER_88_1436 ();
 sg13g2_fill_1 FILLER_88_1441 ();
 sg13g2_fill_4 FILLER_88_1463 ();
 sg13g2_fill_2 FILLER_88_1467 ();
 sg13g2_fill_2 FILLER_88_1474 ();
 sg13g2_fill_1 FILLER_88_1476 ();
 sg13g2_fill_4 FILLER_88_1485 ();
 sg13g2_fill_4 FILLER_88_1498 ();
 sg13g2_fill_1 FILLER_88_1502 ();
 sg13g2_fill_4 FILLER_88_1520 ();
 sg13g2_fill_2 FILLER_88_1524 ();
 sg13g2_fill_1 FILLER_88_1526 ();
 sg13g2_fill_8 FILLER_88_1538 ();
 sg13g2_fill_8 FILLER_88_1546 ();
 sg13g2_fill_8 FILLER_88_1554 ();
 sg13g2_fill_8 FILLER_89_0 ();
 sg13g2_fill_8 FILLER_89_8 ();
 sg13g2_fill_8 FILLER_89_16 ();
 sg13g2_fill_8 FILLER_89_24 ();
 sg13g2_fill_8 FILLER_89_32 ();
 sg13g2_fill_1 FILLER_89_40 ();
 sg13g2_fill_2 FILLER_89_103 ();
 sg13g2_fill_8 FILLER_89_125 ();
 sg13g2_fill_8 FILLER_89_133 ();
 sg13g2_fill_8 FILLER_89_141 ();
 sg13g2_fill_8 FILLER_89_149 ();
 sg13g2_fill_4 FILLER_89_157 ();
 sg13g2_fill_8 FILLER_89_193 ();
 sg13g2_fill_4 FILLER_89_201 ();
 sg13g2_fill_2 FILLER_89_205 ();
 sg13g2_fill_4 FILLER_89_215 ();
 sg13g2_fill_2 FILLER_89_219 ();
 sg13g2_fill_8 FILLER_89_231 ();
 sg13g2_fill_2 FILLER_89_239 ();
 sg13g2_fill_2 FILLER_89_267 ();
 sg13g2_fill_8 FILLER_89_275 ();
 sg13g2_fill_8 FILLER_89_283 ();
 sg13g2_fill_2 FILLER_89_291 ();
 sg13g2_fill_8 FILLER_89_319 ();
 sg13g2_fill_8 FILLER_89_327 ();
 sg13g2_fill_2 FILLER_89_335 ();
 sg13g2_fill_8 FILLER_89_347 ();
 sg13g2_fill_8 FILLER_89_355 ();
 sg13g2_fill_8 FILLER_89_363 ();
 sg13g2_fill_2 FILLER_89_371 ();
 sg13g2_fill_2 FILLER_89_383 ();
 sg13g2_fill_4 FILLER_89_390 ();
 sg13g2_fill_1 FILLER_89_394 ();
 sg13g2_fill_4 FILLER_89_421 ();
 sg13g2_fill_1 FILLER_89_433 ();
 sg13g2_fill_2 FILLER_89_460 ();
 sg13g2_fill_2 FILLER_89_481 ();
 sg13g2_fill_8 FILLER_89_527 ();
 sg13g2_fill_8 FILLER_89_535 ();
 sg13g2_fill_8 FILLER_89_543 ();
 sg13g2_fill_4 FILLER_89_551 ();
 sg13g2_fill_1 FILLER_89_555 ();
 sg13g2_fill_2 FILLER_89_607 ();
 sg13g2_fill_1 FILLER_89_609 ();
 sg13g2_fill_8 FILLER_89_640 ();
 sg13g2_fill_4 FILLER_89_648 ();
 sg13g2_fill_8 FILLER_89_657 ();
 sg13g2_fill_8 FILLER_89_665 ();
 sg13g2_fill_8 FILLER_89_673 ();
 sg13g2_fill_8 FILLER_89_681 ();
 sg13g2_fill_2 FILLER_89_689 ();
 sg13g2_fill_1 FILLER_89_701 ();
 sg13g2_fill_1 FILLER_89_723 ();
 sg13g2_fill_8 FILLER_89_742 ();
 sg13g2_fill_2 FILLER_89_750 ();
 sg13g2_fill_4 FILLER_89_762 ();
 sg13g2_fill_2 FILLER_89_766 ();
 sg13g2_fill_1 FILLER_89_768 ();
 sg13g2_fill_4 FILLER_89_815 ();
 sg13g2_fill_2 FILLER_89_819 ();
 sg13g2_fill_8 FILLER_89_850 ();
 sg13g2_fill_8 FILLER_89_858 ();
 sg13g2_fill_8 FILLER_89_866 ();
 sg13g2_fill_1 FILLER_89_886 ();
 sg13g2_fill_1 FILLER_89_900 ();
 sg13g2_fill_4 FILLER_89_931 ();
 sg13g2_fill_2 FILLER_89_944 ();
 sg13g2_fill_1 FILLER_89_971 ();
 sg13g2_fill_1 FILLER_89_1026 ();
 sg13g2_fill_1 FILLER_89_1050 ();
 sg13g2_fill_1 FILLER_89_1076 ();
 sg13g2_fill_4 FILLER_89_1105 ();
 sg13g2_fill_1 FILLER_89_1119 ();
 sg13g2_fill_8 FILLER_89_1125 ();
 sg13g2_fill_8 FILLER_89_1133 ();
 sg13g2_fill_8 FILLER_89_1141 ();
 sg13g2_fill_2 FILLER_89_1149 ();
 sg13g2_fill_1 FILLER_89_1160 ();
 sg13g2_fill_4 FILLER_89_1165 ();
 sg13g2_fill_2 FILLER_89_1169 ();
 sg13g2_fill_1 FILLER_89_1171 ();
 sg13g2_fill_1 FILLER_89_1177 ();
 sg13g2_fill_8 FILLER_89_1199 ();
 sg13g2_fill_8 FILLER_89_1207 ();
 sg13g2_fill_8 FILLER_89_1241 ();
 sg13g2_fill_4 FILLER_89_1249 ();
 sg13g2_fill_8 FILLER_89_1269 ();
 sg13g2_fill_4 FILLER_89_1319 ();
 sg13g2_fill_2 FILLER_89_1323 ();
 sg13g2_fill_2 FILLER_89_1347 ();
 sg13g2_fill_8 FILLER_89_1365 ();
 sg13g2_fill_8 FILLER_89_1373 ();
 sg13g2_fill_8 FILLER_89_1381 ();
 sg13g2_fill_2 FILLER_89_1389 ();
 sg13g2_fill_4 FILLER_89_1399 ();
 sg13g2_fill_4 FILLER_89_1408 ();
 sg13g2_fill_2 FILLER_89_1412 ();
 sg13g2_fill_8 FILLER_89_1418 ();
 sg13g2_fill_4 FILLER_89_1426 ();
 sg13g2_fill_1 FILLER_89_1430 ();
 sg13g2_fill_4 FILLER_89_1436 ();
 sg13g2_fill_8 FILLER_89_1444 ();
 sg13g2_fill_8 FILLER_89_1452 ();
 sg13g2_fill_4 FILLER_89_1460 ();
 sg13g2_fill_2 FILLER_89_1464 ();
 sg13g2_fill_2 FILLER_89_1472 ();
 sg13g2_fill_1 FILLER_89_1474 ();
 sg13g2_fill_4 FILLER_89_1481 ();
 sg13g2_fill_1 FILLER_89_1490 ();
 sg13g2_fill_1 FILLER_89_1519 ();
 sg13g2_fill_4 FILLER_89_1585 ();
 sg13g2_fill_2 FILLER_89_1589 ();
 sg13g2_fill_1 FILLER_89_1591 ();
 sg13g2_fill_8 FILLER_90_0 ();
 sg13g2_fill_8 FILLER_90_8 ();
 sg13g2_fill_8 FILLER_90_16 ();
 sg13g2_fill_8 FILLER_90_24 ();
 sg13g2_fill_8 FILLER_90_32 ();
 sg13g2_fill_8 FILLER_90_40 ();
 sg13g2_fill_8 FILLER_90_48 ();
 sg13g2_fill_8 FILLER_90_56 ();
 sg13g2_fill_2 FILLER_90_64 ();
 sg13g2_fill_4 FILLER_90_106 ();
 sg13g2_fill_1 FILLER_90_110 ();
 sg13g2_fill_1 FILLER_90_121 ();
 sg13g2_fill_2 FILLER_90_128 ();
 sg13g2_fill_4 FILLER_90_134 ();
 sg13g2_fill_2 FILLER_90_138 ();
 sg13g2_fill_4 FILLER_90_150 ();
 sg13g2_fill_2 FILLER_90_154 ();
 sg13g2_fill_1 FILLER_90_156 ();
 sg13g2_fill_2 FILLER_90_185 ();
 sg13g2_fill_4 FILLER_90_205 ();
 sg13g2_fill_4 FILLER_90_217 ();
 sg13g2_fill_8 FILLER_90_229 ();
 sg13g2_fill_1 FILLER_90_262 ();
 sg13g2_fill_2 FILLER_90_279 ();
 sg13g2_fill_1 FILLER_90_336 ();
 sg13g2_fill_8 FILLER_90_363 ();
 sg13g2_fill_1 FILLER_90_381 ();
 sg13g2_fill_8 FILLER_90_388 ();
 sg13g2_fill_2 FILLER_90_432 ();
 sg13g2_fill_1 FILLER_90_434 ();
 sg13g2_fill_8 FILLER_90_440 ();
 sg13g2_fill_4 FILLER_90_448 ();
 sg13g2_fill_2 FILLER_90_475 ();
 sg13g2_fill_8 FILLER_90_483 ();
 sg13g2_fill_2 FILLER_90_539 ();
 sg13g2_fill_1 FILLER_90_541 ();
 sg13g2_fill_8 FILLER_90_558 ();
 sg13g2_fill_4 FILLER_90_566 ();
 sg13g2_fill_1 FILLER_90_599 ();
 sg13g2_fill_8 FILLER_90_610 ();
 sg13g2_fill_8 FILLER_90_618 ();
 sg13g2_fill_4 FILLER_90_626 ();
 sg13g2_fill_8 FILLER_90_646 ();
 sg13g2_fill_2 FILLER_90_690 ();
 sg13g2_fill_1 FILLER_90_726 ();
 sg13g2_fill_2 FILLER_90_757 ();
 sg13g2_fill_4 FILLER_90_769 ();
 sg13g2_fill_2 FILLER_90_773 ();
 sg13g2_fill_1 FILLER_90_775 ();
 sg13g2_fill_8 FILLER_90_786 ();
 sg13g2_fill_4 FILLER_90_794 ();
 sg13g2_fill_1 FILLER_90_798 ();
 sg13g2_fill_2 FILLER_90_829 ();
 sg13g2_fill_8 FILLER_90_840 ();
 sg13g2_fill_4 FILLER_90_848 ();
 sg13g2_fill_1 FILLER_90_852 ();
 sg13g2_fill_1 FILLER_90_886 ();
 sg13g2_fill_1 FILLER_90_898 ();
 sg13g2_fill_2 FILLER_90_910 ();
 sg13g2_fill_2 FILLER_90_922 ();
 sg13g2_fill_2 FILLER_90_954 ();
 sg13g2_fill_1 FILLER_90_977 ();
 sg13g2_fill_2 FILLER_90_1004 ();
 sg13g2_fill_1 FILLER_90_1020 ();
 sg13g2_fill_2 FILLER_90_1035 ();
 sg13g2_fill_2 FILLER_90_1063 ();
 sg13g2_fill_1 FILLER_90_1110 ();
 sg13g2_fill_4 FILLER_90_1116 ();
 sg13g2_fill_2 FILLER_90_1120 ();
 sg13g2_fill_1 FILLER_90_1122 ();
 sg13g2_fill_4 FILLER_90_1127 ();
 sg13g2_fill_4 FILLER_90_1140 ();
 sg13g2_fill_2 FILLER_90_1150 ();
 sg13g2_fill_8 FILLER_90_1201 ();
 sg13g2_fill_8 FILLER_90_1209 ();
 sg13g2_fill_4 FILLER_90_1217 ();
 sg13g2_fill_2 FILLER_90_1221 ();
 sg13g2_fill_4 FILLER_90_1236 ();
 sg13g2_fill_2 FILLER_90_1240 ();
 sg13g2_fill_8 FILLER_90_1247 ();
 sg13g2_fill_8 FILLER_90_1255 ();
 sg13g2_fill_1 FILLER_90_1263 ();
 sg13g2_fill_1 FILLER_90_1273 ();
 sg13g2_fill_2 FILLER_90_1289 ();
 sg13g2_fill_2 FILLER_90_1298 ();
 sg13g2_fill_2 FILLER_90_1308 ();
 sg13g2_fill_1 FILLER_90_1310 ();
 sg13g2_fill_2 FILLER_90_1321 ();
 sg13g2_fill_2 FILLER_90_1334 ();
 sg13g2_fill_1 FILLER_90_1350 ();
 sg13g2_fill_2 FILLER_90_1369 ();
 sg13g2_fill_1 FILLER_90_1380 ();
 sg13g2_fill_2 FILLER_90_1386 ();
 sg13g2_fill_2 FILLER_90_1403 ();
 sg13g2_fill_4 FILLER_90_1431 ();
 sg13g2_fill_4 FILLER_90_1461 ();
 sg13g2_fill_2 FILLER_90_1465 ();
 sg13g2_fill_1 FILLER_90_1508 ();
 sg13g2_fill_8 FILLER_90_1517 ();
 sg13g2_fill_8 FILLER_90_1525 ();
 sg13g2_fill_1 FILLER_90_1533 ();
 sg13g2_fill_8 FILLER_90_1559 ();
 sg13g2_fill_8 FILLER_90_1567 ();
 sg13g2_fill_8 FILLER_90_1575 ();
 sg13g2_fill_8 FILLER_90_1583 ();
 sg13g2_fill_1 FILLER_90_1591 ();
 sg13g2_fill_8 FILLER_91_0 ();
 sg13g2_fill_8 FILLER_91_8 ();
 sg13g2_fill_8 FILLER_91_16 ();
 sg13g2_fill_8 FILLER_91_24 ();
 sg13g2_fill_8 FILLER_91_32 ();
 sg13g2_fill_1 FILLER_91_40 ();
 sg13g2_fill_4 FILLER_91_67 ();
 sg13g2_fill_2 FILLER_91_71 ();
 sg13g2_fill_4 FILLER_91_83 ();
 sg13g2_fill_2 FILLER_91_87 ();
 sg13g2_fill_1 FILLER_91_89 ();
 sg13g2_fill_8 FILLER_91_132 ();
 sg13g2_fill_1 FILLER_91_140 ();
 sg13g2_fill_4 FILLER_91_167 ();
 sg13g2_fill_2 FILLER_91_171 ();
 sg13g2_fill_2 FILLER_91_187 ();
 sg13g2_fill_4 FILLER_91_215 ();
 sg13g2_fill_1 FILLER_91_219 ();
 sg13g2_fill_2 FILLER_91_274 ();
 sg13g2_fill_1 FILLER_91_276 ();
 sg13g2_fill_8 FILLER_91_287 ();
 sg13g2_fill_8 FILLER_91_295 ();
 sg13g2_fill_2 FILLER_91_303 ();
 sg13g2_fill_2 FILLER_91_315 ();
 sg13g2_fill_4 FILLER_91_342 ();
 sg13g2_fill_2 FILLER_91_372 ();
 sg13g2_fill_1 FILLER_91_374 ();
 sg13g2_fill_8 FILLER_91_398 ();
 sg13g2_fill_8 FILLER_91_406 ();
 sg13g2_fill_8 FILLER_91_414 ();
 sg13g2_fill_8 FILLER_91_422 ();
 sg13g2_fill_4 FILLER_91_430 ();
 sg13g2_fill_1 FILLER_91_434 ();
 sg13g2_fill_8 FILLER_91_484 ();
 sg13g2_fill_2 FILLER_91_492 ();
 sg13g2_fill_1 FILLER_91_494 ();
 sg13g2_fill_2 FILLER_91_508 ();
 sg13g2_fill_2 FILLER_91_546 ();
 sg13g2_fill_1 FILLER_91_574 ();
 sg13g2_fill_4 FILLER_91_585 ();
 sg13g2_fill_1 FILLER_91_589 ();
 sg13g2_fill_1 FILLER_91_600 ();
 sg13g2_fill_2 FILLER_91_619 ();
 sg13g2_fill_2 FILLER_91_629 ();
 sg13g2_fill_4 FILLER_91_647 ();
 sg13g2_fill_4 FILLER_91_687 ();
 sg13g2_fill_1 FILLER_91_691 ();
 sg13g2_fill_1 FILLER_91_696 ();
 sg13g2_fill_8 FILLER_91_723 ();
 sg13g2_fill_4 FILLER_91_731 ();
 sg13g2_fill_8 FILLER_91_740 ();
 sg13g2_fill_1 FILLER_91_748 ();
 sg13g2_fill_8 FILLER_91_814 ();
 sg13g2_fill_2 FILLER_91_822 ();
 sg13g2_fill_1 FILLER_91_824 ();
 sg13g2_fill_2 FILLER_91_867 ();
 sg13g2_fill_2 FILLER_91_903 ();
 sg13g2_fill_1 FILLER_91_905 ();
 sg13g2_fill_4 FILLER_91_913 ();
 sg13g2_fill_1 FILLER_91_917 ();
 sg13g2_fill_8 FILLER_91_937 ();
 sg13g2_fill_8 FILLER_91_945 ();
 sg13g2_fill_1 FILLER_91_953 ();
 sg13g2_fill_2 FILLER_91_964 ();
 sg13g2_fill_1 FILLER_91_976 ();
 sg13g2_fill_2 FILLER_91_1006 ();
 sg13g2_fill_1 FILLER_91_1028 ();
 sg13g2_fill_2 FILLER_91_1034 ();
 sg13g2_fill_2 FILLER_91_1044 ();
 sg13g2_fill_2 FILLER_91_1055 ();
 sg13g2_fill_4 FILLER_91_1090 ();
 sg13g2_fill_1 FILLER_91_1094 ();
 sg13g2_fill_2 FILLER_91_1115 ();
 sg13g2_fill_1 FILLER_91_1117 ();
 sg13g2_fill_8 FILLER_91_1139 ();
 sg13g2_fill_8 FILLER_91_1147 ();
 sg13g2_fill_4 FILLER_91_1155 ();
 sg13g2_fill_8 FILLER_91_1163 ();
 sg13g2_fill_8 FILLER_91_1171 ();
 sg13g2_fill_2 FILLER_91_1179 ();
 sg13g2_fill_8 FILLER_91_1197 ();
 sg13g2_fill_8 FILLER_91_1205 ();
 sg13g2_fill_8 FILLER_91_1213 ();
 sg13g2_fill_8 FILLER_91_1221 ();
 sg13g2_fill_4 FILLER_91_1229 ();
 sg13g2_fill_2 FILLER_91_1271 ();
 sg13g2_fill_1 FILLER_91_1286 ();
 sg13g2_fill_2 FILLER_91_1302 ();
 sg13g2_fill_8 FILLER_91_1319 ();
 sg13g2_fill_4 FILLER_91_1327 ();
 sg13g2_fill_1 FILLER_91_1331 ();
 sg13g2_fill_2 FILLER_91_1337 ();
 sg13g2_fill_1 FILLER_91_1345 ();
 sg13g2_fill_1 FILLER_91_1351 ();
 sg13g2_fill_8 FILLER_91_1361 ();
 sg13g2_fill_4 FILLER_91_1369 ();
 sg13g2_fill_2 FILLER_91_1373 ();
 sg13g2_fill_1 FILLER_91_1375 ();
 sg13g2_fill_4 FILLER_91_1414 ();
 sg13g2_fill_8 FILLER_91_1451 ();
 sg13g2_fill_2 FILLER_91_1459 ();
 sg13g2_fill_1 FILLER_91_1461 ();
 sg13g2_fill_1 FILLER_91_1517 ();
 sg13g2_fill_8 FILLER_91_1522 ();
 sg13g2_fill_8 FILLER_91_1530 ();
 sg13g2_fill_8 FILLER_91_1538 ();
 sg13g2_fill_8 FILLER_91_1546 ();
 sg13g2_fill_8 FILLER_91_1554 ();
 sg13g2_fill_8 FILLER_91_1562 ();
 sg13g2_fill_1 FILLER_91_1570 ();
 sg13g2_fill_8 FILLER_91_1579 ();
 sg13g2_fill_4 FILLER_91_1587 ();
 sg13g2_fill_1 FILLER_91_1591 ();
 sg13g2_fill_8 FILLER_92_0 ();
 sg13g2_fill_8 FILLER_92_8 ();
 sg13g2_fill_8 FILLER_92_16 ();
 sg13g2_fill_8 FILLER_92_24 ();
 sg13g2_fill_1 FILLER_92_32 ();
 sg13g2_fill_4 FILLER_92_69 ();
 sg13g2_fill_2 FILLER_92_73 ();
 sg13g2_fill_8 FILLER_92_91 ();
 sg13g2_fill_8 FILLER_92_99 ();
 sg13g2_fill_8 FILLER_92_107 ();
 sg13g2_fill_8 FILLER_92_115 ();
 sg13g2_fill_4 FILLER_92_123 ();
 sg13g2_fill_2 FILLER_92_127 ();
 sg13g2_fill_8 FILLER_92_142 ();
 sg13g2_fill_8 FILLER_92_150 ();
 sg13g2_fill_8 FILLER_92_158 ();
 sg13g2_fill_8 FILLER_92_166 ();
 sg13g2_fill_8 FILLER_92_174 ();
 sg13g2_fill_8 FILLER_92_191 ();
 sg13g2_fill_8 FILLER_92_199 ();
 sg13g2_fill_4 FILLER_92_207 ();
 sg13g2_fill_2 FILLER_92_211 ();
 sg13g2_fill_8 FILLER_92_229 ();
 sg13g2_fill_8 FILLER_92_250 ();
 sg13g2_fill_4 FILLER_92_263 ();
 sg13g2_fill_8 FILLER_92_282 ();
 sg13g2_fill_8 FILLER_92_290 ();
 sg13g2_fill_4 FILLER_92_298 ();
 sg13g2_fill_2 FILLER_92_302 ();
 sg13g2_fill_1 FILLER_92_304 ();
 sg13g2_fill_2 FILLER_92_326 ();
 sg13g2_fill_1 FILLER_92_328 ();
 sg13g2_fill_8 FILLER_92_349 ();
 sg13g2_fill_8 FILLER_92_357 ();
 sg13g2_fill_8 FILLER_92_365 ();
 sg13g2_fill_8 FILLER_92_373 ();
 sg13g2_fill_4 FILLER_92_381 ();
 sg13g2_fill_2 FILLER_92_385 ();
 sg13g2_fill_1 FILLER_92_387 ();
 sg13g2_fill_2 FILLER_92_395 ();
 sg13g2_fill_4 FILLER_92_417 ();
 sg13g2_fill_2 FILLER_92_421 ();
 sg13g2_fill_1 FILLER_92_423 ();
 sg13g2_fill_4 FILLER_92_460 ();
 sg13g2_fill_2 FILLER_92_464 ();
 sg13g2_fill_1 FILLER_92_466 ();
 sg13g2_fill_2 FILLER_92_475 ();
 sg13g2_fill_8 FILLER_92_503 ();
 sg13g2_fill_2 FILLER_92_511 ();
 sg13g2_fill_8 FILLER_92_523 ();
 sg13g2_fill_8 FILLER_92_531 ();
 sg13g2_fill_2 FILLER_92_539 ();
 sg13g2_fill_1 FILLER_92_541 ();
 sg13g2_fill_8 FILLER_92_552 ();
 sg13g2_fill_4 FILLER_92_560 ();
 sg13g2_fill_2 FILLER_92_564 ();
 sg13g2_fill_1 FILLER_92_566 ();
 sg13g2_fill_8 FILLER_92_593 ();
 sg13g2_fill_8 FILLER_92_601 ();
 sg13g2_fill_1 FILLER_92_614 ();
 sg13g2_fill_8 FILLER_92_619 ();
 sg13g2_fill_8 FILLER_92_627 ();
 sg13g2_fill_2 FILLER_92_635 ();
 sg13g2_fill_4 FILLER_92_648 ();
 sg13g2_fill_2 FILLER_92_652 ();
 sg13g2_fill_1 FILLER_92_654 ();
 sg13g2_fill_8 FILLER_92_680 ();
 sg13g2_fill_8 FILLER_92_688 ();
 sg13g2_fill_8 FILLER_92_696 ();
 sg13g2_fill_2 FILLER_92_704 ();
 sg13g2_fill_4 FILLER_92_711 ();
 sg13g2_fill_2 FILLER_92_715 ();
 sg13g2_fill_1 FILLER_92_717 ();
 sg13g2_fill_8 FILLER_92_736 ();
 sg13g2_fill_4 FILLER_92_744 ();
 sg13g2_fill_1 FILLER_92_748 ();
 sg13g2_fill_8 FILLER_92_754 ();
 sg13g2_fill_8 FILLER_92_762 ();
 sg13g2_fill_8 FILLER_92_770 ();
 sg13g2_fill_8 FILLER_92_778 ();
 sg13g2_fill_1 FILLER_92_786 ();
 sg13g2_fill_2 FILLER_92_813 ();
 sg13g2_fill_1 FILLER_92_815 ();
 sg13g2_fill_8 FILLER_92_828 ();
 sg13g2_fill_2 FILLER_92_876 ();
 sg13g2_fill_1 FILLER_92_883 ();
 sg13g2_fill_1 FILLER_92_897 ();
 sg13g2_fill_4 FILLER_92_933 ();
 sg13g2_fill_2 FILLER_92_937 ();
 sg13g2_fill_8 FILLER_92_944 ();
 sg13g2_fill_1 FILLER_92_952 ();
 sg13g2_fill_1 FILLER_92_1023 ();
 sg13g2_fill_2 FILLER_92_1035 ();
 sg13g2_fill_1 FILLER_92_1062 ();
 sg13g2_fill_1 FILLER_92_1079 ();
 sg13g2_fill_4 FILLER_92_1085 ();
 sg13g2_fill_8 FILLER_92_1097 ();
 sg13g2_fill_8 FILLER_92_1105 ();
 sg13g2_fill_8 FILLER_92_1113 ();
 sg13g2_fill_4 FILLER_92_1121 ();
 sg13g2_fill_4 FILLER_92_1142 ();
 sg13g2_fill_1 FILLER_92_1146 ();
 sg13g2_fill_2 FILLER_92_1151 ();
 sg13g2_fill_8 FILLER_92_1179 ();
 sg13g2_fill_4 FILLER_92_1187 ();
 sg13g2_fill_2 FILLER_92_1191 ();
 sg13g2_fill_1 FILLER_92_1193 ();
 sg13g2_fill_4 FILLER_92_1200 ();
 sg13g2_fill_1 FILLER_92_1213 ();
 sg13g2_fill_8 FILLER_92_1227 ();
 sg13g2_fill_4 FILLER_92_1235 ();
 sg13g2_fill_1 FILLER_92_1239 ();
 sg13g2_fill_4 FILLER_92_1266 ();
 sg13g2_fill_2 FILLER_92_1270 ();
 sg13g2_fill_1 FILLER_92_1272 ();
 sg13g2_fill_2 FILLER_92_1277 ();
 sg13g2_fill_1 FILLER_92_1287 ();
 sg13g2_fill_4 FILLER_92_1292 ();
 sg13g2_fill_2 FILLER_92_1296 ();
 sg13g2_fill_1 FILLER_92_1303 ();
 sg13g2_fill_8 FILLER_92_1309 ();
 sg13g2_fill_2 FILLER_92_1320 ();
 sg13g2_fill_2 FILLER_92_1327 ();
 sg13g2_fill_1 FILLER_92_1329 ();
 sg13g2_fill_8 FILLER_92_1335 ();
 sg13g2_fill_8 FILLER_92_1346 ();
 sg13g2_fill_4 FILLER_92_1354 ();
 sg13g2_fill_2 FILLER_92_1358 ();
 sg13g2_fill_1 FILLER_92_1360 ();
 sg13g2_fill_2 FILLER_92_1365 ();
 sg13g2_fill_8 FILLER_92_1375 ();
 sg13g2_fill_4 FILLER_92_1383 ();
 sg13g2_fill_2 FILLER_92_1387 ();
 sg13g2_fill_1 FILLER_92_1394 ();
 sg13g2_fill_2 FILLER_92_1409 ();
 sg13g2_fill_1 FILLER_92_1411 ();
 sg13g2_fill_2 FILLER_92_1425 ();
 sg13g2_fill_1 FILLER_92_1484 ();
 sg13g2_fill_4 FILLER_92_1490 ();
 sg13g2_fill_8 FILLER_92_1504 ();
 sg13g2_fill_8 FILLER_92_1532 ();
 sg13g2_fill_1 FILLER_92_1540 ();
 sg13g2_fill_4 FILLER_92_1546 ();
 sg13g2_fill_1 FILLER_92_1550 ();
 sg13g2_fill_4 FILLER_92_1556 ();
 sg13g2_fill_2 FILLER_92_1589 ();
 sg13g2_fill_1 FILLER_92_1591 ();
 sg13g2_fill_8 FILLER_93_0 ();
 sg13g2_fill_8 FILLER_93_8 ();
 sg13g2_fill_8 FILLER_93_16 ();
 sg13g2_fill_8 FILLER_93_24 ();
 sg13g2_fill_2 FILLER_93_32 ();
 sg13g2_fill_1 FILLER_93_34 ();
 sg13g2_fill_8 FILLER_93_45 ();
 sg13g2_fill_8 FILLER_93_53 ();
 sg13g2_fill_8 FILLER_93_61 ();
 sg13g2_fill_2 FILLER_93_69 ();
 sg13g2_fill_1 FILLER_93_81 ();
 sg13g2_fill_2 FILLER_93_88 ();
 sg13g2_fill_8 FILLER_93_98 ();
 sg13g2_fill_8 FILLER_93_106 ();
 sg13g2_fill_2 FILLER_93_114 ();
 sg13g2_fill_1 FILLER_93_116 ();
 sg13g2_fill_4 FILLER_93_140 ();
 sg13g2_fill_8 FILLER_93_190 ();
 sg13g2_fill_8 FILLER_93_198 ();
 sg13g2_fill_8 FILLER_93_206 ();
 sg13g2_fill_1 FILLER_93_214 ();
 sg13g2_fill_4 FILLER_93_223 ();
 sg13g2_fill_2 FILLER_93_227 ();
 sg13g2_fill_1 FILLER_93_229 ();
 sg13g2_fill_8 FILLER_93_238 ();
 sg13g2_fill_1 FILLER_93_246 ();
 sg13g2_fill_8 FILLER_93_369 ();
 sg13g2_fill_2 FILLER_93_377 ();
 sg13g2_fill_4 FILLER_93_395 ();
 sg13g2_fill_2 FILLER_93_399 ();
 sg13g2_fill_1 FILLER_93_401 ();
 sg13g2_fill_4 FILLER_93_428 ();
 sg13g2_fill_2 FILLER_93_432 ();
 sg13g2_fill_1 FILLER_93_434 ();
 sg13g2_fill_4 FILLER_93_441 ();
 sg13g2_fill_4 FILLER_93_479 ();
 sg13g2_fill_8 FILLER_93_488 ();
 sg13g2_fill_2 FILLER_93_496 ();
 sg13g2_fill_1 FILLER_93_498 ();
 sg13g2_fill_1 FILLER_93_507 ();
 sg13g2_fill_8 FILLER_93_551 ();
 sg13g2_fill_1 FILLER_93_559 ();
 sg13g2_fill_4 FILLER_93_596 ();
 sg13g2_fill_1 FILLER_93_600 ();
 sg13g2_fill_8 FILLER_93_608 ();
 sg13g2_fill_8 FILLER_93_616 ();
 sg13g2_fill_4 FILLER_93_624 ();
 sg13g2_fill_1 FILLER_93_628 ();
 sg13g2_fill_4 FILLER_93_640 ();
 sg13g2_fill_1 FILLER_93_654 ();
 sg13g2_fill_2 FILLER_93_676 ();
 sg13g2_fill_1 FILLER_93_678 ();
 sg13g2_fill_4 FILLER_93_687 ();
 sg13g2_fill_2 FILLER_93_691 ();
 sg13g2_fill_1 FILLER_93_693 ();
 sg13g2_fill_4 FILLER_93_724 ();
 sg13g2_fill_8 FILLER_93_780 ();
 sg13g2_fill_8 FILLER_93_788 ();
 sg13g2_fill_2 FILLER_93_796 ();
 sg13g2_fill_1 FILLER_93_798 ();
 sg13g2_fill_2 FILLER_93_830 ();
 sg13g2_fill_1 FILLER_93_832 ();
 sg13g2_fill_2 FILLER_93_859 ();
 sg13g2_fill_1 FILLER_93_888 ();
 sg13g2_fill_4 FILLER_93_902 ();
 sg13g2_fill_2 FILLER_93_906 ();
 sg13g2_fill_1 FILLER_93_908 ();
 sg13g2_fill_2 FILLER_93_919 ();
 sg13g2_fill_1 FILLER_93_921 ();
 sg13g2_fill_8 FILLER_93_927 ();
 sg13g2_fill_8 FILLER_93_935 ();
 sg13g2_fill_4 FILLER_93_943 ();
 sg13g2_fill_1 FILLER_93_947 ();
 sg13g2_fill_8 FILLER_93_952 ();
 sg13g2_fill_4 FILLER_93_960 ();
 sg13g2_fill_2 FILLER_93_964 ();
 sg13g2_fill_8 FILLER_93_1005 ();
 sg13g2_fill_8 FILLER_93_1013 ();
 sg13g2_fill_1 FILLER_93_1021 ();
 sg13g2_fill_2 FILLER_93_1034 ();
 sg13g2_fill_1 FILLER_93_1049 ();
 sg13g2_fill_1 FILLER_93_1078 ();
 sg13g2_fill_4 FILLER_93_1087 ();
 sg13g2_fill_8 FILLER_93_1107 ();
 sg13g2_fill_4 FILLER_93_1115 ();
 sg13g2_fill_1 FILLER_93_1127 ();
 sg13g2_fill_8 FILLER_93_1146 ();
 sg13g2_fill_8 FILLER_93_1173 ();
 sg13g2_fill_8 FILLER_93_1181 ();
 sg13g2_fill_2 FILLER_93_1189 ();
 sg13g2_fill_1 FILLER_93_1191 ();
 sg13g2_fill_2 FILLER_93_1210 ();
 sg13g2_fill_2 FILLER_93_1260 ();
 sg13g2_fill_1 FILLER_93_1262 ();
 sg13g2_fill_8 FILLER_93_1273 ();
 sg13g2_fill_8 FILLER_93_1281 ();
 sg13g2_fill_8 FILLER_93_1289 ();
 sg13g2_fill_8 FILLER_93_1297 ();
 sg13g2_fill_1 FILLER_93_1311 ();
 sg13g2_fill_1 FILLER_93_1325 ();
 sg13g2_fill_8 FILLER_93_1345 ();
 sg13g2_fill_2 FILLER_93_1353 ();
 sg13g2_fill_1 FILLER_93_1355 ();
 sg13g2_fill_8 FILLER_93_1383 ();
 sg13g2_fill_2 FILLER_93_1391 ();
 sg13g2_fill_1 FILLER_93_1393 ();
 sg13g2_fill_2 FILLER_93_1406 ();
 sg13g2_fill_1 FILLER_93_1408 ();
 sg13g2_fill_1 FILLER_93_1414 ();
 sg13g2_fill_8 FILLER_93_1446 ();
 sg13g2_fill_8 FILLER_93_1454 ();
 sg13g2_fill_8 FILLER_93_1462 ();
 sg13g2_fill_2 FILLER_93_1482 ();
 sg13g2_fill_1 FILLER_93_1489 ();
 sg13g2_fill_8 FILLER_93_1495 ();
 sg13g2_fill_2 FILLER_93_1503 ();
 sg13g2_fill_2 FILLER_93_1516 ();
 sg13g2_fill_1 FILLER_93_1518 ();
 sg13g2_fill_8 FILLER_93_1525 ();
 sg13g2_fill_2 FILLER_93_1533 ();
 sg13g2_fill_1 FILLER_93_1535 ();
 sg13g2_fill_4 FILLER_93_1558 ();
 sg13g2_fill_2 FILLER_93_1562 ();
 sg13g2_fill_2 FILLER_93_1590 ();
 sg13g2_fill_8 FILLER_94_0 ();
 sg13g2_fill_8 FILLER_94_8 ();
 sg13g2_fill_8 FILLER_94_16 ();
 sg13g2_fill_4 FILLER_94_24 ();
 sg13g2_fill_2 FILLER_94_28 ();
 sg13g2_fill_1 FILLER_94_30 ();
 sg13g2_fill_4 FILLER_94_67 ();
 sg13g2_fill_1 FILLER_94_71 ();
 sg13g2_fill_8 FILLER_94_82 ();
 sg13g2_fill_2 FILLER_94_90 ();
 sg13g2_fill_1 FILLER_94_92 ();
 sg13g2_fill_4 FILLER_94_119 ();
 sg13g2_fill_4 FILLER_94_133 ();
 sg13g2_fill_2 FILLER_94_137 ();
 sg13g2_fill_1 FILLER_94_139 ();
 sg13g2_fill_4 FILLER_94_174 ();
 sg13g2_fill_2 FILLER_94_178 ();
 sg13g2_fill_8 FILLER_94_206 ();
 sg13g2_fill_4 FILLER_94_214 ();
 sg13g2_fill_2 FILLER_94_218 ();
 sg13g2_fill_1 FILLER_94_220 ();
 sg13g2_fill_4 FILLER_94_257 ();
 sg13g2_fill_2 FILLER_94_261 ();
 sg13g2_fill_8 FILLER_94_288 ();
 sg13g2_fill_8 FILLER_94_296 ();
 sg13g2_fill_2 FILLER_94_304 ();
 sg13g2_fill_1 FILLER_94_306 ();
 sg13g2_fill_8 FILLER_94_310 ();
 sg13g2_fill_8 FILLER_94_318 ();
 sg13g2_fill_1 FILLER_94_326 ();
 sg13g2_fill_8 FILLER_94_335 ();
 sg13g2_fill_4 FILLER_94_343 ();
 sg13g2_fill_2 FILLER_94_347 ();
 sg13g2_fill_1 FILLER_94_349 ();
 sg13g2_fill_8 FILLER_94_402 ();
 sg13g2_fill_4 FILLER_94_410 ();
 sg13g2_fill_2 FILLER_94_414 ();
 sg13g2_fill_1 FILLER_94_416 ();
 sg13g2_fill_2 FILLER_94_427 ();
 sg13g2_fill_8 FILLER_94_439 ();
 sg13g2_fill_2 FILLER_94_447 ();
 sg13g2_fill_1 FILLER_94_449 ();
 sg13g2_fill_1 FILLER_94_475 ();
 sg13g2_fill_4 FILLER_94_497 ();
 sg13g2_fill_2 FILLER_94_506 ();
 sg13g2_fill_8 FILLER_94_527 ();
 sg13g2_fill_4 FILLER_94_535 ();
 sg13g2_fill_1 FILLER_94_549 ();
 sg13g2_fill_4 FILLER_94_556 ();
 sg13g2_fill_1 FILLER_94_567 ();
 sg13g2_fill_8 FILLER_94_573 ();
 sg13g2_fill_8 FILLER_94_581 ();
 sg13g2_fill_8 FILLER_94_589 ();
 sg13g2_fill_2 FILLER_94_597 ();
 sg13g2_fill_1 FILLER_94_609 ();
 sg13g2_fill_4 FILLER_94_636 ();
 sg13g2_fill_1 FILLER_94_640 ();
 sg13g2_fill_8 FILLER_94_743 ();
 sg13g2_fill_8 FILLER_94_751 ();
 sg13g2_fill_8 FILLER_94_759 ();
 sg13g2_fill_2 FILLER_94_767 ();
 sg13g2_fill_4 FILLER_94_772 ();
 sg13g2_fill_2 FILLER_94_776 ();
 sg13g2_fill_8 FILLER_94_786 ();
 sg13g2_fill_8 FILLER_94_794 ();
 sg13g2_fill_8 FILLER_94_802 ();
 sg13g2_fill_8 FILLER_94_810 ();
 sg13g2_fill_8 FILLER_94_818 ();
 sg13g2_fill_8 FILLER_94_826 ();
 sg13g2_fill_4 FILLER_94_834 ();
 sg13g2_fill_2 FILLER_94_838 ();
 sg13g2_fill_1 FILLER_94_840 ();
 sg13g2_fill_4 FILLER_94_845 ();
 sg13g2_fill_2 FILLER_94_849 ();
 sg13g2_fill_1 FILLER_94_868 ();
 sg13g2_fill_4 FILLER_94_888 ();
 sg13g2_fill_1 FILLER_94_892 ();
 sg13g2_fill_1 FILLER_94_898 ();
 sg13g2_fill_4 FILLER_94_902 ();
 sg13g2_fill_8 FILLER_94_911 ();
 sg13g2_fill_4 FILLER_94_937 ();
 sg13g2_fill_8 FILLER_94_961 ();
 sg13g2_fill_1 FILLER_94_974 ();
 sg13g2_fill_8 FILLER_94_1012 ();
 sg13g2_fill_2 FILLER_94_1020 ();
 sg13g2_fill_8 FILLER_94_1033 ();
 sg13g2_fill_8 FILLER_94_1041 ();
 sg13g2_fill_4 FILLER_94_1049 ();
 sg13g2_fill_1 FILLER_94_1053 ();
 sg13g2_fill_8 FILLER_94_1057 ();
 sg13g2_fill_8 FILLER_94_1065 ();
 sg13g2_fill_1 FILLER_94_1073 ();
 sg13g2_fill_2 FILLER_94_1083 ();
 sg13g2_fill_1 FILLER_94_1085 ();
 sg13g2_fill_8 FILLER_94_1091 ();
 sg13g2_fill_8 FILLER_94_1099 ();
 sg13g2_fill_8 FILLER_94_1132 ();
 sg13g2_fill_4 FILLER_94_1140 ();
 sg13g2_fill_1 FILLER_94_1144 ();
 sg13g2_fill_4 FILLER_94_1159 ();
 sg13g2_fill_2 FILLER_94_1163 ();
 sg13g2_fill_1 FILLER_94_1165 ();
 sg13g2_fill_1 FILLER_94_1183 ();
 sg13g2_fill_1 FILLER_94_1198 ();
 sg13g2_fill_4 FILLER_94_1233 ();
 sg13g2_fill_2 FILLER_94_1237 ();
 sg13g2_fill_2 FILLER_94_1243 ();
 sg13g2_fill_1 FILLER_94_1245 ();
 sg13g2_fill_1 FILLER_94_1259 ();
 sg13g2_fill_4 FILLER_94_1268 ();
 sg13g2_fill_1 FILLER_94_1272 ();
 sg13g2_fill_2 FILLER_94_1278 ();
 sg13g2_fill_8 FILLER_94_1297 ();
 sg13g2_fill_4 FILLER_94_1305 ();
 sg13g2_fill_4 FILLER_94_1313 ();
 sg13g2_fill_2 FILLER_94_1352 ();
 sg13g2_fill_8 FILLER_94_1374 ();
 sg13g2_fill_2 FILLER_94_1417 ();
 sg13g2_fill_4 FILLER_94_1445 ();
 sg13g2_fill_2 FILLER_94_1449 ();
 sg13g2_fill_2 FILLER_94_1474 ();
 sg13g2_fill_4 FILLER_94_1505 ();
 sg13g2_fill_4 FILLER_94_1531 ();
 sg13g2_fill_4 FILLER_94_1543 ();
 sg13g2_fill_8 FILLER_94_1570 ();
 sg13g2_fill_8 FILLER_94_1578 ();
 sg13g2_fill_4 FILLER_94_1586 ();
 sg13g2_fill_2 FILLER_94_1590 ();
 sg13g2_fill_8 FILLER_95_0 ();
 sg13g2_fill_8 FILLER_95_8 ();
 sg13g2_fill_8 FILLER_95_16 ();
 sg13g2_fill_4 FILLER_95_24 ();
 sg13g2_fill_2 FILLER_95_28 ();
 sg13g2_fill_4 FILLER_95_71 ();
 sg13g2_fill_1 FILLER_95_75 ();
 sg13g2_fill_2 FILLER_95_84 ();
 sg13g2_fill_1 FILLER_95_86 ();
 sg13g2_fill_1 FILLER_95_123 ();
 sg13g2_fill_8 FILLER_95_140 ();
 sg13g2_fill_8 FILLER_95_148 ();
 sg13g2_fill_4 FILLER_95_156 ();
 sg13g2_fill_2 FILLER_95_160 ();
 sg13g2_fill_4 FILLER_95_172 ();
 sg13g2_fill_2 FILLER_95_176 ();
 sg13g2_fill_1 FILLER_95_178 ();
 sg13g2_fill_8 FILLER_95_189 ();
 sg13g2_fill_2 FILLER_95_197 ();
 sg13g2_fill_1 FILLER_95_199 ();
 sg13g2_fill_4 FILLER_95_221 ();
 sg13g2_fill_1 FILLER_95_225 ();
 sg13g2_fill_8 FILLER_95_236 ();
 sg13g2_fill_4 FILLER_95_244 ();
 sg13g2_fill_4 FILLER_95_302 ();
 sg13g2_fill_1 FILLER_95_306 ();
 sg13g2_fill_8 FILLER_95_333 ();
 sg13g2_fill_8 FILLER_95_341 ();
 sg13g2_fill_8 FILLER_95_349 ();
 sg13g2_fill_8 FILLER_95_357 ();
 sg13g2_fill_8 FILLER_95_365 ();
 sg13g2_fill_8 FILLER_95_373 ();
 sg13g2_fill_4 FILLER_95_381 ();
 sg13g2_fill_8 FILLER_95_395 ();
 sg13g2_fill_4 FILLER_95_403 ();
 sg13g2_fill_4 FILLER_95_427 ();
 sg13g2_fill_2 FILLER_95_431 ();
 sg13g2_fill_8 FILLER_95_484 ();
 sg13g2_fill_4 FILLER_95_492 ();
 sg13g2_fill_1 FILLER_95_496 ();
 sg13g2_fill_1 FILLER_95_510 ();
 sg13g2_fill_4 FILLER_95_561 ();
 sg13g2_fill_4 FILLER_95_570 ();
 sg13g2_fill_1 FILLER_95_578 ();
 sg13g2_fill_8 FILLER_95_588 ();
 sg13g2_fill_4 FILLER_95_596 ();
 sg13g2_fill_4 FILLER_95_616 ();
 sg13g2_fill_2 FILLER_95_620 ();
 sg13g2_fill_1 FILLER_95_622 ();
 sg13g2_fill_8 FILLER_95_633 ();
 sg13g2_fill_4 FILLER_95_641 ();
 sg13g2_fill_2 FILLER_95_645 ();
 sg13g2_fill_1 FILLER_95_647 ();
 sg13g2_fill_8 FILLER_95_656 ();
 sg13g2_fill_4 FILLER_95_664 ();
 sg13g2_fill_1 FILLER_95_668 ();
 sg13g2_fill_8 FILLER_95_695 ();
 sg13g2_fill_8 FILLER_95_703 ();
 sg13g2_fill_8 FILLER_95_711 ();
 sg13g2_fill_4 FILLER_95_719 ();
 sg13g2_fill_8 FILLER_95_733 ();
 sg13g2_fill_1 FILLER_95_779 ();
 sg13g2_fill_4 FILLER_95_788 ();
 sg13g2_fill_1 FILLER_95_792 ();
 sg13g2_fill_4 FILLER_95_810 ();
 sg13g2_fill_2 FILLER_95_814 ();
 sg13g2_fill_8 FILLER_95_826 ();
 sg13g2_fill_2 FILLER_95_834 ();
 sg13g2_fill_1 FILLER_95_836 ();
 sg13g2_fill_8 FILLER_95_852 ();
 sg13g2_fill_4 FILLER_95_860 ();
 sg13g2_fill_1 FILLER_95_864 ();
 sg13g2_fill_2 FILLER_95_872 ();
 sg13g2_fill_1 FILLER_95_874 ();
 sg13g2_fill_4 FILLER_95_882 ();
 sg13g2_fill_1 FILLER_95_886 ();
 sg13g2_fill_1 FILLER_95_901 ();
 sg13g2_fill_4 FILLER_95_927 ();
 sg13g2_fill_1 FILLER_95_931 ();
 sg13g2_fill_8 FILLER_95_954 ();
 sg13g2_fill_2 FILLER_95_962 ();
 sg13g2_fill_1 FILLER_95_964 ();
 sg13g2_fill_2 FILLER_95_975 ();
 sg13g2_fill_4 FILLER_95_1030 ();
 sg13g2_fill_4 FILLER_95_1054 ();
 sg13g2_fill_1 FILLER_95_1058 ();
 sg13g2_fill_2 FILLER_95_1064 ();
 sg13g2_fill_1 FILLER_95_1074 ();
 sg13g2_fill_1 FILLER_95_1085 ();
 sg13g2_fill_8 FILLER_95_1096 ();
 sg13g2_fill_2 FILLER_95_1114 ();
 sg13g2_fill_4 FILLER_95_1121 ();
 sg13g2_fill_1 FILLER_95_1125 ();
 sg13g2_fill_2 FILLER_95_1149 ();
 sg13g2_fill_1 FILLER_95_1151 ();
 sg13g2_fill_8 FILLER_95_1160 ();
 sg13g2_fill_8 FILLER_95_1168 ();
 sg13g2_fill_8 FILLER_95_1176 ();
 sg13g2_fill_8 FILLER_95_1184 ();
 sg13g2_fill_2 FILLER_95_1192 ();
 sg13g2_fill_2 FILLER_95_1199 ();
 sg13g2_fill_8 FILLER_95_1206 ();
 sg13g2_fill_2 FILLER_95_1214 ();
 sg13g2_fill_8 FILLER_95_1220 ();
 sg13g2_fill_1 FILLER_95_1228 ();
 sg13g2_fill_8 FILLER_95_1261 ();
 sg13g2_fill_2 FILLER_95_1269 ();
 sg13g2_fill_1 FILLER_95_1271 ();
 sg13g2_fill_4 FILLER_95_1290 ();
 sg13g2_fill_2 FILLER_95_1294 ();
 sg13g2_fill_1 FILLER_95_1296 ();
 sg13g2_fill_2 FILLER_95_1302 ();
 sg13g2_fill_1 FILLER_95_1304 ();
 sg13g2_fill_1 FILLER_95_1310 ();
 sg13g2_fill_1 FILLER_95_1325 ();
 sg13g2_fill_8 FILLER_95_1330 ();
 sg13g2_fill_2 FILLER_95_1338 ();
 sg13g2_fill_2 FILLER_95_1359 ();
 sg13g2_fill_1 FILLER_95_1361 ();
 sg13g2_fill_1 FILLER_95_1370 ();
 sg13g2_fill_2 FILLER_95_1391 ();
 sg13g2_fill_1 FILLER_95_1393 ();
 sg13g2_fill_2 FILLER_95_1402 ();
 sg13g2_fill_1 FILLER_95_1404 ();
 sg13g2_fill_1 FILLER_95_1414 ();
 sg13g2_fill_8 FILLER_95_1428 ();
 sg13g2_fill_8 FILLER_95_1436 ();
 sg13g2_fill_8 FILLER_95_1444 ();
 sg13g2_fill_8 FILLER_95_1452 ();
 sg13g2_fill_4 FILLER_95_1460 ();
 sg13g2_fill_1 FILLER_95_1464 ();
 sg13g2_fill_2 FILLER_95_1471 ();
 sg13g2_fill_1 FILLER_95_1473 ();
 sg13g2_fill_8 FILLER_95_1499 ();
 sg13g2_fill_8 FILLER_95_1507 ();
 sg13g2_fill_1 FILLER_95_1515 ();
 sg13g2_fill_2 FILLER_95_1521 ();
 sg13g2_fill_1 FILLER_95_1523 ();
 sg13g2_fill_8 FILLER_95_1529 ();
 sg13g2_fill_2 FILLER_95_1537 ();
 sg13g2_fill_4 FILLER_95_1558 ();
 sg13g2_fill_8 FILLER_96_0 ();
 sg13g2_fill_8 FILLER_96_8 ();
 sg13g2_fill_8 FILLER_96_16 ();
 sg13g2_fill_8 FILLER_96_24 ();
 sg13g2_fill_8 FILLER_96_32 ();
 sg13g2_fill_8 FILLER_96_40 ();
 sg13g2_fill_8 FILLER_96_48 ();
 sg13g2_fill_8 FILLER_96_56 ();
 sg13g2_fill_8 FILLER_96_64 ();
 sg13g2_fill_4 FILLER_96_82 ();
 sg13g2_fill_8 FILLER_96_96 ();
 sg13g2_fill_1 FILLER_96_149 ();
 sg13g2_fill_1 FILLER_96_175 ();
 sg13g2_fill_4 FILLER_96_223 ();
 sg13g2_fill_1 FILLER_96_227 ();
 sg13g2_fill_8 FILLER_96_254 ();
 sg13g2_fill_1 FILLER_96_262 ();
 sg13g2_fill_8 FILLER_96_288 ();
 sg13g2_fill_8 FILLER_96_296 ();
 sg13g2_fill_2 FILLER_96_304 ();
 sg13g2_fill_1 FILLER_96_306 ();
 sg13g2_fill_8 FILLER_96_346 ();
 sg13g2_fill_8 FILLER_96_354 ();
 sg13g2_fill_8 FILLER_96_372 ();
 sg13g2_fill_4 FILLER_96_380 ();
 sg13g2_fill_2 FILLER_96_384 ();
 sg13g2_fill_1 FILLER_96_396 ();
 sg13g2_fill_1 FILLER_96_439 ();
 sg13g2_fill_4 FILLER_96_501 ();
 sg13g2_fill_1 FILLER_96_513 ();
 sg13g2_fill_8 FILLER_96_519 ();
 sg13g2_fill_8 FILLER_96_527 ();
 sg13g2_fill_8 FILLER_96_535 ();
 sg13g2_fill_8 FILLER_96_543 ();
 sg13g2_fill_8 FILLER_96_551 ();
 sg13g2_fill_8 FILLER_96_559 ();
 sg13g2_fill_8 FILLER_96_567 ();
 sg13g2_fill_4 FILLER_96_575 ();
 sg13g2_fill_1 FILLER_96_579 ();
 sg13g2_fill_4 FILLER_96_587 ();
 sg13g2_fill_2 FILLER_96_591 ();
 sg13g2_fill_1 FILLER_96_593 ();
 sg13g2_fill_2 FILLER_96_630 ();
 sg13g2_fill_8 FILLER_96_653 ();
 sg13g2_fill_8 FILLER_96_661 ();
 sg13g2_fill_8 FILLER_96_693 ();
 sg13g2_fill_8 FILLER_96_701 ();
 sg13g2_fill_8 FILLER_96_709 ();
 sg13g2_fill_4 FILLER_96_717 ();
 sg13g2_fill_1 FILLER_96_721 ();
 sg13g2_fill_4 FILLER_96_782 ();
 sg13g2_fill_4 FILLER_96_812 ();
 sg13g2_fill_2 FILLER_96_834 ();
 sg13g2_fill_2 FILLER_96_840 ();
 sg13g2_fill_1 FILLER_96_842 ();
 sg13g2_fill_1 FILLER_96_885 ();
 sg13g2_fill_1 FILLER_96_917 ();
 sg13g2_fill_8 FILLER_96_924 ();
 sg13g2_fill_4 FILLER_96_937 ();
 sg13g2_fill_1 FILLER_96_941 ();
 sg13g2_fill_4 FILLER_96_946 ();
 sg13g2_fill_2 FILLER_96_950 ();
 sg13g2_fill_4 FILLER_96_956 ();
 sg13g2_fill_4 FILLER_96_1026 ();
 sg13g2_fill_2 FILLER_96_1078 ();
 sg13g2_fill_1 FILLER_96_1080 ();
 sg13g2_fill_1 FILLER_96_1085 ();
 sg13g2_fill_1 FILLER_96_1090 ();
 sg13g2_fill_8 FILLER_96_1096 ();
 sg13g2_fill_4 FILLER_96_1104 ();
 sg13g2_fill_1 FILLER_96_1113 ();
 sg13g2_fill_8 FILLER_96_1119 ();
 sg13g2_fill_8 FILLER_96_1127 ();
 sg13g2_fill_8 FILLER_96_1135 ();
 sg13g2_fill_4 FILLER_96_1167 ();
 sg13g2_fill_2 FILLER_96_1171 ();
 sg13g2_fill_1 FILLER_96_1173 ();
 sg13g2_fill_1 FILLER_96_1198 ();
 sg13g2_fill_1 FILLER_96_1204 ();
 sg13g2_fill_4 FILLER_96_1215 ();
 sg13g2_fill_2 FILLER_96_1219 ();
 sg13g2_fill_1 FILLER_96_1221 ();
 sg13g2_fill_2 FILLER_96_1237 ();
 sg13g2_fill_1 FILLER_96_1239 ();
 sg13g2_fill_8 FILLER_96_1248 ();
 sg13g2_fill_8 FILLER_96_1256 ();
 sg13g2_fill_8 FILLER_96_1264 ();
 sg13g2_fill_4 FILLER_96_1272 ();
 sg13g2_fill_2 FILLER_96_1285 ();
 sg13g2_fill_1 FILLER_96_1287 ();
 sg13g2_fill_4 FILLER_96_1293 ();
 sg13g2_fill_2 FILLER_96_1297 ();
 sg13g2_fill_8 FILLER_96_1323 ();
 sg13g2_fill_2 FILLER_96_1331 ();
 sg13g2_fill_1 FILLER_96_1333 ();
 sg13g2_fill_1 FILLER_96_1344 ();
 sg13g2_fill_1 FILLER_96_1360 ();
 sg13g2_fill_1 FILLER_96_1384 ();
 sg13g2_fill_8 FILLER_96_1389 ();
 sg13g2_fill_8 FILLER_96_1497 ();
 sg13g2_fill_2 FILLER_96_1515 ();
 sg13g2_fill_1 FILLER_96_1517 ();
 sg13g2_fill_4 FILLER_96_1529 ();
 sg13g2_fill_2 FILLER_96_1533 ();
 sg13g2_fill_1 FILLER_96_1535 ();
 sg13g2_fill_8 FILLER_96_1547 ();
 sg13g2_fill_8 FILLER_96_1555 ();
 sg13g2_fill_8 FILLER_96_1563 ();
 sg13g2_fill_4 FILLER_96_1571 ();
 sg13g2_fill_2 FILLER_96_1575 ();
 sg13g2_fill_2 FILLER_96_1590 ();
 sg13g2_fill_8 FILLER_97_0 ();
 sg13g2_fill_8 FILLER_97_8 ();
 sg13g2_fill_8 FILLER_97_16 ();
 sg13g2_fill_8 FILLER_97_24 ();
 sg13g2_fill_8 FILLER_97_32 ();
 sg13g2_fill_8 FILLER_97_40 ();
 sg13g2_fill_2 FILLER_97_48 ();
 sg13g2_fill_8 FILLER_97_84 ();
 sg13g2_fill_8 FILLER_97_92 ();
 sg13g2_fill_2 FILLER_97_100 ();
 sg13g2_fill_8 FILLER_97_107 ();
 sg13g2_fill_8 FILLER_97_115 ();
 sg13g2_fill_2 FILLER_97_123 ();
 sg13g2_fill_1 FILLER_97_135 ();
 sg13g2_fill_8 FILLER_97_180 ();
 sg13g2_fill_8 FILLER_97_188 ();
 sg13g2_fill_2 FILLER_97_196 ();
 sg13g2_fill_1 FILLER_97_198 ();
 sg13g2_fill_2 FILLER_97_209 ();
 sg13g2_fill_8 FILLER_97_227 ();
 sg13g2_fill_4 FILLER_97_235 ();
 sg13g2_fill_1 FILLER_97_239 ();
 sg13g2_fill_8 FILLER_97_313 ();
 sg13g2_fill_2 FILLER_97_321 ();
 sg13g2_fill_2 FILLER_97_333 ();
 sg13g2_fill_1 FILLER_97_335 ();
 sg13g2_fill_4 FILLER_97_362 ();
 sg13g2_fill_8 FILLER_97_392 ();
 sg13g2_fill_8 FILLER_97_400 ();
 sg13g2_fill_1 FILLER_97_408 ();
 sg13g2_fill_2 FILLER_97_420 ();
 sg13g2_fill_8 FILLER_97_428 ();
 sg13g2_fill_8 FILLER_97_436 ();
 sg13g2_fill_4 FILLER_97_470 ();
 sg13g2_fill_2 FILLER_97_474 ();
 sg13g2_fill_1 FILLER_97_476 ();
 sg13g2_fill_8 FILLER_97_502 ();
 sg13g2_fill_8 FILLER_97_510 ();
 sg13g2_fill_8 FILLER_97_518 ();
 sg13g2_fill_8 FILLER_97_526 ();
 sg13g2_fill_4 FILLER_97_534 ();
 sg13g2_fill_2 FILLER_97_538 ();
 sg13g2_fill_1 FILLER_97_540 ();
 sg13g2_fill_4 FILLER_97_551 ();
 sg13g2_fill_2 FILLER_97_555 ();
 sg13g2_fill_1 FILLER_97_557 ();
 sg13g2_fill_4 FILLER_97_574 ();
 sg13g2_fill_4 FILLER_97_588 ();
 sg13g2_fill_2 FILLER_97_592 ();
 sg13g2_fill_4 FILLER_97_599 ();
 sg13g2_fill_1 FILLER_97_603 ();
 sg13g2_fill_8 FILLER_97_614 ();
 sg13g2_fill_4 FILLER_97_622 ();
 sg13g2_fill_1 FILLER_97_626 ();
 sg13g2_fill_4 FILLER_97_633 ();
 sg13g2_fill_2 FILLER_97_637 ();
 sg13g2_fill_1 FILLER_97_639 ();
 sg13g2_fill_2 FILLER_97_676 ();
 sg13g2_fill_4 FILLER_97_688 ();
 sg13g2_fill_2 FILLER_97_692 ();
 sg13g2_fill_1 FILLER_97_694 ();
 sg13g2_fill_8 FILLER_97_721 ();
 sg13g2_fill_8 FILLER_97_729 ();
 sg13g2_fill_8 FILLER_97_737 ();
 sg13g2_fill_8 FILLER_97_745 ();
 sg13g2_fill_8 FILLER_97_753 ();
 sg13g2_fill_1 FILLER_97_761 ();
 sg13g2_fill_8 FILLER_97_772 ();
 sg13g2_fill_8 FILLER_97_780 ();
 sg13g2_fill_2 FILLER_97_788 ();
 sg13g2_fill_4 FILLER_97_839 ();
 sg13g2_fill_1 FILLER_97_843 ();
 sg13g2_fill_8 FILLER_97_852 ();
 sg13g2_fill_8 FILLER_97_860 ();
 sg13g2_fill_1 FILLER_97_868 ();
 sg13g2_fill_4 FILLER_97_882 ();
 sg13g2_fill_2 FILLER_97_894 ();
 sg13g2_fill_8 FILLER_97_900 ();
 sg13g2_fill_4 FILLER_97_908 ();
 sg13g2_fill_2 FILLER_97_915 ();
 sg13g2_fill_1 FILLER_97_917 ();
 sg13g2_fill_4 FILLER_97_934 ();
 sg13g2_fill_2 FILLER_97_944 ();
 sg13g2_fill_1 FILLER_97_946 ();
 sg13g2_fill_1 FILLER_97_952 ();
 sg13g2_fill_8 FILLER_97_957 ();
 sg13g2_fill_2 FILLER_97_965 ();
 sg13g2_fill_1 FILLER_97_967 ();
 sg13g2_fill_1 FILLER_97_976 ();
 sg13g2_fill_8 FILLER_97_994 ();
 sg13g2_fill_4 FILLER_97_1002 ();
 sg13g2_fill_1 FILLER_97_1006 ();
 sg13g2_fill_4 FILLER_97_1035 ();
 sg13g2_fill_8 FILLER_97_1045 ();
 sg13g2_fill_4 FILLER_97_1053 ();
 sg13g2_fill_1 FILLER_97_1080 ();
 sg13g2_fill_4 FILLER_97_1113 ();
 sg13g2_fill_8 FILLER_97_1122 ();
 sg13g2_fill_8 FILLER_97_1138 ();
 sg13g2_fill_8 FILLER_97_1146 ();
 sg13g2_fill_8 FILLER_97_1154 ();
 sg13g2_fill_2 FILLER_97_1162 ();
 sg13g2_fill_1 FILLER_97_1164 ();
 sg13g2_fill_4 FILLER_97_1173 ();
 sg13g2_fill_2 FILLER_97_1177 ();
 sg13g2_fill_8 FILLER_97_1195 ();
 sg13g2_fill_1 FILLER_97_1203 ();
 sg13g2_fill_8 FILLER_97_1208 ();
 sg13g2_fill_8 FILLER_97_1221 ();
 sg13g2_fill_4 FILLER_97_1229 ();
 sg13g2_fill_2 FILLER_97_1233 ();
 sg13g2_fill_8 FILLER_97_1246 ();
 sg13g2_fill_2 FILLER_97_1254 ();
 sg13g2_fill_1 FILLER_97_1256 ();
 sg13g2_fill_2 FILLER_97_1262 ();
 sg13g2_fill_1 FILLER_97_1264 ();
 sg13g2_fill_8 FILLER_97_1286 ();
 sg13g2_fill_2 FILLER_97_1294 ();
 sg13g2_fill_1 FILLER_97_1296 ();
 sg13g2_fill_1 FILLER_97_1301 ();
 sg13g2_fill_8 FILLER_97_1316 ();
 sg13g2_fill_4 FILLER_97_1324 ();
 sg13g2_fill_1 FILLER_97_1328 ();
 sg13g2_fill_8 FILLER_97_1340 ();
 sg13g2_fill_2 FILLER_97_1348 ();
 sg13g2_fill_1 FILLER_97_1350 ();
 sg13g2_fill_4 FILLER_97_1356 ();
 sg13g2_fill_2 FILLER_97_1360 ();
 sg13g2_fill_1 FILLER_97_1362 ();
 sg13g2_fill_4 FILLER_97_1366 ();
 sg13g2_fill_8 FILLER_97_1384 ();
 sg13g2_fill_8 FILLER_97_1392 ();
 sg13g2_fill_1 FILLER_97_1404 ();
 sg13g2_fill_8 FILLER_97_1408 ();
 sg13g2_fill_4 FILLER_97_1416 ();
 sg13g2_fill_2 FILLER_97_1420 ();
 sg13g2_fill_1 FILLER_97_1422 ();
 sg13g2_fill_4 FILLER_97_1427 ();
 sg13g2_fill_8 FILLER_97_1452 ();
 sg13g2_fill_1 FILLER_97_1460 ();
 sg13g2_fill_4 FILLER_97_1494 ();
 sg13g2_fill_2 FILLER_97_1498 ();
 sg13g2_fill_8 FILLER_97_1526 ();
 sg13g2_fill_2 FILLER_97_1534 ();
 sg13g2_fill_4 FILLER_97_1540 ();
 sg13g2_fill_1 FILLER_97_1544 ();
 sg13g2_fill_4 FILLER_97_1587 ();
 sg13g2_fill_1 FILLER_97_1591 ();
 sg13g2_fill_8 FILLER_98_0 ();
 sg13g2_fill_8 FILLER_98_8 ();
 sg13g2_fill_8 FILLER_98_16 ();
 sg13g2_fill_8 FILLER_98_24 ();
 sg13g2_fill_8 FILLER_98_32 ();
 sg13g2_fill_8 FILLER_98_40 ();
 sg13g2_fill_4 FILLER_98_48 ();
 sg13g2_fill_2 FILLER_98_52 ();
 sg13g2_fill_1 FILLER_98_54 ();
 sg13g2_fill_8 FILLER_98_65 ();
 sg13g2_fill_8 FILLER_98_125 ();
 sg13g2_fill_8 FILLER_98_133 ();
 sg13g2_fill_2 FILLER_98_141 ();
 sg13g2_fill_1 FILLER_98_143 ();
 sg13g2_fill_2 FILLER_98_148 ();
 sg13g2_fill_1 FILLER_98_161 ();
 sg13g2_fill_4 FILLER_98_167 ();
 sg13g2_fill_1 FILLER_98_171 ();
 sg13g2_fill_2 FILLER_98_198 ();
 sg13g2_fill_8 FILLER_98_226 ();
 sg13g2_fill_1 FILLER_98_234 ();
 sg13g2_fill_8 FILLER_98_270 ();
 sg13g2_fill_8 FILLER_98_278 ();
 sg13g2_fill_2 FILLER_98_286 ();
 sg13g2_fill_8 FILLER_98_327 ();
 sg13g2_fill_4 FILLER_98_335 ();
 sg13g2_fill_2 FILLER_98_339 ();
 sg13g2_fill_4 FILLER_98_362 ();
 sg13g2_fill_2 FILLER_98_366 ();
 sg13g2_fill_1 FILLER_98_394 ();
 sg13g2_fill_2 FILLER_98_400 ();
 sg13g2_fill_2 FILLER_98_427 ();
 sg13g2_fill_4 FILLER_98_434 ();
 sg13g2_fill_8 FILLER_98_447 ();
 sg13g2_fill_8 FILLER_98_455 ();
 sg13g2_fill_8 FILLER_98_463 ();
 sg13g2_fill_4 FILLER_98_471 ();
 sg13g2_fill_8 FILLER_98_491 ();
 sg13g2_fill_4 FILLER_98_499 ();
 sg13g2_fill_2 FILLER_98_503 ();
 sg13g2_fill_1 FILLER_98_577 ();
 sg13g2_fill_8 FILLER_98_604 ();
 sg13g2_fill_2 FILLER_98_638 ();
 sg13g2_fill_1 FILLER_98_640 ();
 sg13g2_fill_8 FILLER_98_649 ();
 sg13g2_fill_4 FILLER_98_657 ();
 sg13g2_fill_2 FILLER_98_661 ();
 sg13g2_fill_4 FILLER_98_671 ();
 sg13g2_fill_1 FILLER_98_675 ();
 sg13g2_fill_2 FILLER_98_696 ();
 sg13g2_fill_4 FILLER_98_794 ();
 sg13g2_fill_2 FILLER_98_804 ();
 sg13g2_fill_1 FILLER_98_806 ();
 sg13g2_fill_4 FILLER_98_812 ();
 sg13g2_fill_1 FILLER_98_816 ();
 sg13g2_fill_4 FILLER_98_821 ();
 sg13g2_fill_2 FILLER_98_830 ();
 sg13g2_fill_4 FILLER_98_859 ();
 sg13g2_fill_1 FILLER_98_863 ();
 sg13g2_fill_8 FILLER_98_878 ();
 sg13g2_fill_8 FILLER_98_886 ();
 sg13g2_fill_2 FILLER_98_894 ();
 sg13g2_fill_4 FILLER_98_906 ();
 sg13g2_fill_2 FILLER_98_910 ();
 sg13g2_fill_8 FILLER_98_916 ();
 sg13g2_fill_8 FILLER_98_924 ();
 sg13g2_fill_4 FILLER_98_932 ();
 sg13g2_fill_1 FILLER_98_936 ();
 sg13g2_fill_2 FILLER_98_941 ();
 sg13g2_fill_1 FILLER_98_957 ();
 sg13g2_fill_2 FILLER_98_961 ();
 sg13g2_fill_1 FILLER_98_963 ();
 sg13g2_fill_4 FILLER_98_989 ();
 sg13g2_fill_2 FILLER_98_993 ();
 sg13g2_fill_1 FILLER_98_995 ();
 sg13g2_fill_2 FILLER_98_1001 ();
 sg13g2_fill_1 FILLER_98_1006 ();
 sg13g2_fill_2 FILLER_98_1017 ();
 sg13g2_fill_8 FILLER_98_1027 ();
 sg13g2_fill_2 FILLER_98_1035 ();
 sg13g2_fill_1 FILLER_98_1037 ();
 sg13g2_fill_8 FILLER_98_1044 ();
 sg13g2_fill_8 FILLER_98_1052 ();
 sg13g2_fill_4 FILLER_98_1060 ();
 sg13g2_fill_1 FILLER_98_1064 ();
 sg13g2_fill_2 FILLER_98_1075 ();
 sg13g2_fill_1 FILLER_98_1077 ();
 sg13g2_fill_4 FILLER_98_1081 ();
 sg13g2_fill_2 FILLER_98_1085 ();
 sg13g2_fill_8 FILLER_98_1098 ();
 sg13g2_fill_2 FILLER_98_1114 ();
 sg13g2_fill_1 FILLER_98_1116 ();
 sg13g2_fill_4 FILLER_98_1135 ();
 sg13g2_fill_2 FILLER_98_1139 ();
 sg13g2_fill_2 FILLER_98_1146 ();
 sg13g2_fill_8 FILLER_98_1156 ();
 sg13g2_fill_1 FILLER_98_1164 ();
 sg13g2_fill_8 FILLER_98_1175 ();
 sg13g2_fill_8 FILLER_98_1183 ();
 sg13g2_fill_8 FILLER_98_1197 ();
 sg13g2_fill_4 FILLER_98_1205 ();
 sg13g2_fill_1 FILLER_98_1209 ();
 sg13g2_fill_2 FILLER_98_1215 ();
 sg13g2_fill_8 FILLER_98_1222 ();
 sg13g2_fill_8 FILLER_98_1230 ();
 sg13g2_fill_4 FILLER_98_1238 ();
 sg13g2_fill_1 FILLER_98_1242 ();
 sg13g2_fill_4 FILLER_98_1256 ();
 sg13g2_fill_4 FILLER_98_1264 ();
 sg13g2_fill_1 FILLER_98_1268 ();
 sg13g2_fill_2 FILLER_98_1273 ();
 sg13g2_fill_8 FILLER_98_1281 ();
 sg13g2_fill_8 FILLER_98_1289 ();
 sg13g2_fill_4 FILLER_98_1297 ();
 sg13g2_fill_8 FILLER_98_1304 ();
 sg13g2_fill_8 FILLER_98_1312 ();
 sg13g2_fill_8 FILLER_98_1320 ();
 sg13g2_fill_2 FILLER_98_1328 ();
 sg13g2_fill_1 FILLER_98_1330 ();
 sg13g2_fill_4 FILLER_98_1335 ();
 sg13g2_fill_1 FILLER_98_1339 ();
 sg13g2_fill_8 FILLER_98_1344 ();
 sg13g2_fill_8 FILLER_98_1352 ();
 sg13g2_fill_8 FILLER_98_1360 ();
 sg13g2_fill_1 FILLER_98_1368 ();
 sg13g2_fill_8 FILLER_98_1373 ();
 sg13g2_fill_8 FILLER_98_1381 ();
 sg13g2_fill_2 FILLER_98_1389 ();
 sg13g2_fill_1 FILLER_98_1391 ();
 sg13g2_fill_1 FILLER_98_1397 ();
 sg13g2_fill_2 FILLER_98_1403 ();
 sg13g2_fill_2 FILLER_98_1408 ();
 sg13g2_fill_8 FILLER_98_1441 ();
 sg13g2_fill_4 FILLER_98_1449 ();
 sg13g2_fill_2 FILLER_98_1453 ();
 sg13g2_fill_1 FILLER_98_1455 ();
 sg13g2_fill_2 FILLER_98_1486 ();
 sg13g2_fill_2 FILLER_98_1500 ();
 sg13g2_fill_8 FILLER_98_1512 ();
 sg13g2_fill_2 FILLER_98_1520 ();
 sg13g2_fill_1 FILLER_98_1522 ();
 sg13g2_fill_2 FILLER_98_1529 ();
 sg13g2_fill_1 FILLER_98_1531 ();
 sg13g2_fill_2 FILLER_98_1546 ();
 sg13g2_fill_4 FILLER_98_1553 ();
 sg13g2_fill_2 FILLER_98_1557 ();
 sg13g2_fill_4 FILLER_98_1563 ();
 sg13g2_fill_8 FILLER_98_1572 ();
 sg13g2_fill_8 FILLER_98_1580 ();
 sg13g2_fill_4 FILLER_98_1588 ();
 sg13g2_fill_8 FILLER_99_0 ();
 sg13g2_fill_8 FILLER_99_8 ();
 sg13g2_fill_8 FILLER_99_16 ();
 sg13g2_fill_8 FILLER_99_24 ();
 sg13g2_fill_8 FILLER_99_32 ();
 sg13g2_fill_8 FILLER_99_40 ();
 sg13g2_fill_8 FILLER_99_48 ();
 sg13g2_fill_8 FILLER_99_56 ();
 sg13g2_fill_4 FILLER_99_64 ();
 sg13g2_fill_2 FILLER_99_68 ();
 sg13g2_fill_2 FILLER_99_105 ();
 sg13g2_fill_4 FILLER_99_117 ();
 sg13g2_fill_8 FILLER_99_137 ();
 sg13g2_fill_8 FILLER_99_145 ();
 sg13g2_fill_8 FILLER_99_153 ();
 sg13g2_fill_4 FILLER_99_161 ();
 sg13g2_fill_2 FILLER_99_165 ();
 sg13g2_fill_8 FILLER_99_177 ();
 sg13g2_fill_8 FILLER_99_185 ();
 sg13g2_fill_2 FILLER_99_193 ();
 sg13g2_fill_4 FILLER_99_224 ();
 sg13g2_fill_4 FILLER_99_238 ();
 sg13g2_fill_2 FILLER_99_267 ();
 sg13g2_fill_2 FILLER_99_313 ();
 sg13g2_fill_8 FILLER_99_351 ();
 sg13g2_fill_8 FILLER_99_359 ();
 sg13g2_fill_8 FILLER_99_367 ();
 sg13g2_fill_2 FILLER_99_375 ();
 sg13g2_fill_1 FILLER_99_377 ();
 sg13g2_fill_1 FILLER_99_396 ();
 sg13g2_fill_2 FILLER_99_438 ();
 sg13g2_fill_8 FILLER_99_458 ();
 sg13g2_fill_1 FILLER_99_466 ();
 sg13g2_fill_4 FILLER_99_477 ();
 sg13g2_fill_1 FILLER_99_481 ();
 sg13g2_fill_4 FILLER_99_492 ();
 sg13g2_fill_2 FILLER_99_532 ();
 sg13g2_fill_1 FILLER_99_534 ();
 sg13g2_fill_8 FILLER_99_560 ();
 sg13g2_fill_4 FILLER_99_568 ();
 sg13g2_fill_2 FILLER_99_572 ();
 sg13g2_fill_4 FILLER_99_580 ();
 sg13g2_fill_8 FILLER_99_589 ();
 sg13g2_fill_4 FILLER_99_597 ();
 sg13g2_fill_1 FILLER_99_601 ();
 sg13g2_fill_8 FILLER_99_612 ();
 sg13g2_fill_4 FILLER_99_620 ();
 sg13g2_fill_1 FILLER_99_624 ();
 sg13g2_fill_2 FILLER_99_635 ();
 sg13g2_fill_1 FILLER_99_637 ();
 sg13g2_fill_1 FILLER_99_643 ();
 sg13g2_fill_8 FILLER_99_652 ();
 sg13g2_fill_4 FILLER_99_660 ();
 sg13g2_fill_2 FILLER_99_664 ();
 sg13g2_fill_1 FILLER_99_666 ();
 sg13g2_fill_8 FILLER_99_672 ();
 sg13g2_fill_8 FILLER_99_680 ();
 sg13g2_fill_4 FILLER_99_688 ();
 sg13g2_fill_2 FILLER_99_692 ();
 sg13g2_fill_1 FILLER_99_694 ();
 sg13g2_fill_8 FILLER_99_724 ();
 sg13g2_fill_8 FILLER_99_732 ();
 sg13g2_fill_8 FILLER_99_740 ();
 sg13g2_fill_8 FILLER_99_748 ();
 sg13g2_fill_8 FILLER_99_756 ();
 sg13g2_fill_8 FILLER_99_764 ();
 sg13g2_fill_8 FILLER_99_772 ();
 sg13g2_fill_4 FILLER_99_785 ();
 sg13g2_fill_2 FILLER_99_789 ();
 sg13g2_fill_1 FILLER_99_791 ();
 sg13g2_fill_1 FILLER_99_805 ();
 sg13g2_fill_2 FILLER_99_816 ();
 sg13g2_fill_1 FILLER_99_848 ();
 sg13g2_fill_4 FILLER_99_854 ();
 sg13g2_fill_8 FILLER_99_880 ();
 sg13g2_fill_2 FILLER_99_888 ();
 sg13g2_fill_1 FILLER_99_940 ();
 sg13g2_fill_1 FILLER_99_944 ();
 sg13g2_fill_4 FILLER_99_955 ();
 sg13g2_fill_1 FILLER_99_959 ();
 sg13g2_fill_4 FILLER_99_984 ();
 sg13g2_fill_4 FILLER_99_996 ();
 sg13g2_fill_2 FILLER_99_1000 ();
 sg13g2_fill_1 FILLER_99_1002 ();
 sg13g2_fill_2 FILLER_99_1043 ();
 sg13g2_fill_1 FILLER_99_1045 ();
 sg13g2_fill_8 FILLER_99_1059 ();
 sg13g2_fill_8 FILLER_99_1067 ();
 sg13g2_fill_2 FILLER_99_1075 ();
 sg13g2_fill_1 FILLER_99_1077 ();
 sg13g2_fill_8 FILLER_99_1096 ();
 sg13g2_fill_4 FILLER_99_1104 ();
 sg13g2_fill_1 FILLER_99_1108 ();
 sg13g2_fill_2 FILLER_99_1114 ();
 sg13g2_fill_1 FILLER_99_1116 ();
 sg13g2_fill_1 FILLER_99_1130 ();
 sg13g2_fill_1 FILLER_99_1136 ();
 sg13g2_fill_4 FILLER_99_1143 ();
 sg13g2_fill_1 FILLER_99_1147 ();
 sg13g2_fill_8 FILLER_99_1194 ();
 sg13g2_fill_2 FILLER_99_1202 ();
 sg13g2_fill_2 FILLER_99_1235 ();
 sg13g2_fill_1 FILLER_99_1264 ();
 sg13g2_fill_4 FILLER_99_1270 ();
 sg13g2_fill_1 FILLER_99_1274 ();
 sg13g2_fill_8 FILLER_99_1280 ();
 sg13g2_fill_4 FILLER_99_1310 ();
 sg13g2_fill_2 FILLER_99_1333 ();
 sg13g2_fill_4 FILLER_99_1343 ();
 sg13g2_fill_2 FILLER_99_1355 ();
 sg13g2_fill_1 FILLER_99_1357 ();
 sg13g2_fill_4 FILLER_99_1379 ();
 sg13g2_fill_4 FILLER_99_1410 ();
 sg13g2_fill_2 FILLER_99_1414 ();
 sg13g2_fill_4 FILLER_99_1420 ();
 sg13g2_fill_2 FILLER_99_1424 ();
 sg13g2_fill_8 FILLER_99_1430 ();
 sg13g2_fill_4 FILLER_99_1438 ();
 sg13g2_fill_2 FILLER_99_1442 ();
 sg13g2_fill_4 FILLER_99_1474 ();
 sg13g2_fill_4 FILLER_99_1517 ();
 sg13g2_fill_8 FILLER_99_1533 ();
 sg13g2_fill_8 FILLER_99_1541 ();
 sg13g2_fill_2 FILLER_99_1549 ();
 sg13g2_fill_1 FILLER_99_1551 ();
 sg13g2_fill_8 FILLER_100_0 ();
 sg13g2_fill_8 FILLER_100_8 ();
 sg13g2_fill_8 FILLER_100_16 ();
 sg13g2_fill_8 FILLER_100_24 ();
 sg13g2_fill_8 FILLER_100_32 ();
 sg13g2_fill_8 FILLER_100_40 ();
 sg13g2_fill_8 FILLER_100_48 ();
 sg13g2_fill_2 FILLER_100_56 ();
 sg13g2_fill_1 FILLER_100_58 ();
 sg13g2_fill_8 FILLER_100_69 ();
 sg13g2_fill_2 FILLER_100_77 ();
 sg13g2_fill_1 FILLER_100_79 ();
 sg13g2_fill_2 FILLER_100_83 ();
 sg13g2_fill_1 FILLER_100_111 ();
 sg13g2_fill_4 FILLER_100_132 ();
 sg13g2_fill_8 FILLER_100_150 ();
 sg13g2_fill_4 FILLER_100_158 ();
 sg13g2_fill_2 FILLER_100_162 ();
 sg13g2_fill_1 FILLER_100_164 ();
 sg13g2_fill_8 FILLER_100_175 ();
 sg13g2_fill_8 FILLER_100_183 ();
 sg13g2_fill_4 FILLER_100_191 ();
 sg13g2_fill_1 FILLER_100_195 ();
 sg13g2_fill_8 FILLER_100_217 ();
 sg13g2_fill_4 FILLER_100_225 ();
 sg13g2_fill_8 FILLER_100_276 ();
 sg13g2_fill_8 FILLER_100_284 ();
 sg13g2_fill_8 FILLER_100_292 ();
 sg13g2_fill_8 FILLER_100_300 ();
 sg13g2_fill_1 FILLER_100_308 ();
 sg13g2_fill_8 FILLER_100_317 ();
 sg13g2_fill_4 FILLER_100_325 ();
 sg13g2_fill_1 FILLER_100_329 ();
 sg13g2_fill_8 FILLER_100_366 ();
 sg13g2_fill_8 FILLER_100_374 ();
 sg13g2_fill_4 FILLER_100_382 ();
 sg13g2_fill_2 FILLER_100_386 ();
 sg13g2_fill_1 FILLER_100_388 ();
 sg13g2_fill_4 FILLER_100_397 ();
 sg13g2_fill_1 FILLER_100_401 ();
 sg13g2_fill_2 FILLER_100_427 ();
 sg13g2_fill_8 FILLER_100_489 ();
 sg13g2_fill_4 FILLER_100_497 ();
 sg13g2_fill_2 FILLER_100_501 ();
 sg13g2_fill_8 FILLER_100_511 ();
 sg13g2_fill_1 FILLER_100_519 ();
 sg13g2_fill_8 FILLER_100_546 ();
 sg13g2_fill_1 FILLER_100_554 ();
 sg13g2_fill_4 FILLER_100_575 ();
 sg13g2_fill_2 FILLER_100_579 ();
 sg13g2_fill_2 FILLER_100_595 ();
 sg13g2_fill_1 FILLER_100_597 ();
 sg13g2_fill_2 FILLER_100_634 ();
 sg13g2_fill_1 FILLER_100_636 ();
 sg13g2_fill_4 FILLER_100_653 ();
 sg13g2_fill_8 FILLER_100_678 ();
 sg13g2_fill_8 FILLER_100_686 ();
 sg13g2_fill_8 FILLER_100_694 ();
 sg13g2_fill_2 FILLER_100_702 ();
 sg13g2_fill_4 FILLER_100_730 ();
 sg13g2_fill_1 FILLER_100_734 ();
 sg13g2_fill_8 FILLER_100_743 ();
 sg13g2_fill_2 FILLER_100_785 ();
 sg13g2_fill_1 FILLER_100_787 ();
 sg13g2_fill_1 FILLER_100_800 ();
 sg13g2_fill_2 FILLER_100_811 ();
 sg13g2_fill_8 FILLER_100_847 ();
 sg13g2_fill_8 FILLER_100_855 ();
 sg13g2_fill_8 FILLER_100_863 ();
 sg13g2_fill_2 FILLER_100_871 ();
 sg13g2_fill_1 FILLER_100_873 ();
 sg13g2_fill_4 FILLER_100_886 ();
 sg13g2_fill_2 FILLER_100_890 ();
 sg13g2_fill_1 FILLER_100_892 ();
 sg13g2_fill_2 FILLER_100_898 ();
 sg13g2_fill_2 FILLER_100_909 ();
 sg13g2_fill_8 FILLER_100_919 ();
 sg13g2_fill_8 FILLER_100_932 ();
 sg13g2_fill_8 FILLER_100_940 ();
 sg13g2_fill_4 FILLER_100_948 ();
 sg13g2_fill_8 FILLER_100_956 ();
 sg13g2_fill_8 FILLER_100_964 ();
 sg13g2_fill_8 FILLER_100_972 ();
 sg13g2_fill_4 FILLER_100_980 ();
 sg13g2_fill_2 FILLER_100_984 ();
 sg13g2_fill_1 FILLER_100_986 ();
 sg13g2_fill_4 FILLER_100_992 ();
 sg13g2_fill_8 FILLER_100_1004 ();
 sg13g2_fill_8 FILLER_100_1012 ();
 sg13g2_fill_1 FILLER_100_1020 ();
 sg13g2_fill_8 FILLER_100_1025 ();
 sg13g2_fill_1 FILLER_100_1040 ();
 sg13g2_fill_2 FILLER_100_1051 ();
 sg13g2_fill_8 FILLER_100_1064 ();
 sg13g2_fill_4 FILLER_100_1072 ();
 sg13g2_fill_2 FILLER_100_1084 ();
 sg13g2_fill_8 FILLER_100_1091 ();
 sg13g2_fill_2 FILLER_100_1099 ();
 sg13g2_fill_4 FILLER_100_1106 ();
 sg13g2_fill_8 FILLER_100_1115 ();
 sg13g2_fill_8 FILLER_100_1123 ();
 sg13g2_fill_1 FILLER_100_1131 ();
 sg13g2_fill_2 FILLER_100_1156 ();
 sg13g2_fill_1 FILLER_100_1158 ();
 sg13g2_fill_4 FILLER_100_1164 ();
 sg13g2_fill_1 FILLER_100_1168 ();
 sg13g2_fill_8 FILLER_100_1174 ();
 sg13g2_fill_2 FILLER_100_1182 ();
 sg13g2_fill_1 FILLER_100_1184 ();
 sg13g2_fill_8 FILLER_100_1204 ();
 sg13g2_fill_4 FILLER_100_1212 ();
 sg13g2_fill_1 FILLER_100_1216 ();
 sg13g2_fill_2 FILLER_100_1235 ();
 sg13g2_fill_1 FILLER_100_1237 ();
 sg13g2_fill_4 FILLER_100_1254 ();
 sg13g2_fill_2 FILLER_100_1258 ();
 sg13g2_fill_1 FILLER_100_1260 ();
 sg13g2_fill_2 FILLER_100_1269 ();
 sg13g2_fill_1 FILLER_100_1335 ();
 sg13g2_fill_4 FILLER_100_1384 ();
 sg13g2_fill_2 FILLER_100_1388 ();
 sg13g2_fill_1 FILLER_100_1390 ();
 sg13g2_fill_4 FILLER_100_1403 ();
 sg13g2_fill_2 FILLER_100_1407 ();
 sg13g2_fill_1 FILLER_100_1409 ();
 sg13g2_fill_2 FILLER_100_1441 ();
 sg13g2_fill_4 FILLER_100_1503 ();
 sg13g2_fill_1 FILLER_100_1507 ();
 sg13g2_fill_2 FILLER_100_1514 ();
 sg13g2_fill_8 FILLER_100_1526 ();
 sg13g2_fill_2 FILLER_100_1534 ();
 sg13g2_fill_2 FILLER_100_1554 ();
 sg13g2_fill_4 FILLER_100_1572 ();
 sg13g2_fill_2 FILLER_100_1576 ();
 sg13g2_fill_1 FILLER_100_1578 ();
 sg13g2_fill_4 FILLER_100_1587 ();
 sg13g2_fill_1 FILLER_100_1591 ();
 sg13g2_fill_8 FILLER_101_0 ();
 sg13g2_fill_8 FILLER_101_8 ();
 sg13g2_fill_8 FILLER_101_16 ();
 sg13g2_fill_8 FILLER_101_24 ();
 sg13g2_fill_8 FILLER_101_32 ();
 sg13g2_fill_8 FILLER_101_40 ();
 sg13g2_fill_4 FILLER_101_48 ();
 sg13g2_fill_2 FILLER_101_52 ();
 sg13g2_fill_8 FILLER_101_90 ();
 sg13g2_fill_8 FILLER_101_98 ();
 sg13g2_fill_4 FILLER_101_106 ();
 sg13g2_fill_2 FILLER_101_110 ();
 sg13g2_fill_1 FILLER_101_112 ();
 sg13g2_fill_8 FILLER_101_123 ();
 sg13g2_fill_4 FILLER_101_139 ();
 sg13g2_fill_1 FILLER_101_143 ();
 sg13g2_fill_1 FILLER_101_170 ();
 sg13g2_fill_8 FILLER_101_207 ();
 sg13g2_fill_8 FILLER_101_215 ();
 sg13g2_fill_1 FILLER_101_223 ();
 sg13g2_fill_8 FILLER_101_232 ();
 sg13g2_fill_8 FILLER_101_240 ();
 sg13g2_fill_8 FILLER_101_248 ();
 sg13g2_fill_8 FILLER_101_256 ();
 sg13g2_fill_8 FILLER_101_264 ();
 sg13g2_fill_4 FILLER_101_308 ();
 sg13g2_fill_2 FILLER_101_312 ();
 sg13g2_fill_8 FILLER_101_339 ();
 sg13g2_fill_8 FILLER_101_347 ();
 sg13g2_fill_1 FILLER_101_355 ();
 sg13g2_fill_2 FILLER_101_396 ();
 sg13g2_fill_1 FILLER_101_398 ();
 sg13g2_fill_4 FILLER_101_460 ();
 sg13g2_fill_1 FILLER_101_464 ();
 sg13g2_fill_4 FILLER_101_468 ();
 sg13g2_fill_2 FILLER_101_472 ();
 sg13g2_fill_1 FILLER_101_474 ();
 sg13g2_fill_8 FILLER_101_517 ();
 sg13g2_fill_8 FILLER_101_588 ();
 sg13g2_fill_8 FILLER_101_602 ();
 sg13g2_fill_8 FILLER_101_610 ();
 sg13g2_fill_1 FILLER_101_618 ();
 sg13g2_fill_8 FILLER_101_647 ();
 sg13g2_fill_8 FILLER_101_666 ();
 sg13g2_fill_1 FILLER_101_674 ();
 sg13g2_fill_4 FILLER_101_711 ();
 sg13g2_fill_8 FILLER_101_751 ();
 sg13g2_fill_2 FILLER_101_759 ();
 sg13g2_fill_1 FILLER_101_761 ();
 sg13g2_fill_2 FILLER_101_768 ();
 sg13g2_fill_2 FILLER_101_779 ();
 sg13g2_fill_1 FILLER_101_781 ();
 sg13g2_fill_1 FILLER_101_791 ();
 sg13g2_fill_2 FILLER_101_801 ();
 sg13g2_fill_1 FILLER_101_803 ();
 sg13g2_fill_2 FILLER_101_855 ();
 sg13g2_fill_1 FILLER_101_857 ();
 sg13g2_fill_2 FILLER_101_871 ();
 sg13g2_fill_1 FILLER_101_873 ();
 sg13g2_fill_8 FILLER_101_885 ();
 sg13g2_fill_4 FILLER_101_893 ();
 sg13g2_fill_1 FILLER_101_897 ();
 sg13g2_fill_8 FILLER_101_919 ();
 sg13g2_fill_8 FILLER_101_927 ();
 sg13g2_fill_4 FILLER_101_935 ();
 sg13g2_fill_2 FILLER_101_943 ();
 sg13g2_fill_1 FILLER_101_945 ();
 sg13g2_fill_8 FILLER_101_950 ();
 sg13g2_fill_4 FILLER_101_958 ();
 sg13g2_fill_2 FILLER_101_962 ();
 sg13g2_fill_1 FILLER_101_964 ();
 sg13g2_fill_8 FILLER_101_970 ();
 sg13g2_fill_8 FILLER_101_978 ();
 sg13g2_fill_8 FILLER_101_986 ();
 sg13g2_fill_8 FILLER_101_994 ();
 sg13g2_fill_8 FILLER_101_1011 ();
 sg13g2_fill_4 FILLER_101_1019 ();
 sg13g2_fill_2 FILLER_101_1049 ();
 sg13g2_fill_4 FILLER_101_1056 ();
 sg13g2_fill_2 FILLER_101_1065 ();
 sg13g2_fill_4 FILLER_101_1090 ();
 sg13g2_fill_2 FILLER_101_1112 ();
 sg13g2_fill_1 FILLER_101_1119 ();
 sg13g2_fill_8 FILLER_101_1134 ();
 sg13g2_fill_8 FILLER_101_1142 ();
 sg13g2_fill_4 FILLER_101_1150 ();
 sg13g2_fill_8 FILLER_101_1159 ();
 sg13g2_fill_1 FILLER_101_1167 ();
 sg13g2_fill_8 FILLER_101_1176 ();
 sg13g2_fill_8 FILLER_101_1184 ();
 sg13g2_fill_1 FILLER_101_1197 ();
 sg13g2_fill_4 FILLER_101_1208 ();
 sg13g2_fill_1 FILLER_101_1212 ();
 sg13g2_fill_8 FILLER_101_1242 ();
 sg13g2_fill_2 FILLER_101_1250 ();
 sg13g2_fill_1 FILLER_101_1252 ();
 sg13g2_fill_8 FILLER_101_1256 ();
 sg13g2_fill_4 FILLER_101_1264 ();
 sg13g2_fill_2 FILLER_101_1268 ();
 sg13g2_fill_4 FILLER_101_1283 ();
 sg13g2_fill_2 FILLER_101_1287 ();
 sg13g2_fill_1 FILLER_101_1289 ();
 sg13g2_fill_2 FILLER_101_1295 ();
 sg13g2_fill_2 FILLER_101_1306 ();
 sg13g2_fill_1 FILLER_101_1308 ();
 sg13g2_fill_1 FILLER_101_1316 ();
 sg13g2_fill_8 FILLER_101_1329 ();
 sg13g2_fill_8 FILLER_101_1358 ();
 sg13g2_fill_2 FILLER_101_1366 ();
 sg13g2_fill_8 FILLER_101_1384 ();
 sg13g2_fill_8 FILLER_101_1392 ();
 sg13g2_fill_8 FILLER_101_1400 ();
 sg13g2_fill_4 FILLER_101_1408 ();
 sg13g2_fill_2 FILLER_101_1412 ();
 sg13g2_fill_4 FILLER_101_1419 ();
 sg13g2_fill_2 FILLER_101_1423 ();
 sg13g2_fill_1 FILLER_101_1425 ();
 sg13g2_fill_8 FILLER_101_1451 ();
 sg13g2_fill_1 FILLER_101_1459 ();
 sg13g2_fill_1 FILLER_101_1472 ();
 sg13g2_fill_8 FILLER_101_1477 ();
 sg13g2_fill_8 FILLER_101_1485 ();
 sg13g2_fill_8 FILLER_101_1493 ();
 sg13g2_fill_2 FILLER_101_1501 ();
 sg13g2_fill_1 FILLER_101_1503 ();
 sg13g2_fill_8 FILLER_101_1518 ();
 sg13g2_fill_2 FILLER_101_1526 ();
 sg13g2_fill_2 FILLER_101_1590 ();
 sg13g2_fill_8 FILLER_102_0 ();
 sg13g2_fill_8 FILLER_102_8 ();
 sg13g2_fill_8 FILLER_102_16 ();
 sg13g2_fill_8 FILLER_102_24 ();
 sg13g2_fill_8 FILLER_102_32 ();
 sg13g2_fill_8 FILLER_102_40 ();
 sg13g2_fill_8 FILLER_102_48 ();
 sg13g2_fill_8 FILLER_102_56 ();
 sg13g2_fill_8 FILLER_102_90 ();
 sg13g2_fill_1 FILLER_102_98 ();
 sg13g2_fill_8 FILLER_102_109 ();
 sg13g2_fill_1 FILLER_102_117 ();
 sg13g2_fill_8 FILLER_102_140 ();
 sg13g2_fill_8 FILLER_102_148 ();
 sg13g2_fill_2 FILLER_102_166 ();
 sg13g2_fill_1 FILLER_102_168 ();
 sg13g2_fill_1 FILLER_102_172 ();
 sg13g2_fill_8 FILLER_102_199 ();
 sg13g2_fill_8 FILLER_102_207 ();
 sg13g2_fill_8 FILLER_102_215 ();
 sg13g2_fill_1 FILLER_102_223 ();
 sg13g2_fill_8 FILLER_102_229 ();
 sg13g2_fill_8 FILLER_102_250 ();
 sg13g2_fill_2 FILLER_102_258 ();
 sg13g2_fill_4 FILLER_102_270 ();
 sg13g2_fill_2 FILLER_102_274 ();
 sg13g2_fill_1 FILLER_102_276 ();
 sg13g2_fill_8 FILLER_102_287 ();
 sg13g2_fill_8 FILLER_102_295 ();
 sg13g2_fill_8 FILLER_102_303 ();
 sg13g2_fill_1 FILLER_102_311 ();
 sg13g2_fill_4 FILLER_102_317 ();
 sg13g2_fill_1 FILLER_102_321 ();
 sg13g2_fill_8 FILLER_102_330 ();
 sg13g2_fill_8 FILLER_102_338 ();
 sg13g2_fill_2 FILLER_102_374 ();
 sg13g2_fill_4 FILLER_102_386 ();
 sg13g2_fill_4 FILLER_102_403 ();
 sg13g2_fill_1 FILLER_102_407 ();
 sg13g2_fill_4 FILLER_102_444 ();
 sg13g2_fill_1 FILLER_102_448 ();
 sg13g2_fill_4 FILLER_102_507 ();
 sg13g2_fill_2 FILLER_102_511 ();
 sg13g2_fill_1 FILLER_102_513 ();
 sg13g2_fill_8 FILLER_102_524 ();
 sg13g2_fill_8 FILLER_102_532 ();
 sg13g2_fill_8 FILLER_102_540 ();
 sg13g2_fill_8 FILLER_102_548 ();
 sg13g2_fill_2 FILLER_102_556 ();
 sg13g2_fill_1 FILLER_102_558 ();
 sg13g2_fill_8 FILLER_102_569 ();
 sg13g2_fill_1 FILLER_102_577 ();
 sg13g2_fill_2 FILLER_102_612 ();
 sg13g2_fill_1 FILLER_102_614 ();
 sg13g2_fill_8 FILLER_102_641 ();
 sg13g2_fill_8 FILLER_102_649 ();
 sg13g2_fill_1 FILLER_102_657 ();
 sg13g2_fill_4 FILLER_102_668 ();
 sg13g2_fill_2 FILLER_102_672 ();
 sg13g2_fill_4 FILLER_102_684 ();
 sg13g2_fill_1 FILLER_102_688 ();
 sg13g2_fill_4 FILLER_102_699 ();
 sg13g2_fill_2 FILLER_102_703 ();
 sg13g2_fill_1 FILLER_102_705 ();
 sg13g2_fill_4 FILLER_102_711 ();
 sg13g2_fill_1 FILLER_102_725 ();
 sg13g2_fill_1 FILLER_102_752 ();
 sg13g2_fill_1 FILLER_102_799 ();
 sg13g2_fill_2 FILLER_102_815 ();
 sg13g2_fill_2 FILLER_102_842 ();
 sg13g2_fill_1 FILLER_102_844 ();
 sg13g2_fill_4 FILLER_102_853 ();
 sg13g2_fill_2 FILLER_102_857 ();
 sg13g2_fill_8 FILLER_102_863 ();
 sg13g2_fill_8 FILLER_102_871 ();
 sg13g2_fill_8 FILLER_102_879 ();
 sg13g2_fill_2 FILLER_102_887 ();
 sg13g2_fill_2 FILLER_102_904 ();
 sg13g2_fill_4 FILLER_102_968 ();
 sg13g2_fill_2 FILLER_102_972 ();
 sg13g2_fill_2 FILLER_102_982 ();
 sg13g2_fill_1 FILLER_102_998 ();
 sg13g2_fill_1 FILLER_102_1022 ();
 sg13g2_fill_1 FILLER_102_1047 ();
 sg13g2_fill_8 FILLER_102_1056 ();
 sg13g2_fill_1 FILLER_102_1064 ();
 sg13g2_fill_4 FILLER_102_1095 ();
 sg13g2_fill_2 FILLER_102_1099 ();
 sg13g2_fill_8 FILLER_102_1106 ();
 sg13g2_fill_4 FILLER_102_1114 ();
 sg13g2_fill_1 FILLER_102_1118 ();
 sg13g2_fill_4 FILLER_102_1124 ();
 sg13g2_fill_2 FILLER_102_1128 ();
 sg13g2_fill_1 FILLER_102_1130 ();
 sg13g2_fill_4 FILLER_102_1138 ();
 sg13g2_fill_8 FILLER_102_1146 ();
 sg13g2_fill_8 FILLER_102_1159 ();
 sg13g2_fill_2 FILLER_102_1167 ();
 sg13g2_fill_2 FILLER_102_1174 ();
 sg13g2_fill_2 FILLER_102_1181 ();
 sg13g2_fill_1 FILLER_102_1203 ();
 sg13g2_fill_4 FILLER_102_1210 ();
 sg13g2_fill_2 FILLER_102_1214 ();
 sg13g2_fill_1 FILLER_102_1216 ();
 sg13g2_fill_8 FILLER_102_1235 ();
 sg13g2_fill_8 FILLER_102_1250 ();
 sg13g2_fill_2 FILLER_102_1258 ();
 sg13g2_fill_1 FILLER_102_1260 ();
 sg13g2_fill_4 FILLER_102_1265 ();
 sg13g2_fill_1 FILLER_102_1269 ();
 sg13g2_fill_8 FILLER_102_1279 ();
 sg13g2_fill_1 FILLER_102_1287 ();
 sg13g2_fill_8 FILLER_102_1291 ();
 sg13g2_fill_4 FILLER_102_1299 ();
 sg13g2_fill_8 FILLER_102_1309 ();
 sg13g2_fill_8 FILLER_102_1317 ();
 sg13g2_fill_8 FILLER_102_1325 ();
 sg13g2_fill_8 FILLER_102_1333 ();
 sg13g2_fill_2 FILLER_102_1341 ();
 sg13g2_fill_8 FILLER_102_1347 ();
 sg13g2_fill_8 FILLER_102_1355 ();
 sg13g2_fill_8 FILLER_102_1363 ();
 sg13g2_fill_1 FILLER_102_1371 ();
 sg13g2_fill_1 FILLER_102_1388 ();
 sg13g2_fill_2 FILLER_102_1394 ();
 sg13g2_fill_2 FILLER_102_1404 ();
 sg13g2_fill_1 FILLER_102_1406 ();
 sg13g2_fill_8 FILLER_102_1425 ();
 sg13g2_fill_1 FILLER_102_1433 ();
 sg13g2_fill_2 FILLER_102_1442 ();
 sg13g2_fill_8 FILLER_102_1454 ();
 sg13g2_fill_2 FILLER_102_1462 ();
 sg13g2_fill_1 FILLER_102_1464 ();
 sg13g2_fill_8 FILLER_102_1478 ();
 sg13g2_fill_2 FILLER_102_1486 ();
 sg13g2_fill_1 FILLER_102_1488 ();
 sg13g2_fill_4 FILLER_102_1497 ();
 sg13g2_fill_8 FILLER_102_1527 ();
 sg13g2_fill_8 FILLER_102_1535 ();
 sg13g2_fill_2 FILLER_102_1557 ();
 sg13g2_fill_2 FILLER_102_1572 ();
 sg13g2_fill_8 FILLER_102_1582 ();
 sg13g2_fill_2 FILLER_102_1590 ();
 sg13g2_fill_8 FILLER_103_0 ();
 sg13g2_fill_8 FILLER_103_8 ();
 sg13g2_fill_8 FILLER_103_16 ();
 sg13g2_fill_8 FILLER_103_24 ();
 sg13g2_fill_8 FILLER_103_32 ();
 sg13g2_fill_8 FILLER_103_40 ();
 sg13g2_fill_8 FILLER_103_48 ();
 sg13g2_fill_8 FILLER_103_56 ();
 sg13g2_fill_8 FILLER_103_64 ();
 sg13g2_fill_8 FILLER_103_72 ();
 sg13g2_fill_4 FILLER_103_80 ();
 sg13g2_fill_1 FILLER_103_84 ();
 sg13g2_fill_1 FILLER_103_111 ();
 sg13g2_fill_1 FILLER_103_168 ();
 sg13g2_fill_8 FILLER_103_194 ();
 sg13g2_fill_8 FILLER_103_202 ();
 sg13g2_fill_4 FILLER_103_210 ();
 sg13g2_fill_2 FILLER_103_214 ();
 sg13g2_fill_8 FILLER_103_266 ();
 sg13g2_fill_1 FILLER_103_310 ();
 sg13g2_fill_4 FILLER_103_355 ();
 sg13g2_fill_2 FILLER_103_359 ();
 sg13g2_fill_1 FILLER_103_361 ();
 sg13g2_fill_8 FILLER_103_411 ();
 sg13g2_fill_8 FILLER_103_419 ();
 sg13g2_fill_8 FILLER_103_427 ();
 sg13g2_fill_8 FILLER_103_435 ();
 sg13g2_fill_8 FILLER_103_443 ();
 sg13g2_fill_4 FILLER_103_451 ();
 sg13g2_fill_8 FILLER_103_463 ();
 sg13g2_fill_2 FILLER_103_471 ();
 sg13g2_fill_1 FILLER_103_473 ();
 sg13g2_fill_8 FILLER_103_496 ();
 sg13g2_fill_4 FILLER_103_504 ();
 sg13g2_fill_2 FILLER_103_508 ();
 sg13g2_fill_8 FILLER_103_526 ();
 sg13g2_fill_8 FILLER_103_534 ();
 sg13g2_fill_8 FILLER_103_542 ();
 sg13g2_fill_8 FILLER_103_550 ();
 sg13g2_fill_1 FILLER_103_568 ();
 sg13g2_fill_8 FILLER_103_577 ();
 sg13g2_fill_8 FILLER_103_585 ();
 sg13g2_fill_4 FILLER_103_593 ();
 sg13g2_fill_2 FILLER_103_597 ();
 sg13g2_fill_8 FILLER_103_619 ();
 sg13g2_fill_2 FILLER_103_627 ();
 sg13g2_fill_1 FILLER_103_629 ();
 sg13g2_fill_4 FILLER_103_656 ();
 sg13g2_fill_1 FILLER_103_660 ();
 sg13g2_fill_4 FILLER_103_687 ();
 sg13g2_fill_2 FILLER_103_691 ();
 sg13g2_fill_8 FILLER_103_711 ();
 sg13g2_fill_8 FILLER_103_719 ();
 sg13g2_fill_8 FILLER_103_727 ();
 sg13g2_fill_8 FILLER_103_735 ();
 sg13g2_fill_8 FILLER_103_743 ();
 sg13g2_fill_4 FILLER_103_751 ();
 sg13g2_fill_2 FILLER_103_755 ();
 sg13g2_fill_8 FILLER_103_792 ();
 sg13g2_fill_2 FILLER_103_812 ();
 sg13g2_fill_2 FILLER_103_820 ();
 sg13g2_fill_4 FILLER_103_847 ();
 sg13g2_fill_1 FILLER_103_851 ();
 sg13g2_fill_2 FILLER_103_891 ();
 sg13g2_fill_1 FILLER_103_910 ();
 sg13g2_fill_4 FILLER_103_965 ();
 sg13g2_fill_1 FILLER_103_994 ();
 sg13g2_fill_4 FILLER_103_1002 ();
 sg13g2_fill_2 FILLER_103_1006 ();
 sg13g2_fill_2 FILLER_103_1013 ();
 sg13g2_fill_1 FILLER_103_1035 ();
 sg13g2_fill_2 FILLER_103_1049 ();
 sg13g2_fill_8 FILLER_103_1056 ();
 sg13g2_fill_8 FILLER_103_1064 ();
 sg13g2_fill_2 FILLER_103_1072 ();
 sg13g2_fill_1 FILLER_103_1074 ();
 sg13g2_fill_8 FILLER_103_1085 ();
 sg13g2_fill_8 FILLER_103_1093 ();
 sg13g2_fill_2 FILLER_103_1101 ();
 sg13g2_fill_1 FILLER_103_1103 ();
 sg13g2_fill_2 FILLER_103_1109 ();
 sg13g2_fill_1 FILLER_103_1111 ();
 sg13g2_fill_2 FILLER_103_1122 ();
 sg13g2_fill_1 FILLER_103_1124 ();
 sg13g2_fill_2 FILLER_103_1147 ();
 sg13g2_fill_1 FILLER_103_1171 ();
 sg13g2_fill_2 FILLER_103_1182 ();
 sg13g2_fill_8 FILLER_103_1207 ();
 sg13g2_fill_4 FILLER_103_1215 ();
 sg13g2_fill_2 FILLER_103_1219 ();
 sg13g2_fill_1 FILLER_103_1221 ();
 sg13g2_fill_8 FILLER_103_1226 ();
 sg13g2_fill_8 FILLER_103_1234 ();
 sg13g2_fill_2 FILLER_103_1242 ();
 sg13g2_fill_4 FILLER_103_1275 ();
 sg13g2_fill_2 FILLER_103_1279 ();
 sg13g2_fill_8 FILLER_103_1302 ();
 sg13g2_fill_4 FILLER_103_1310 ();
 sg13g2_fill_2 FILLER_103_1314 ();
 sg13g2_fill_1 FILLER_103_1316 ();
 sg13g2_fill_4 FILLER_103_1322 ();
 sg13g2_fill_2 FILLER_103_1326 ();
 sg13g2_fill_1 FILLER_103_1328 ();
 sg13g2_fill_4 FILLER_103_1371 ();
 sg13g2_fill_2 FILLER_103_1375 ();
 sg13g2_fill_1 FILLER_103_1377 ();
 sg13g2_fill_2 FILLER_103_1385 ();
 sg13g2_fill_1 FILLER_103_1387 ();
 sg13g2_fill_8 FILLER_103_1400 ();
 sg13g2_fill_1 FILLER_103_1448 ();
 sg13g2_fill_2 FILLER_103_1475 ();
 sg13g2_fill_2 FILLER_103_1527 ();
 sg13g2_fill_1 FILLER_103_1529 ();
 sg13g2_fill_4 FILLER_103_1534 ();
 sg13g2_fill_8 FILLER_103_1544 ();
 sg13g2_fill_4 FILLER_103_1561 ();
 sg13g2_fill_1 FILLER_103_1565 ();
 sg13g2_fill_8 FILLER_104_0 ();
 sg13g2_fill_8 FILLER_104_8 ();
 sg13g2_fill_8 FILLER_104_16 ();
 sg13g2_fill_8 FILLER_104_24 ();
 sg13g2_fill_8 FILLER_104_32 ();
 sg13g2_fill_8 FILLER_104_40 ();
 sg13g2_fill_8 FILLER_104_48 ();
 sg13g2_fill_8 FILLER_104_56 ();
 sg13g2_fill_8 FILLER_104_64 ();
 sg13g2_fill_8 FILLER_104_72 ();
 sg13g2_fill_8 FILLER_104_80 ();
 sg13g2_fill_8 FILLER_104_88 ();
 sg13g2_fill_8 FILLER_104_96 ();
 sg13g2_fill_8 FILLER_104_104 ();
 sg13g2_fill_8 FILLER_104_112 ();
 sg13g2_fill_8 FILLER_104_120 ();
 sg13g2_fill_1 FILLER_104_128 ();
 sg13g2_fill_8 FILLER_104_139 ();
 sg13g2_fill_8 FILLER_104_147 ();
 sg13g2_fill_8 FILLER_104_155 ();
 sg13g2_fill_4 FILLER_104_163 ();
 sg13g2_fill_2 FILLER_104_167 ();
 sg13g2_fill_2 FILLER_104_174 ();
 sg13g2_fill_1 FILLER_104_176 ();
 sg13g2_fill_2 FILLER_104_195 ();
 sg13g2_fill_1 FILLER_104_197 ();
 sg13g2_fill_4 FILLER_104_219 ();
 sg13g2_fill_4 FILLER_104_244 ();
 sg13g2_fill_2 FILLER_104_248 ();
 sg13g2_fill_1 FILLER_104_250 ();
 sg13g2_fill_8 FILLER_104_259 ();
 sg13g2_fill_8 FILLER_104_293 ();
 sg13g2_fill_1 FILLER_104_301 ();
 sg13g2_fill_2 FILLER_104_307 ();
 sg13g2_fill_2 FILLER_104_324 ();
 sg13g2_fill_1 FILLER_104_326 ();
 sg13g2_fill_4 FILLER_104_358 ();
 sg13g2_fill_1 FILLER_104_372 ();
 sg13g2_fill_8 FILLER_104_383 ();
 sg13g2_fill_8 FILLER_104_391 ();
 sg13g2_fill_8 FILLER_104_399 ();
 sg13g2_fill_1 FILLER_104_407 ();
 sg13g2_fill_8 FILLER_104_418 ();
 sg13g2_fill_8 FILLER_104_426 ();
 sg13g2_fill_8 FILLER_104_434 ();
 sg13g2_fill_4 FILLER_104_442 ();
 sg13g2_fill_4 FILLER_104_467 ();
 sg13g2_fill_2 FILLER_104_471 ();
 sg13g2_fill_1 FILLER_104_473 ();
 sg13g2_fill_2 FILLER_104_502 ();
 sg13g2_fill_1 FILLER_104_504 ();
 sg13g2_fill_1 FILLER_104_510 ();
 sg13g2_fill_4 FILLER_104_521 ();
 sg13g2_fill_4 FILLER_104_587 ();
 sg13g2_fill_8 FILLER_104_595 ();
 sg13g2_fill_8 FILLER_104_603 ();
 sg13g2_fill_8 FILLER_104_615 ();
 sg13g2_fill_4 FILLER_104_623 ();
 sg13g2_fill_1 FILLER_104_627 ();
 sg13g2_fill_8 FILLER_104_638 ();
 sg13g2_fill_8 FILLER_104_646 ();
 sg13g2_fill_1 FILLER_104_654 ();
 sg13g2_fill_8 FILLER_104_665 ();
 sg13g2_fill_8 FILLER_104_673 ();
 sg13g2_fill_4 FILLER_104_681 ();
 sg13g2_fill_1 FILLER_104_685 ();
 sg13g2_fill_8 FILLER_104_696 ();
 sg13g2_fill_8 FILLER_104_704 ();
 sg13g2_fill_8 FILLER_104_738 ();
 sg13g2_fill_4 FILLER_104_746 ();
 sg13g2_fill_1 FILLER_104_750 ();
 sg13g2_fill_4 FILLER_104_767 ();
 sg13g2_fill_2 FILLER_104_804 ();
 sg13g2_fill_1 FILLER_104_806 ();
 sg13g2_fill_1 FILLER_104_828 ();
 sg13g2_fill_2 FILLER_104_834 ();
 sg13g2_fill_1 FILLER_104_836 ();
 sg13g2_fill_2 FILLER_104_878 ();
 sg13g2_fill_1 FILLER_104_880 ();
 sg13g2_fill_1 FILLER_104_907 ();
 sg13g2_fill_4 FILLER_104_944 ();
 sg13g2_fill_2 FILLER_104_948 ();
 sg13g2_fill_8 FILLER_104_958 ();
 sg13g2_fill_4 FILLER_104_966 ();
 sg13g2_fill_2 FILLER_104_970 ();
 sg13g2_fill_1 FILLER_104_972 ();
 sg13g2_fill_4 FILLER_104_982 ();
 sg13g2_fill_1 FILLER_104_986 ();
 sg13g2_fill_8 FILLER_104_992 ();
 sg13g2_fill_8 FILLER_104_1000 ();
 sg13g2_fill_8 FILLER_104_1008 ();
 sg13g2_fill_8 FILLER_104_1016 ();
 sg13g2_fill_2 FILLER_104_1024 ();
 sg13g2_fill_1 FILLER_104_1026 ();
 sg13g2_fill_4 FILLER_104_1031 ();
 sg13g2_fill_1 FILLER_104_1035 ();
 sg13g2_fill_2 FILLER_104_1042 ();
 sg13g2_fill_2 FILLER_104_1048 ();
 sg13g2_fill_1 FILLER_104_1050 ();
 sg13g2_fill_8 FILLER_104_1057 ();
 sg13g2_fill_4 FILLER_104_1065 ();
 sg13g2_fill_2 FILLER_104_1069 ();
 sg13g2_fill_2 FILLER_104_1076 ();
 sg13g2_fill_8 FILLER_104_1081 ();
 sg13g2_fill_4 FILLER_104_1089 ();
 sg13g2_fill_1 FILLER_104_1093 ();
 sg13g2_fill_2 FILLER_104_1102 ();
 sg13g2_fill_1 FILLER_104_1104 ();
 sg13g2_fill_1 FILLER_104_1110 ();
 sg13g2_fill_8 FILLER_104_1121 ();
 sg13g2_fill_2 FILLER_104_1129 ();
 sg13g2_fill_4 FILLER_104_1134 ();
 sg13g2_fill_1 FILLER_104_1138 ();
 sg13g2_fill_1 FILLER_104_1144 ();
 sg13g2_fill_2 FILLER_104_1158 ();
 sg13g2_fill_1 FILLER_104_1160 ();
 sg13g2_fill_8 FILLER_104_1177 ();
 sg13g2_fill_4 FILLER_104_1185 ();
 sg13g2_fill_2 FILLER_104_1189 ();
 sg13g2_fill_8 FILLER_104_1196 ();
 sg13g2_fill_8 FILLER_104_1204 ();
 sg13g2_fill_4 FILLER_104_1212 ();
 sg13g2_fill_2 FILLER_104_1216 ();
 sg13g2_fill_4 FILLER_104_1227 ();
 sg13g2_fill_2 FILLER_104_1231 ();
 sg13g2_fill_1 FILLER_104_1233 ();
 sg13g2_fill_4 FILLER_104_1241 ();
 sg13g2_fill_2 FILLER_104_1245 ();
 sg13g2_fill_1 FILLER_104_1247 ();
 sg13g2_fill_2 FILLER_104_1263 ();
 sg13g2_fill_1 FILLER_104_1270 ();
 sg13g2_fill_1 FILLER_104_1280 ();
 sg13g2_fill_8 FILLER_104_1303 ();
 sg13g2_fill_2 FILLER_104_1311 ();
 sg13g2_fill_4 FILLER_104_1333 ();
 sg13g2_fill_1 FILLER_104_1337 ();
 sg13g2_fill_2 FILLER_104_1343 ();
 sg13g2_fill_1 FILLER_104_1345 ();
 sg13g2_fill_8 FILLER_104_1402 ();
 sg13g2_fill_2 FILLER_104_1410 ();
 sg13g2_fill_4 FILLER_104_1417 ();
 sg13g2_fill_2 FILLER_104_1421 ();
 sg13g2_fill_8 FILLER_104_1427 ();
 sg13g2_fill_4 FILLER_104_1435 ();
 sg13g2_fill_2 FILLER_104_1439 ();
 sg13g2_fill_2 FILLER_104_1446 ();
 sg13g2_fill_8 FILLER_104_1457 ();
 sg13g2_fill_8 FILLER_104_1476 ();
 sg13g2_fill_4 FILLER_104_1484 ();
 sg13g2_fill_2 FILLER_104_1488 ();
 sg13g2_fill_8 FILLER_104_1499 ();
 sg13g2_fill_1 FILLER_104_1507 ();
 sg13g2_fill_2 FILLER_104_1512 ();
 sg13g2_fill_4 FILLER_104_1540 ();
 sg13g2_fill_4 FILLER_104_1570 ();
 sg13g2_fill_1 FILLER_104_1574 ();
 sg13g2_fill_8 FILLER_104_1580 ();
 sg13g2_fill_4 FILLER_104_1588 ();
 sg13g2_fill_8 FILLER_105_0 ();
 sg13g2_fill_8 FILLER_105_8 ();
 sg13g2_fill_8 FILLER_105_16 ();
 sg13g2_fill_8 FILLER_105_24 ();
 sg13g2_fill_8 FILLER_105_32 ();
 sg13g2_fill_8 FILLER_105_40 ();
 sg13g2_fill_8 FILLER_105_48 ();
 sg13g2_fill_8 FILLER_105_56 ();
 sg13g2_fill_8 FILLER_105_64 ();
 sg13g2_fill_8 FILLER_105_72 ();
 sg13g2_fill_8 FILLER_105_80 ();
 sg13g2_fill_8 FILLER_105_88 ();
 sg13g2_fill_8 FILLER_105_96 ();
 sg13g2_fill_2 FILLER_105_104 ();
 sg13g2_fill_1 FILLER_105_126 ();
 sg13g2_fill_8 FILLER_105_132 ();
 sg13g2_fill_1 FILLER_105_140 ();
 sg13g2_fill_4 FILLER_105_149 ();
 sg13g2_fill_1 FILLER_105_153 ();
 sg13g2_fill_4 FILLER_105_170 ();
 sg13g2_fill_1 FILLER_105_174 ();
 sg13g2_fill_8 FILLER_105_285 ();
 sg13g2_fill_8 FILLER_105_330 ();
 sg13g2_fill_4 FILLER_105_338 ();
 sg13g2_fill_2 FILLER_105_342 ();
 sg13g2_fill_1 FILLER_105_344 ();
 sg13g2_fill_4 FILLER_105_371 ();
 sg13g2_fill_2 FILLER_105_375 ();
 sg13g2_fill_1 FILLER_105_377 ();
 sg13g2_fill_1 FILLER_105_404 ();
 sg13g2_fill_2 FILLER_105_439 ();
 sg13g2_fill_1 FILLER_105_441 ();
 sg13g2_fill_1 FILLER_105_452 ();
 sg13g2_fill_2 FILLER_105_460 ();
 sg13g2_fill_1 FILLER_105_462 ();
 sg13g2_fill_1 FILLER_105_468 ();
 sg13g2_fill_2 FILLER_105_480 ();
 sg13g2_fill_4 FILLER_105_487 ();
 sg13g2_fill_1 FILLER_105_491 ();
 sg13g2_fill_4 FILLER_105_526 ();
 sg13g2_fill_4 FILLER_105_546 ();
 sg13g2_fill_4 FILLER_105_558 ();
 sg13g2_fill_2 FILLER_105_562 ();
 sg13g2_fill_1 FILLER_105_572 ();
 sg13g2_fill_8 FILLER_105_618 ();
 sg13g2_fill_8 FILLER_105_626 ();
 sg13g2_fill_2 FILLER_105_634 ();
 sg13g2_fill_2 FILLER_105_660 ();
 sg13g2_fill_1 FILLER_105_662 ();
 sg13g2_fill_4 FILLER_105_668 ();
 sg13g2_fill_2 FILLER_105_672 ();
 sg13g2_fill_4 FILLER_105_682 ();
 sg13g2_fill_1 FILLER_105_686 ();
 sg13g2_fill_4 FILLER_105_717 ();
 sg13g2_fill_4 FILLER_105_747 ();
 sg13g2_fill_2 FILLER_105_751 ();
 sg13g2_fill_1 FILLER_105_753 ();
 sg13g2_fill_8 FILLER_105_767 ();
 sg13g2_fill_8 FILLER_105_775 ();
 sg13g2_fill_8 FILLER_105_787 ();
 sg13g2_fill_8 FILLER_105_795 ();
 sg13g2_fill_8 FILLER_105_803 ();
 sg13g2_fill_8 FILLER_105_811 ();
 sg13g2_fill_4 FILLER_105_819 ();
 sg13g2_fill_1 FILLER_105_823 ();
 sg13g2_fill_8 FILLER_105_827 ();
 sg13g2_fill_8 FILLER_105_835 ();
 sg13g2_fill_8 FILLER_105_843 ();
 sg13g2_fill_1 FILLER_105_851 ();
 sg13g2_fill_2 FILLER_105_877 ();
 sg13g2_fill_8 FILLER_105_884 ();
 sg13g2_fill_4 FILLER_105_892 ();
 sg13g2_fill_2 FILLER_105_896 ();
 sg13g2_fill_1 FILLER_105_898 ();
 sg13g2_fill_2 FILLER_105_912 ();
 sg13g2_fill_8 FILLER_105_924 ();
 sg13g2_fill_8 FILLER_105_932 ();
 sg13g2_fill_8 FILLER_105_940 ();
 sg13g2_fill_2 FILLER_105_948 ();
 sg13g2_fill_1 FILLER_105_950 ();
 sg13g2_fill_8 FILLER_105_959 ();
 sg13g2_fill_4 FILLER_105_967 ();
 sg13g2_fill_1 FILLER_105_971 ();
 sg13g2_fill_8 FILLER_105_982 ();
 sg13g2_fill_4 FILLER_105_990 ();
 sg13g2_fill_2 FILLER_105_994 ();
 sg13g2_fill_4 FILLER_105_1016 ();
 sg13g2_fill_2 FILLER_105_1020 ();
 sg13g2_fill_1 FILLER_105_1047 ();
 sg13g2_fill_2 FILLER_105_1054 ();
 sg13g2_fill_1 FILLER_105_1056 ();
 sg13g2_fill_1 FILLER_105_1063 ();
 sg13g2_fill_2 FILLER_105_1082 ();
 sg13g2_fill_1 FILLER_105_1084 ();
 sg13g2_fill_4 FILLER_105_1105 ();
 sg13g2_fill_1 FILLER_105_1109 ();
 sg13g2_fill_8 FILLER_105_1114 ();
 sg13g2_fill_4 FILLER_105_1122 ();
 sg13g2_fill_2 FILLER_105_1126 ();
 sg13g2_fill_8 FILLER_105_1133 ();
 sg13g2_fill_4 FILLER_105_1141 ();
 sg13g2_fill_1 FILLER_105_1145 ();
 sg13g2_fill_1 FILLER_105_1162 ();
 sg13g2_fill_8 FILLER_105_1167 ();
 sg13g2_fill_2 FILLER_105_1175 ();
 sg13g2_fill_1 FILLER_105_1184 ();
 sg13g2_fill_2 FILLER_105_1205 ();
 sg13g2_fill_1 FILLER_105_1207 ();
 sg13g2_fill_1 FILLER_105_1236 ();
 sg13g2_fill_8 FILLER_105_1242 ();
 sg13g2_fill_4 FILLER_105_1250 ();
 sg13g2_fill_2 FILLER_105_1254 ();
 sg13g2_fill_1 FILLER_105_1256 ();
 sg13g2_fill_1 FILLER_105_1262 ();
 sg13g2_fill_8 FILLER_105_1268 ();
 sg13g2_fill_8 FILLER_105_1276 ();
 sg13g2_fill_4 FILLER_105_1284 ();
 sg13g2_fill_2 FILLER_105_1293 ();
 sg13g2_fill_8 FILLER_105_1301 ();
 sg13g2_fill_2 FILLER_105_1309 ();
 sg13g2_fill_1 FILLER_105_1311 ();
 sg13g2_fill_8 FILLER_105_1317 ();
 sg13g2_fill_4 FILLER_105_1325 ();
 sg13g2_fill_1 FILLER_105_1329 ();
 sg13g2_fill_8 FILLER_105_1347 ();
 sg13g2_fill_1 FILLER_105_1355 ();
 sg13g2_fill_4 FILLER_105_1375 ();
 sg13g2_fill_2 FILLER_105_1379 ();
 sg13g2_fill_2 FILLER_105_1390 ();
 sg13g2_fill_1 FILLER_105_1392 ();
 sg13g2_fill_4 FILLER_105_1398 ();
 sg13g2_fill_8 FILLER_105_1417 ();
 sg13g2_fill_8 FILLER_105_1425 ();
 sg13g2_fill_8 FILLER_105_1433 ();
 sg13g2_fill_4 FILLER_105_1441 ();
 sg13g2_fill_8 FILLER_105_1467 ();
 sg13g2_fill_8 FILLER_105_1475 ();
 sg13g2_fill_8 FILLER_105_1483 ();
 sg13g2_fill_1 FILLER_105_1491 ();
 sg13g2_fill_2 FILLER_105_1507 ();
 sg13g2_fill_1 FILLER_105_1509 ();
 sg13g2_fill_2 FILLER_105_1518 ();
 sg13g2_fill_1 FILLER_105_1520 ();
 sg13g2_fill_8 FILLER_105_1524 ();
 sg13g2_fill_8 FILLER_105_1532 ();
 sg13g2_fill_8 FILLER_105_1540 ();
 sg13g2_fill_2 FILLER_105_1548 ();
 sg13g2_fill_2 FILLER_105_1564 ();
 sg13g2_fill_8 FILLER_106_0 ();
 sg13g2_fill_8 FILLER_106_8 ();
 sg13g2_fill_8 FILLER_106_16 ();
 sg13g2_fill_8 FILLER_106_24 ();
 sg13g2_fill_8 FILLER_106_32 ();
 sg13g2_fill_8 FILLER_106_40 ();
 sg13g2_fill_8 FILLER_106_48 ();
 sg13g2_fill_8 FILLER_106_56 ();
 sg13g2_fill_8 FILLER_106_64 ();
 sg13g2_fill_4 FILLER_106_72 ();
 sg13g2_fill_8 FILLER_106_110 ();
 sg13g2_fill_4 FILLER_106_134 ();
 sg13g2_fill_4 FILLER_106_148 ();
 sg13g2_fill_2 FILLER_106_152 ();
 sg13g2_fill_8 FILLER_106_167 ();
 sg13g2_fill_2 FILLER_106_175 ();
 sg13g2_fill_4 FILLER_106_187 ();
 sg13g2_fill_8 FILLER_106_201 ();
 sg13g2_fill_4 FILLER_106_209 ();
 sg13g2_fill_2 FILLER_106_213 ();
 sg13g2_fill_1 FILLER_106_215 ();
 sg13g2_fill_8 FILLER_106_250 ();
 sg13g2_fill_2 FILLER_106_258 ();
 sg13g2_fill_1 FILLER_106_260 ();
 sg13g2_fill_8 FILLER_106_271 ();
 sg13g2_fill_8 FILLER_106_279 ();
 sg13g2_fill_8 FILLER_106_287 ();
 sg13g2_fill_1 FILLER_106_295 ();
 sg13g2_fill_8 FILLER_106_306 ();
 sg13g2_fill_8 FILLER_106_314 ();
 sg13g2_fill_8 FILLER_106_322 ();
 sg13g2_fill_4 FILLER_106_330 ();
 sg13g2_fill_8 FILLER_106_345 ();
 sg13g2_fill_8 FILLER_106_353 ();
 sg13g2_fill_2 FILLER_106_361 ();
 sg13g2_fill_8 FILLER_106_373 ();
 sg13g2_fill_8 FILLER_106_381 ();
 sg13g2_fill_8 FILLER_106_409 ();
 sg13g2_fill_2 FILLER_106_417 ();
 sg13g2_fill_2 FILLER_106_469 ();
 sg13g2_fill_1 FILLER_106_481 ();
 sg13g2_fill_8 FILLER_106_487 ();
 sg13g2_fill_8 FILLER_106_495 ();
 sg13g2_fill_8 FILLER_106_503 ();
 sg13g2_fill_8 FILLER_106_511 ();
 sg13g2_fill_4 FILLER_106_519 ();
 sg13g2_fill_2 FILLER_106_523 ();
 sg13g2_fill_1 FILLER_106_525 ();
 sg13g2_fill_2 FILLER_106_536 ();
 sg13g2_fill_4 FILLER_106_544 ();
 sg13g2_fill_2 FILLER_106_548 ();
 sg13g2_fill_1 FILLER_106_550 ();
 sg13g2_fill_8 FILLER_106_587 ();
 sg13g2_fill_8 FILLER_106_595 ();
 sg13g2_fill_8 FILLER_106_603 ();
 sg13g2_fill_4 FILLER_106_611 ();
 sg13g2_fill_1 FILLER_106_615 ();
 sg13g2_fill_4 FILLER_106_642 ();
 sg13g2_fill_1 FILLER_106_678 ();
 sg13g2_fill_8 FILLER_106_699 ();
 sg13g2_fill_8 FILLER_106_707 ();
 sg13g2_fill_4 FILLER_106_715 ();
 sg13g2_fill_2 FILLER_106_719 ();
 sg13g2_fill_1 FILLER_106_721 ();
 sg13g2_fill_4 FILLER_106_748 ();
 sg13g2_fill_1 FILLER_106_752 ();
 sg13g2_fill_2 FILLER_106_756 ();
 sg13g2_fill_2 FILLER_106_766 ();
 sg13g2_fill_8 FILLER_106_801 ();
 sg13g2_fill_8 FILLER_106_809 ();
 sg13g2_fill_8 FILLER_106_817 ();
 sg13g2_fill_8 FILLER_106_825 ();
 sg13g2_fill_8 FILLER_106_833 ();
 sg13g2_fill_2 FILLER_106_841 ();
 sg13g2_fill_1 FILLER_106_843 ();
 sg13g2_fill_8 FILLER_106_888 ();
 sg13g2_fill_8 FILLER_106_900 ();
 sg13g2_fill_2 FILLER_106_908 ();
 sg13g2_fill_1 FILLER_106_910 ();
 sg13g2_fill_2 FILLER_106_968 ();
 sg13g2_fill_1 FILLER_106_1014 ();
 sg13g2_fill_1 FILLER_106_1020 ();
 sg13g2_fill_1 FILLER_106_1026 ();
 sg13g2_fill_1 FILLER_106_1035 ();
 sg13g2_fill_1 FILLER_106_1042 ();
 sg13g2_fill_8 FILLER_106_1058 ();
 sg13g2_fill_1 FILLER_106_1066 ();
 sg13g2_fill_4 FILLER_106_1077 ();
 sg13g2_fill_1 FILLER_106_1081 ();
 sg13g2_fill_4 FILLER_106_1100 ();
 sg13g2_fill_8 FILLER_106_1137 ();
 sg13g2_fill_2 FILLER_106_1145 ();
 sg13g2_fill_4 FILLER_106_1152 ();
 sg13g2_fill_2 FILLER_106_1164 ();
 sg13g2_fill_1 FILLER_106_1166 ();
 sg13g2_fill_2 FILLER_106_1177 ();
 sg13g2_fill_2 FILLER_106_1209 ();
 sg13g2_fill_1 FILLER_106_1215 ();
 sg13g2_fill_1 FILLER_106_1220 ();
 sg13g2_fill_4 FILLER_106_1227 ();
 sg13g2_fill_4 FILLER_106_1235 ();
 sg13g2_fill_2 FILLER_106_1249 ();
 sg13g2_fill_4 FILLER_106_1270 ();
 sg13g2_fill_2 FILLER_106_1274 ();
 sg13g2_fill_1 FILLER_106_1276 ();
 sg13g2_fill_8 FILLER_106_1282 ();
 sg13g2_fill_8 FILLER_106_1290 ();
 sg13g2_fill_8 FILLER_106_1298 ();
 sg13g2_fill_8 FILLER_106_1306 ();
 sg13g2_fill_4 FILLER_106_1314 ();
 sg13g2_fill_1 FILLER_106_1318 ();
 sg13g2_fill_2 FILLER_106_1340 ();
 sg13g2_fill_8 FILLER_106_1351 ();
 sg13g2_fill_8 FILLER_106_1359 ();
 sg13g2_fill_8 FILLER_106_1367 ();
 sg13g2_fill_4 FILLER_106_1375 ();
 sg13g2_fill_2 FILLER_106_1379 ();
 sg13g2_fill_1 FILLER_106_1381 ();
 sg13g2_fill_2 FILLER_106_1395 ();
 sg13g2_fill_8 FILLER_106_1411 ();
 sg13g2_fill_2 FILLER_106_1419 ();
 sg13g2_fill_1 FILLER_106_1421 ();
 sg13g2_fill_4 FILLER_106_1430 ();
 sg13g2_fill_2 FILLER_106_1434 ();
 sg13g2_fill_2 FILLER_106_1502 ();
 sg13g2_fill_8 FILLER_106_1528 ();
 sg13g2_fill_4 FILLER_106_1536 ();
 sg13g2_fill_1 FILLER_106_1540 ();
 sg13g2_fill_4 FILLER_106_1546 ();
 sg13g2_fill_2 FILLER_106_1550 ();
 sg13g2_fill_1 FILLER_106_1552 ();
 sg13g2_fill_2 FILLER_106_1562 ();
 sg13g2_fill_1 FILLER_106_1564 ();
 sg13g2_fill_8 FILLER_106_1570 ();
 sg13g2_fill_8 FILLER_106_1578 ();
 sg13g2_fill_4 FILLER_106_1586 ();
 sg13g2_fill_2 FILLER_106_1590 ();
 sg13g2_fill_8 FILLER_107_0 ();
 sg13g2_fill_8 FILLER_107_8 ();
 sg13g2_fill_8 FILLER_107_16 ();
 sg13g2_fill_8 FILLER_107_24 ();
 sg13g2_fill_8 FILLER_107_32 ();
 sg13g2_fill_8 FILLER_107_40 ();
 sg13g2_fill_8 FILLER_107_48 ();
 sg13g2_fill_8 FILLER_107_56 ();
 sg13g2_fill_8 FILLER_107_64 ();
 sg13g2_fill_8 FILLER_107_72 ();
 sg13g2_fill_8 FILLER_107_116 ();
 sg13g2_fill_4 FILLER_107_135 ();
 sg13g2_fill_1 FILLER_107_139 ();
 sg13g2_fill_8 FILLER_107_166 ();
 sg13g2_fill_2 FILLER_107_174 ();
 sg13g2_fill_1 FILLER_107_176 ();
 sg13g2_fill_8 FILLER_107_203 ();
 sg13g2_fill_8 FILLER_107_211 ();
 sg13g2_fill_8 FILLER_107_219 ();
 sg13g2_fill_8 FILLER_107_227 ();
 sg13g2_fill_1 FILLER_107_235 ();
 sg13g2_fill_1 FILLER_107_261 ();
 sg13g2_fill_8 FILLER_107_270 ();
 sg13g2_fill_1 FILLER_107_278 ();
 sg13g2_fill_4 FILLER_107_322 ();
 sg13g2_fill_2 FILLER_107_326 ();
 sg13g2_fill_1 FILLER_107_333 ();
 sg13g2_fill_8 FILLER_107_338 ();
 sg13g2_fill_2 FILLER_107_346 ();
 sg13g2_fill_2 FILLER_107_374 ();
 sg13g2_fill_8 FILLER_107_381 ();
 sg13g2_fill_8 FILLER_107_389 ();
 sg13g2_fill_4 FILLER_107_397 ();
 sg13g2_fill_2 FILLER_107_401 ();
 sg13g2_fill_1 FILLER_107_403 ();
 sg13g2_fill_8 FILLER_107_422 ();
 sg13g2_fill_8 FILLER_107_430 ();
 sg13g2_fill_8 FILLER_107_438 ();
 sg13g2_fill_8 FILLER_107_446 ();
 sg13g2_fill_8 FILLER_107_454 ();
 sg13g2_fill_8 FILLER_107_462 ();
 sg13g2_fill_4 FILLER_107_497 ();
 sg13g2_fill_1 FILLER_107_501 ();
 sg13g2_fill_8 FILLER_107_520 ();
 sg13g2_fill_4 FILLER_107_528 ();
 sg13g2_fill_2 FILLER_107_532 ();
 sg13g2_fill_4 FILLER_107_546 ();
 sg13g2_fill_8 FILLER_107_558 ();
 sg13g2_fill_1 FILLER_107_566 ();
 sg13g2_fill_8 FILLER_107_593 ();
 sg13g2_fill_1 FILLER_107_647 ();
 sg13g2_fill_8 FILLER_107_683 ();
 sg13g2_fill_1 FILLER_107_691 ();
 sg13g2_fill_8 FILLER_107_697 ();
 sg13g2_fill_2 FILLER_107_705 ();
 sg13g2_fill_1 FILLER_107_707 ();
 sg13g2_fill_8 FILLER_107_718 ();
 sg13g2_fill_8 FILLER_107_726 ();
 sg13g2_fill_8 FILLER_107_734 ();
 sg13g2_fill_8 FILLER_107_742 ();
 sg13g2_fill_8 FILLER_107_761 ();
 sg13g2_fill_8 FILLER_107_769 ();
 sg13g2_fill_4 FILLER_107_777 ();
 sg13g2_fill_1 FILLER_107_781 ();
 sg13g2_fill_2 FILLER_107_799 ();
 sg13g2_fill_1 FILLER_107_801 ();
 sg13g2_fill_4 FILLER_107_818 ();
 sg13g2_fill_1 FILLER_107_863 ();
 sg13g2_fill_8 FILLER_107_890 ();
 sg13g2_fill_4 FILLER_107_898 ();
 sg13g2_fill_8 FILLER_107_912 ();
 sg13g2_fill_8 FILLER_107_920 ();
 sg13g2_fill_4 FILLER_107_928 ();
 sg13g2_fill_2 FILLER_107_932 ();
 sg13g2_fill_2 FILLER_107_949 ();
 sg13g2_fill_1 FILLER_107_951 ();
 sg13g2_fill_2 FILLER_107_965 ();
 sg13g2_fill_2 FILLER_107_977 ();
 sg13g2_fill_4 FILLER_107_985 ();
 sg13g2_fill_4 FILLER_107_992 ();
 sg13g2_fill_4 FILLER_107_1036 ();
 sg13g2_fill_1 FILLER_107_1040 ();
 sg13g2_fill_1 FILLER_107_1054 ();
 sg13g2_fill_8 FILLER_107_1061 ();
 sg13g2_fill_8 FILLER_107_1074 ();
 sg13g2_fill_8 FILLER_107_1082 ();
 sg13g2_fill_2 FILLER_107_1090 ();
 sg13g2_fill_1 FILLER_107_1092 ();
 sg13g2_fill_2 FILLER_107_1108 ();
 sg13g2_fill_1 FILLER_107_1110 ();
 sg13g2_fill_4 FILLER_107_1131 ();
 sg13g2_fill_2 FILLER_107_1148 ();
 sg13g2_fill_8 FILLER_107_1165 ();
 sg13g2_fill_4 FILLER_107_1186 ();
 sg13g2_fill_8 FILLER_107_1200 ();
 sg13g2_fill_8 FILLER_107_1227 ();
 sg13g2_fill_2 FILLER_107_1235 ();
 sg13g2_fill_1 FILLER_107_1242 ();
 sg13g2_fill_8 FILLER_107_1263 ();
 sg13g2_fill_2 FILLER_107_1271 ();
 sg13g2_fill_1 FILLER_107_1299 ();
 sg13g2_fill_4 FILLER_107_1313 ();
 sg13g2_fill_1 FILLER_107_1317 ();
 sg13g2_fill_2 FILLER_107_1328 ();
 sg13g2_fill_1 FILLER_107_1330 ();
 sg13g2_fill_1 FILLER_107_1336 ();
 sg13g2_fill_2 FILLER_107_1350 ();
 sg13g2_fill_8 FILLER_107_1360 ();
 sg13g2_fill_1 FILLER_107_1368 ();
 sg13g2_fill_2 FILLER_107_1373 ();
 sg13g2_fill_1 FILLER_107_1375 ();
 sg13g2_fill_2 FILLER_107_1384 ();
 sg13g2_fill_1 FILLER_107_1386 ();
 sg13g2_fill_2 FILLER_107_1391 ();
 sg13g2_fill_8 FILLER_107_1398 ();
 sg13g2_fill_8 FILLER_107_1406 ();
 sg13g2_fill_4 FILLER_107_1414 ();
 sg13g2_fill_1 FILLER_107_1444 ();
 sg13g2_fill_8 FILLER_107_1470 ();
 sg13g2_fill_8 FILLER_107_1478 ();
 sg13g2_fill_8 FILLER_107_1486 ();
 sg13g2_fill_8 FILLER_107_1494 ();
 sg13g2_fill_2 FILLER_107_1514 ();
 sg13g2_fill_8 FILLER_107_1536 ();
 sg13g2_fill_1 FILLER_107_1544 ();
 sg13g2_fill_2 FILLER_107_1556 ();
 sg13g2_fill_2 FILLER_107_1563 ();
 sg13g2_fill_1 FILLER_107_1565 ();
 sg13g2_fill_8 FILLER_108_0 ();
 sg13g2_fill_8 FILLER_108_8 ();
 sg13g2_fill_8 FILLER_108_16 ();
 sg13g2_fill_2 FILLER_108_24 ();
 sg13g2_fill_1 FILLER_108_26 ();
 sg13g2_fill_8 FILLER_108_37 ();
 sg13g2_fill_8 FILLER_108_45 ();
 sg13g2_fill_1 FILLER_108_53 ();
 sg13g2_fill_8 FILLER_108_80 ();
 sg13g2_fill_8 FILLER_108_88 ();
 sg13g2_fill_4 FILLER_108_106 ();
 sg13g2_fill_2 FILLER_108_110 ();
 sg13g2_fill_1 FILLER_108_112 ();
 sg13g2_fill_8 FILLER_108_123 ();
 sg13g2_fill_8 FILLER_108_131 ();
 sg13g2_fill_4 FILLER_108_139 ();
 sg13g2_fill_1 FILLER_108_143 ();
 sg13g2_fill_8 FILLER_108_149 ();
 sg13g2_fill_8 FILLER_108_157 ();
 sg13g2_fill_1 FILLER_108_165 ();
 sg13g2_fill_8 FILLER_108_174 ();
 sg13g2_fill_8 FILLER_108_182 ();
 sg13g2_fill_8 FILLER_108_190 ();
 sg13g2_fill_4 FILLER_108_224 ();
 sg13g2_fill_2 FILLER_108_228 ();
 sg13g2_fill_1 FILLER_108_230 ();
 sg13g2_fill_1 FILLER_108_267 ();
 sg13g2_fill_4 FILLER_108_294 ();
 sg13g2_fill_1 FILLER_108_298 ();
 sg13g2_fill_8 FILLER_108_350 ();
 sg13g2_fill_8 FILLER_108_358 ();
 sg13g2_fill_8 FILLER_108_366 ();
 sg13g2_fill_1 FILLER_108_374 ();
 sg13g2_fill_8 FILLER_108_380 ();
 sg13g2_fill_1 FILLER_108_388 ();
 sg13g2_fill_8 FILLER_108_403 ();
 sg13g2_fill_4 FILLER_108_411 ();
 sg13g2_fill_1 FILLER_108_415 ();
 sg13g2_fill_8 FILLER_108_444 ();
 sg13g2_fill_2 FILLER_108_452 ();
 sg13g2_fill_1 FILLER_108_454 ();
 sg13g2_fill_4 FILLER_108_471 ();
 sg13g2_fill_2 FILLER_108_475 ();
 sg13g2_fill_1 FILLER_108_552 ();
 sg13g2_fill_8 FILLER_108_576 ();
 sg13g2_fill_8 FILLER_108_584 ();
 sg13g2_fill_4 FILLER_108_592 ();
 sg13g2_fill_2 FILLER_108_606 ();
 sg13g2_fill_8 FILLER_108_618 ();
 sg13g2_fill_8 FILLER_108_626 ();
 sg13g2_fill_2 FILLER_108_634 ();
 sg13g2_fill_2 FILLER_108_646 ();
 sg13g2_fill_2 FILLER_108_674 ();
 sg13g2_fill_1 FILLER_108_676 ();
 sg13g2_fill_8 FILLER_108_687 ();
 sg13g2_fill_4 FILLER_108_695 ();
 sg13g2_fill_1 FILLER_108_699 ();
 sg13g2_fill_2 FILLER_108_715 ();
 sg13g2_fill_2 FILLER_108_743 ();
 sg13g2_fill_4 FILLER_108_780 ();
 sg13g2_fill_1 FILLER_108_784 ();
 sg13g2_fill_1 FILLER_108_790 ();
 sg13g2_fill_2 FILLER_108_796 ();
 sg13g2_fill_1 FILLER_108_798 ();
 sg13g2_fill_1 FILLER_108_809 ();
 sg13g2_fill_8 FILLER_108_814 ();
 sg13g2_fill_8 FILLER_108_822 ();
 sg13g2_fill_8 FILLER_108_830 ();
 sg13g2_fill_2 FILLER_108_838 ();
 sg13g2_fill_1 FILLER_108_840 ();
 sg13g2_fill_2 FILLER_108_851 ();
 sg13g2_fill_4 FILLER_108_864 ();
 sg13g2_fill_8 FILLER_108_871 ();
 sg13g2_fill_2 FILLER_108_879 ();
 sg13g2_fill_1 FILLER_108_881 ();
 sg13g2_fill_2 FILLER_108_886 ();
 sg13g2_fill_1 FILLER_108_888 ();
 sg13g2_fill_4 FILLER_108_894 ();
 sg13g2_fill_8 FILLER_108_917 ();
 sg13g2_fill_8 FILLER_108_925 ();
 sg13g2_fill_8 FILLER_108_933 ();
 sg13g2_fill_8 FILLER_108_941 ();
 sg13g2_fill_8 FILLER_108_949 ();
 sg13g2_fill_4 FILLER_108_957 ();
 sg13g2_fill_8 FILLER_108_971 ();
 sg13g2_fill_8 FILLER_108_985 ();
 sg13g2_fill_8 FILLER_108_993 ();
 sg13g2_fill_8 FILLER_108_1001 ();
 sg13g2_fill_1 FILLER_108_1009 ();
 sg13g2_fill_8 FILLER_108_1016 ();
 sg13g2_fill_4 FILLER_108_1024 ();
 sg13g2_fill_8 FILLER_108_1031 ();
 sg13g2_fill_4 FILLER_108_1039 ();
 sg13g2_fill_2 FILLER_108_1043 ();
 sg13g2_fill_1 FILLER_108_1045 ();
 sg13g2_fill_2 FILLER_108_1056 ();
 sg13g2_fill_8 FILLER_108_1074 ();
 sg13g2_fill_8 FILLER_108_1082 ();
 sg13g2_fill_1 FILLER_108_1090 ();
 sg13g2_fill_2 FILLER_108_1096 ();
 sg13g2_fill_1 FILLER_108_1111 ();
 sg13g2_fill_2 FILLER_108_1117 ();
 sg13g2_fill_8 FILLER_108_1124 ();
 sg13g2_fill_8 FILLER_108_1132 ();
 sg13g2_fill_2 FILLER_108_1140 ();
 sg13g2_fill_8 FILLER_108_1146 ();
 sg13g2_fill_4 FILLER_108_1158 ();
 sg13g2_fill_2 FILLER_108_1162 ();
 sg13g2_fill_8 FILLER_108_1186 ();
 sg13g2_fill_8 FILLER_108_1194 ();
 sg13g2_fill_4 FILLER_108_1202 ();
 sg13g2_fill_1 FILLER_108_1206 ();
 sg13g2_fill_8 FILLER_108_1233 ();
 sg13g2_fill_2 FILLER_108_1241 ();
 sg13g2_fill_1 FILLER_108_1243 ();
 sg13g2_fill_2 FILLER_108_1264 ();
 sg13g2_fill_1 FILLER_108_1266 ();
 sg13g2_fill_4 FILLER_108_1273 ();
 sg13g2_fill_2 FILLER_108_1277 ();
 sg13g2_fill_2 FILLER_108_1288 ();
 sg13g2_fill_1 FILLER_108_1290 ();
 sg13g2_fill_1 FILLER_108_1321 ();
 sg13g2_fill_1 FILLER_108_1326 ();
 sg13g2_fill_8 FILLER_108_1348 ();
 sg13g2_fill_2 FILLER_108_1356 ();
 sg13g2_fill_2 FILLER_108_1383 ();
 sg13g2_fill_2 FILLER_108_1388 ();
 sg13g2_fill_1 FILLER_108_1390 ();
 sg13g2_fill_8 FILLER_108_1399 ();
 sg13g2_fill_4 FILLER_108_1407 ();
 sg13g2_fill_4 FILLER_108_1416 ();
 sg13g2_fill_2 FILLER_108_1420 ();
 sg13g2_fill_4 FILLER_108_1430 ();
 sg13g2_fill_1 FILLER_108_1434 ();
 sg13g2_fill_2 FILLER_108_1440 ();
 sg13g2_fill_1 FILLER_108_1461 ();
 sg13g2_fill_4 FILLER_108_1470 ();
 sg13g2_fill_1 FILLER_108_1474 ();
 sg13g2_fill_8 FILLER_108_1501 ();
 sg13g2_fill_4 FILLER_108_1509 ();
 sg13g2_fill_2 FILLER_108_1513 ();
 sg13g2_fill_1 FILLER_108_1515 ();
 sg13g2_fill_2 FILLER_108_1521 ();
 sg13g2_fill_8 FILLER_108_1528 ();
 sg13g2_fill_2 FILLER_108_1536 ();
 sg13g2_fill_8 FILLER_108_1543 ();
 sg13g2_fill_2 FILLER_108_1561 ();
 sg13g2_fill_1 FILLER_108_1563 ();
 sg13g2_fill_8 FILLER_108_1573 ();
 sg13g2_fill_8 FILLER_108_1581 ();
 sg13g2_fill_2 FILLER_108_1589 ();
 sg13g2_fill_1 FILLER_108_1591 ();
 sg13g2_fill_4 FILLER_109_0 ();
 sg13g2_fill_1 FILLER_109_4 ();
 sg13g2_fill_8 FILLER_109_15 ();
 sg13g2_fill_2 FILLER_109_55 ();
 sg13g2_fill_2 FILLER_109_113 ();
 sg13g2_fill_4 FILLER_109_135 ();
 sg13g2_fill_8 FILLER_109_189 ();
 sg13g2_fill_4 FILLER_109_197 ();
 sg13g2_fill_1 FILLER_109_201 ();
 sg13g2_fill_8 FILLER_109_247 ();
 sg13g2_fill_2 FILLER_109_255 ();
 sg13g2_fill_1 FILLER_109_257 ();
 sg13g2_fill_8 FILLER_109_287 ();
 sg13g2_fill_8 FILLER_109_295 ();
 sg13g2_fill_8 FILLER_109_303 ();
 sg13g2_fill_8 FILLER_109_311 ();
 sg13g2_fill_8 FILLER_109_335 ();
 sg13g2_fill_8 FILLER_109_343 ();
 sg13g2_fill_8 FILLER_109_351 ();
 sg13g2_fill_4 FILLER_109_359 ();
 sg13g2_fill_1 FILLER_109_363 ();
 sg13g2_fill_8 FILLER_109_404 ();
 sg13g2_fill_8 FILLER_109_412 ();
 sg13g2_fill_4 FILLER_109_433 ();
 sg13g2_fill_8 FILLER_109_488 ();
 sg13g2_fill_8 FILLER_109_496 ();
 sg13g2_fill_2 FILLER_109_504 ();
 sg13g2_fill_8 FILLER_109_519 ();
 sg13g2_fill_8 FILLER_109_527 ();
 sg13g2_fill_8 FILLER_109_535 ();
 sg13g2_fill_2 FILLER_109_543 ();
 sg13g2_fill_1 FILLER_109_545 ();
 sg13g2_fill_8 FILLER_109_554 ();
 sg13g2_fill_4 FILLER_109_562 ();
 sg13g2_fill_4 FILLER_109_592 ();
 sg13g2_fill_4 FILLER_109_606 ();
 sg13g2_fill_2 FILLER_109_610 ();
 sg13g2_fill_1 FILLER_109_612 ();
 sg13g2_fill_1 FILLER_109_628 ();
 sg13g2_fill_8 FILLER_109_642 ();
 sg13g2_fill_8 FILLER_109_650 ();
 sg13g2_fill_8 FILLER_109_658 ();
 sg13g2_fill_8 FILLER_109_666 ();
 sg13g2_fill_4 FILLER_109_674 ();
 sg13g2_fill_1 FILLER_109_678 ();
 sg13g2_fill_2 FILLER_109_684 ();
 sg13g2_fill_4 FILLER_109_699 ();
 sg13g2_fill_8 FILLER_109_723 ();
 sg13g2_fill_2 FILLER_109_760 ();
 sg13g2_fill_1 FILLER_109_762 ();
 sg13g2_fill_1 FILLER_109_773 ();
 sg13g2_fill_4 FILLER_109_784 ();
 sg13g2_fill_2 FILLER_109_793 ();
 sg13g2_fill_1 FILLER_109_795 ();
 sg13g2_fill_2 FILLER_109_823 ();
 sg13g2_fill_1 FILLER_109_825 ();
 sg13g2_fill_8 FILLER_109_842 ();
 sg13g2_fill_2 FILLER_109_850 ();
 sg13g2_fill_1 FILLER_109_852 ();
 sg13g2_fill_8 FILLER_109_858 ();
 sg13g2_fill_4 FILLER_109_866 ();
 sg13g2_fill_8 FILLER_109_879 ();
 sg13g2_fill_4 FILLER_109_887 ();
 sg13g2_fill_2 FILLER_109_896 ();
 sg13g2_fill_1 FILLER_109_898 ();
 sg13g2_fill_8 FILLER_109_912 ();
 sg13g2_fill_8 FILLER_109_937 ();
 sg13g2_fill_4 FILLER_109_945 ();
 sg13g2_fill_1 FILLER_109_949 ();
 sg13g2_fill_8 FILLER_109_958 ();
 sg13g2_fill_8 FILLER_109_966 ();
 sg13g2_fill_2 FILLER_109_992 ();
 sg13g2_fill_2 FILLER_109_1016 ();
 sg13g2_fill_1 FILLER_109_1018 ();
 sg13g2_fill_2 FILLER_109_1022 ();
 sg13g2_fill_4 FILLER_109_1037 ();
 sg13g2_fill_1 FILLER_109_1041 ();
 sg13g2_fill_1 FILLER_109_1054 ();
 sg13g2_fill_8 FILLER_109_1063 ();
 sg13g2_fill_2 FILLER_109_1083 ();
 sg13g2_fill_1 FILLER_109_1085 ();
 sg13g2_fill_2 FILLER_109_1098 ();
 sg13g2_fill_1 FILLER_109_1100 ();
 sg13g2_fill_2 FILLER_109_1109 ();
 sg13g2_fill_1 FILLER_109_1111 ();
 sg13g2_fill_8 FILLER_109_1130 ();
 sg13g2_fill_8 FILLER_109_1160 ();
 sg13g2_fill_1 FILLER_109_1185 ();
 sg13g2_fill_8 FILLER_109_1197 ();
 sg13g2_fill_8 FILLER_109_1205 ();
 sg13g2_fill_2 FILLER_109_1213 ();
 sg13g2_fill_1 FILLER_109_1215 ();
 sg13g2_fill_8 FILLER_109_1234 ();
 sg13g2_fill_4 FILLER_109_1247 ();
 sg13g2_fill_1 FILLER_109_1251 ();
 sg13g2_fill_8 FILLER_109_1266 ();
 sg13g2_fill_1 FILLER_109_1274 ();
 sg13g2_fill_1 FILLER_109_1287 ();
 sg13g2_fill_8 FILLER_109_1293 ();
 sg13g2_fill_1 FILLER_109_1301 ();
 sg13g2_fill_2 FILLER_109_1306 ();
 sg13g2_fill_8 FILLER_109_1322 ();
 sg13g2_fill_8 FILLER_109_1330 ();
 sg13g2_fill_2 FILLER_109_1338 ();
 sg13g2_fill_4 FILLER_109_1350 ();
 sg13g2_fill_2 FILLER_109_1354 ();
 sg13g2_fill_1 FILLER_109_1368 ();
 sg13g2_fill_1 FILLER_109_1386 ();
 sg13g2_fill_8 FILLER_109_1441 ();
 sg13g2_fill_4 FILLER_109_1449 ();
 sg13g2_fill_2 FILLER_109_1453 ();
 sg13g2_fill_1 FILLER_109_1455 ();
 sg13g2_fill_8 FILLER_109_1487 ();
 sg13g2_fill_4 FILLER_109_1495 ();
 sg13g2_fill_1 FILLER_109_1499 ();
 sg13g2_fill_8 FILLER_109_1525 ();
 sg13g2_fill_8 FILLER_109_1533 ();
 sg13g2_fill_2 FILLER_109_1564 ();
 sg13g2_fill_1 FILLER_109_1591 ();
 sg13g2_fill_4 FILLER_110_0 ();
 sg13g2_fill_2 FILLER_110_4 ();
 sg13g2_fill_1 FILLER_110_32 ();
 sg13g2_fill_8 FILLER_110_71 ();
 sg13g2_fill_8 FILLER_110_79 ();
 sg13g2_fill_4 FILLER_110_87 ();
 sg13g2_fill_1 FILLER_110_91 ();
 sg13g2_fill_1 FILLER_110_164 ();
 sg13g2_fill_8 FILLER_110_175 ();
 sg13g2_fill_4 FILLER_110_183 ();
 sg13g2_fill_2 FILLER_110_187 ();
 sg13g2_fill_1 FILLER_110_189 ();
 sg13g2_fill_2 FILLER_110_200 ();
 sg13g2_fill_4 FILLER_110_223 ();
 sg13g2_fill_1 FILLER_110_227 ();
 sg13g2_fill_8 FILLER_110_233 ();
 sg13g2_fill_8 FILLER_110_241 ();
 sg13g2_fill_2 FILLER_110_249 ();
 sg13g2_fill_1 FILLER_110_251 ();
 sg13g2_fill_8 FILLER_110_277 ();
 sg13g2_fill_8 FILLER_110_285 ();
 sg13g2_fill_8 FILLER_110_293 ();
 sg13g2_fill_8 FILLER_110_301 ();
 sg13g2_fill_8 FILLER_110_309 ();
 sg13g2_fill_8 FILLER_110_317 ();
 sg13g2_fill_4 FILLER_110_325 ();
 sg13g2_fill_2 FILLER_110_329 ();
 sg13g2_fill_4 FILLER_110_339 ();
 sg13g2_fill_1 FILLER_110_343 ();
 sg13g2_fill_1 FILLER_110_359 ();
 sg13g2_fill_2 FILLER_110_370 ();
 sg13g2_fill_1 FILLER_110_372 ();
 sg13g2_fill_4 FILLER_110_381 ();
 sg13g2_fill_1 FILLER_110_385 ();
 sg13g2_fill_4 FILLER_110_412 ();
 sg13g2_fill_4 FILLER_110_446 ();
 sg13g2_fill_2 FILLER_110_450 ();
 sg13g2_fill_1 FILLER_110_452 ();
 sg13g2_fill_8 FILLER_110_489 ();
 sg13g2_fill_8 FILLER_110_497 ();
 sg13g2_fill_8 FILLER_110_505 ();
 sg13g2_fill_8 FILLER_110_535 ();
 sg13g2_fill_2 FILLER_110_543 ();
 sg13g2_fill_1 FILLER_110_545 ();
 sg13g2_fill_4 FILLER_110_554 ();
 sg13g2_fill_2 FILLER_110_558 ();
 sg13g2_fill_8 FILLER_110_570 ();
 sg13g2_fill_2 FILLER_110_604 ();
 sg13g2_fill_1 FILLER_110_622 ();
 sg13g2_fill_8 FILLER_110_649 ();
 sg13g2_fill_4 FILLER_110_657 ();
 sg13g2_fill_2 FILLER_110_661 ();
 sg13g2_fill_4 FILLER_110_679 ();
 sg13g2_fill_1 FILLER_110_683 ();
 sg13g2_fill_8 FILLER_110_694 ();
 sg13g2_fill_8 FILLER_110_702 ();
 sg13g2_fill_8 FILLER_110_710 ();
 sg13g2_fill_2 FILLER_110_718 ();
 sg13g2_fill_1 FILLER_110_720 ();
 sg13g2_fill_8 FILLER_110_731 ();
 sg13g2_fill_8 FILLER_110_739 ();
 sg13g2_fill_2 FILLER_110_771 ();
 sg13g2_fill_1 FILLER_110_788 ();
 sg13g2_fill_4 FILLER_110_803 ();
 sg13g2_fill_1 FILLER_110_836 ();
 sg13g2_fill_2 FILLER_110_847 ();
 sg13g2_fill_8 FILLER_110_857 ();
 sg13g2_fill_8 FILLER_110_865 ();
 sg13g2_fill_4 FILLER_110_873 ();
 sg13g2_fill_1 FILLER_110_877 ();
 sg13g2_fill_8 FILLER_110_888 ();
 sg13g2_fill_8 FILLER_110_896 ();
 sg13g2_fill_2 FILLER_110_904 ();
 sg13g2_fill_2 FILLER_110_912 ();
 sg13g2_fill_1 FILLER_110_914 ();
 sg13g2_fill_2 FILLER_110_938 ();
 sg13g2_fill_4 FILLER_110_969 ();
 sg13g2_fill_1 FILLER_110_1023 ();
 sg13g2_fill_2 FILLER_110_1030 ();
 sg13g2_fill_1 FILLER_110_1032 ();
 sg13g2_fill_1 FILLER_110_1041 ();
 sg13g2_fill_2 FILLER_110_1055 ();
 sg13g2_fill_1 FILLER_110_1076 ();
 sg13g2_fill_8 FILLER_110_1089 ();
 sg13g2_fill_8 FILLER_110_1097 ();
 sg13g2_fill_8 FILLER_110_1105 ();
 sg13g2_fill_8 FILLER_110_1113 ();
 sg13g2_fill_8 FILLER_110_1121 ();
 sg13g2_fill_8 FILLER_110_1129 ();
 sg13g2_fill_4 FILLER_110_1137 ();
 sg13g2_fill_1 FILLER_110_1141 ();
 sg13g2_fill_4 FILLER_110_1206 ();
 sg13g2_fill_2 FILLER_110_1210 ();
 sg13g2_fill_4 FILLER_110_1230 ();
 sg13g2_fill_1 FILLER_110_1234 ();
 sg13g2_fill_8 FILLER_110_1239 ();
 sg13g2_fill_8 FILLER_110_1247 ();
 sg13g2_fill_4 FILLER_110_1255 ();
 sg13g2_fill_2 FILLER_110_1259 ();
 sg13g2_fill_2 FILLER_110_1269 ();
 sg13g2_fill_2 FILLER_110_1282 ();
 sg13g2_fill_1 FILLER_110_1284 ();
 sg13g2_fill_8 FILLER_110_1301 ();
 sg13g2_fill_1 FILLER_110_1309 ();
 sg13g2_fill_8 FILLER_110_1329 ();
 sg13g2_fill_1 FILLER_110_1337 ();
 sg13g2_fill_4 FILLER_110_1353 ();
 sg13g2_fill_2 FILLER_110_1357 ();
 sg13g2_fill_1 FILLER_110_1359 ();
 sg13g2_fill_4 FILLER_110_1373 ();
 sg13g2_fill_1 FILLER_110_1377 ();
 sg13g2_fill_2 FILLER_110_1385 ();
 sg13g2_fill_8 FILLER_110_1400 ();
 sg13g2_fill_8 FILLER_110_1408 ();
 sg13g2_fill_8 FILLER_110_1416 ();
 sg13g2_fill_8 FILLER_110_1424 ();
 sg13g2_fill_8 FILLER_110_1432 ();
 sg13g2_fill_4 FILLER_110_1440 ();
 sg13g2_fill_1 FILLER_110_1444 ();
 sg13g2_fill_2 FILLER_110_1450 ();
 sg13g2_fill_1 FILLER_110_1452 ();
 sg13g2_fill_8 FILLER_110_1472 ();
 sg13g2_fill_8 FILLER_110_1480 ();
 sg13g2_fill_8 FILLER_110_1488 ();
 sg13g2_fill_4 FILLER_110_1496 ();
 sg13g2_fill_2 FILLER_110_1500 ();
 sg13g2_fill_2 FILLER_110_1535 ();
 sg13g2_fill_8 FILLER_110_1579 ();
 sg13g2_fill_4 FILLER_110_1587 ();
 sg13g2_fill_1 FILLER_110_1591 ();
 sg13g2_fill_2 FILLER_111_0 ();
 sg13g2_fill_1 FILLER_111_2 ();
 sg13g2_fill_8 FILLER_111_44 ();
 sg13g2_fill_8 FILLER_111_72 ();
 sg13g2_fill_2 FILLER_111_80 ();
 sg13g2_fill_1 FILLER_111_82 ();
 sg13g2_fill_4 FILLER_111_88 ();
 sg13g2_fill_2 FILLER_111_92 ();
 sg13g2_fill_2 FILLER_111_97 ();
 sg13g2_fill_1 FILLER_111_107 ();
 sg13g2_fill_8 FILLER_111_133 ();
 sg13g2_fill_8 FILLER_111_141 ();
 sg13g2_fill_4 FILLER_111_149 ();
 sg13g2_fill_1 FILLER_111_153 ();
 sg13g2_fill_8 FILLER_111_206 ();
 sg13g2_fill_4 FILLER_111_214 ();
 sg13g2_fill_2 FILLER_111_218 ();
 sg13g2_fill_1 FILLER_111_220 ();
 sg13g2_fill_1 FILLER_111_265 ();
 sg13g2_fill_2 FILLER_111_342 ();
 sg13g2_fill_8 FILLER_111_386 ();
 sg13g2_fill_4 FILLER_111_394 ();
 sg13g2_fill_1 FILLER_111_398 ();
 sg13g2_fill_8 FILLER_111_409 ();
 sg13g2_fill_4 FILLER_111_417 ();
 sg13g2_fill_8 FILLER_111_451 ();
 sg13g2_fill_2 FILLER_111_459 ();
 sg13g2_fill_2 FILLER_111_506 ();
 sg13g2_fill_1 FILLER_111_508 ();
 sg13g2_fill_8 FILLER_111_518 ();
 sg13g2_fill_4 FILLER_111_526 ();
 sg13g2_fill_2 FILLER_111_530 ();
 sg13g2_fill_8 FILLER_111_558 ();
 sg13g2_fill_8 FILLER_111_566 ();
 sg13g2_fill_8 FILLER_111_574 ();
 sg13g2_fill_8 FILLER_111_622 ();
 sg13g2_fill_4 FILLER_111_630 ();
 sg13g2_fill_1 FILLER_111_634 ();
 sg13g2_fill_2 FILLER_111_645 ();
 sg13g2_fill_1 FILLER_111_647 ();
 sg13g2_fill_4 FILLER_111_656 ();
 sg13g2_fill_2 FILLER_111_660 ();
 sg13g2_fill_4 FILLER_111_679 ();
 sg13g2_fill_1 FILLER_111_683 ();
 sg13g2_fill_4 FILLER_111_710 ();
 sg13g2_fill_8 FILLER_111_740 ();
 sg13g2_fill_4 FILLER_111_748 ();
 sg13g2_fill_2 FILLER_111_752 ();
 sg13g2_fill_8 FILLER_111_789 ();
 sg13g2_fill_8 FILLER_111_797 ();
 sg13g2_fill_8 FILLER_111_805 ();
 sg13g2_fill_8 FILLER_111_817 ();
 sg13g2_fill_2 FILLER_111_825 ();
 sg13g2_fill_4 FILLER_111_832 ();
 sg13g2_fill_1 FILLER_111_836 ();
 sg13g2_fill_4 FILLER_111_842 ();
 sg13g2_fill_2 FILLER_111_846 ();
 sg13g2_fill_1 FILLER_111_848 ();
 sg13g2_fill_1 FILLER_111_885 ();
 sg13g2_fill_8 FILLER_111_897 ();
 sg13g2_fill_1 FILLER_111_905 ();
 sg13g2_fill_8 FILLER_111_941 ();
 sg13g2_fill_2 FILLER_111_949 ();
 sg13g2_fill_1 FILLER_111_951 ();
 sg13g2_fill_2 FILLER_111_961 ();
 sg13g2_fill_1 FILLER_111_963 ();
 sg13g2_fill_4 FILLER_111_981 ();
 sg13g2_fill_2 FILLER_111_993 ();
 sg13g2_fill_2 FILLER_111_1014 ();
 sg13g2_fill_1 FILLER_111_1016 ();
 sg13g2_fill_2 FILLER_111_1022 ();
 sg13g2_fill_1 FILLER_111_1033 ();
 sg13g2_fill_1 FILLER_111_1053 ();
 sg13g2_fill_8 FILLER_111_1062 ();
 sg13g2_fill_2 FILLER_111_1070 ();
 sg13g2_fill_2 FILLER_111_1086 ();
 sg13g2_fill_1 FILLER_111_1088 ();
 sg13g2_fill_8 FILLER_111_1121 ();
 sg13g2_fill_8 FILLER_111_1129 ();
 sg13g2_fill_8 FILLER_111_1153 ();
 sg13g2_fill_1 FILLER_111_1161 ();
 sg13g2_fill_8 FILLER_111_1170 ();
 sg13g2_fill_2 FILLER_111_1196 ();
 sg13g2_fill_8 FILLER_111_1206 ();
 sg13g2_fill_1 FILLER_111_1214 ();
 sg13g2_fill_8 FILLER_111_1225 ();
 sg13g2_fill_4 FILLER_111_1233 ();
 sg13g2_fill_2 FILLER_111_1237 ();
 sg13g2_fill_8 FILLER_111_1249 ();
 sg13g2_fill_2 FILLER_111_1277 ();
 sg13g2_fill_1 FILLER_111_1279 ();
 sg13g2_fill_2 FILLER_111_1285 ();
 sg13g2_fill_1 FILLER_111_1287 ();
 sg13g2_fill_8 FILLER_111_1299 ();
 sg13g2_fill_1 FILLER_111_1307 ();
 sg13g2_fill_2 FILLER_111_1316 ();
 sg13g2_fill_1 FILLER_111_1334 ();
 sg13g2_fill_4 FILLER_111_1354 ();
 sg13g2_fill_1 FILLER_111_1358 ();
 sg13g2_fill_8 FILLER_111_1362 ();
 sg13g2_fill_8 FILLER_111_1370 ();
 sg13g2_fill_8 FILLER_111_1378 ();
 sg13g2_fill_8 FILLER_111_1386 ();
 sg13g2_fill_8 FILLER_111_1394 ();
 sg13g2_fill_8 FILLER_111_1402 ();
 sg13g2_fill_8 FILLER_111_1410 ();
 sg13g2_fill_2 FILLER_111_1418 ();
 sg13g2_fill_1 FILLER_111_1420 ();
 sg13g2_fill_2 FILLER_111_1447 ();
 sg13g2_fill_2 FILLER_111_1455 ();
 sg13g2_fill_1 FILLER_111_1457 ();
 sg13g2_fill_4 FILLER_111_1466 ();
 sg13g2_fill_1 FILLER_111_1470 ();
 sg13g2_fill_8 FILLER_111_1506 ();
 sg13g2_fill_4 FILLER_111_1514 ();
 sg13g2_fill_2 FILLER_111_1518 ();
 sg13g2_fill_8 FILLER_111_1525 ();
 sg13g2_fill_4 FILLER_111_1533 ();
 sg13g2_fill_1 FILLER_111_1537 ();
 sg13g2_fill_4 FILLER_112_0 ();
 sg13g2_fill_8 FILLER_112_14 ();
 sg13g2_fill_8 FILLER_112_22 ();
 sg13g2_fill_1 FILLER_112_30 ();
 sg13g2_fill_2 FILLER_112_83 ();
 sg13g2_fill_1 FILLER_112_85 ();
 sg13g2_fill_1 FILLER_112_102 ();
 sg13g2_fill_4 FILLER_112_132 ();
 sg13g2_fill_1 FILLER_112_136 ();
 sg13g2_fill_8 FILLER_112_153 ();
 sg13g2_fill_4 FILLER_112_161 ();
 sg13g2_fill_2 FILLER_112_165 ();
 sg13g2_fill_4 FILLER_112_197 ();
 sg13g2_fill_2 FILLER_112_201 ();
 sg13g2_fill_8 FILLER_112_213 ();
 sg13g2_fill_4 FILLER_112_221 ();
 sg13g2_fill_2 FILLER_112_225 ();
 sg13g2_fill_1 FILLER_112_227 ();
 sg13g2_fill_4 FILLER_112_233 ();
 sg13g2_fill_2 FILLER_112_237 ();
 sg13g2_fill_1 FILLER_112_239 ();
 sg13g2_fill_2 FILLER_112_250 ();
 sg13g2_fill_8 FILLER_112_277 ();
 sg13g2_fill_2 FILLER_112_285 ();
 sg13g2_fill_8 FILLER_112_322 ();
 sg13g2_fill_8 FILLER_112_330 ();
 sg13g2_fill_4 FILLER_112_338 ();
 sg13g2_fill_8 FILLER_112_363 ();
 sg13g2_fill_1 FILLER_112_371 ();
 sg13g2_fill_8 FILLER_112_376 ();
 sg13g2_fill_8 FILLER_112_384 ();
 sg13g2_fill_2 FILLER_112_392 ();
 sg13g2_fill_4 FILLER_112_418 ();
 sg13g2_fill_8 FILLER_112_429 ();
 sg13g2_fill_2 FILLER_112_437 ();
 sg13g2_fill_1 FILLER_112_439 ();
 sg13g2_fill_8 FILLER_112_456 ();
 sg13g2_fill_2 FILLER_112_464 ();
 sg13g2_fill_4 FILLER_112_476 ();
 sg13g2_fill_1 FILLER_112_480 ();
 sg13g2_fill_8 FILLER_112_486 ();
 sg13g2_fill_4 FILLER_112_494 ();
 sg13g2_fill_1 FILLER_112_498 ();
 sg13g2_fill_1 FILLER_112_507 ();
 sg13g2_fill_2 FILLER_112_524 ();
 sg13g2_fill_1 FILLER_112_526 ();
 sg13g2_fill_4 FILLER_112_545 ();
 sg13g2_fill_2 FILLER_112_549 ();
 sg13g2_fill_2 FILLER_112_559 ();
 sg13g2_fill_8 FILLER_112_565 ();
 sg13g2_fill_8 FILLER_112_573 ();
 sg13g2_fill_8 FILLER_112_581 ();
 sg13g2_fill_8 FILLER_112_589 ();
 sg13g2_fill_2 FILLER_112_597 ();
 sg13g2_fill_1 FILLER_112_599 ();
 sg13g2_fill_4 FILLER_112_607 ();
 sg13g2_fill_4 FILLER_112_647 ();
 sg13g2_fill_4 FILLER_112_655 ();
 sg13g2_fill_2 FILLER_112_659 ();
 sg13g2_fill_1 FILLER_112_697 ();
 sg13g2_fill_1 FILLER_112_718 ();
 sg13g2_fill_8 FILLER_112_760 ();
 sg13g2_fill_2 FILLER_112_768 ();
 sg13g2_fill_2 FILLER_112_777 ();
 sg13g2_fill_1 FILLER_112_779 ();
 sg13g2_fill_8 FILLER_112_789 ();
 sg13g2_fill_2 FILLER_112_797 ();
 sg13g2_fill_2 FILLER_112_816 ();
 sg13g2_fill_2 FILLER_112_823 ();
 sg13g2_fill_2 FILLER_112_830 ();
 sg13g2_fill_4 FILLER_112_842 ();
 sg13g2_fill_2 FILLER_112_846 ();
 sg13g2_fill_1 FILLER_112_848 ();
 sg13g2_fill_8 FILLER_112_860 ();
 sg13g2_fill_4 FILLER_112_868 ();
 sg13g2_fill_8 FILLER_112_895 ();
 sg13g2_fill_2 FILLER_112_911 ();
 sg13g2_fill_4 FILLER_112_918 ();
 sg13g2_fill_2 FILLER_112_922 ();
 sg13g2_fill_8 FILLER_112_933 ();
 sg13g2_fill_1 FILLER_112_941 ();
 sg13g2_fill_2 FILLER_112_951 ();
 sg13g2_fill_2 FILLER_112_993 ();
 sg13g2_fill_2 FILLER_112_1000 ();
 sg13g2_fill_1 FILLER_112_1002 ();
 sg13g2_fill_4 FILLER_112_1008 ();
 sg13g2_fill_2 FILLER_112_1012 ();
 sg13g2_fill_8 FILLER_112_1020 ();
 sg13g2_fill_8 FILLER_112_1028 ();
 sg13g2_fill_8 FILLER_112_1046 ();
 sg13g2_fill_8 FILLER_112_1054 ();
 sg13g2_fill_8 FILLER_112_1062 ();
 sg13g2_fill_2 FILLER_112_1070 ();
 sg13g2_fill_8 FILLER_112_1087 ();
 sg13g2_fill_8 FILLER_112_1095 ();
 sg13g2_fill_4 FILLER_112_1108 ();
 sg13g2_fill_2 FILLER_112_1112 ();
 sg13g2_fill_1 FILLER_112_1114 ();
 sg13g2_fill_4 FILLER_112_1132 ();
 sg13g2_fill_8 FILLER_112_1141 ();
 sg13g2_fill_4 FILLER_112_1149 ();
 sg13g2_fill_4 FILLER_112_1158 ();
 sg13g2_fill_1 FILLER_112_1162 ();
 sg13g2_fill_8 FILLER_112_1171 ();
 sg13g2_fill_8 FILLER_112_1179 ();
 sg13g2_fill_8 FILLER_112_1187 ();
 sg13g2_fill_8 FILLER_112_1195 ();
 sg13g2_fill_8 FILLER_112_1203 ();
 sg13g2_fill_4 FILLER_112_1211 ();
 sg13g2_fill_2 FILLER_112_1215 ();
 sg13g2_fill_1 FILLER_112_1217 ();
 sg13g2_fill_2 FILLER_112_1224 ();
 sg13g2_fill_4 FILLER_112_1234 ();
 sg13g2_fill_2 FILLER_112_1238 ();
 sg13g2_fill_1 FILLER_112_1240 ();
 sg13g2_fill_4 FILLER_112_1245 ();
 sg13g2_fill_4 FILLER_112_1257 ();
 sg13g2_fill_1 FILLER_112_1261 ();
 sg13g2_fill_2 FILLER_112_1266 ();
 sg13g2_fill_1 FILLER_112_1268 ();
 sg13g2_fill_8 FILLER_112_1274 ();
 sg13g2_fill_4 FILLER_112_1282 ();
 sg13g2_fill_1 FILLER_112_1286 ();
 sg13g2_fill_4 FILLER_112_1296 ();
 sg13g2_fill_8 FILLER_112_1304 ();
 sg13g2_fill_1 FILLER_112_1312 ();
 sg13g2_fill_2 FILLER_112_1317 ();
 sg13g2_fill_1 FILLER_112_1319 ();
 sg13g2_fill_8 FILLER_112_1325 ();
 sg13g2_fill_2 FILLER_112_1333 ();
 sg13g2_fill_1 FILLER_112_1339 ();
 sg13g2_fill_8 FILLER_112_1349 ();
 sg13g2_fill_4 FILLER_112_1357 ();
 sg13g2_fill_1 FILLER_112_1371 ();
 sg13g2_fill_4 FILLER_112_1438 ();
 sg13g2_fill_2 FILLER_112_1442 ();
 sg13g2_fill_1 FILLER_112_1444 ();
 sg13g2_fill_4 FILLER_112_1450 ();
 sg13g2_fill_8 FILLER_112_1458 ();
 sg13g2_fill_4 FILLER_112_1466 ();
 sg13g2_fill_1 FILLER_112_1470 ();
 sg13g2_fill_2 FILLER_112_1476 ();
 sg13g2_fill_1 FILLER_112_1478 ();
 sg13g2_fill_1 FILLER_112_1484 ();
 sg13g2_fill_2 FILLER_112_1511 ();
 sg13g2_fill_8 FILLER_112_1539 ();
 sg13g2_fill_1 FILLER_112_1547 ();
 sg13g2_fill_1 FILLER_112_1577 ();
 sg13g2_fill_2 FILLER_112_1589 ();
 sg13g2_fill_1 FILLER_112_1591 ();
 sg13g2_fill_4 FILLER_113_0 ();
 sg13g2_fill_1 FILLER_113_4 ();
 sg13g2_fill_4 FILLER_113_15 ();
 sg13g2_fill_8 FILLER_113_54 ();
 sg13g2_fill_4 FILLER_113_62 ();
 sg13g2_fill_1 FILLER_113_66 ();
 sg13g2_fill_2 FILLER_113_89 ();
 sg13g2_fill_1 FILLER_113_91 ();
 sg13g2_fill_8 FILLER_113_146 ();
 sg13g2_fill_8 FILLER_113_154 ();
 sg13g2_fill_8 FILLER_113_162 ();
 sg13g2_fill_8 FILLER_113_170 ();
 sg13g2_fill_4 FILLER_113_178 ();
 sg13g2_fill_2 FILLER_113_182 ();
 sg13g2_fill_8 FILLER_113_192 ();
 sg13g2_fill_4 FILLER_113_200 ();
 sg13g2_fill_1 FILLER_113_204 ();
 sg13g2_fill_8 FILLER_113_239 ();
 sg13g2_fill_1 FILLER_113_247 ();
 sg13g2_fill_8 FILLER_113_274 ();
 sg13g2_fill_8 FILLER_113_282 ();
 sg13g2_fill_2 FILLER_113_290 ();
 sg13g2_fill_1 FILLER_113_306 ();
 sg13g2_fill_8 FILLER_113_328 ();
 sg13g2_fill_4 FILLER_113_336 ();
 sg13g2_fill_2 FILLER_113_340 ();
 sg13g2_fill_4 FILLER_113_352 ();
 sg13g2_fill_1 FILLER_113_356 ();
 sg13g2_fill_4 FILLER_113_403 ();
 sg13g2_fill_4 FILLER_113_425 ();
 sg13g2_fill_8 FILLER_113_437 ();
 sg13g2_fill_1 FILLER_113_445 ();
 sg13g2_fill_8 FILLER_113_454 ();
 sg13g2_fill_8 FILLER_113_462 ();
 sg13g2_fill_8 FILLER_113_474 ();
 sg13g2_fill_8 FILLER_113_482 ();
 sg13g2_fill_4 FILLER_113_498 ();
 sg13g2_fill_8 FILLER_113_507 ();
 sg13g2_fill_4 FILLER_113_515 ();
 sg13g2_fill_8 FILLER_113_527 ();
 sg13g2_fill_8 FILLER_113_543 ();
 sg13g2_fill_8 FILLER_113_551 ();
 sg13g2_fill_1 FILLER_113_559 ();
 sg13g2_fill_8 FILLER_113_576 ();
 sg13g2_fill_4 FILLER_113_592 ();
 sg13g2_fill_1 FILLER_113_596 ();
 sg13g2_fill_8 FILLER_113_611 ();
 sg13g2_fill_8 FILLER_113_619 ();
 sg13g2_fill_2 FILLER_113_643 ();
 sg13g2_fill_8 FILLER_113_653 ();
 sg13g2_fill_1 FILLER_113_661 ();
 sg13g2_fill_8 FILLER_113_667 ();
 sg13g2_fill_8 FILLER_113_675 ();
 sg13g2_fill_8 FILLER_113_683 ();
 sg13g2_fill_8 FILLER_113_691 ();
 sg13g2_fill_1 FILLER_113_699 ();
 sg13g2_fill_4 FILLER_113_710 ();
 sg13g2_fill_2 FILLER_113_747 ();
 sg13g2_fill_1 FILLER_113_749 ();
 sg13g2_fill_1 FILLER_113_788 ();
 sg13g2_fill_2 FILLER_113_817 ();
 sg13g2_fill_1 FILLER_113_829 ();
 sg13g2_fill_1 FILLER_113_842 ();
 sg13g2_fill_1 FILLER_113_854 ();
 sg13g2_fill_1 FILLER_113_863 ();
 sg13g2_fill_8 FILLER_113_872 ();
 sg13g2_fill_4 FILLER_113_883 ();
 sg13g2_fill_2 FILLER_113_887 ();
 sg13g2_fill_1 FILLER_113_905 ();
 sg13g2_fill_8 FILLER_113_919 ();
 sg13g2_fill_1 FILLER_113_932 ();
 sg13g2_fill_1 FILLER_113_963 ();
 sg13g2_fill_8 FILLER_113_978 ();
 sg13g2_fill_8 FILLER_113_986 ();
 sg13g2_fill_8 FILLER_113_994 ();
 sg13g2_fill_8 FILLER_113_1002 ();
 sg13g2_fill_1 FILLER_113_1010 ();
 sg13g2_fill_2 FILLER_113_1020 ();
 sg13g2_fill_1 FILLER_113_1028 ();
 sg13g2_fill_1 FILLER_113_1034 ();
 sg13g2_fill_4 FILLER_113_1055 ();
 sg13g2_fill_4 FILLER_113_1080 ();
 sg13g2_fill_2 FILLER_113_1084 ();
 sg13g2_fill_1 FILLER_113_1086 ();
 sg13g2_fill_2 FILLER_113_1092 ();
 sg13g2_fill_1 FILLER_113_1094 ();
 sg13g2_fill_2 FILLER_113_1100 ();
 sg13g2_fill_1 FILLER_113_1102 ();
 sg13g2_fill_4 FILLER_113_1118 ();
 sg13g2_fill_1 FILLER_113_1122 ();
 sg13g2_fill_4 FILLER_113_1128 ();
 sg13g2_fill_2 FILLER_113_1132 ();
 sg13g2_fill_2 FILLER_113_1147 ();
 sg13g2_fill_1 FILLER_113_1149 ();
 sg13g2_fill_4 FILLER_113_1158 ();
 sg13g2_fill_2 FILLER_113_1162 ();
 sg13g2_fill_4 FILLER_113_1172 ();
 sg13g2_fill_1 FILLER_113_1192 ();
 sg13g2_fill_2 FILLER_113_1218 ();
 sg13g2_fill_1 FILLER_113_1220 ();
 sg13g2_fill_2 FILLER_113_1257 ();
 sg13g2_fill_8 FILLER_113_1266 ();
 sg13g2_fill_8 FILLER_113_1279 ();
 sg13g2_fill_2 FILLER_113_1287 ();
 sg13g2_fill_1 FILLER_113_1289 ();
 sg13g2_fill_4 FILLER_113_1297 ();
 sg13g2_fill_8 FILLER_113_1328 ();
 sg13g2_fill_8 FILLER_113_1336 ();
 sg13g2_fill_2 FILLER_113_1344 ();
 sg13g2_fill_4 FILLER_113_1349 ();
 sg13g2_fill_8 FILLER_113_1373 ();
 sg13g2_fill_1 FILLER_113_1381 ();
 sg13g2_fill_8 FILLER_113_1408 ();
 sg13g2_fill_4 FILLER_113_1416 ();
 sg13g2_fill_4 FILLER_113_1429 ();
 sg13g2_fill_2 FILLER_113_1433 ();
 sg13g2_fill_8 FILLER_113_1445 ();
 sg13g2_fill_2 FILLER_113_1500 ();
 sg13g2_fill_1 FILLER_113_1502 ();
 sg13g2_fill_2 FILLER_113_1531 ();
 sg13g2_fill_1 FILLER_113_1533 ();
 sg13g2_fill_2 FILLER_113_1560 ();
 sg13g2_fill_4 FILLER_113_1572 ();
 sg13g2_fill_1 FILLER_113_1576 ();
 sg13g2_fill_4 FILLER_113_1588 ();
 sg13g2_fill_4 FILLER_114_0 ();
 sg13g2_fill_1 FILLER_114_4 ();
 sg13g2_fill_4 FILLER_114_31 ();
 sg13g2_fill_4 FILLER_114_61 ();
 sg13g2_fill_2 FILLER_114_65 ();
 sg13g2_fill_1 FILLER_114_67 ();
 sg13g2_fill_4 FILLER_114_73 ();
 sg13g2_fill_1 FILLER_114_77 ();
 sg13g2_fill_4 FILLER_114_90 ();
 sg13g2_fill_2 FILLER_114_94 ();
 sg13g2_fill_1 FILLER_114_96 ();
 sg13g2_fill_4 FILLER_114_133 ();
 sg13g2_fill_2 FILLER_114_137 ();
 sg13g2_fill_1 FILLER_114_191 ();
 sg13g2_fill_8 FILLER_114_196 ();
 sg13g2_fill_8 FILLER_114_204 ();
 sg13g2_fill_8 FILLER_114_212 ();
 sg13g2_fill_2 FILLER_114_220 ();
 sg13g2_fill_1 FILLER_114_222 ();
 sg13g2_fill_8 FILLER_114_260 ();
 sg13g2_fill_4 FILLER_114_346 ();
 sg13g2_fill_2 FILLER_114_350 ();
 sg13g2_fill_2 FILLER_114_365 ();
 sg13g2_fill_8 FILLER_114_401 ();
 sg13g2_fill_8 FILLER_114_409 ();
 sg13g2_fill_1 FILLER_114_417 ();
 sg13g2_fill_1 FILLER_114_431 ();
 sg13g2_fill_2 FILLER_114_464 ();
 sg13g2_fill_1 FILLER_114_466 ();
 sg13g2_fill_1 FILLER_114_481 ();
 sg13g2_fill_1 FILLER_114_486 ();
 sg13g2_fill_8 FILLER_114_495 ();
 sg13g2_fill_4 FILLER_114_511 ();
 sg13g2_fill_1 FILLER_114_515 ();
 sg13g2_fill_4 FILLER_114_524 ();
 sg13g2_fill_2 FILLER_114_554 ();
 sg13g2_fill_1 FILLER_114_572 ();
 sg13g2_fill_2 FILLER_114_594 ();
 sg13g2_fill_1 FILLER_114_596 ();
 sg13g2_fill_4 FILLER_114_633 ();
 sg13g2_fill_2 FILLER_114_637 ();
 sg13g2_fill_8 FILLER_114_649 ();
 sg13g2_fill_4 FILLER_114_657 ();
 sg13g2_fill_1 FILLER_114_661 ();
 sg13g2_fill_8 FILLER_114_672 ();
 sg13g2_fill_2 FILLER_114_680 ();
 sg13g2_fill_1 FILLER_114_682 ();
 sg13g2_fill_8 FILLER_114_689 ();
 sg13g2_fill_4 FILLER_114_697 ();
 sg13g2_fill_2 FILLER_114_701 ();
 sg13g2_fill_2 FILLER_114_721 ();
 sg13g2_fill_2 FILLER_114_749 ();
 sg13g2_fill_8 FILLER_114_759 ();
 sg13g2_fill_8 FILLER_114_767 ();
 sg13g2_fill_4 FILLER_114_784 ();
 sg13g2_fill_2 FILLER_114_788 ();
 sg13g2_fill_1 FILLER_114_790 ();
 sg13g2_fill_2 FILLER_114_800 ();
 sg13g2_fill_2 FILLER_114_811 ();
 sg13g2_fill_4 FILLER_114_817 ();
 sg13g2_fill_8 FILLER_114_869 ();
 sg13g2_fill_4 FILLER_114_877 ();
 sg13g2_fill_1 FILLER_114_881 ();
 sg13g2_fill_8 FILLER_114_886 ();
 sg13g2_fill_8 FILLER_114_894 ();
 sg13g2_fill_2 FILLER_114_902 ();
 sg13g2_fill_4 FILLER_114_908 ();
 sg13g2_fill_2 FILLER_114_912 ();
 sg13g2_fill_8 FILLER_114_925 ();
 sg13g2_fill_1 FILLER_114_933 ();
 sg13g2_fill_1 FILLER_114_976 ();
 sg13g2_fill_4 FILLER_114_981 ();
 sg13g2_fill_2 FILLER_114_985 ();
 sg13g2_fill_1 FILLER_114_987 ();
 sg13g2_fill_8 FILLER_114_1014 ();
 sg13g2_fill_8 FILLER_114_1022 ();
 sg13g2_fill_8 FILLER_114_1030 ();
 sg13g2_fill_8 FILLER_114_1043 ();
 sg13g2_fill_8 FILLER_114_1051 ();
 sg13g2_fill_4 FILLER_114_1059 ();
 sg13g2_fill_2 FILLER_114_1063 ();
 sg13g2_fill_2 FILLER_114_1068 ();
 sg13g2_fill_4 FILLER_114_1075 ();
 sg13g2_fill_2 FILLER_114_1079 ();
 sg13g2_fill_1 FILLER_114_1081 ();
 sg13g2_fill_4 FILLER_114_1097 ();
 sg13g2_fill_1 FILLER_114_1111 ();
 sg13g2_fill_2 FILLER_114_1122 ();
 sg13g2_fill_1 FILLER_114_1124 ();
 sg13g2_fill_1 FILLER_114_1130 ();
 sg13g2_fill_8 FILLER_114_1148 ();
 sg13g2_fill_2 FILLER_114_1156 ();
 sg13g2_fill_1 FILLER_114_1158 ();
 sg13g2_fill_4 FILLER_114_1164 ();
 sg13g2_fill_2 FILLER_114_1168 ();
 sg13g2_fill_8 FILLER_114_1180 ();
 sg13g2_fill_8 FILLER_114_1188 ();
 sg13g2_fill_8 FILLER_114_1196 ();
 sg13g2_fill_8 FILLER_114_1204 ();
 sg13g2_fill_8 FILLER_114_1212 ();
 sg13g2_fill_4 FILLER_114_1220 ();
 sg13g2_fill_1 FILLER_114_1224 ();
 sg13g2_fill_8 FILLER_114_1235 ();
 sg13g2_fill_1 FILLER_114_1243 ();
 sg13g2_fill_1 FILLER_114_1261 ();
 sg13g2_fill_8 FILLER_114_1266 ();
 sg13g2_fill_1 FILLER_114_1274 ();
 sg13g2_fill_1 FILLER_114_1293 ();
 sg13g2_fill_2 FILLER_114_1299 ();
 sg13g2_fill_8 FILLER_114_1312 ();
 sg13g2_fill_8 FILLER_114_1320 ();
 sg13g2_fill_8 FILLER_114_1384 ();
 sg13g2_fill_8 FILLER_114_1392 ();
 sg13g2_fill_4 FILLER_114_1410 ();
 sg13g2_fill_2 FILLER_114_1414 ();
 sg13g2_fill_4 FILLER_114_1447 ();
 sg13g2_fill_8 FILLER_114_1495 ();
 sg13g2_fill_4 FILLER_114_1503 ();
 sg13g2_fill_2 FILLER_114_1507 ();
 sg13g2_fill_8 FILLER_114_1540 ();
 sg13g2_fill_4 FILLER_114_1548 ();
 sg13g2_fill_2 FILLER_114_1552 ();
 sg13g2_fill_1 FILLER_114_1576 ();
 sg13g2_fill_4 FILLER_114_1588 ();
 sg13g2_fill_4 FILLER_115_0 ();
 sg13g2_fill_8 FILLER_115_14 ();
 sg13g2_fill_2 FILLER_115_22 ();
 sg13g2_fill_1 FILLER_115_24 ();
 sg13g2_fill_8 FILLER_115_47 ();
 sg13g2_fill_4 FILLER_115_55 ();
 sg13g2_fill_2 FILLER_115_59 ();
 sg13g2_fill_1 FILLER_115_61 ();
 sg13g2_fill_8 FILLER_115_83 ();
 sg13g2_fill_4 FILLER_115_91 ();
 sg13g2_fill_2 FILLER_115_99 ();
 sg13g2_fill_4 FILLER_115_109 ();
 sg13g2_fill_2 FILLER_115_113 ();
 sg13g2_fill_1 FILLER_115_115 ();
 sg13g2_fill_4 FILLER_115_124 ();
 sg13g2_fill_1 FILLER_115_128 ();
 sg13g2_fill_8 FILLER_115_137 ();
 sg13g2_fill_4 FILLER_115_145 ();
 sg13g2_fill_8 FILLER_115_175 ();
 sg13g2_fill_8 FILLER_115_240 ();
 sg13g2_fill_8 FILLER_115_248 ();
 sg13g2_fill_8 FILLER_115_256 ();
 sg13g2_fill_4 FILLER_115_264 ();
 sg13g2_fill_1 FILLER_115_268 ();
 sg13g2_fill_1 FILLER_115_279 ();
 sg13g2_fill_4 FILLER_115_288 ();
 sg13g2_fill_1 FILLER_115_292 ();
 sg13g2_fill_8 FILLER_115_303 ();
 sg13g2_fill_4 FILLER_115_311 ();
 sg13g2_fill_1 FILLER_115_315 ();
 sg13g2_fill_8 FILLER_115_326 ();
 sg13g2_fill_8 FILLER_115_344 ();
 sg13g2_fill_4 FILLER_115_352 ();
 sg13g2_fill_1 FILLER_115_356 ();
 sg13g2_fill_8 FILLER_115_418 ();
 sg13g2_fill_8 FILLER_115_426 ();
 sg13g2_fill_1 FILLER_115_434 ();
 sg13g2_fill_4 FILLER_115_440 ();
 sg13g2_fill_2 FILLER_115_444 ();
 sg13g2_fill_4 FILLER_115_450 ();
 sg13g2_fill_4 FILLER_115_458 ();
 sg13g2_fill_2 FILLER_115_462 ();
 sg13g2_fill_2 FILLER_115_472 ();
 sg13g2_fill_4 FILLER_115_504 ();
 sg13g2_fill_2 FILLER_115_508 ();
 sg13g2_fill_8 FILLER_115_518 ();
 sg13g2_fill_8 FILLER_115_526 ();
 sg13g2_fill_4 FILLER_115_534 ();
 sg13g2_fill_2 FILLER_115_538 ();
 sg13g2_fill_1 FILLER_115_540 ();
 sg13g2_fill_8 FILLER_115_573 ();
 sg13g2_fill_8 FILLER_115_581 ();
 sg13g2_fill_8 FILLER_115_589 ();
 sg13g2_fill_4 FILLER_115_633 ();
 sg13g2_fill_2 FILLER_115_637 ();
 sg13g2_fill_1 FILLER_115_639 ();
 sg13g2_fill_4 FILLER_115_686 ();
 sg13g2_fill_2 FILLER_115_690 ();
 sg13g2_fill_1 FILLER_115_692 ();
 sg13g2_fill_8 FILLER_115_698 ();
 sg13g2_fill_4 FILLER_115_706 ();
 sg13g2_fill_2 FILLER_115_710 ();
 sg13g2_fill_1 FILLER_115_722 ();
 sg13g2_fill_8 FILLER_115_749 ();
 sg13g2_fill_8 FILLER_115_757 ();
 sg13g2_fill_4 FILLER_115_765 ();
 sg13g2_fill_1 FILLER_115_769 ();
 sg13g2_fill_1 FILLER_115_801 ();
 sg13g2_fill_4 FILLER_115_824 ();
 sg13g2_fill_1 FILLER_115_838 ();
 sg13g2_fill_8 FILLER_115_869 ();
 sg13g2_fill_1 FILLER_115_877 ();
 sg13g2_fill_2 FILLER_115_915 ();
 sg13g2_fill_1 FILLER_115_917 ();
 sg13g2_fill_2 FILLER_115_942 ();
 sg13g2_fill_4 FILLER_115_972 ();
 sg13g2_fill_2 FILLER_115_976 ();
 sg13g2_fill_1 FILLER_115_978 ();
 sg13g2_fill_8 FILLER_115_1000 ();
 sg13g2_fill_4 FILLER_115_1008 ();
 sg13g2_fill_2 FILLER_115_1012 ();
 sg13g2_fill_2 FILLER_115_1038 ();
 sg13g2_fill_4 FILLER_115_1045 ();
 sg13g2_fill_8 FILLER_115_1056 ();
 sg13g2_fill_4 FILLER_115_1064 ();
 sg13g2_fill_2 FILLER_115_1068 ();
 sg13g2_fill_8 FILLER_115_1086 ();
 sg13g2_fill_1 FILLER_115_1094 ();
 sg13g2_fill_8 FILLER_115_1103 ();
 sg13g2_fill_4 FILLER_115_1111 ();
 sg13g2_fill_2 FILLER_115_1115 ();
 sg13g2_fill_8 FILLER_115_1122 ();
 sg13g2_fill_8 FILLER_115_1130 ();
 sg13g2_fill_8 FILLER_115_1138 ();
 sg13g2_fill_2 FILLER_115_1146 ();
 sg13g2_fill_8 FILLER_115_1182 ();
 sg13g2_fill_4 FILLER_115_1190 ();
 sg13g2_fill_2 FILLER_115_1194 ();
 sg13g2_fill_4 FILLER_115_1200 ();
 sg13g2_fill_2 FILLER_115_1204 ();
 sg13g2_fill_4 FILLER_115_1211 ();
 sg13g2_fill_1 FILLER_115_1215 ();
 sg13g2_fill_4 FILLER_115_1221 ();
 sg13g2_fill_4 FILLER_115_1238 ();
 sg13g2_fill_2 FILLER_115_1242 ();
 sg13g2_fill_4 FILLER_115_1249 ();
 sg13g2_fill_1 FILLER_115_1253 ();
 sg13g2_fill_2 FILLER_115_1260 ();
 sg13g2_fill_1 FILLER_115_1262 ();
 sg13g2_fill_2 FILLER_115_1276 ();
 sg13g2_fill_1 FILLER_115_1288 ();
 sg13g2_fill_4 FILLER_115_1294 ();
 sg13g2_fill_2 FILLER_115_1298 ();
 sg13g2_fill_4 FILLER_115_1308 ();
 sg13g2_fill_1 FILLER_115_1312 ();
 sg13g2_fill_8 FILLER_115_1349 ();
 sg13g2_fill_8 FILLER_115_1357 ();
 sg13g2_fill_2 FILLER_115_1365 ();
 sg13g2_fill_2 FILLER_115_1372 ();
 sg13g2_fill_8 FILLER_115_1378 ();
 sg13g2_fill_4 FILLER_115_1386 ();
 sg13g2_fill_2 FILLER_115_1390 ();
 sg13g2_fill_1 FILLER_115_1392 ();
 sg13g2_fill_2 FILLER_115_1399 ();
 sg13g2_fill_1 FILLER_115_1401 ();
 sg13g2_fill_2 FILLER_115_1427 ();
 sg13g2_fill_1 FILLER_115_1429 ();
 sg13g2_fill_8 FILLER_115_1439 ();
 sg13g2_fill_4 FILLER_115_1447 ();
 sg13g2_fill_1 FILLER_115_1451 ();
 sg13g2_fill_8 FILLER_115_1461 ();
 sg13g2_fill_2 FILLER_115_1469 ();
 sg13g2_fill_8 FILLER_115_1500 ();
 sg13g2_fill_4 FILLER_115_1508 ();
 sg13g2_fill_2 FILLER_115_1512 ();
 sg13g2_fill_2 FILLER_115_1519 ();
 sg13g2_fill_1 FILLER_115_1521 ();
 sg13g2_fill_8 FILLER_115_1532 ();
 sg13g2_fill_8 FILLER_115_1540 ();
 sg13g2_fill_8 FILLER_115_1548 ();
 sg13g2_fill_4 FILLER_115_1556 ();
 sg13g2_fill_4 FILLER_115_1573 ();
 sg13g2_fill_4 FILLER_115_1588 ();
 sg13g2_fill_1 FILLER_116_26 ();
 sg13g2_fill_4 FILLER_116_42 ();
 sg13g2_fill_4 FILLER_116_59 ();
 sg13g2_fill_2 FILLER_116_95 ();
 sg13g2_fill_1 FILLER_116_97 ();
 sg13g2_fill_1 FILLER_116_111 ();
 sg13g2_fill_8 FILLER_116_122 ();
 sg13g2_fill_2 FILLER_116_130 ();
 sg13g2_fill_1 FILLER_116_132 ();
 sg13g2_fill_4 FILLER_116_143 ();
 sg13g2_fill_2 FILLER_116_157 ();
 sg13g2_fill_1 FILLER_116_159 ();
 sg13g2_fill_4 FILLER_116_168 ();
 sg13g2_fill_1 FILLER_116_172 ();
 sg13g2_fill_8 FILLER_116_194 ();
 sg13g2_fill_8 FILLER_116_202 ();
 sg13g2_fill_2 FILLER_116_210 ();
 sg13g2_fill_8 FILLER_116_233 ();
 sg13g2_fill_2 FILLER_116_241 ();
 sg13g2_fill_8 FILLER_116_287 ();
 sg13g2_fill_8 FILLER_116_357 ();
 sg13g2_fill_8 FILLER_116_365 ();
 sg13g2_fill_4 FILLER_116_373 ();
 sg13g2_fill_8 FILLER_116_439 ();
 sg13g2_fill_8 FILLER_116_447 ();
 sg13g2_fill_1 FILLER_116_455 ();
 sg13g2_fill_4 FILLER_116_464 ();
 sg13g2_fill_2 FILLER_116_468 ();
 sg13g2_fill_8 FILLER_116_478 ();
 sg13g2_fill_2 FILLER_116_486 ();
 sg13g2_fill_1 FILLER_116_488 ();
 sg13g2_fill_8 FILLER_116_525 ();
 sg13g2_fill_2 FILLER_116_533 ();
 sg13g2_fill_2 FILLER_116_545 ();
 sg13g2_fill_1 FILLER_116_547 ();
 sg13g2_fill_2 FILLER_116_554 ();
 sg13g2_fill_4 FILLER_116_592 ();
 sg13g2_fill_2 FILLER_116_596 ();
 sg13g2_fill_8 FILLER_116_608 ();
 sg13g2_fill_8 FILLER_116_616 ();
 sg13g2_fill_8 FILLER_116_624 ();
 sg13g2_fill_8 FILLER_116_632 ();
 sg13g2_fill_8 FILLER_116_640 ();
 sg13g2_fill_8 FILLER_116_648 ();
 sg13g2_fill_1 FILLER_116_656 ();
 sg13g2_fill_8 FILLER_116_667 ();
 sg13g2_fill_2 FILLER_116_711 ();
 sg13g2_fill_2 FILLER_116_723 ();
 sg13g2_fill_4 FILLER_116_751 ();
 sg13g2_fill_8 FILLER_116_768 ();
 sg13g2_fill_1 FILLER_116_776 ();
 sg13g2_fill_8 FILLER_116_787 ();
 sg13g2_fill_8 FILLER_116_795 ();
 sg13g2_fill_8 FILLER_116_803 ();
 sg13g2_fill_8 FILLER_116_811 ();
 sg13g2_fill_2 FILLER_116_819 ();
 sg13g2_fill_8 FILLER_116_833 ();
 sg13g2_fill_2 FILLER_116_841 ();
 sg13g2_fill_1 FILLER_116_843 ();
 sg13g2_fill_4 FILLER_116_850 ();
 sg13g2_fill_2 FILLER_116_854 ();
 sg13g2_fill_1 FILLER_116_856 ();
 sg13g2_fill_1 FILLER_116_926 ();
 sg13g2_fill_1 FILLER_116_953 ();
 sg13g2_fill_2 FILLER_116_958 ();
 sg13g2_fill_4 FILLER_116_970 ();
 sg13g2_fill_2 FILLER_116_978 ();
 sg13g2_fill_2 FILLER_116_989 ();
 sg13g2_fill_1 FILLER_116_991 ();
 sg13g2_fill_2 FILLER_116_1001 ();
 sg13g2_fill_2 FILLER_116_1010 ();
 sg13g2_fill_1 FILLER_116_1012 ();
 sg13g2_fill_2 FILLER_116_1039 ();
 sg13g2_fill_4 FILLER_116_1058 ();
 sg13g2_fill_2 FILLER_116_1062 ();
 sg13g2_fill_1 FILLER_116_1064 ();
 sg13g2_fill_8 FILLER_116_1081 ();
 sg13g2_fill_1 FILLER_116_1089 ();
 sg13g2_fill_4 FILLER_116_1095 ();
 sg13g2_fill_2 FILLER_116_1099 ();
 sg13g2_fill_1 FILLER_116_1109 ();
 sg13g2_fill_2 FILLER_116_1122 ();
 sg13g2_fill_8 FILLER_116_1134 ();
 sg13g2_fill_2 FILLER_116_1142 ();
 sg13g2_fill_1 FILLER_116_1144 ();
 sg13g2_fill_4 FILLER_116_1148 ();
 sg13g2_fill_4 FILLER_116_1175 ();
 sg13g2_fill_2 FILLER_116_1179 ();
 sg13g2_fill_1 FILLER_116_1181 ();
 sg13g2_fill_4 FILLER_116_1244 ();
 sg13g2_fill_8 FILLER_116_1252 ();
 sg13g2_fill_8 FILLER_116_1260 ();
 sg13g2_fill_8 FILLER_116_1268 ();
 sg13g2_fill_8 FILLER_116_1276 ();
 sg13g2_fill_4 FILLER_116_1284 ();
 sg13g2_fill_2 FILLER_116_1288 ();
 sg13g2_fill_1 FILLER_116_1290 ();
 sg13g2_fill_8 FILLER_116_1317 ();
 sg13g2_fill_2 FILLER_116_1325 ();
 sg13g2_fill_8 FILLER_116_1330 ();
 sg13g2_fill_8 FILLER_116_1338 ();
 sg13g2_fill_4 FILLER_116_1346 ();
 sg13g2_fill_1 FILLER_116_1350 ();
 sg13g2_fill_4 FILLER_116_1359 ();
 sg13g2_fill_1 FILLER_116_1363 ();
 sg13g2_fill_2 FILLER_116_1417 ();
 sg13g2_fill_1 FILLER_116_1419 ();
 sg13g2_fill_2 FILLER_116_1429 ();
 sg13g2_fill_8 FILLER_116_1439 ();
 sg13g2_fill_2 FILLER_116_1447 ();
 sg13g2_fill_1 FILLER_116_1449 ();
 sg13g2_fill_4 FILLER_116_1462 ();
 sg13g2_fill_4 FILLER_116_1517 ();
 sg13g2_fill_8 FILLER_116_1553 ();
 sg13g2_fill_2 FILLER_116_1561 ();
 sg13g2_fill_4 FILLER_116_1568 ();
 sg13g2_fill_2 FILLER_116_1572 ();
 sg13g2_fill_1 FILLER_116_1574 ();
 sg13g2_fill_8 FILLER_116_1580 ();
 sg13g2_fill_4 FILLER_116_1588 ();
 sg13g2_fill_8 FILLER_117_0 ();
 sg13g2_fill_8 FILLER_117_8 ();
 sg13g2_fill_2 FILLER_117_16 ();
 sg13g2_fill_1 FILLER_117_18 ();
 sg13g2_fill_2 FILLER_117_47 ();
 sg13g2_fill_2 FILLER_117_54 ();
 sg13g2_fill_1 FILLER_117_56 ();
 sg13g2_fill_8 FILLER_117_63 ();
 sg13g2_fill_2 FILLER_117_71 ();
 sg13g2_fill_8 FILLER_117_76 ();
 sg13g2_fill_4 FILLER_117_84 ();
 sg13g2_fill_2 FILLER_117_98 ();
 sg13g2_fill_2 FILLER_117_116 ();
 sg13g2_fill_8 FILLER_117_167 ();
 sg13g2_fill_8 FILLER_117_196 ();
 sg13g2_fill_8 FILLER_117_204 ();
 sg13g2_fill_8 FILLER_117_212 ();
 sg13g2_fill_2 FILLER_117_220 ();
 sg13g2_fill_4 FILLER_117_258 ();
 sg13g2_fill_1 FILLER_117_287 ();
 sg13g2_fill_8 FILLER_117_296 ();
 sg13g2_fill_8 FILLER_117_304 ();
 sg13g2_fill_8 FILLER_117_312 ();
 sg13g2_fill_8 FILLER_117_320 ();
 sg13g2_fill_8 FILLER_117_328 ();
 sg13g2_fill_8 FILLER_117_336 ();
 sg13g2_fill_8 FILLER_117_344 ();
 sg13g2_fill_4 FILLER_117_352 ();
 sg13g2_fill_2 FILLER_117_356 ();
 sg13g2_fill_8 FILLER_117_384 ();
 sg13g2_fill_8 FILLER_117_392 ();
 sg13g2_fill_8 FILLER_117_400 ();
 sg13g2_fill_8 FILLER_117_408 ();
 sg13g2_fill_2 FILLER_117_416 ();
 sg13g2_fill_1 FILLER_117_418 ();
 sg13g2_fill_4 FILLER_117_424 ();
 sg13g2_fill_8 FILLER_117_446 ();
 sg13g2_fill_4 FILLER_117_454 ();
 sg13g2_fill_2 FILLER_117_468 ();
 sg13g2_fill_1 FILLER_117_470 ();
 sg13g2_fill_4 FILLER_117_475 ();
 sg13g2_fill_2 FILLER_117_479 ();
 sg13g2_fill_1 FILLER_117_481 ();
 sg13g2_fill_8 FILLER_117_490 ();
 sg13g2_fill_8 FILLER_117_498 ();
 sg13g2_fill_8 FILLER_117_506 ();
 sg13g2_fill_4 FILLER_117_514 ();
 sg13g2_fill_1 FILLER_117_518 ();
 sg13g2_fill_1 FILLER_117_545 ();
 sg13g2_fill_8 FILLER_117_563 ();
 sg13g2_fill_8 FILLER_117_571 ();
 sg13g2_fill_8 FILLER_117_579 ();
 sg13g2_fill_4 FILLER_117_587 ();
 sg13g2_fill_8 FILLER_117_599 ();
 sg13g2_fill_8 FILLER_117_607 ();
 sg13g2_fill_1 FILLER_117_615 ();
 sg13g2_fill_4 FILLER_117_624 ();
 sg13g2_fill_2 FILLER_117_628 ();
 sg13g2_fill_4 FILLER_117_655 ();
 sg13g2_fill_1 FILLER_117_659 ();
 sg13g2_fill_4 FILLER_117_670 ();
 sg13g2_fill_2 FILLER_117_674 ();
 sg13g2_fill_1 FILLER_117_676 ();
 sg13g2_fill_8 FILLER_117_703 ();
 sg13g2_fill_8 FILLER_117_711 ();
 sg13g2_fill_8 FILLER_117_719 ();
 sg13g2_fill_8 FILLER_117_727 ();
 sg13g2_fill_8 FILLER_117_735 ();
 sg13g2_fill_8 FILLER_117_743 ();
 sg13g2_fill_4 FILLER_117_751 ();
 sg13g2_fill_2 FILLER_117_755 ();
 sg13g2_fill_1 FILLER_117_757 ();
 sg13g2_fill_8 FILLER_117_766 ();
 sg13g2_fill_8 FILLER_117_774 ();
 sg13g2_fill_8 FILLER_117_812 ();
 sg13g2_fill_4 FILLER_117_820 ();
 sg13g2_fill_2 FILLER_117_824 ();
 sg13g2_fill_8 FILLER_117_834 ();
 sg13g2_fill_8 FILLER_117_842 ();
 sg13g2_fill_8 FILLER_117_850 ();
 sg13g2_fill_8 FILLER_117_858 ();
 sg13g2_fill_8 FILLER_117_866 ();
 sg13g2_fill_8 FILLER_117_874 ();
 sg13g2_fill_2 FILLER_117_890 ();
 sg13g2_fill_1 FILLER_117_892 ();
 sg13g2_fill_2 FILLER_117_908 ();
 sg13g2_fill_8 FILLER_117_915 ();
 sg13g2_fill_4 FILLER_117_923 ();
 sg13g2_fill_1 FILLER_117_927 ();
 sg13g2_fill_2 FILLER_117_934 ();
 sg13g2_fill_2 FILLER_117_945 ();
 sg13g2_fill_8 FILLER_117_970 ();
 sg13g2_fill_4 FILLER_117_978 ();
 sg13g2_fill_8 FILLER_117_996 ();
 sg13g2_fill_8 FILLER_117_1004 ();
 sg13g2_fill_4 FILLER_117_1012 ();
 sg13g2_fill_8 FILLER_117_1033 ();
 sg13g2_fill_4 FILLER_117_1041 ();
 sg13g2_fill_2 FILLER_117_1045 ();
 sg13g2_fill_4 FILLER_117_1055 ();
 sg13g2_fill_1 FILLER_117_1059 ();
 sg13g2_fill_8 FILLER_117_1065 ();
 sg13g2_fill_4 FILLER_117_1073 ();
 sg13g2_fill_1 FILLER_117_1098 ();
 sg13g2_fill_8 FILLER_117_1104 ();
 sg13g2_fill_4 FILLER_117_1112 ();
 sg13g2_fill_1 FILLER_117_1116 ();
 sg13g2_fill_2 FILLER_117_1127 ();
 sg13g2_fill_1 FILLER_117_1129 ();
 sg13g2_fill_2 FILLER_117_1134 ();
 sg13g2_fill_8 FILLER_117_1149 ();
 sg13g2_fill_8 FILLER_117_1157 ();
 sg13g2_fill_8 FILLER_117_1165 ();
 sg13g2_fill_2 FILLER_117_1173 ();
 sg13g2_fill_1 FILLER_117_1175 ();
 sg13g2_fill_4 FILLER_117_1193 ();
 sg13g2_fill_2 FILLER_117_1197 ();
 sg13g2_fill_1 FILLER_117_1199 ();
 sg13g2_fill_2 FILLER_117_1210 ();
 sg13g2_fill_2 FILLER_117_1237 ();
 sg13g2_fill_1 FILLER_117_1239 ();
 sg13g2_fill_4 FILLER_117_1269 ();
 sg13g2_fill_4 FILLER_117_1283 ();
 sg13g2_fill_1 FILLER_117_1287 ();
 sg13g2_fill_4 FILLER_117_1301 ();
 sg13g2_fill_1 FILLER_117_1305 ();
 sg13g2_fill_4 FILLER_117_1340 ();
 sg13g2_fill_2 FILLER_117_1344 ();
 sg13g2_fill_8 FILLER_117_1367 ();
 sg13g2_fill_8 FILLER_117_1375 ();
 sg13g2_fill_8 FILLER_117_1383 ();
 sg13g2_fill_2 FILLER_117_1391 ();
 sg13g2_fill_1 FILLER_117_1393 ();
 sg13g2_fill_4 FILLER_117_1405 ();
 sg13g2_fill_1 FILLER_117_1409 ();
 sg13g2_fill_1 FILLER_117_1415 ();
 sg13g2_fill_8 FILLER_117_1452 ();
 sg13g2_fill_4 FILLER_117_1460 ();
 sg13g2_fill_2 FILLER_117_1464 ();
 sg13g2_fill_2 FILLER_117_1476 ();
 sg13g2_fill_8 FILLER_117_1509 ();
 sg13g2_fill_1 FILLER_117_1517 ();
 sg13g2_fill_8 FILLER_117_1536 ();
 sg13g2_fill_8 FILLER_117_1544 ();
 sg13g2_fill_4 FILLER_117_1552 ();
 sg13g2_fill_2 FILLER_117_1589 ();
 sg13g2_fill_1 FILLER_117_1591 ();
 sg13g2_fill_4 FILLER_118_0 ();
 sg13g2_fill_1 FILLER_118_4 ();
 sg13g2_fill_1 FILLER_118_13 ();
 sg13g2_fill_2 FILLER_118_20 ();
 sg13g2_fill_8 FILLER_118_36 ();
 sg13g2_fill_8 FILLER_118_44 ();
 sg13g2_fill_8 FILLER_118_52 ();
 sg13g2_fill_4 FILLER_118_60 ();
 sg13g2_fill_1 FILLER_118_64 ();
 sg13g2_fill_1 FILLER_118_71 ();
 sg13g2_fill_4 FILLER_118_78 ();
 sg13g2_fill_1 FILLER_118_88 ();
 sg13g2_fill_8 FILLER_118_94 ();
 sg13g2_fill_8 FILLER_118_102 ();
 sg13g2_fill_8 FILLER_118_110 ();
 sg13g2_fill_2 FILLER_118_118 ();
 sg13g2_fill_8 FILLER_118_126 ();
 sg13g2_fill_4 FILLER_118_134 ();
 sg13g2_fill_1 FILLER_118_138 ();
 sg13g2_fill_1 FILLER_118_158 ();
 sg13g2_fill_2 FILLER_118_185 ();
 sg13g2_fill_1 FILLER_118_187 ();
 sg13g2_fill_2 FILLER_118_206 ();
 sg13g2_fill_1 FILLER_118_208 ();
 sg13g2_fill_8 FILLER_118_219 ();
 sg13g2_fill_8 FILLER_118_227 ();
 sg13g2_fill_4 FILLER_118_235 ();
 sg13g2_fill_8 FILLER_118_244 ();
 sg13g2_fill_2 FILLER_118_252 ();
 sg13g2_fill_2 FILLER_118_275 ();
 sg13g2_fill_1 FILLER_118_277 ();
 sg13g2_fill_4 FILLER_118_294 ();
 sg13g2_fill_4 FILLER_118_314 ();
 sg13g2_fill_1 FILLER_118_318 ();
 sg13g2_fill_2 FILLER_118_327 ();
 sg13g2_fill_1 FILLER_118_337 ();
 sg13g2_fill_4 FILLER_118_346 ();
 sg13g2_fill_2 FILLER_118_364 ();
 sg13g2_fill_2 FILLER_118_371 ();
 sg13g2_fill_1 FILLER_118_373 ();
 sg13g2_fill_4 FILLER_118_383 ();
 sg13g2_fill_2 FILLER_118_387 ();
 sg13g2_fill_1 FILLER_118_389 ();
 sg13g2_fill_8 FILLER_118_400 ();
 sg13g2_fill_2 FILLER_118_408 ();
 sg13g2_fill_4 FILLER_118_425 ();
 sg13g2_fill_2 FILLER_118_429 ();
 sg13g2_fill_1 FILLER_118_431 ();
 sg13g2_fill_2 FILLER_118_447 ();
 sg13g2_fill_1 FILLER_118_449 ();
 sg13g2_fill_4 FILLER_118_470 ();
 sg13g2_fill_2 FILLER_118_478 ();
 sg13g2_fill_4 FILLER_118_488 ();
 sg13g2_fill_8 FILLER_118_500 ();
 sg13g2_fill_4 FILLER_118_518 ();
 sg13g2_fill_2 FILLER_118_522 ();
 sg13g2_fill_1 FILLER_118_572 ();
 sg13g2_fill_8 FILLER_118_583 ();
 sg13g2_fill_1 FILLER_118_591 ();
 sg13g2_fill_8 FILLER_118_602 ();
 sg13g2_fill_8 FILLER_118_610 ();
 sg13g2_fill_1 FILLER_118_618 ();
 sg13g2_fill_2 FILLER_118_629 ();
 sg13g2_fill_2 FILLER_118_676 ();
 sg13g2_fill_1 FILLER_118_678 ();
 sg13g2_fill_1 FILLER_118_696 ();
 sg13g2_fill_2 FILLER_118_707 ();
 sg13g2_fill_1 FILLER_118_709 ();
 sg13g2_fill_8 FILLER_118_720 ();
 sg13g2_fill_8 FILLER_118_728 ();
 sg13g2_fill_8 FILLER_118_736 ();
 sg13g2_fill_8 FILLER_118_744 ();
 sg13g2_fill_8 FILLER_118_777 ();
 sg13g2_fill_8 FILLER_118_785 ();
 sg13g2_fill_8 FILLER_118_793 ();
 sg13g2_fill_8 FILLER_118_815 ();
 sg13g2_fill_4 FILLER_118_823 ();
 sg13g2_fill_2 FILLER_118_827 ();
 sg13g2_fill_1 FILLER_118_829 ();
 sg13g2_fill_8 FILLER_118_870 ();
 sg13g2_fill_8 FILLER_118_878 ();
 sg13g2_fill_8 FILLER_118_886 ();
 sg13g2_fill_8 FILLER_118_894 ();
 sg13g2_fill_8 FILLER_118_902 ();
 sg13g2_fill_1 FILLER_118_910 ();
 sg13g2_fill_2 FILLER_118_926 ();
 sg13g2_fill_1 FILLER_118_928 ();
 sg13g2_fill_1 FILLER_118_966 ();
 sg13g2_fill_2 FILLER_118_982 ();
 sg13g2_fill_8 FILLER_118_1004 ();
 sg13g2_fill_8 FILLER_118_1012 ();
 sg13g2_fill_8 FILLER_118_1020 ();
 sg13g2_fill_8 FILLER_118_1028 ();
 sg13g2_fill_2 FILLER_118_1036 ();
 sg13g2_fill_4 FILLER_118_1047 ();
 sg13g2_fill_2 FILLER_118_1051 ();
 sg13g2_fill_4 FILLER_118_1071 ();
 sg13g2_fill_2 FILLER_118_1075 ();
 sg13g2_fill_2 FILLER_118_1082 ();
 sg13g2_fill_2 FILLER_118_1096 ();
 sg13g2_fill_1 FILLER_118_1098 ();
 sg13g2_fill_2 FILLER_118_1122 ();
 sg13g2_fill_1 FILLER_118_1124 ();
 sg13g2_fill_4 FILLER_118_1131 ();
 sg13g2_fill_2 FILLER_118_1135 ();
 sg13g2_fill_4 FILLER_118_1155 ();
 sg13g2_fill_2 FILLER_118_1159 ();
 sg13g2_fill_4 FILLER_118_1174 ();
 sg13g2_fill_4 FILLER_118_1182 ();
 sg13g2_fill_2 FILLER_118_1194 ();
 sg13g2_fill_8 FILLER_118_1201 ();
 sg13g2_fill_4 FILLER_118_1209 ();
 sg13g2_fill_8 FILLER_118_1291 ();
 sg13g2_fill_2 FILLER_118_1311 ();
 sg13g2_fill_1 FILLER_118_1343 ();
 sg13g2_fill_8 FILLER_118_1348 ();
 sg13g2_fill_8 FILLER_118_1356 ();
 sg13g2_fill_4 FILLER_118_1370 ();
 sg13g2_fill_2 FILLER_118_1374 ();
 sg13g2_fill_8 FILLER_118_1393 ();
 sg13g2_fill_2 FILLER_118_1401 ();
 sg13g2_fill_1 FILLER_118_1403 ();
 sg13g2_fill_2 FILLER_118_1411 ();
 sg13g2_fill_1 FILLER_118_1413 ();
 sg13g2_fill_1 FILLER_118_1470 ();
 sg13g2_fill_4 FILLER_118_1476 ();
 sg13g2_fill_8 FILLER_118_1484 ();
 sg13g2_fill_8 FILLER_118_1492 ();
 sg13g2_fill_8 FILLER_118_1500 ();
 sg13g2_fill_8 FILLER_118_1508 ();
 sg13g2_fill_8 FILLER_118_1516 ();
 sg13g2_fill_4 FILLER_118_1524 ();
 sg13g2_fill_2 FILLER_118_1551 ();
 sg13g2_fill_2 FILLER_118_1575 ();
 sg13g2_fill_1 FILLER_118_1577 ();
 sg13g2_fill_2 FILLER_118_1589 ();
 sg13g2_fill_1 FILLER_118_1591 ();
 sg13g2_fill_8 FILLER_119_0 ();
 sg13g2_fill_4 FILLER_119_8 ();
 sg13g2_fill_4 FILLER_119_38 ();
 sg13g2_fill_8 FILLER_119_47 ();
 sg13g2_fill_8 FILLER_119_87 ();
 sg13g2_fill_2 FILLER_119_95 ();
 sg13g2_fill_2 FILLER_119_102 ();
 sg13g2_fill_1 FILLER_119_117 ();
 sg13g2_fill_8 FILLER_119_122 ();
 sg13g2_fill_4 FILLER_119_130 ();
 sg13g2_fill_2 FILLER_119_134 ();
 sg13g2_fill_1 FILLER_119_136 ();
 sg13g2_fill_2 FILLER_119_147 ();
 sg13g2_fill_8 FILLER_119_184 ();
 sg13g2_fill_4 FILLER_119_223 ();
 sg13g2_fill_8 FILLER_119_235 ();
 sg13g2_fill_4 FILLER_119_243 ();
 sg13g2_fill_1 FILLER_119_247 ();
 sg13g2_fill_4 FILLER_119_272 ();
 sg13g2_fill_2 FILLER_119_276 ();
 sg13g2_fill_1 FILLER_119_278 ();
 sg13g2_fill_2 FILLER_119_295 ();
 sg13g2_fill_1 FILLER_119_297 ();
 sg13g2_fill_8 FILLER_119_306 ();
 sg13g2_fill_4 FILLER_119_314 ();
 sg13g2_fill_1 FILLER_119_318 ();
 sg13g2_fill_8 FILLER_119_327 ();
 sg13g2_fill_4 FILLER_119_348 ();
 sg13g2_fill_2 FILLER_119_352 ();
 sg13g2_fill_2 FILLER_119_365 ();
 sg13g2_fill_4 FILLER_119_384 ();
 sg13g2_fill_2 FILLER_119_388 ();
 sg13g2_fill_4 FILLER_119_416 ();
 sg13g2_fill_2 FILLER_119_420 ();
 sg13g2_fill_8 FILLER_119_433 ();
 sg13g2_fill_8 FILLER_119_441 ();
 sg13g2_fill_2 FILLER_119_449 ();
 sg13g2_fill_4 FILLER_119_470 ();
 sg13g2_fill_4 FILLER_119_494 ();
 sg13g2_fill_2 FILLER_119_498 ();
 sg13g2_fill_1 FILLER_119_500 ();
 sg13g2_fill_2 FILLER_119_517 ();
 sg13g2_fill_1 FILLER_119_519 ();
 sg13g2_fill_4 FILLER_119_530 ();
 sg13g2_fill_1 FILLER_119_534 ();
 sg13g2_fill_2 FILLER_119_555 ();
 sg13g2_fill_1 FILLER_119_557 ();
 sg13g2_fill_2 FILLER_119_584 ();
 sg13g2_fill_1 FILLER_119_586 ();
 sg13g2_fill_1 FILLER_119_593 ();
 sg13g2_fill_8 FILLER_119_636 ();
 sg13g2_fill_8 FILLER_119_644 ();
 sg13g2_fill_2 FILLER_119_652 ();
 sg13g2_fill_2 FILLER_119_697 ();
 sg13g2_fill_8 FILLER_119_751 ();
 sg13g2_fill_1 FILLER_119_767 ();
 sg13g2_fill_1 FILLER_119_798 ();
 sg13g2_fill_8 FILLER_119_838 ();
 sg13g2_fill_8 FILLER_119_846 ();
 sg13g2_fill_8 FILLER_119_854 ();
 sg13g2_fill_4 FILLER_119_862 ();
 sg13g2_fill_2 FILLER_119_879 ();
 sg13g2_fill_1 FILLER_119_881 ();
 sg13g2_fill_2 FILLER_119_892 ();
 sg13g2_fill_1 FILLER_119_894 ();
 sg13g2_fill_8 FILLER_119_906 ();
 sg13g2_fill_2 FILLER_119_914 ();
 sg13g2_fill_8 FILLER_119_925 ();
 sg13g2_fill_8 FILLER_119_933 ();
 sg13g2_fill_2 FILLER_119_941 ();
 sg13g2_fill_1 FILLER_119_943 ();
 sg13g2_fill_2 FILLER_119_957 ();
 sg13g2_fill_2 FILLER_119_966 ();
 sg13g2_fill_8 FILLER_119_979 ();
 sg13g2_fill_8 FILLER_119_987 ();
 sg13g2_fill_2 FILLER_119_995 ();
 sg13g2_fill_4 FILLER_119_1002 ();
 sg13g2_fill_2 FILLER_119_1006 ();
 sg13g2_fill_1 FILLER_119_1008 ();
 sg13g2_fill_8 FILLER_119_1020 ();
 sg13g2_fill_2 FILLER_119_1028 ();
 sg13g2_fill_1 FILLER_119_1030 ();
 sg13g2_fill_8 FILLER_119_1038 ();
 sg13g2_fill_2 FILLER_119_1046 ();
 sg13g2_fill_1 FILLER_119_1048 ();
 sg13g2_fill_8 FILLER_119_1057 ();
 sg13g2_fill_4 FILLER_119_1065 ();
 sg13g2_fill_2 FILLER_119_1069 ();
 sg13g2_fill_4 FILLER_119_1078 ();
 sg13g2_fill_2 FILLER_119_1087 ();
 sg13g2_fill_1 FILLER_119_1089 ();
 sg13g2_fill_4 FILLER_119_1099 ();
 sg13g2_fill_1 FILLER_119_1103 ();
 sg13g2_fill_2 FILLER_119_1109 ();
 sg13g2_fill_4 FILLER_119_1132 ();
 sg13g2_fill_1 FILLER_119_1136 ();
 sg13g2_fill_2 FILLER_119_1141 ();
 sg13g2_fill_1 FILLER_119_1143 ();
 sg13g2_fill_8 FILLER_119_1148 ();
 sg13g2_fill_2 FILLER_119_1181 ();
 sg13g2_fill_1 FILLER_119_1183 ();
 sg13g2_fill_4 FILLER_119_1189 ();
 sg13g2_fill_1 FILLER_119_1219 ();
 sg13g2_fill_8 FILLER_119_1229 ();
 sg13g2_fill_8 FILLER_119_1237 ();
 sg13g2_fill_2 FILLER_119_1245 ();
 sg13g2_fill_8 FILLER_119_1251 ();
 sg13g2_fill_1 FILLER_119_1259 ();
 sg13g2_fill_2 FILLER_119_1304 ();
 sg13g2_fill_2 FILLER_119_1317 ();
 sg13g2_fill_1 FILLER_119_1324 ();
 sg13g2_fill_4 FILLER_119_1351 ();
 sg13g2_fill_1 FILLER_119_1355 ();
 sg13g2_fill_4 FILLER_119_1364 ();
 sg13g2_fill_1 FILLER_119_1381 ();
 sg13g2_fill_2 FILLER_119_1400 ();
 sg13g2_fill_1 FILLER_119_1402 ();
 sg13g2_fill_1 FILLER_119_1433 ();
 sg13g2_fill_2 FILLER_119_1448 ();
 sg13g2_fill_1 FILLER_119_1450 ();
 sg13g2_fill_2 FILLER_119_1460 ();
 sg13g2_fill_1 FILLER_119_1462 ();
 sg13g2_fill_2 FILLER_119_1468 ();
 sg13g2_fill_1 FILLER_119_1470 ();
 sg13g2_fill_1 FILLER_119_1523 ();
 sg13g2_fill_8 FILLER_119_1555 ();
 sg13g2_fill_4 FILLER_119_1563 ();
 sg13g2_fill_1 FILLER_119_1567 ();
 sg13g2_fill_4 FILLER_119_1587 ();
 sg13g2_fill_1 FILLER_119_1591 ();
 sg13g2_fill_8 FILLER_120_0 ();
 sg13g2_fill_8 FILLER_120_8 ();
 sg13g2_fill_4 FILLER_120_16 ();
 sg13g2_fill_1 FILLER_120_20 ();
 sg13g2_fill_2 FILLER_120_24 ();
 sg13g2_fill_8 FILLER_120_42 ();
 sg13g2_fill_8 FILLER_120_50 ();
 sg13g2_fill_1 FILLER_120_58 ();
 sg13g2_fill_1 FILLER_120_68 ();
 sg13g2_fill_4 FILLER_120_100 ();
 sg13g2_fill_2 FILLER_120_112 ();
 sg13g2_fill_1 FILLER_120_114 ();
 sg13g2_fill_4 FILLER_120_155 ();
 sg13g2_fill_2 FILLER_120_159 ();
 sg13g2_fill_8 FILLER_120_187 ();
 sg13g2_fill_1 FILLER_120_195 ();
 sg13g2_fill_8 FILLER_120_204 ();
 sg13g2_fill_2 FILLER_120_212 ();
 sg13g2_fill_2 FILLER_120_240 ();
 sg13g2_fill_8 FILLER_120_252 ();
 sg13g2_fill_8 FILLER_120_260 ();
 sg13g2_fill_8 FILLER_120_268 ();
 sg13g2_fill_8 FILLER_120_276 ();
 sg13g2_fill_4 FILLER_120_284 ();
 sg13g2_fill_2 FILLER_120_288 ();
 sg13g2_fill_4 FILLER_120_298 ();
 sg13g2_fill_1 FILLER_120_302 ();
 sg13g2_fill_4 FILLER_120_311 ();
 sg13g2_fill_4 FILLER_120_323 ();
 sg13g2_fill_2 FILLER_120_327 ();
 sg13g2_fill_1 FILLER_120_329 ();
 sg13g2_fill_8 FILLER_120_338 ();
 sg13g2_fill_4 FILLER_120_346 ();
 sg13g2_fill_1 FILLER_120_350 ();
 sg13g2_fill_2 FILLER_120_362 ();
 sg13g2_fill_1 FILLER_120_364 ();
 sg13g2_fill_8 FILLER_120_378 ();
 sg13g2_fill_8 FILLER_120_386 ();
 sg13g2_fill_8 FILLER_120_394 ();
 sg13g2_fill_4 FILLER_120_402 ();
 sg13g2_fill_1 FILLER_120_406 ();
 sg13g2_fill_4 FILLER_120_418 ();
 sg13g2_fill_2 FILLER_120_430 ();
 sg13g2_fill_1 FILLER_120_432 ();
 sg13g2_fill_1 FILLER_120_457 ();
 sg13g2_fill_1 FILLER_120_464 ();
 sg13g2_fill_2 FILLER_120_470 ();
 sg13g2_fill_8 FILLER_120_485 ();
 sg13g2_fill_8 FILLER_120_507 ();
 sg13g2_fill_8 FILLER_120_515 ();
 sg13g2_fill_8 FILLER_120_523 ();
 sg13g2_fill_4 FILLER_120_531 ();
 sg13g2_fill_2 FILLER_120_535 ();
 sg13g2_fill_1 FILLER_120_537 ();
 sg13g2_fill_1 FILLER_120_543 ();
 sg13g2_fill_8 FILLER_120_548 ();
 sg13g2_fill_8 FILLER_120_556 ();
 sg13g2_fill_8 FILLER_120_564 ();
 sg13g2_fill_4 FILLER_120_588 ();
 sg13g2_fill_2 FILLER_120_592 ();
 sg13g2_fill_8 FILLER_120_630 ();
 sg13g2_fill_2 FILLER_120_656 ();
 sg13g2_fill_8 FILLER_120_675 ();
 sg13g2_fill_8 FILLER_120_683 ();
 sg13g2_fill_8 FILLER_120_691 ();
 sg13g2_fill_8 FILLER_120_699 ();
 sg13g2_fill_4 FILLER_120_707 ();
 sg13g2_fill_4 FILLER_120_721 ();
 sg13g2_fill_8 FILLER_120_751 ();
 sg13g2_fill_4 FILLER_120_759 ();
 sg13g2_fill_2 FILLER_120_763 ();
 sg13g2_fill_1 FILLER_120_765 ();
 sg13g2_fill_2 FILLER_120_771 ();
 sg13g2_fill_8 FILLER_120_776 ();
 sg13g2_fill_8 FILLER_120_784 ();
 sg13g2_fill_8 FILLER_120_792 ();
 sg13g2_fill_8 FILLER_120_800 ();
 sg13g2_fill_1 FILLER_120_808 ();
 sg13g2_fill_8 FILLER_120_814 ();
 sg13g2_fill_2 FILLER_120_822 ();
 sg13g2_fill_1 FILLER_120_824 ();
 sg13g2_fill_4 FILLER_120_869 ();
 sg13g2_fill_8 FILLER_120_883 ();
 sg13g2_fill_4 FILLER_120_891 ();
 sg13g2_fill_8 FILLER_120_913 ();
 sg13g2_fill_2 FILLER_120_921 ();
 sg13g2_fill_8 FILLER_120_929 ();
 sg13g2_fill_2 FILLER_120_937 ();
 sg13g2_fill_1 FILLER_120_939 ();
 sg13g2_fill_1 FILLER_120_966 ();
 sg13g2_fill_8 FILLER_120_972 ();
 sg13g2_fill_8 FILLER_120_980 ();
 sg13g2_fill_1 FILLER_120_988 ();
 sg13g2_fill_2 FILLER_120_1001 ();
 sg13g2_fill_1 FILLER_120_1003 ();
 sg13g2_fill_2 FILLER_120_1022 ();
 sg13g2_fill_2 FILLER_120_1039 ();
 sg13g2_fill_1 FILLER_120_1041 ();
 sg13g2_fill_8 FILLER_120_1066 ();
 sg13g2_fill_8 FILLER_120_1090 ();
 sg13g2_fill_8 FILLER_120_1098 ();
 sg13g2_fill_4 FILLER_120_1106 ();
 sg13g2_fill_2 FILLER_120_1110 ();
 sg13g2_fill_1 FILLER_120_1112 ();
 sg13g2_fill_2 FILLER_120_1138 ();
 sg13g2_fill_1 FILLER_120_1140 ();
 sg13g2_fill_2 FILLER_120_1146 ();
 sg13g2_fill_1 FILLER_120_1148 ();
 sg13g2_fill_4 FILLER_120_1162 ();
 sg13g2_fill_2 FILLER_120_1166 ();
 sg13g2_fill_2 FILLER_120_1176 ();
 sg13g2_fill_8 FILLER_120_1183 ();
 sg13g2_fill_8 FILLER_120_1191 ();
 sg13g2_fill_4 FILLER_120_1199 ();
 sg13g2_fill_1 FILLER_120_1203 ();
 sg13g2_fill_4 FILLER_120_1208 ();
 sg13g2_fill_2 FILLER_120_1212 ();
 sg13g2_fill_1 FILLER_120_1214 ();
 sg13g2_fill_1 FILLER_120_1220 ();
 sg13g2_fill_1 FILLER_120_1254 ();
 sg13g2_fill_4 FILLER_120_1260 ();
 sg13g2_fill_1 FILLER_120_1306 ();
 sg13g2_fill_1 FILLER_120_1316 ();
 sg13g2_fill_1 FILLER_120_1349 ();
 sg13g2_fill_8 FILLER_120_1355 ();
 sg13g2_fill_2 FILLER_120_1363 ();
 sg13g2_fill_1 FILLER_120_1365 ();
 sg13g2_fill_2 FILLER_120_1379 ();
 sg13g2_fill_4 FILLER_120_1394 ();
 sg13g2_fill_1 FILLER_120_1398 ();
 sg13g2_fill_8 FILLER_120_1404 ();
 sg13g2_fill_8 FILLER_120_1412 ();
 sg13g2_fill_1 FILLER_120_1452 ();
 sg13g2_fill_1 FILLER_120_1463 ();
 sg13g2_fill_4 FILLER_120_1473 ();
 sg13g2_fill_8 FILLER_120_1486 ();
 sg13g2_fill_8 FILLER_120_1494 ();
 sg13g2_fill_8 FILLER_120_1502 ();
 sg13g2_fill_4 FILLER_120_1510 ();
 sg13g2_fill_2 FILLER_120_1514 ();
 sg13g2_fill_2 FILLER_120_1521 ();
 sg13g2_fill_1 FILLER_120_1527 ();
 sg13g2_fill_8 FILLER_120_1532 ();
 sg13g2_fill_8 FILLER_120_1540 ();
 sg13g2_fill_2 FILLER_120_1548 ();
 sg13g2_fill_2 FILLER_120_1572 ();
 sg13g2_fill_4 FILLER_120_1585 ();
 sg13g2_fill_2 FILLER_120_1589 ();
 sg13g2_fill_1 FILLER_120_1591 ();
 sg13g2_fill_4 FILLER_121_0 ();
 sg13g2_fill_4 FILLER_121_14 ();
 sg13g2_fill_2 FILLER_121_18 ();
 sg13g2_fill_2 FILLER_121_28 ();
 sg13g2_fill_4 FILLER_121_35 ();
 sg13g2_fill_2 FILLER_121_39 ();
 sg13g2_fill_1 FILLER_121_41 ();
 sg13g2_fill_8 FILLER_121_47 ();
 sg13g2_fill_8 FILLER_121_55 ();
 sg13g2_fill_1 FILLER_121_69 ();
 sg13g2_fill_2 FILLER_121_73 ();
 sg13g2_fill_1 FILLER_121_75 ();
 sg13g2_fill_8 FILLER_121_96 ();
 sg13g2_fill_4 FILLER_121_104 ();
 sg13g2_fill_1 FILLER_121_108 ();
 sg13g2_fill_8 FILLER_121_114 ();
 sg13g2_fill_8 FILLER_121_132 ();
 sg13g2_fill_4 FILLER_121_140 ();
 sg13g2_fill_1 FILLER_121_154 ();
 sg13g2_fill_4 FILLER_121_160 ();
 sg13g2_fill_1 FILLER_121_164 ();
 sg13g2_fill_8 FILLER_121_175 ();
 sg13g2_fill_4 FILLER_121_183 ();
 sg13g2_fill_2 FILLER_121_187 ();
 sg13g2_fill_8 FILLER_121_210 ();
 sg13g2_fill_8 FILLER_121_218 ();
 sg13g2_fill_8 FILLER_121_226 ();
 sg13g2_fill_4 FILLER_121_234 ();
 sg13g2_fill_2 FILLER_121_238 ();
 sg13g2_fill_2 FILLER_121_266 ();
 sg13g2_fill_1 FILLER_121_268 ();
 sg13g2_fill_2 FILLER_121_305 ();
 sg13g2_fill_1 FILLER_121_307 ();
 sg13g2_fill_4 FILLER_121_316 ();
 sg13g2_fill_2 FILLER_121_320 ();
 sg13g2_fill_8 FILLER_121_330 ();
 sg13g2_fill_4 FILLER_121_338 ();
 sg13g2_fill_1 FILLER_121_342 ();
 sg13g2_fill_8 FILLER_121_360 ();
 sg13g2_fill_1 FILLER_121_368 ();
 sg13g2_fill_1 FILLER_121_415 ();
 sg13g2_fill_4 FILLER_121_426 ();
 sg13g2_fill_2 FILLER_121_448 ();
 sg13g2_fill_1 FILLER_121_464 ();
 sg13g2_fill_8 FILLER_121_494 ();
 sg13g2_fill_8 FILLER_121_502 ();
 sg13g2_fill_2 FILLER_121_510 ();
 sg13g2_fill_2 FILLER_121_548 ();
 sg13g2_fill_1 FILLER_121_550 ();
 sg13g2_fill_8 FILLER_121_577 ();
 sg13g2_fill_8 FILLER_121_585 ();
 sg13g2_fill_8 FILLER_121_593 ();
 sg13g2_fill_8 FILLER_121_601 ();
 sg13g2_fill_8 FILLER_121_609 ();
 sg13g2_fill_8 FILLER_121_617 ();
 sg13g2_fill_4 FILLER_121_625 ();
 sg13g2_fill_2 FILLER_121_629 ();
 sg13g2_fill_1 FILLER_121_639 ();
 sg13g2_fill_8 FILLER_121_676 ();
 sg13g2_fill_8 FILLER_121_684 ();
 sg13g2_fill_8 FILLER_121_692 ();
 sg13g2_fill_8 FILLER_121_700 ();
 sg13g2_fill_8 FILLER_121_708 ();
 sg13g2_fill_8 FILLER_121_716 ();
 sg13g2_fill_8 FILLER_121_724 ();
 sg13g2_fill_8 FILLER_121_732 ();
 sg13g2_fill_4 FILLER_121_740 ();
 sg13g2_fill_1 FILLER_121_744 ();
 sg13g2_fill_8 FILLER_121_770 ();
 sg13g2_fill_8 FILLER_121_778 ();
 sg13g2_fill_2 FILLER_121_786 ();
 sg13g2_fill_8 FILLER_121_813 ();
 sg13g2_fill_8 FILLER_121_821 ();
 sg13g2_fill_1 FILLER_121_829 ();
 sg13g2_fill_1 FILLER_121_850 ();
 sg13g2_fill_4 FILLER_121_894 ();
 sg13g2_fill_2 FILLER_121_898 ();
 sg13g2_fill_1 FILLER_121_900 ();
 sg13g2_fill_4 FILLER_121_925 ();
 sg13g2_fill_2 FILLER_121_929 ();
 sg13g2_fill_1 FILLER_121_931 ();
 sg13g2_fill_4 FILLER_121_940 ();
 sg13g2_fill_1 FILLER_121_944 ();
 sg13g2_fill_1 FILLER_121_959 ();
 sg13g2_fill_8 FILLER_121_965 ();
 sg13g2_fill_8 FILLER_121_973 ();
 sg13g2_fill_8 FILLER_121_981 ();
 sg13g2_fill_4 FILLER_121_989 ();
 sg13g2_fill_2 FILLER_121_993 ();
 sg13g2_fill_1 FILLER_121_995 ();
 sg13g2_fill_1 FILLER_121_1008 ();
 sg13g2_fill_4 FILLER_121_1027 ();
 sg13g2_fill_1 FILLER_121_1031 ();
 sg13g2_fill_8 FILLER_121_1037 ();
 sg13g2_fill_4 FILLER_121_1045 ();
 sg13g2_fill_1 FILLER_121_1049 ();
 sg13g2_fill_4 FILLER_121_1067 ();
 sg13g2_fill_2 FILLER_121_1071 ();
 sg13g2_fill_1 FILLER_121_1073 ();
 sg13g2_fill_2 FILLER_121_1093 ();
 sg13g2_fill_1 FILLER_121_1100 ();
 sg13g2_fill_1 FILLER_121_1113 ();
 sg13g2_fill_1 FILLER_121_1143 ();
 sg13g2_fill_2 FILLER_121_1156 ();
 sg13g2_fill_4 FILLER_121_1168 ();
 sg13g2_fill_2 FILLER_121_1172 ();
 sg13g2_fill_8 FILLER_121_1204 ();
 sg13g2_fill_2 FILLER_121_1212 ();
 sg13g2_fill_1 FILLER_121_1214 ();
 sg13g2_fill_1 FILLER_121_1221 ();
 sg13g2_fill_4 FILLER_121_1233 ();
 sg13g2_fill_2 FILLER_121_1237 ();
 sg13g2_fill_1 FILLER_121_1239 ();
 sg13g2_fill_4 FILLER_121_1248 ();
 sg13g2_fill_2 FILLER_121_1252 ();
 sg13g2_fill_1 FILLER_121_1254 ();
 sg13g2_fill_8 FILLER_121_1264 ();
 sg13g2_fill_2 FILLER_121_1284 ();
 sg13g2_fill_1 FILLER_121_1306 ();
 sg13g2_fill_2 FILLER_121_1322 ();
 sg13g2_fill_1 FILLER_121_1354 ();
 sg13g2_fill_2 FILLER_121_1365 ();
 sg13g2_fill_1 FILLER_121_1367 ();
 sg13g2_fill_2 FILLER_121_1380 ();
 sg13g2_fill_1 FILLER_121_1382 ();
 sg13g2_fill_2 FILLER_121_1389 ();
 sg13g2_fill_4 FILLER_121_1396 ();
 sg13g2_fill_4 FILLER_121_1405 ();
 sg13g2_fill_1 FILLER_121_1409 ();
 sg13g2_fill_4 FILLER_121_1415 ();
 sg13g2_fill_1 FILLER_121_1419 ();
 sg13g2_fill_8 FILLER_121_1424 ();
 sg13g2_fill_8 FILLER_121_1432 ();
 sg13g2_fill_4 FILLER_121_1440 ();
 sg13g2_fill_8 FILLER_121_1454 ();
 sg13g2_fill_2 FILLER_121_1462 ();
 sg13g2_fill_8 FILLER_121_1469 ();
 sg13g2_fill_4 FILLER_121_1477 ();
 sg13g2_fill_1 FILLER_121_1481 ();
 sg13g2_fill_4 FILLER_121_1486 ();
 sg13g2_fill_8 FILLER_121_1541 ();
 sg13g2_fill_1 FILLER_121_1549 ();
 sg13g2_fill_8 FILLER_121_1561 ();
 sg13g2_fill_2 FILLER_121_1569 ();
 sg13g2_fill_1 FILLER_121_1571 ();
 sg13g2_fill_8 FILLER_121_1580 ();
 sg13g2_fill_4 FILLER_121_1588 ();
 sg13g2_fill_1 FILLER_122_26 ();
 sg13g2_fill_1 FILLER_122_36 ();
 sg13g2_fill_8 FILLER_122_52 ();
 sg13g2_fill_8 FILLER_122_60 ();
 sg13g2_fill_2 FILLER_122_68 ();
 sg13g2_fill_2 FILLER_122_87 ();
 sg13g2_fill_2 FILLER_122_99 ();
 sg13g2_fill_8 FILLER_122_119 ();
 sg13g2_fill_8 FILLER_122_127 ();
 sg13g2_fill_8 FILLER_122_135 ();
 sg13g2_fill_4 FILLER_122_143 ();
 sg13g2_fill_1 FILLER_122_213 ();
 sg13g2_fill_8 FILLER_122_229 ();
 sg13g2_fill_2 FILLER_122_237 ();
 sg13g2_fill_8 FILLER_122_249 ();
 sg13g2_fill_4 FILLER_122_257 ();
 sg13g2_fill_1 FILLER_122_261 ();
 sg13g2_fill_8 FILLER_122_283 ();
 sg13g2_fill_8 FILLER_122_291 ();
 sg13g2_fill_1 FILLER_122_299 ();
 sg13g2_fill_4 FILLER_122_305 ();
 sg13g2_fill_1 FILLER_122_309 ();
 sg13g2_fill_1 FILLER_122_333 ();
 sg13g2_fill_8 FILLER_122_360 ();
 sg13g2_fill_2 FILLER_122_368 ();
 sg13g2_fill_1 FILLER_122_370 ();
 sg13g2_fill_4 FILLER_122_402 ();
 sg13g2_fill_2 FILLER_122_406 ();
 sg13g2_fill_1 FILLER_122_408 ();
 sg13g2_fill_2 FILLER_122_419 ();
 sg13g2_fill_8 FILLER_122_426 ();
 sg13g2_fill_2 FILLER_122_434 ();
 sg13g2_fill_1 FILLER_122_436 ();
 sg13g2_fill_8 FILLER_122_449 ();
 sg13g2_fill_8 FILLER_122_457 ();
 sg13g2_fill_8 FILLER_122_465 ();
 sg13g2_fill_8 FILLER_122_473 ();
 sg13g2_fill_8 FILLER_122_481 ();
 sg13g2_fill_4 FILLER_122_489 ();
 sg13g2_fill_1 FILLER_122_493 ();
 sg13g2_fill_4 FILLER_122_520 ();
 sg13g2_fill_4 FILLER_122_534 ();
 sg13g2_fill_1 FILLER_122_542 ();
 sg13g2_fill_8 FILLER_122_553 ();
 sg13g2_fill_1 FILLER_122_561 ();
 sg13g2_fill_2 FILLER_122_567 ();
 sg13g2_fill_8 FILLER_122_595 ();
 sg13g2_fill_8 FILLER_122_603 ();
 sg13g2_fill_8 FILLER_122_611 ();
 sg13g2_fill_2 FILLER_122_619 ();
 sg13g2_fill_1 FILLER_122_626 ();
 sg13g2_fill_4 FILLER_122_632 ();
 sg13g2_fill_1 FILLER_122_641 ();
 sg13g2_fill_8 FILLER_122_658 ();
 sg13g2_fill_8 FILLER_122_666 ();
 sg13g2_fill_2 FILLER_122_674 ();
 sg13g2_fill_1 FILLER_122_676 ();
 sg13g2_fill_2 FILLER_122_747 ();
 sg13g2_fill_1 FILLER_122_816 ();
 sg13g2_fill_8 FILLER_122_825 ();
 sg13g2_fill_4 FILLER_122_833 ();
 sg13g2_fill_2 FILLER_122_837 ();
 sg13g2_fill_1 FILLER_122_839 ();
 sg13g2_fill_4 FILLER_122_848 ();
 sg13g2_fill_2 FILLER_122_893 ();
 sg13g2_fill_8 FILLER_122_912 ();
 sg13g2_fill_8 FILLER_122_920 ();
 sg13g2_fill_2 FILLER_122_928 ();
 sg13g2_fill_4 FILLER_122_942 ();
 sg13g2_fill_1 FILLER_122_946 ();
 sg13g2_fill_1 FILLER_122_970 ();
 sg13g2_fill_1 FILLER_122_977 ();
 sg13g2_fill_8 FILLER_122_983 ();
 sg13g2_fill_4 FILLER_122_991 ();
 sg13g2_fill_1 FILLER_122_995 ();
 sg13g2_fill_4 FILLER_122_1003 ();
 sg13g2_fill_4 FILLER_122_1013 ();
 sg13g2_fill_2 FILLER_122_1044 ();
 sg13g2_fill_1 FILLER_122_1046 ();
 sg13g2_fill_1 FILLER_122_1054 ();
 sg13g2_fill_4 FILLER_122_1059 ();
 sg13g2_fill_1 FILLER_122_1063 ();
 sg13g2_fill_8 FILLER_122_1079 ();
 sg13g2_fill_2 FILLER_122_1087 ();
 sg13g2_fill_1 FILLER_122_1089 ();
 sg13g2_fill_2 FILLER_122_1096 ();
 sg13g2_fill_8 FILLER_122_1101 ();
 sg13g2_fill_2 FILLER_122_1148 ();
 sg13g2_fill_8 FILLER_122_1158 ();
 sg13g2_fill_8 FILLER_122_1166 ();
 sg13g2_fill_8 FILLER_122_1179 ();
 sg13g2_fill_8 FILLER_122_1187 ();
 sg13g2_fill_8 FILLER_122_1195 ();
 sg13g2_fill_4 FILLER_122_1203 ();
 sg13g2_fill_2 FILLER_122_1207 ();
 sg13g2_fill_2 FILLER_122_1212 ();
 sg13g2_fill_1 FILLER_122_1232 ();
 sg13g2_fill_1 FILLER_122_1242 ();
 sg13g2_fill_2 FILLER_122_1274 ();
 sg13g2_fill_1 FILLER_122_1279 ();
 sg13g2_fill_1 FILLER_122_1291 ();
 sg13g2_fill_2 FILLER_122_1318 ();
 sg13g2_fill_1 FILLER_122_1358 ();
 sg13g2_fill_4 FILLER_122_1373 ();
 sg13g2_fill_1 FILLER_122_1386 ();
 sg13g2_fill_1 FILLER_122_1402 ();
 sg13g2_fill_8 FILLER_122_1447 ();
 sg13g2_fill_4 FILLER_122_1455 ();
 sg13g2_fill_2 FILLER_122_1459 ();
 sg13g2_fill_1 FILLER_122_1461 ();
 sg13g2_fill_4 FILLER_122_1472 ();
 sg13g2_fill_2 FILLER_122_1476 ();
 sg13g2_fill_8 FILLER_122_1483 ();
 sg13g2_fill_2 FILLER_122_1491 ();
 sg13g2_fill_1 FILLER_122_1493 ();
 sg13g2_fill_8 FILLER_122_1549 ();
 sg13g2_fill_8 FILLER_122_1557 ();
 sg13g2_fill_8 FILLER_122_1565 ();
 sg13g2_fill_2 FILLER_122_1573 ();
 sg13g2_fill_1 FILLER_122_1575 ();
 sg13g2_fill_4 FILLER_122_1587 ();
 sg13g2_fill_1 FILLER_122_1591 ();
 sg13g2_fill_8 FILLER_123_0 ();
 sg13g2_fill_2 FILLER_123_8 ();
 sg13g2_fill_1 FILLER_123_10 ();
 sg13g2_fill_2 FILLER_123_34 ();
 sg13g2_fill_2 FILLER_123_42 ();
 sg13g2_fill_1 FILLER_123_44 ();
 sg13g2_fill_2 FILLER_123_65 ();
 sg13g2_fill_1 FILLER_123_67 ();
 sg13g2_fill_8 FILLER_123_86 ();
 sg13g2_fill_4 FILLER_123_94 ();
 sg13g2_fill_2 FILLER_123_98 ();
 sg13g2_fill_1 FILLER_123_100 ();
 sg13g2_fill_4 FILLER_123_121 ();
 sg13g2_fill_8 FILLER_123_151 ();
 sg13g2_fill_8 FILLER_123_159 ();
 sg13g2_fill_1 FILLER_123_167 ();
 sg13g2_fill_8 FILLER_123_176 ();
 sg13g2_fill_8 FILLER_123_184 ();
 sg13g2_fill_8 FILLER_123_192 ();
 sg13g2_fill_8 FILLER_123_200 ();
 sg13g2_fill_4 FILLER_123_208 ();
 sg13g2_fill_1 FILLER_123_212 ();
 sg13g2_fill_4 FILLER_123_286 ();
 sg13g2_fill_8 FILLER_123_307 ();
 sg13g2_fill_8 FILLER_123_315 ();
 sg13g2_fill_4 FILLER_123_323 ();
 sg13g2_fill_2 FILLER_123_327 ();
 sg13g2_fill_8 FILLER_123_334 ();
 sg13g2_fill_8 FILLER_123_342 ();
 sg13g2_fill_8 FILLER_123_350 ();
 sg13g2_fill_8 FILLER_123_358 ();
 sg13g2_fill_4 FILLER_123_366 ();
 sg13g2_fill_2 FILLER_123_370 ();
 sg13g2_fill_4 FILLER_123_421 ();
 sg13g2_fill_2 FILLER_123_425 ();
 sg13g2_fill_1 FILLER_123_427 ();
 sg13g2_fill_2 FILLER_123_441 ();
 sg13g2_fill_8 FILLER_123_449 ();
 sg13g2_fill_8 FILLER_123_457 ();
 sg13g2_fill_4 FILLER_123_475 ();
 sg13g2_fill_1 FILLER_123_479 ();
 sg13g2_fill_8 FILLER_123_501 ();
 sg13g2_fill_4 FILLER_123_509 ();
 sg13g2_fill_2 FILLER_123_513 ();
 sg13g2_fill_1 FILLER_123_515 ();
 sg13g2_fill_8 FILLER_123_526 ();
 sg13g2_fill_4 FILLER_123_534 ();
 sg13g2_fill_2 FILLER_123_538 ();
 sg13g2_fill_8 FILLER_123_550 ();
 sg13g2_fill_8 FILLER_123_558 ();
 sg13g2_fill_2 FILLER_123_566 ();
 sg13g2_fill_1 FILLER_123_568 ();
 sg13g2_fill_2 FILLER_123_579 ();
 sg13g2_fill_8 FILLER_123_625 ();
 sg13g2_fill_8 FILLER_123_633 ();
 sg13g2_fill_8 FILLER_123_641 ();
 sg13g2_fill_4 FILLER_123_649 ();
 sg13g2_fill_8 FILLER_123_689 ();
 sg13g2_fill_1 FILLER_123_697 ();
 sg13g2_fill_4 FILLER_123_774 ();
 sg13g2_fill_1 FILLER_123_778 ();
 sg13g2_fill_4 FILLER_123_795 ();
 sg13g2_fill_2 FILLER_123_799 ();
 sg13g2_fill_1 FILLER_123_843 ();
 sg13g2_fill_8 FILLER_123_852 ();
 sg13g2_fill_2 FILLER_123_860 ();
 sg13g2_fill_1 FILLER_123_862 ();
 sg13g2_fill_2 FILLER_123_921 ();
 sg13g2_fill_2 FILLER_123_966 ();
 sg13g2_fill_4 FILLER_123_984 ();
 sg13g2_fill_2 FILLER_123_1000 ();
 sg13g2_fill_1 FILLER_123_1017 ();
 sg13g2_fill_8 FILLER_123_1028 ();
 sg13g2_fill_4 FILLER_123_1053 ();
 sg13g2_fill_2 FILLER_123_1057 ();
 sg13g2_fill_4 FILLER_123_1069 ();
 sg13g2_fill_2 FILLER_123_1073 ();
 sg13g2_fill_1 FILLER_123_1075 ();
 sg13g2_fill_4 FILLER_123_1080 ();
 sg13g2_fill_2 FILLER_123_1084 ();
 sg13g2_fill_1 FILLER_123_1086 ();
 sg13g2_fill_2 FILLER_123_1091 ();
 sg13g2_fill_8 FILLER_123_1103 ();
 sg13g2_fill_4 FILLER_123_1137 ();
 sg13g2_fill_4 FILLER_123_1168 ();
 sg13g2_fill_1 FILLER_123_1177 ();
 sg13g2_fill_4 FILLER_123_1183 ();
 sg13g2_fill_2 FILLER_123_1187 ();
 sg13g2_fill_1 FILLER_123_1221 ();
 sg13g2_fill_8 FILLER_123_1248 ();
 sg13g2_fill_4 FILLER_123_1256 ();
 sg13g2_fill_1 FILLER_123_1260 ();
 sg13g2_fill_4 FILLER_123_1266 ();
 sg13g2_fill_2 FILLER_123_1288 ();
 sg13g2_fill_8 FILLER_123_1354 ();
 sg13g2_fill_8 FILLER_123_1362 ();
 sg13g2_fill_8 FILLER_123_1375 ();
 sg13g2_fill_8 FILLER_123_1383 ();
 sg13g2_fill_4 FILLER_123_1391 ();
 sg13g2_fill_2 FILLER_123_1395 ();
 sg13g2_fill_1 FILLER_123_1397 ();
 sg13g2_fill_8 FILLER_123_1403 ();
 sg13g2_fill_8 FILLER_123_1411 ();
 sg13g2_fill_8 FILLER_123_1419 ();
 sg13g2_fill_4 FILLER_123_1427 ();
 sg13g2_fill_2 FILLER_123_1431 ();
 sg13g2_fill_1 FILLER_123_1433 ();
 sg13g2_fill_2 FILLER_123_1439 ();
 sg13g2_fill_1 FILLER_123_1441 ();
 sg13g2_fill_2 FILLER_123_1446 ();
 sg13g2_fill_8 FILLER_123_1453 ();
 sg13g2_fill_1 FILLER_123_1475 ();
 sg13g2_fill_2 FILLER_123_1489 ();
 sg13g2_fill_8 FILLER_123_1533 ();
 sg13g2_fill_8 FILLER_123_1541 ();
 sg13g2_fill_2 FILLER_123_1549 ();
 sg13g2_fill_2 FILLER_123_1573 ();
 sg13g2_fill_4 FILLER_123_1586 ();
 sg13g2_fill_2 FILLER_123_1590 ();
 sg13g2_fill_8 FILLER_124_0 ();
 sg13g2_fill_4 FILLER_124_8 ();
 sg13g2_fill_2 FILLER_124_12 ();
 sg13g2_fill_8 FILLER_124_55 ();
 sg13g2_fill_4 FILLER_124_63 ();
 sg13g2_fill_2 FILLER_124_67 ();
 sg13g2_fill_2 FILLER_124_73 ();
 sg13g2_fill_8 FILLER_124_82 ();
 sg13g2_fill_1 FILLER_124_90 ();
 sg13g2_fill_8 FILLER_124_101 ();
 sg13g2_fill_1 FILLER_124_109 ();
 sg13g2_fill_8 FILLER_124_115 ();
 sg13g2_fill_8 FILLER_124_123 ();
 sg13g2_fill_4 FILLER_124_131 ();
 sg13g2_fill_2 FILLER_124_135 ();
 sg13g2_fill_8 FILLER_124_142 ();
 sg13g2_fill_8 FILLER_124_150 ();
 sg13g2_fill_1 FILLER_124_158 ();
 sg13g2_fill_8 FILLER_124_167 ();
 sg13g2_fill_8 FILLER_124_175 ();
 sg13g2_fill_1 FILLER_124_228 ();
 sg13g2_fill_8 FILLER_124_240 ();
 sg13g2_fill_8 FILLER_124_248 ();
 sg13g2_fill_8 FILLER_124_256 ();
 sg13g2_fill_8 FILLER_124_264 ();
 sg13g2_fill_2 FILLER_124_272 ();
 sg13g2_fill_2 FILLER_124_312 ();
 sg13g2_fill_1 FILLER_124_314 ();
 sg13g2_fill_8 FILLER_124_333 ();
 sg13g2_fill_8 FILLER_124_341 ();
 sg13g2_fill_2 FILLER_124_359 ();
 sg13g2_fill_1 FILLER_124_361 ();
 sg13g2_fill_8 FILLER_124_388 ();
 sg13g2_fill_1 FILLER_124_396 ();
 sg13g2_fill_8 FILLER_124_407 ();
 sg13g2_fill_4 FILLER_124_415 ();
 sg13g2_fill_2 FILLER_124_419 ();
 sg13g2_fill_1 FILLER_124_421 ();
 sg13g2_fill_8 FILLER_124_427 ();
 sg13g2_fill_4 FILLER_124_435 ();
 sg13g2_fill_1 FILLER_124_478 ();
 sg13g2_fill_2 FILLER_124_515 ();
 sg13g2_fill_1 FILLER_124_517 ();
 sg13g2_fill_4 FILLER_124_528 ();
 sg13g2_fill_2 FILLER_124_532 ();
 sg13g2_fill_1 FILLER_124_539 ();
 sg13g2_fill_8 FILLER_124_550 ();
 sg13g2_fill_4 FILLER_124_558 ();
 sg13g2_fill_8 FILLER_124_592 ();
 sg13g2_fill_1 FILLER_124_600 ();
 sg13g2_fill_8 FILLER_124_627 ();
 sg13g2_fill_4 FILLER_124_635 ();
 sg13g2_fill_1 FILLER_124_639 ();
 sg13g2_fill_8 FILLER_124_653 ();
 sg13g2_fill_8 FILLER_124_661 ();
 sg13g2_fill_8 FILLER_124_669 ();
 sg13g2_fill_8 FILLER_124_677 ();
 sg13g2_fill_8 FILLER_124_685 ();
 sg13g2_fill_1 FILLER_124_693 ();
 sg13g2_fill_8 FILLER_124_725 ();
 sg13g2_fill_8 FILLER_124_733 ();
 sg13g2_fill_8 FILLER_124_741 ();
 sg13g2_fill_8 FILLER_124_749 ();
 sg13g2_fill_2 FILLER_124_757 ();
 sg13g2_fill_1 FILLER_124_759 ();
 sg13g2_fill_8 FILLER_124_771 ();
 sg13g2_fill_8 FILLER_124_779 ();
 sg13g2_fill_4 FILLER_124_787 ();
 sg13g2_fill_1 FILLER_124_791 ();
 sg13g2_fill_4 FILLER_124_817 ();
 sg13g2_fill_2 FILLER_124_821 ();
 sg13g2_fill_4 FILLER_124_861 ();
 sg13g2_fill_1 FILLER_124_865 ();
 sg13g2_fill_8 FILLER_124_906 ();
 sg13g2_fill_2 FILLER_124_914 ();
 sg13g2_fill_4 FILLER_124_945 ();
 sg13g2_fill_1 FILLER_124_949 ();
 sg13g2_fill_2 FILLER_124_978 ();
 sg13g2_fill_1 FILLER_124_980 ();
 sg13g2_fill_8 FILLER_124_986 ();
 sg13g2_fill_4 FILLER_124_994 ();
 sg13g2_fill_1 FILLER_124_998 ();
 sg13g2_fill_4 FILLER_124_1009 ();
 sg13g2_fill_1 FILLER_124_1013 ();
 sg13g2_fill_2 FILLER_124_1022 ();
 sg13g2_fill_1 FILLER_124_1024 ();
 sg13g2_fill_8 FILLER_124_1038 ();
 sg13g2_fill_4 FILLER_124_1046 ();
 sg13g2_fill_1 FILLER_124_1050 ();
 sg13g2_fill_2 FILLER_124_1069 ();
 sg13g2_fill_4 FILLER_124_1102 ();
 sg13g2_fill_2 FILLER_124_1106 ();
 sg13g2_fill_4 FILLER_124_1117 ();
 sg13g2_fill_1 FILLER_124_1121 ();
 sg13g2_fill_2 FILLER_124_1126 ();
 sg13g2_fill_2 FILLER_124_1141 ();
 sg13g2_fill_1 FILLER_124_1143 ();
 sg13g2_fill_4 FILLER_124_1169 ();
 sg13g2_fill_1 FILLER_124_1173 ();
 sg13g2_fill_2 FILLER_124_1183 ();
 sg13g2_fill_2 FILLER_124_1205 ();
 sg13g2_fill_2 FILLER_124_1250 ();
 sg13g2_fill_4 FILLER_124_1261 ();
 sg13g2_fill_1 FILLER_124_1265 ();
 sg13g2_fill_2 FILLER_124_1274 ();
 sg13g2_fill_8 FILLER_124_1339 ();
 sg13g2_fill_1 FILLER_124_1347 ();
 sg13g2_fill_2 FILLER_124_1358 ();
 sg13g2_fill_8 FILLER_124_1370 ();
 sg13g2_fill_8 FILLER_124_1378 ();
 sg13g2_fill_2 FILLER_124_1386 ();
 sg13g2_fill_1 FILLER_124_1388 ();
 sg13g2_fill_4 FILLER_124_1393 ();
 sg13g2_fill_2 FILLER_124_1397 ();
 sg13g2_fill_4 FILLER_124_1404 ();
 sg13g2_fill_2 FILLER_124_1408 ();
 sg13g2_fill_1 FILLER_124_1410 ();
 sg13g2_fill_4 FILLER_124_1429 ();
 sg13g2_fill_2 FILLER_124_1433 ();
 sg13g2_fill_1 FILLER_124_1435 ();
 sg13g2_fill_2 FILLER_124_1467 ();
 sg13g2_fill_8 FILLER_124_1495 ();
 sg13g2_fill_8 FILLER_124_1503 ();
 sg13g2_fill_4 FILLER_124_1511 ();
 sg13g2_fill_2 FILLER_124_1515 ();
 sg13g2_fill_1 FILLER_124_1517 ();
 sg13g2_fill_8 FILLER_124_1522 ();
 sg13g2_fill_8 FILLER_124_1530 ();
 sg13g2_fill_8 FILLER_124_1538 ();
 sg13g2_fill_2 FILLER_124_1546 ();
 sg13g2_fill_4 FILLER_125_0 ();
 sg13g2_fill_8 FILLER_125_14 ();
 sg13g2_fill_4 FILLER_125_25 ();
 sg13g2_fill_2 FILLER_125_29 ();
 sg13g2_fill_1 FILLER_125_31 ();
 sg13g2_fill_8 FILLER_125_40 ();
 sg13g2_fill_4 FILLER_125_48 ();
 sg13g2_fill_1 FILLER_125_52 ();
 sg13g2_fill_4 FILLER_125_57 ();
 sg13g2_fill_2 FILLER_125_61 ();
 sg13g2_fill_4 FILLER_125_68 ();
 sg13g2_fill_8 FILLER_125_76 ();
 sg13g2_fill_2 FILLER_125_108 ();
 sg13g2_fill_2 FILLER_125_120 ();
 sg13g2_fill_1 FILLER_125_122 ();
 sg13g2_fill_1 FILLER_125_127 ();
 sg13g2_fill_4 FILLER_125_132 ();
 sg13g2_fill_2 FILLER_125_136 ();
 sg13g2_fill_8 FILLER_125_147 ();
 sg13g2_fill_1 FILLER_125_155 ();
 sg13g2_fill_1 FILLER_125_166 ();
 sg13g2_fill_4 FILLER_125_193 ();
 sg13g2_fill_2 FILLER_125_197 ();
 sg13g2_fill_1 FILLER_125_225 ();
 sg13g2_fill_8 FILLER_125_268 ();
 sg13g2_fill_4 FILLER_125_276 ();
 sg13g2_fill_2 FILLER_125_280 ();
 sg13g2_fill_1 FILLER_125_282 ();
 sg13g2_fill_4 FILLER_125_288 ();
 sg13g2_fill_4 FILLER_125_394 ();
 sg13g2_fill_2 FILLER_125_398 ();
 sg13g2_fill_1 FILLER_125_400 ();
 sg13g2_fill_1 FILLER_125_427 ();
 sg13g2_fill_8 FILLER_125_435 ();
 sg13g2_fill_8 FILLER_125_443 ();
 sg13g2_fill_8 FILLER_125_451 ();
 sg13g2_fill_4 FILLER_125_459 ();
 sg13g2_fill_2 FILLER_125_463 ();
 sg13g2_fill_2 FILLER_125_526 ();
 sg13g2_fill_2 FILLER_125_534 ();
 sg13g2_fill_2 FILLER_125_578 ();
 sg13g2_fill_1 FILLER_125_580 ();
 sg13g2_fill_2 FILLER_125_611 ();
 sg13g2_fill_1 FILLER_125_613 ();
 sg13g2_fill_1 FILLER_125_622 ();
 sg13g2_fill_4 FILLER_125_631 ();
 sg13g2_fill_1 FILLER_125_635 ();
 sg13g2_fill_2 FILLER_125_657 ();
 sg13g2_fill_1 FILLER_125_659 ();
 sg13g2_fill_4 FILLER_125_696 ();
 sg13g2_fill_2 FILLER_125_700 ();
 sg13g2_fill_8 FILLER_125_727 ();
 sg13g2_fill_8 FILLER_125_735 ();
 sg13g2_fill_8 FILLER_125_743 ();
 sg13g2_fill_1 FILLER_125_751 ();
 sg13g2_fill_8 FILLER_125_790 ();
 sg13g2_fill_8 FILLER_125_798 ();
 sg13g2_fill_4 FILLER_125_806 ();
 sg13g2_fill_2 FILLER_125_810 ();
 sg13g2_fill_1 FILLER_125_851 ();
 sg13g2_fill_2 FILLER_125_860 ();
 sg13g2_fill_8 FILLER_125_867 ();
 sg13g2_fill_4 FILLER_125_875 ();
 sg13g2_fill_2 FILLER_125_879 ();
 sg13g2_fill_1 FILLER_125_881 ();
 sg13g2_fill_8 FILLER_125_887 ();
 sg13g2_fill_8 FILLER_125_895 ();
 sg13g2_fill_8 FILLER_125_903 ();
 sg13g2_fill_1 FILLER_125_911 ();
 sg13g2_fill_4 FILLER_125_922 ();
 sg13g2_fill_2 FILLER_125_926 ();
 sg13g2_fill_2 FILLER_125_938 ();
 sg13g2_fill_1 FILLER_125_940 ();
 sg13g2_fill_4 FILLER_125_954 ();
 sg13g2_fill_2 FILLER_125_958 ();
 sg13g2_fill_1 FILLER_125_960 ();
 sg13g2_fill_8 FILLER_125_970 ();
 sg13g2_fill_1 FILLER_125_978 ();
 sg13g2_fill_8 FILLER_125_985 ();
 sg13g2_fill_4 FILLER_125_993 ();
 sg13g2_fill_2 FILLER_125_997 ();
 sg13g2_fill_8 FILLER_125_1013 ();
 sg13g2_fill_1 FILLER_125_1021 ();
 sg13g2_fill_8 FILLER_125_1030 ();
 sg13g2_fill_4 FILLER_125_1038 ();
 sg13g2_fill_2 FILLER_125_1042 ();
 sg13g2_fill_1 FILLER_125_1044 ();
 sg13g2_fill_8 FILLER_125_1053 ();
 sg13g2_fill_1 FILLER_125_1061 ();
 sg13g2_fill_2 FILLER_125_1075 ();
 sg13g2_fill_8 FILLER_125_1082 ();
 sg13g2_fill_4 FILLER_125_1090 ();
 sg13g2_fill_2 FILLER_125_1099 ();
 sg13g2_fill_8 FILLER_125_1120 ();
 sg13g2_fill_8 FILLER_125_1128 ();
 sg13g2_fill_1 FILLER_125_1136 ();
 sg13g2_fill_4 FILLER_125_1141 ();
 sg13g2_fill_2 FILLER_125_1145 ();
 sg13g2_fill_2 FILLER_125_1152 ();
 sg13g2_fill_2 FILLER_125_1184 ();
 sg13g2_fill_8 FILLER_125_1191 ();
 sg13g2_fill_2 FILLER_125_1199 ();
 sg13g2_fill_1 FILLER_125_1201 ();
 sg13g2_fill_2 FILLER_125_1230 ();
 sg13g2_fill_1 FILLER_125_1232 ();
 sg13g2_fill_2 FILLER_125_1241 ();
 sg13g2_fill_1 FILLER_125_1243 ();
 sg13g2_fill_4 FILLER_125_1247 ();
 sg13g2_fill_8 FILLER_125_1255 ();
 sg13g2_fill_8 FILLER_125_1263 ();
 sg13g2_fill_4 FILLER_125_1271 ();
 sg13g2_fill_1 FILLER_125_1275 ();
 sg13g2_fill_4 FILLER_125_1285 ();
 sg13g2_fill_8 FILLER_125_1294 ();
 sg13g2_fill_8 FILLER_125_1302 ();
 sg13g2_fill_8 FILLER_125_1310 ();
 sg13g2_fill_8 FILLER_125_1318 ();
 sg13g2_fill_4 FILLER_125_1326 ();
 sg13g2_fill_4 FILLER_125_1343 ();
 sg13g2_fill_2 FILLER_125_1347 ();
 sg13g2_fill_1 FILLER_125_1349 ();
 sg13g2_fill_1 FILLER_125_1359 ();
 sg13g2_fill_2 FILLER_125_1370 ();
 sg13g2_fill_1 FILLER_125_1372 ();
 sg13g2_fill_1 FILLER_125_1393 ();
 sg13g2_fill_8 FILLER_125_1409 ();
 sg13g2_fill_2 FILLER_125_1417 ();
 sg13g2_fill_1 FILLER_125_1419 ();
 sg13g2_fill_2 FILLER_125_1469 ();
 sg13g2_fill_8 FILLER_125_1510 ();
 sg13g2_fill_4 FILLER_125_1518 ();
 sg13g2_fill_2 FILLER_125_1522 ();
 sg13g2_fill_8 FILLER_125_1550 ();
 sg13g2_fill_8 FILLER_125_1558 ();
 sg13g2_fill_4 FILLER_125_1566 ();
 sg13g2_fill_2 FILLER_125_1570 ();
 sg13g2_fill_1 FILLER_125_1572 ();
 sg13g2_fill_8 FILLER_125_1584 ();
 sg13g2_fill_8 FILLER_126_30 ();
 sg13g2_fill_2 FILLER_126_47 ();
 sg13g2_fill_2 FILLER_126_54 ();
 sg13g2_fill_1 FILLER_126_56 ();
 sg13g2_fill_1 FILLER_126_83 ();
 sg13g2_fill_4 FILLER_126_93 ();
 sg13g2_fill_8 FILLER_126_102 ();
 sg13g2_fill_2 FILLER_126_110 ();
 sg13g2_fill_1 FILLER_126_112 ();
 sg13g2_fill_1 FILLER_126_139 ();
 sg13g2_fill_8 FILLER_126_166 ();
 sg13g2_fill_8 FILLER_126_174 ();
 sg13g2_fill_8 FILLER_126_182 ();
 sg13g2_fill_8 FILLER_126_190 ();
 sg13g2_fill_8 FILLER_126_198 ();
 sg13g2_fill_8 FILLER_126_206 ();
 sg13g2_fill_8 FILLER_126_239 ();
 sg13g2_fill_4 FILLER_126_247 ();
 sg13g2_fill_2 FILLER_126_251 ();
 sg13g2_fill_1 FILLER_126_289 ();
 sg13g2_fill_2 FILLER_126_301 ();
 sg13g2_fill_8 FILLER_126_338 ();
 sg13g2_fill_4 FILLER_126_346 ();
 sg13g2_fill_1 FILLER_126_350 ();
 sg13g2_fill_8 FILLER_126_371 ();
 sg13g2_fill_8 FILLER_126_379 ();
 sg13g2_fill_8 FILLER_126_387 ();
 sg13g2_fill_8 FILLER_126_395 ();
 sg13g2_fill_4 FILLER_126_413 ();
 sg13g2_fill_1 FILLER_126_417 ();
 sg13g2_fill_4 FILLER_126_469 ();
 sg13g2_fill_2 FILLER_126_473 ();
 sg13g2_fill_1 FILLER_126_475 ();
 sg13g2_fill_4 FILLER_126_528 ();
 sg13g2_fill_1 FILLER_126_532 ();
 sg13g2_fill_2 FILLER_126_542 ();
 sg13g2_fill_1 FILLER_126_544 ();
 sg13g2_fill_2 FILLER_126_551 ();
 sg13g2_fill_2 FILLER_126_561 ();
 sg13g2_fill_1 FILLER_126_563 ();
 sg13g2_fill_2 FILLER_126_567 ();
 sg13g2_fill_1 FILLER_126_569 ();
 sg13g2_fill_8 FILLER_126_596 ();
 sg13g2_fill_4 FILLER_126_604 ();
 sg13g2_fill_2 FILLER_126_638 ();
 sg13g2_fill_1 FILLER_126_640 ();
 sg13g2_fill_4 FILLER_126_657 ();
 sg13g2_fill_1 FILLER_126_661 ();
 sg13g2_fill_8 FILLER_126_672 ();
 sg13g2_fill_2 FILLER_126_680 ();
 sg13g2_fill_1 FILLER_126_723 ();
 sg13g2_fill_4 FILLER_126_755 ();
 sg13g2_fill_8 FILLER_126_767 ();
 sg13g2_fill_4 FILLER_126_775 ();
 sg13g2_fill_1 FILLER_126_779 ();
 sg13g2_fill_2 FILLER_126_805 ();
 sg13g2_fill_8 FILLER_126_817 ();
 sg13g2_fill_2 FILLER_126_825 ();
 sg13g2_fill_1 FILLER_126_827 ();
 sg13g2_fill_4 FILLER_126_894 ();
 sg13g2_fill_1 FILLER_126_898 ();
 sg13g2_fill_4 FILLER_126_925 ();
 sg13g2_fill_2 FILLER_126_929 ();
 sg13g2_fill_1 FILLER_126_931 ();
 sg13g2_fill_2 FILLER_126_944 ();
 sg13g2_fill_1 FILLER_126_946 ();
 sg13g2_fill_2 FILLER_126_965 ();
 sg13g2_fill_1 FILLER_126_967 ();
 sg13g2_fill_8 FILLER_126_973 ();
 sg13g2_fill_8 FILLER_126_981 ();
 sg13g2_fill_8 FILLER_126_989 ();
 sg13g2_fill_1 FILLER_126_997 ();
 sg13g2_fill_1 FILLER_126_1007 ();
 sg13g2_fill_4 FILLER_126_1022 ();
 sg13g2_fill_8 FILLER_126_1043 ();
 sg13g2_fill_4 FILLER_126_1051 ();
 sg13g2_fill_8 FILLER_126_1063 ();
 sg13g2_fill_8 FILLER_126_1071 ();
 sg13g2_fill_4 FILLER_126_1079 ();
 sg13g2_fill_2 FILLER_126_1083 ();
 sg13g2_fill_8 FILLER_126_1094 ();
 sg13g2_fill_8 FILLER_126_1112 ();
 sg13g2_fill_8 FILLER_126_1120 ();
 sg13g2_fill_2 FILLER_126_1128 ();
 sg13g2_fill_1 FILLER_126_1130 ();
 sg13g2_fill_2 FILLER_126_1135 ();
 sg13g2_fill_1 FILLER_126_1137 ();
 sg13g2_fill_2 FILLER_126_1169 ();
 sg13g2_fill_2 FILLER_126_1186 ();
 sg13g2_fill_8 FILLER_126_1200 ();
 sg13g2_fill_2 FILLER_126_1208 ();
 sg13g2_fill_1 FILLER_126_1210 ();
 sg13g2_fill_1 FILLER_126_1224 ();
 sg13g2_fill_1 FILLER_126_1243 ();
 sg13g2_fill_2 FILLER_126_1247 ();
 sg13g2_fill_8 FILLER_126_1279 ();
 sg13g2_fill_1 FILLER_126_1287 ();
 sg13g2_fill_8 FILLER_126_1294 ();
 sg13g2_fill_8 FILLER_126_1311 ();
 sg13g2_fill_2 FILLER_126_1319 ();
 sg13g2_fill_8 FILLER_126_1324 ();
 sg13g2_fill_4 FILLER_126_1332 ();
 sg13g2_fill_2 FILLER_126_1336 ();
 sg13g2_fill_1 FILLER_126_1338 ();
 sg13g2_fill_8 FILLER_126_1358 ();
 sg13g2_fill_2 FILLER_126_1366 ();
 sg13g2_fill_1 FILLER_126_1368 ();
 sg13g2_fill_1 FILLER_126_1381 ();
 sg13g2_fill_1 FILLER_126_1413 ();
 sg13g2_fill_4 FILLER_126_1428 ();
 sg13g2_fill_2 FILLER_126_1432 ();
 sg13g2_fill_2 FILLER_126_1453 ();
 sg13g2_fill_8 FILLER_126_1512 ();
 sg13g2_fill_8 FILLER_126_1520 ();
 sg13g2_fill_4 FILLER_126_1528 ();
 sg13g2_fill_2 FILLER_126_1532 ();
 sg13g2_fill_2 FILLER_126_1542 ();
 sg13g2_fill_8 FILLER_126_1555 ();
 sg13g2_fill_8 FILLER_126_1563 ();
 sg13g2_fill_4 FILLER_126_1571 ();
 sg13g2_fill_1 FILLER_126_1575 ();
 sg13g2_fill_4 FILLER_126_1587 ();
 sg13g2_fill_1 FILLER_126_1591 ();
 sg13g2_fill_8 FILLER_127_0 ();
 sg13g2_fill_8 FILLER_127_8 ();
 sg13g2_fill_8 FILLER_127_16 ();
 sg13g2_fill_8 FILLER_127_41 ();
 sg13g2_fill_2 FILLER_127_49 ();
 sg13g2_fill_8 FILLER_127_56 ();
 sg13g2_fill_2 FILLER_127_64 ();
 sg13g2_fill_4 FILLER_127_70 ();
 sg13g2_fill_4 FILLER_127_78 ();
 sg13g2_fill_8 FILLER_127_86 ();
 sg13g2_fill_2 FILLER_127_94 ();
 sg13g2_fill_1 FILLER_127_96 ();
 sg13g2_fill_8 FILLER_127_107 ();
 sg13g2_fill_2 FILLER_127_115 ();
 sg13g2_fill_4 FILLER_127_121 ();
 sg13g2_fill_1 FILLER_127_125 ();
 sg13g2_fill_2 FILLER_127_130 ();
 sg13g2_fill_1 FILLER_127_132 ();
 sg13g2_fill_4 FILLER_127_143 ();
 sg13g2_fill_1 FILLER_127_147 ();
 sg13g2_fill_2 FILLER_127_152 ();
 sg13g2_fill_1 FILLER_127_154 ();
 sg13g2_fill_4 FILLER_127_160 ();
 sg13g2_fill_1 FILLER_127_164 ();
 sg13g2_fill_2 FILLER_127_217 ();
 sg13g2_fill_2 FILLER_127_228 ();
 sg13g2_fill_4 FILLER_127_238 ();
 sg13g2_fill_1 FILLER_127_242 ();
 sg13g2_fill_8 FILLER_127_253 ();
 sg13g2_fill_8 FILLER_127_261 ();
 sg13g2_fill_8 FILLER_127_269 ();
 sg13g2_fill_1 FILLER_127_277 ();
 sg13g2_fill_8 FILLER_127_310 ();
 sg13g2_fill_1 FILLER_127_318 ();
 sg13g2_fill_8 FILLER_127_340 ();
 sg13g2_fill_4 FILLER_127_348 ();
 sg13g2_fill_2 FILLER_127_383 ();
 sg13g2_fill_8 FILLER_127_395 ();
 sg13g2_fill_8 FILLER_127_403 ();
 sg13g2_fill_8 FILLER_127_411 ();
 sg13g2_fill_2 FILLER_127_419 ();
 sg13g2_fill_2 FILLER_127_440 ();
 sg13g2_fill_1 FILLER_127_442 ();
 sg13g2_fill_8 FILLER_127_469 ();
 sg13g2_fill_8 FILLER_127_477 ();
 sg13g2_fill_8 FILLER_127_485 ();
 sg13g2_fill_8 FILLER_127_493 ();
 sg13g2_fill_8 FILLER_127_501 ();
 sg13g2_fill_8 FILLER_127_509 ();
 sg13g2_fill_8 FILLER_127_517 ();
 sg13g2_fill_8 FILLER_127_525 ();
 sg13g2_fill_2 FILLER_127_533 ();
 sg13g2_fill_8 FILLER_127_545 ();
 sg13g2_fill_8 FILLER_127_553 ();
 sg13g2_fill_2 FILLER_127_561 ();
 sg13g2_fill_1 FILLER_127_563 ();
 sg13g2_fill_1 FILLER_127_589 ();
 sg13g2_fill_2 FILLER_127_639 ();
 sg13g2_fill_1 FILLER_127_651 ();
 sg13g2_fill_2 FILLER_127_704 ();
 sg13g2_fill_1 FILLER_127_706 ();
 sg13g2_fill_1 FILLER_127_717 ();
 sg13g2_fill_4 FILLER_127_744 ();
 sg13g2_fill_1 FILLER_127_748 ();
 sg13g2_fill_8 FILLER_127_781 ();
 sg13g2_fill_8 FILLER_127_804 ();
 sg13g2_fill_8 FILLER_127_812 ();
 sg13g2_fill_8 FILLER_127_820 ();
 sg13g2_fill_8 FILLER_127_838 ();
 sg13g2_fill_8 FILLER_127_846 ();
 sg13g2_fill_8 FILLER_127_854 ();
 sg13g2_fill_8 FILLER_127_862 ();
 sg13g2_fill_8 FILLER_127_870 ();
 sg13g2_fill_8 FILLER_127_878 ();
 sg13g2_fill_4 FILLER_127_886 ();
 sg13g2_fill_2 FILLER_127_890 ();
 sg13g2_fill_4 FILLER_127_933 ();
 sg13g2_fill_2 FILLER_127_937 ();
 sg13g2_fill_1 FILLER_127_939 ();
 sg13g2_fill_1 FILLER_127_952 ();
 sg13g2_fill_2 FILLER_127_964 ();
 sg13g2_fill_2 FILLER_127_972 ();
 sg13g2_fill_1 FILLER_127_974 ();
 sg13g2_fill_2 FILLER_127_980 ();
 sg13g2_fill_4 FILLER_127_995 ();
 sg13g2_fill_2 FILLER_127_999 ();
 sg13g2_fill_1 FILLER_127_1001 ();
 sg13g2_fill_2 FILLER_127_1028 ();
 sg13g2_fill_1 FILLER_127_1030 ();
 sg13g2_fill_4 FILLER_127_1047 ();
 sg13g2_fill_2 FILLER_127_1051 ();
 sg13g2_fill_1 FILLER_127_1053 ();
 sg13g2_fill_1 FILLER_127_1075 ();
 sg13g2_fill_2 FILLER_127_1097 ();
 sg13g2_fill_8 FILLER_127_1104 ();
 sg13g2_fill_4 FILLER_127_1112 ();
 sg13g2_fill_2 FILLER_127_1116 ();
 sg13g2_fill_8 FILLER_127_1145 ();
 sg13g2_fill_4 FILLER_127_1153 ();
 sg13g2_fill_4 FILLER_127_1167 ();
 sg13g2_fill_1 FILLER_127_1171 ();
 sg13g2_fill_8 FILLER_127_1190 ();
 sg13g2_fill_1 FILLER_127_1213 ();
 sg13g2_fill_4 FILLER_127_1224 ();
 sg13g2_fill_8 FILLER_127_1233 ();
 sg13g2_fill_2 FILLER_127_1241 ();
 sg13g2_fill_1 FILLER_127_1243 ();
 sg13g2_fill_8 FILLER_127_1257 ();
 sg13g2_fill_8 FILLER_127_1265 ();
 sg13g2_fill_1 FILLER_127_1273 ();
 sg13g2_fill_4 FILLER_127_1292 ();
 sg13g2_fill_2 FILLER_127_1296 ();
 sg13g2_fill_1 FILLER_127_1298 ();
 sg13g2_fill_1 FILLER_127_1338 ();
 sg13g2_fill_2 FILLER_127_1344 ();
 sg13g2_fill_1 FILLER_127_1363 ();
 sg13g2_fill_2 FILLER_127_1388 ();
 sg13g2_fill_8 FILLER_127_1400 ();
 sg13g2_fill_4 FILLER_127_1408 ();
 sg13g2_fill_2 FILLER_127_1412 ();
 sg13g2_fill_1 FILLER_127_1414 ();
 sg13g2_fill_2 FILLER_127_1420 ();
 sg13g2_fill_1 FILLER_127_1426 ();
 sg13g2_fill_4 FILLER_127_1436 ();
 sg13g2_fill_1 FILLER_127_1440 ();
 sg13g2_fill_2 FILLER_127_1449 ();
 sg13g2_fill_1 FILLER_127_1456 ();
 sg13g2_fill_2 FILLER_127_1487 ();
 sg13g2_fill_1 FILLER_127_1489 ();
 sg13g2_fill_1 FILLER_127_1516 ();
 sg13g2_fill_4 FILLER_127_1522 ();
 sg13g2_fill_2 FILLER_127_1526 ();
 sg13g2_fill_1 FILLER_127_1528 ();
 sg13g2_fill_2 FILLER_127_1554 ();
 sg13g2_fill_8 FILLER_127_1567 ();
 sg13g2_fill_2 FILLER_127_1575 ();
 sg13g2_fill_4 FILLER_127_1588 ();
 sg13g2_fill_4 FILLER_128_0 ();
 sg13g2_fill_2 FILLER_128_4 ();
 sg13g2_fill_4 FILLER_128_11 ();
 sg13g2_fill_2 FILLER_128_15 ();
 sg13g2_fill_8 FILLER_128_37 ();
 sg13g2_fill_2 FILLER_128_45 ();
 sg13g2_fill_4 FILLER_128_51 ();
 sg13g2_fill_2 FILLER_128_55 ();
 sg13g2_fill_8 FILLER_128_62 ();
 sg13g2_fill_8 FILLER_128_70 ();
 sg13g2_fill_8 FILLER_128_78 ();
 sg13g2_fill_1 FILLER_128_86 ();
 sg13g2_fill_1 FILLER_128_95 ();
 sg13g2_fill_4 FILLER_128_105 ();
 sg13g2_fill_2 FILLER_128_109 ();
 sg13g2_fill_1 FILLER_128_137 ();
 sg13g2_fill_8 FILLER_128_184 ();
 sg13g2_fill_8 FILLER_128_192 ();
 sg13g2_fill_4 FILLER_128_200 ();
 sg13g2_fill_1 FILLER_128_204 ();
 sg13g2_fill_2 FILLER_128_215 ();
 sg13g2_fill_1 FILLER_128_217 ();
 sg13g2_fill_2 FILLER_128_239 ();
 sg13g2_fill_1 FILLER_128_241 ();
 sg13g2_fill_8 FILLER_128_268 ();
 sg13g2_fill_8 FILLER_128_286 ();
 sg13g2_fill_4 FILLER_128_294 ();
 sg13g2_fill_1 FILLER_128_298 ();
 sg13g2_fill_4 FILLER_128_325 ();
 sg13g2_fill_2 FILLER_128_329 ();
 sg13g2_fill_1 FILLER_128_331 ();
 sg13g2_fill_2 FILLER_128_364 ();
 sg13g2_fill_2 FILLER_128_418 ();
 sg13g2_fill_1 FILLER_128_420 ();
 sg13g2_fill_8 FILLER_128_452 ();
 sg13g2_fill_1 FILLER_128_460 ();
 sg13g2_fill_8 FILLER_128_471 ();
 sg13g2_fill_4 FILLER_128_479 ();
 sg13g2_fill_8 FILLER_128_493 ();
 sg13g2_fill_4 FILLER_128_501 ();
 sg13g2_fill_2 FILLER_128_505 ();
 sg13g2_fill_1 FILLER_128_507 ();
 sg13g2_fill_2 FILLER_128_556 ();
 sg13g2_fill_8 FILLER_128_593 ();
 sg13g2_fill_8 FILLER_128_601 ();
 sg13g2_fill_4 FILLER_128_609 ();
 sg13g2_fill_2 FILLER_128_613 ();
 sg13g2_fill_1 FILLER_128_615 ();
 sg13g2_fill_8 FILLER_128_621 ();
 sg13g2_fill_4 FILLER_128_629 ();
 sg13g2_fill_2 FILLER_128_633 ();
 sg13g2_fill_8 FILLER_128_640 ();
 sg13g2_fill_8 FILLER_128_648 ();
 sg13g2_fill_1 FILLER_128_656 ();
 sg13g2_fill_8 FILLER_128_673 ();
 sg13g2_fill_8 FILLER_128_681 ();
 sg13g2_fill_8 FILLER_128_689 ();
 sg13g2_fill_8 FILLER_128_697 ();
 sg13g2_fill_8 FILLER_128_705 ();
 sg13g2_fill_8 FILLER_128_713 ();
 sg13g2_fill_8 FILLER_128_721 ();
 sg13g2_fill_8 FILLER_128_729 ();
 sg13g2_fill_4 FILLER_128_737 ();
 sg13g2_fill_2 FILLER_128_741 ();
 sg13g2_fill_8 FILLER_128_768 ();
 sg13g2_fill_8 FILLER_128_776 ();
 sg13g2_fill_8 FILLER_128_784 ();
 sg13g2_fill_8 FILLER_128_792 ();
 sg13g2_fill_2 FILLER_128_800 ();
 sg13g2_fill_1 FILLER_128_802 ();
 sg13g2_fill_4 FILLER_128_811 ();
 sg13g2_fill_2 FILLER_128_823 ();
 sg13g2_fill_8 FILLER_128_851 ();
 sg13g2_fill_1 FILLER_128_859 ();
 sg13g2_fill_4 FILLER_128_870 ();
 sg13g2_fill_2 FILLER_128_874 ();
 sg13g2_fill_1 FILLER_128_876 ();
 sg13g2_fill_8 FILLER_128_887 ();
 sg13g2_fill_8 FILLER_128_895 ();
 sg13g2_fill_2 FILLER_128_903 ();
 sg13g2_fill_1 FILLER_128_905 ();
 sg13g2_fill_2 FILLER_128_927 ();
 sg13g2_fill_8 FILLER_128_934 ();
 sg13g2_fill_2 FILLER_128_942 ();
 sg13g2_fill_1 FILLER_128_944 ();
 sg13g2_fill_2 FILLER_128_971 ();
 sg13g2_fill_1 FILLER_128_980 ();
 sg13g2_fill_8 FILLER_128_996 ();
 sg13g2_fill_8 FILLER_128_1004 ();
 sg13g2_fill_1 FILLER_128_1012 ();
 sg13g2_fill_4 FILLER_128_1018 ();
 sg13g2_fill_1 FILLER_128_1022 ();
 sg13g2_fill_2 FILLER_128_1028 ();
 sg13g2_fill_4 FILLER_128_1043 ();
 sg13g2_fill_2 FILLER_128_1047 ();
 sg13g2_fill_8 FILLER_128_1052 ();
 sg13g2_fill_2 FILLER_128_1060 ();
 sg13g2_fill_1 FILLER_128_1062 ();
 sg13g2_fill_2 FILLER_128_1069 ();
 sg13g2_fill_8 FILLER_128_1076 ();
 sg13g2_fill_1 FILLER_128_1084 ();
 sg13g2_fill_2 FILLER_128_1091 ();
 sg13g2_fill_1 FILLER_128_1093 ();
 sg13g2_fill_1 FILLER_128_1107 ();
 sg13g2_fill_2 FILLER_128_1114 ();
 sg13g2_fill_1 FILLER_128_1116 ();
 sg13g2_fill_4 FILLER_128_1147 ();
 sg13g2_fill_8 FILLER_128_1160 ();
 sg13g2_fill_8 FILLER_128_1168 ();
 sg13g2_fill_1 FILLER_128_1176 ();
 sg13g2_fill_2 FILLER_128_1182 ();
 sg13g2_fill_8 FILLER_128_1196 ();
 sg13g2_fill_8 FILLER_128_1204 ();
 sg13g2_fill_2 FILLER_128_1212 ();
 sg13g2_fill_8 FILLER_128_1225 ();
 sg13g2_fill_4 FILLER_128_1238 ();
 sg13g2_fill_2 FILLER_128_1242 ();
 sg13g2_fill_8 FILLER_128_1256 ();
 sg13g2_fill_8 FILLER_128_1269 ();
 sg13g2_fill_2 FILLER_128_1277 ();
 sg13g2_fill_8 FILLER_128_1284 ();
 sg13g2_fill_8 FILLER_128_1292 ();
 sg13g2_fill_2 FILLER_128_1300 ();
 sg13g2_fill_1 FILLER_128_1307 ();
 sg13g2_fill_4 FILLER_128_1314 ();
 sg13g2_fill_1 FILLER_128_1318 ();
 sg13g2_fill_2 FILLER_128_1324 ();
 sg13g2_fill_1 FILLER_128_1326 ();
 sg13g2_fill_1 FILLER_128_1342 ();
 sg13g2_fill_1 FILLER_128_1365 ();
 sg13g2_fill_4 FILLER_128_1377 ();
 sg13g2_fill_2 FILLER_128_1381 ();
 sg13g2_fill_1 FILLER_128_1383 ();
 sg13g2_fill_2 FILLER_128_1396 ();
 sg13g2_fill_1 FILLER_128_1398 ();
 sg13g2_fill_2 FILLER_128_1403 ();
 sg13g2_fill_1 FILLER_128_1405 ();
 sg13g2_fill_1 FILLER_128_1422 ();
 sg13g2_fill_2 FILLER_128_1427 ();
 sg13g2_fill_1 FILLER_128_1521 ();
 sg13g2_fill_2 FILLER_128_1589 ();
 sg13g2_fill_1 FILLER_128_1591 ();
 sg13g2_fill_4 FILLER_129_0 ();
 sg13g2_fill_1 FILLER_129_4 ();
 sg13g2_fill_1 FILLER_129_50 ();
 sg13g2_fill_2 FILLER_129_84 ();
 sg13g2_fill_2 FILLER_129_92 ();
 sg13g2_fill_1 FILLER_129_99 ();
 sg13g2_fill_8 FILLER_129_110 ();
 sg13g2_fill_8 FILLER_129_118 ();
 sg13g2_fill_1 FILLER_129_126 ();
 sg13g2_fill_8 FILLER_129_131 ();
 sg13g2_fill_8 FILLER_129_139 ();
 sg13g2_fill_4 FILLER_129_147 ();
 sg13g2_fill_1 FILLER_129_151 ();
 sg13g2_fill_1 FILLER_129_195 ();
 sg13g2_fill_4 FILLER_129_243 ();
 sg13g2_fill_2 FILLER_129_247 ();
 sg13g2_fill_4 FILLER_129_259 ();
 sg13g2_fill_2 FILLER_129_263 ();
 sg13g2_fill_1 FILLER_129_265 ();
 sg13g2_fill_8 FILLER_129_287 ();
 sg13g2_fill_4 FILLER_129_295 ();
 sg13g2_fill_2 FILLER_129_299 ();
 sg13g2_fill_1 FILLER_129_301 ();
 sg13g2_fill_8 FILLER_129_312 ();
 sg13g2_fill_4 FILLER_129_320 ();
 sg13g2_fill_4 FILLER_129_345 ();
 sg13g2_fill_2 FILLER_129_349 ();
 sg13g2_fill_1 FILLER_129_351 ();
 sg13g2_fill_2 FILLER_129_375 ();
 sg13g2_fill_4 FILLER_129_387 ();
 sg13g2_fill_8 FILLER_129_447 ();
 sg13g2_fill_2 FILLER_129_455 ();
 sg13g2_fill_1 FILLER_129_457 ();
 sg13g2_fill_8 FILLER_129_468 ();
 sg13g2_fill_4 FILLER_129_476 ();
 sg13g2_fill_2 FILLER_129_480 ();
 sg13g2_fill_1 FILLER_129_482 ();
 sg13g2_fill_8 FILLER_129_509 ();
 sg13g2_fill_8 FILLER_129_517 ();
 sg13g2_fill_4 FILLER_129_525 ();
 sg13g2_fill_1 FILLER_129_529 ();
 sg13g2_fill_2 FILLER_129_576 ();
 sg13g2_fill_1 FILLER_129_578 ();
 sg13g2_fill_2 FILLER_129_597 ();
 sg13g2_fill_1 FILLER_129_599 ();
 sg13g2_fill_8 FILLER_129_606 ();
 sg13g2_fill_4 FILLER_129_614 ();
 sg13g2_fill_2 FILLER_129_618 ();
 sg13g2_fill_1 FILLER_129_620 ();
 sg13g2_fill_4 FILLER_129_655 ();
 sg13g2_fill_2 FILLER_129_659 ();
 sg13g2_fill_1 FILLER_129_661 ();
 sg13g2_fill_2 FILLER_129_672 ();
 sg13g2_fill_1 FILLER_129_674 ();
 sg13g2_fill_8 FILLER_129_711 ();
 sg13g2_fill_2 FILLER_129_729 ();
 sg13g2_fill_2 FILLER_129_760 ();
 sg13g2_fill_1 FILLER_129_762 ();
 sg13g2_fill_8 FILLER_129_771 ();
 sg13g2_fill_1 FILLER_129_779 ();
 sg13g2_fill_8 FILLER_129_806 ();
 sg13g2_fill_4 FILLER_129_814 ();
 sg13g2_fill_1 FILLER_129_818 ();
 sg13g2_fill_8 FILLER_129_829 ();
 sg13g2_fill_8 FILLER_129_837 ();
 sg13g2_fill_1 FILLER_129_845 ();
 sg13g2_fill_8 FILLER_129_902 ();
 sg13g2_fill_8 FILLER_129_910 ();
 sg13g2_fill_2 FILLER_129_918 ();
 sg13g2_fill_8 FILLER_129_925 ();
 sg13g2_fill_1 FILLER_129_933 ();
 sg13g2_fill_1 FILLER_129_943 ();
 sg13g2_fill_4 FILLER_129_948 ();
 sg13g2_fill_1 FILLER_129_952 ();
 sg13g2_fill_8 FILLER_129_970 ();
 sg13g2_fill_1 FILLER_129_978 ();
 sg13g2_fill_8 FILLER_129_985 ();
 sg13g2_fill_4 FILLER_129_993 ();
 sg13g2_fill_2 FILLER_129_997 ();
 sg13g2_fill_1 FILLER_129_999 ();
 sg13g2_fill_2 FILLER_129_1009 ();
 sg13g2_fill_1 FILLER_129_1011 ();
 sg13g2_fill_8 FILLER_129_1032 ();
 sg13g2_fill_4 FILLER_129_1040 ();
 sg13g2_fill_2 FILLER_129_1044 ();
 sg13g2_fill_1 FILLER_129_1052 ();
 sg13g2_fill_8 FILLER_129_1067 ();
 sg13g2_fill_4 FILLER_129_1075 ();
 sg13g2_fill_2 FILLER_129_1079 ();
 sg13g2_fill_1 FILLER_129_1087 ();
 sg13g2_fill_4 FILLER_129_1106 ();
 sg13g2_fill_1 FILLER_129_1110 ();
 sg13g2_fill_8 FILLER_129_1117 ();
 sg13g2_fill_8 FILLER_129_1125 ();
 sg13g2_fill_8 FILLER_129_1133 ();
 sg13g2_fill_8 FILLER_129_1141 ();
 sg13g2_fill_8 FILLER_129_1149 ();
 sg13g2_fill_4 FILLER_129_1157 ();
 sg13g2_fill_2 FILLER_129_1161 ();
 sg13g2_fill_1 FILLER_129_1163 ();
 sg13g2_fill_8 FILLER_129_1173 ();
 sg13g2_fill_1 FILLER_129_1181 ();
 sg13g2_fill_8 FILLER_129_1188 ();
 sg13g2_fill_1 FILLER_129_1196 ();
 sg13g2_fill_2 FILLER_129_1227 ();
 sg13g2_fill_2 FILLER_129_1259 ();
 sg13g2_fill_1 FILLER_129_1261 ();
 sg13g2_fill_2 FILLER_129_1292 ();
 sg13g2_fill_1 FILLER_129_1299 ();
 sg13g2_fill_1 FILLER_129_1305 ();
 sg13g2_fill_8 FILLER_129_1311 ();
 sg13g2_fill_2 FILLER_129_1319 ();
 sg13g2_fill_1 FILLER_129_1321 ();
 sg13g2_fill_1 FILLER_129_1332 ();
 sg13g2_fill_1 FILLER_129_1339 ();
 sg13g2_fill_2 FILLER_129_1375 ();
 sg13g2_fill_1 FILLER_129_1377 ();
 sg13g2_fill_1 FILLER_129_1386 ();
 sg13g2_fill_8 FILLER_129_1416 ();
 sg13g2_fill_2 FILLER_129_1448 ();
 sg13g2_fill_2 FILLER_129_1465 ();
 sg13g2_fill_4 FILLER_129_1472 ();
 sg13g2_fill_1 FILLER_129_1476 ();
 sg13g2_fill_8 FILLER_129_1486 ();
 sg13g2_fill_8 FILLER_129_1494 ();
 sg13g2_fill_1 FILLER_129_1502 ();
 sg13g2_fill_1 FILLER_129_1556 ();
 sg13g2_fill_8 FILLER_129_1567 ();
 sg13g2_fill_4 FILLER_129_1586 ();
 sg13g2_fill_2 FILLER_129_1590 ();
 sg13g2_fill_4 FILLER_130_0 ();
 sg13g2_fill_2 FILLER_130_67 ();
 sg13g2_fill_8 FILLER_130_81 ();
 sg13g2_fill_2 FILLER_130_89 ();
 sg13g2_fill_1 FILLER_130_91 ();
 sg13g2_fill_8 FILLER_130_102 ();
 sg13g2_fill_4 FILLER_130_110 ();
 sg13g2_fill_2 FILLER_130_114 ();
 sg13g2_fill_2 FILLER_130_145 ();
 sg13g2_fill_1 FILLER_130_147 ();
 sg13g2_fill_8 FILLER_130_182 ();
 sg13g2_fill_8 FILLER_130_190 ();
 sg13g2_fill_8 FILLER_130_198 ();
 sg13g2_fill_8 FILLER_130_206 ();
 sg13g2_fill_4 FILLER_130_214 ();
 sg13g2_fill_2 FILLER_130_218 ();
 sg13g2_fill_1 FILLER_130_220 ();
 sg13g2_fill_4 FILLER_130_231 ();
 sg13g2_fill_2 FILLER_130_243 ();
 sg13g2_fill_1 FILLER_130_245 ();
 sg13g2_fill_2 FILLER_130_300 ();
 sg13g2_fill_1 FILLER_130_302 ();
 sg13g2_fill_8 FILLER_130_329 ();
 sg13g2_fill_8 FILLER_130_337 ();
 sg13g2_fill_8 FILLER_130_345 ();
 sg13g2_fill_4 FILLER_130_353 ();
 sg13g2_fill_2 FILLER_130_357 ();
 sg13g2_fill_8 FILLER_130_395 ();
 sg13g2_fill_8 FILLER_130_403 ();
 sg13g2_fill_8 FILLER_130_411 ();
 sg13g2_fill_8 FILLER_130_419 ();
 sg13g2_fill_4 FILLER_130_427 ();
 sg13g2_fill_1 FILLER_130_431 ();
 sg13g2_fill_8 FILLER_130_442 ();
 sg13g2_fill_8 FILLER_130_450 ();
 sg13g2_fill_8 FILLER_130_458 ();
 sg13g2_fill_2 FILLER_130_466 ();
 sg13g2_fill_1 FILLER_130_486 ();
 sg13g2_fill_2 FILLER_130_497 ();
 sg13g2_fill_4 FILLER_130_507 ();
 sg13g2_fill_1 FILLER_130_521 ();
 sg13g2_fill_8 FILLER_130_549 ();
 sg13g2_fill_8 FILLER_130_557 ();
 sg13g2_fill_8 FILLER_130_565 ();
 sg13g2_fill_4 FILLER_130_573 ();
 sg13g2_fill_1 FILLER_130_582 ();
 sg13g2_fill_8 FILLER_130_603 ();
 sg13g2_fill_8 FILLER_130_611 ();
 sg13g2_fill_4 FILLER_130_619 ();
 sg13g2_fill_2 FILLER_130_623 ();
 sg13g2_fill_1 FILLER_130_625 ();
 sg13g2_fill_8 FILLER_130_636 ();
 sg13g2_fill_4 FILLER_130_644 ();
 sg13g2_fill_1 FILLER_130_648 ();
 sg13g2_fill_8 FILLER_130_669 ();
 sg13g2_fill_4 FILLER_130_677 ();
 sg13g2_fill_2 FILLER_130_681 ();
 sg13g2_fill_4 FILLER_130_709 ();
 sg13g2_fill_2 FILLER_130_713 ();
 sg13g2_fill_1 FILLER_130_715 ();
 sg13g2_fill_1 FILLER_130_742 ();
 sg13g2_fill_8 FILLER_130_751 ();
 sg13g2_fill_2 FILLER_130_759 ();
 sg13g2_fill_2 FILLER_130_782 ();
 sg13g2_fill_4 FILLER_130_840 ();
 sg13g2_fill_1 FILLER_130_844 ();
 sg13g2_fill_4 FILLER_130_861 ();
 sg13g2_fill_1 FILLER_130_865 ();
 sg13g2_fill_4 FILLER_130_871 ();
 sg13g2_fill_1 FILLER_130_875 ();
 sg13g2_fill_8 FILLER_130_882 ();
 sg13g2_fill_8 FILLER_130_890 ();
 sg13g2_fill_2 FILLER_130_898 ();
 sg13g2_fill_2 FILLER_130_906 ();
 sg13g2_fill_1 FILLER_130_908 ();
 sg13g2_fill_8 FILLER_130_918 ();
 sg13g2_fill_1 FILLER_130_926 ();
 sg13g2_fill_8 FILLER_130_936 ();
 sg13g2_fill_2 FILLER_130_944 ();
 sg13g2_fill_1 FILLER_130_946 ();
 sg13g2_fill_8 FILLER_130_951 ();
 sg13g2_fill_8 FILLER_130_959 ();
 sg13g2_fill_1 FILLER_130_967 ();
 sg13g2_fill_8 FILLER_130_973 ();
 sg13g2_fill_4 FILLER_130_981 ();
 sg13g2_fill_1 FILLER_130_985 ();
 sg13g2_fill_1 FILLER_130_998 ();
 sg13g2_fill_1 FILLER_130_1003 ();
 sg13g2_fill_1 FILLER_130_1034 ();
 sg13g2_fill_2 FILLER_130_1055 ();
 sg13g2_fill_1 FILLER_130_1061 ();
 sg13g2_fill_1 FILLER_130_1066 ();
 sg13g2_fill_8 FILLER_130_1077 ();
 sg13g2_fill_4 FILLER_130_1085 ();
 sg13g2_fill_2 FILLER_130_1089 ();
 sg13g2_fill_2 FILLER_130_1100 ();
 sg13g2_fill_1 FILLER_130_1102 ();
 sg13g2_fill_1 FILLER_130_1111 ();
 sg13g2_fill_8 FILLER_130_1124 ();
 sg13g2_fill_2 FILLER_130_1146 ();
 sg13g2_fill_8 FILLER_130_1178 ();
 sg13g2_fill_2 FILLER_130_1186 ();
 sg13g2_fill_1 FILLER_130_1188 ();
 sg13g2_fill_4 FILLER_130_1205 ();
 sg13g2_fill_2 FILLER_130_1209 ();
 sg13g2_fill_8 FILLER_130_1219 ();
 sg13g2_fill_8 FILLER_130_1236 ();
 sg13g2_fill_2 FILLER_130_1258 ();
 sg13g2_fill_1 FILLER_130_1260 ();
 sg13g2_fill_8 FILLER_130_1266 ();
 sg13g2_fill_4 FILLER_130_1274 ();
 sg13g2_fill_4 FILLER_130_1314 ();
 sg13g2_fill_2 FILLER_130_1318 ();
 sg13g2_fill_1 FILLER_130_1320 ();
 sg13g2_fill_4 FILLER_130_1326 ();
 sg13g2_fill_2 FILLER_130_1330 ();
 sg13g2_fill_1 FILLER_130_1332 ();
 sg13g2_fill_1 FILLER_130_1346 ();
 sg13g2_fill_1 FILLER_130_1372 ();
 sg13g2_fill_2 FILLER_130_1378 ();
 sg13g2_fill_2 FILLER_130_1387 ();
 sg13g2_fill_1 FILLER_130_1389 ();
 sg13g2_fill_4 FILLER_130_1395 ();
 sg13g2_fill_2 FILLER_130_1399 ();
 sg13g2_fill_8 FILLER_130_1405 ();
 sg13g2_fill_4 FILLER_130_1413 ();
 sg13g2_fill_2 FILLER_130_1417 ();
 sg13g2_fill_1 FILLER_130_1429 ();
 sg13g2_fill_4 FILLER_130_1455 ();
 sg13g2_fill_2 FILLER_130_1459 ();
 sg13g2_fill_2 FILLER_130_1466 ();
 sg13g2_fill_1 FILLER_130_1468 ();
 sg13g2_fill_8 FILLER_130_1500 ();
 sg13g2_fill_4 FILLER_130_1508 ();
 sg13g2_fill_2 FILLER_130_1512 ();
 sg13g2_fill_1 FILLER_130_1514 ();
 sg13g2_fill_4 FILLER_130_1528 ();
 sg13g2_fill_1 FILLER_130_1532 ();
 sg13g2_fill_1 FILLER_130_1543 ();
 sg13g2_fill_8 FILLER_130_1557 ();
 sg13g2_fill_1 FILLER_130_1565 ();
 sg13g2_fill_4 FILLER_130_1588 ();
 sg13g2_fill_2 FILLER_131_34 ();
 sg13g2_fill_8 FILLER_131_41 ();
 sg13g2_fill_8 FILLER_131_49 ();
 sg13g2_fill_2 FILLER_131_57 ();
 sg13g2_fill_1 FILLER_131_59 ();
 sg13g2_fill_1 FILLER_131_71 ();
 sg13g2_fill_4 FILLER_131_78 ();
 sg13g2_fill_2 FILLER_131_82 ();
 sg13g2_fill_1 FILLER_131_84 ();
 sg13g2_fill_2 FILLER_131_91 ();
 sg13g2_fill_1 FILLER_131_101 ();
 sg13g2_fill_8 FILLER_131_112 ();
 sg13g2_fill_8 FILLER_131_120 ();
 sg13g2_fill_4 FILLER_131_128 ();
 sg13g2_fill_1 FILLER_131_132 ();
 sg13g2_fill_4 FILLER_131_180 ();
 sg13g2_fill_2 FILLER_131_205 ();
 sg13g2_fill_1 FILLER_131_207 ();
 sg13g2_fill_4 FILLER_131_218 ();
 sg13g2_fill_1 FILLER_131_222 ();
 sg13g2_fill_2 FILLER_131_275 ();
 sg13g2_fill_1 FILLER_131_277 ();
 sg13g2_fill_2 FILLER_131_302 ();
 sg13g2_fill_1 FILLER_131_304 ();
 sg13g2_fill_8 FILLER_131_315 ();
 sg13g2_fill_8 FILLER_131_323 ();
 sg13g2_fill_1 FILLER_131_331 ();
 sg13g2_fill_2 FILLER_131_374 ();
 sg13g2_fill_1 FILLER_131_376 ();
 sg13g2_fill_4 FILLER_131_429 ();
 sg13g2_fill_4 FILLER_131_469 ();
 sg13g2_fill_8 FILLER_131_478 ();
 sg13g2_fill_2 FILLER_131_486 ();
 sg13g2_fill_8 FILLER_131_514 ();
 sg13g2_fill_1 FILLER_131_522 ();
 sg13g2_fill_4 FILLER_131_533 ();
 sg13g2_fill_4 FILLER_131_583 ();
 sg13g2_fill_1 FILLER_131_587 ();
 sg13g2_fill_8 FILLER_131_624 ();
 sg13g2_fill_8 FILLER_131_632 ();
 sg13g2_fill_8 FILLER_131_640 ();
 sg13g2_fill_1 FILLER_131_648 ();
 sg13g2_fill_8 FILLER_131_661 ();
 sg13g2_fill_4 FILLER_131_669 ();
 sg13g2_fill_1 FILLER_131_673 ();
 sg13g2_fill_8 FILLER_131_684 ();
 sg13g2_fill_8 FILLER_131_692 ();
 sg13g2_fill_8 FILLER_131_700 ();
 sg13g2_fill_1 FILLER_131_708 ();
 sg13g2_fill_4 FILLER_131_719 ();
 sg13g2_fill_2 FILLER_131_723 ();
 sg13g2_fill_1 FILLER_131_725 ();
 sg13g2_fill_8 FILLER_131_792 ();
 sg13g2_fill_8 FILLER_131_800 ();
 sg13g2_fill_8 FILLER_131_808 ();
 sg13g2_fill_4 FILLER_131_816 ();
 sg13g2_fill_2 FILLER_131_820 ();
 sg13g2_fill_1 FILLER_131_822 ();
 sg13g2_fill_8 FILLER_131_833 ();
 sg13g2_fill_1 FILLER_131_841 ();
 sg13g2_fill_8 FILLER_131_867 ();
 sg13g2_fill_8 FILLER_131_875 ();
 sg13g2_fill_1 FILLER_131_883 ();
 sg13g2_fill_4 FILLER_131_894 ();
 sg13g2_fill_1 FILLER_131_898 ();
 sg13g2_fill_8 FILLER_131_921 ();
 sg13g2_fill_1 FILLER_131_943 ();
 sg13g2_fill_4 FILLER_131_978 ();
 sg13g2_fill_8 FILLER_131_989 ();
 sg13g2_fill_1 FILLER_131_997 ();
 sg13g2_fill_8 FILLER_131_1006 ();
 sg13g2_fill_2 FILLER_131_1014 ();
 sg13g2_fill_1 FILLER_131_1016 ();
 sg13g2_fill_8 FILLER_131_1032 ();
 sg13g2_fill_4 FILLER_131_1040 ();
 sg13g2_fill_8 FILLER_131_1049 ();
 sg13g2_fill_8 FILLER_131_1057 ();
 sg13g2_fill_8 FILLER_131_1069 ();
 sg13g2_fill_1 FILLER_131_1077 ();
 sg13g2_fill_1 FILLER_131_1082 ();
 sg13g2_fill_1 FILLER_131_1093 ();
 sg13g2_fill_2 FILLER_131_1115 ();
 sg13g2_fill_1 FILLER_131_1117 ();
 sg13g2_fill_8 FILLER_131_1161 ();
 sg13g2_fill_4 FILLER_131_1169 ();
 sg13g2_fill_2 FILLER_131_1173 ();
 sg13g2_fill_8 FILLER_131_1185 ();
 sg13g2_fill_8 FILLER_131_1213 ();
 sg13g2_fill_8 FILLER_131_1221 ();
 sg13g2_fill_4 FILLER_131_1229 ();
 sg13g2_fill_1 FILLER_131_1233 ();
 sg13g2_fill_2 FILLER_131_1276 ();
 sg13g2_fill_2 FILLER_131_1283 ();
 sg13g2_fill_1 FILLER_131_1285 ();
 sg13g2_fill_2 FILLER_131_1327 ();
 sg13g2_fill_1 FILLER_131_1346 ();
 sg13g2_fill_2 FILLER_131_1375 ();
 sg13g2_fill_1 FILLER_131_1377 ();
 sg13g2_fill_1 FILLER_131_1383 ();
 sg13g2_fill_2 FILLER_131_1399 ();
 sg13g2_fill_1 FILLER_131_1401 ();
 sg13g2_fill_4 FILLER_131_1414 ();
 sg13g2_fill_2 FILLER_131_1418 ();
 sg13g2_fill_1 FILLER_131_1429 ();
 sg13g2_fill_2 FILLER_131_1465 ();
 sg13g2_fill_1 FILLER_131_1467 ();
 sg13g2_fill_2 FILLER_131_1494 ();
 sg13g2_fill_1 FILLER_131_1496 ();
 sg13g2_fill_2 FILLER_131_1512 ();
 sg13g2_fill_1 FILLER_131_1535 ();
 sg13g2_fill_1 FILLER_131_1547 ();
 sg13g2_fill_2 FILLER_131_1574 ();
 sg13g2_fill_1 FILLER_131_1576 ();
 sg13g2_fill_4 FILLER_131_1588 ();
 sg13g2_fill_8 FILLER_132_0 ();
 sg13g2_fill_4 FILLER_132_8 ();
 sg13g2_fill_2 FILLER_132_12 ();
 sg13g2_fill_4 FILLER_132_30 ();
 sg13g2_fill_2 FILLER_132_34 ();
 sg13g2_fill_8 FILLER_132_50 ();
 sg13g2_fill_4 FILLER_132_58 ();
 sg13g2_fill_1 FILLER_132_62 ();
 sg13g2_fill_2 FILLER_132_68 ();
 sg13g2_fill_1 FILLER_132_70 ();
 sg13g2_fill_2 FILLER_132_88 ();
 sg13g2_fill_1 FILLER_132_96 ();
 sg13g2_fill_4 FILLER_132_133 ();
 sg13g2_fill_1 FILLER_132_137 ();
 sg13g2_fill_8 FILLER_132_141 ();
 sg13g2_fill_8 FILLER_132_149 ();
 sg13g2_fill_2 FILLER_132_157 ();
 sg13g2_fill_8 FILLER_132_185 ();
 sg13g2_fill_8 FILLER_132_193 ();
 sg13g2_fill_2 FILLER_132_201 ();
 sg13g2_fill_4 FILLER_132_229 ();
 sg13g2_fill_2 FILLER_132_233 ();
 sg13g2_fill_1 FILLER_132_235 ();
 sg13g2_fill_8 FILLER_132_244 ();
 sg13g2_fill_8 FILLER_132_252 ();
 sg13g2_fill_8 FILLER_132_260 ();
 sg13g2_fill_8 FILLER_132_268 ();
 sg13g2_fill_8 FILLER_132_276 ();
 sg13g2_fill_8 FILLER_132_284 ();
 sg13g2_fill_8 FILLER_132_292 ();
 sg13g2_fill_8 FILLER_132_300 ();
 sg13g2_fill_8 FILLER_132_308 ();
 sg13g2_fill_8 FILLER_132_316 ();
 sg13g2_fill_8 FILLER_132_324 ();
 sg13g2_fill_4 FILLER_132_332 ();
 sg13g2_fill_8 FILLER_132_346 ();
 sg13g2_fill_8 FILLER_132_354 ();
 sg13g2_fill_8 FILLER_132_362 ();
 sg13g2_fill_8 FILLER_132_370 ();
 sg13g2_fill_8 FILLER_132_378 ();
 sg13g2_fill_8 FILLER_132_386 ();
 sg13g2_fill_1 FILLER_132_394 ();
 sg13g2_fill_4 FILLER_132_431 ();
 sg13g2_fill_2 FILLER_132_435 ();
 sg13g2_fill_4 FILLER_132_472 ();
 sg13g2_fill_1 FILLER_132_476 ();
 sg13g2_fill_8 FILLER_132_485 ();
 sg13g2_fill_8 FILLER_132_493 ();
 sg13g2_fill_2 FILLER_132_501 ();
 sg13g2_fill_1 FILLER_132_503 ();
 sg13g2_fill_8 FILLER_132_514 ();
 sg13g2_fill_4 FILLER_132_522 ();
 sg13g2_fill_2 FILLER_132_526 ();
 sg13g2_fill_1 FILLER_132_528 ();
 sg13g2_fill_8 FILLER_132_546 ();
 sg13g2_fill_8 FILLER_132_554 ();
 sg13g2_fill_8 FILLER_132_562 ();
 sg13g2_fill_2 FILLER_132_570 ();
 sg13g2_fill_8 FILLER_132_598 ();
 sg13g2_fill_4 FILLER_132_606 ();
 sg13g2_fill_2 FILLER_132_610 ();
 sg13g2_fill_1 FILLER_132_612 ();
 sg13g2_fill_2 FILLER_132_639 ();
 sg13g2_fill_1 FILLER_132_641 ();
 sg13g2_fill_2 FILLER_132_663 ();
 sg13g2_fill_8 FILLER_132_675 ();
 sg13g2_fill_1 FILLER_132_683 ();
 sg13g2_fill_2 FILLER_132_710 ();
 sg13g2_fill_4 FILLER_132_747 ();
 sg13g2_fill_1 FILLER_132_751 ();
 sg13g2_fill_8 FILLER_132_757 ();
 sg13g2_fill_1 FILLER_132_765 ();
 sg13g2_fill_1 FILLER_132_827 ();
 sg13g2_fill_1 FILLER_132_889 ();
 sg13g2_fill_8 FILLER_132_900 ();
 sg13g2_fill_4 FILLER_132_908 ();
 sg13g2_fill_1 FILLER_132_912 ();
 sg13g2_fill_1 FILLER_132_937 ();
 sg13g2_fill_8 FILLER_132_947 ();
 sg13g2_fill_8 FILLER_132_955 ();
 sg13g2_fill_2 FILLER_132_963 ();
 sg13g2_fill_1 FILLER_132_965 ();
 sg13g2_fill_8 FILLER_132_973 ();
 sg13g2_fill_2 FILLER_132_981 ();
 sg13g2_fill_8 FILLER_132_1008 ();
 sg13g2_fill_8 FILLER_132_1016 ();
 sg13g2_fill_8 FILLER_132_1024 ();
 sg13g2_fill_8 FILLER_132_1032 ();
 sg13g2_fill_8 FILLER_132_1040 ();
 sg13g2_fill_2 FILLER_132_1054 ();
 sg13g2_fill_2 FILLER_132_1075 ();
 sg13g2_fill_2 FILLER_132_1081 ();
 sg13g2_fill_1 FILLER_132_1133 ();
 sg13g2_fill_8 FILLER_132_1143 ();
 sg13g2_fill_1 FILLER_132_1151 ();
 sg13g2_fill_8 FILLER_132_1186 ();
 sg13g2_fill_2 FILLER_132_1194 ();
 sg13g2_fill_1 FILLER_132_1196 ();
 sg13g2_fill_2 FILLER_132_1227 ();
 sg13g2_fill_2 FILLER_132_1234 ();
 sg13g2_fill_1 FILLER_132_1236 ();
 sg13g2_fill_2 FILLER_132_1242 ();
 sg13g2_fill_4 FILLER_132_1285 ();
 sg13g2_fill_2 FILLER_132_1301 ();
 sg13g2_fill_2 FILLER_132_1316 ();
 sg13g2_fill_2 FILLER_132_1322 ();
 sg13g2_fill_8 FILLER_132_1329 ();
 sg13g2_fill_2 FILLER_132_1337 ();
 sg13g2_fill_1 FILLER_132_1352 ();
 sg13g2_fill_2 FILLER_132_1358 ();
 sg13g2_fill_4 FILLER_132_1370 ();
 sg13g2_fill_2 FILLER_132_1379 ();
 sg13g2_fill_2 FILLER_132_1399 ();
 sg13g2_fill_1 FILLER_132_1401 ();
 sg13g2_fill_4 FILLER_132_1417 ();
 sg13g2_fill_2 FILLER_132_1421 ();
 sg13g2_fill_8 FILLER_132_1428 ();
 sg13g2_fill_2 FILLER_132_1440 ();
 sg13g2_fill_1 FILLER_132_1446 ();
 sg13g2_fill_8 FILLER_132_1452 ();
 sg13g2_fill_4 FILLER_132_1460 ();
 sg13g2_fill_2 FILLER_132_1464 ();
 sg13g2_fill_1 FILLER_132_1466 ();
 sg13g2_fill_8 FILLER_132_1480 ();
 sg13g2_fill_8 FILLER_132_1488 ();
 sg13g2_fill_8 FILLER_132_1496 ();
 sg13g2_fill_4 FILLER_132_1509 ();
 sg13g2_fill_4 FILLER_132_1587 ();
 sg13g2_fill_1 FILLER_132_1591 ();
 sg13g2_fill_4 FILLER_133_0 ();
 sg13g2_fill_8 FILLER_133_14 ();
 sg13g2_fill_4 FILLER_133_22 ();
 sg13g2_fill_2 FILLER_133_26 ();
 sg13g2_fill_4 FILLER_133_43 ();
 sg13g2_fill_1 FILLER_133_47 ();
 sg13g2_fill_2 FILLER_133_58 ();
 sg13g2_fill_4 FILLER_133_74 ();
 sg13g2_fill_2 FILLER_133_78 ();
 sg13g2_fill_2 FILLER_133_101 ();
 sg13g2_fill_8 FILLER_133_113 ();
 sg13g2_fill_4 FILLER_133_121 ();
 sg13g2_fill_1 FILLER_133_125 ();
 sg13g2_fill_8 FILLER_133_146 ();
 sg13g2_fill_4 FILLER_133_154 ();
 sg13g2_fill_1 FILLER_133_158 ();
 sg13g2_fill_8 FILLER_133_164 ();
 sg13g2_fill_1 FILLER_133_172 ();
 sg13g2_fill_8 FILLER_133_204 ();
 sg13g2_fill_8 FILLER_133_212 ();
 sg13g2_fill_8 FILLER_133_220 ();
 sg13g2_fill_8 FILLER_133_228 ();
 sg13g2_fill_8 FILLER_133_236 ();
 sg13g2_fill_4 FILLER_133_244 ();
 sg13g2_fill_8 FILLER_133_274 ();
 sg13g2_fill_2 FILLER_133_282 ();
 sg13g2_fill_8 FILLER_133_289 ();
 sg13g2_fill_4 FILLER_133_297 ();
 sg13g2_fill_1 FILLER_133_301 ();
 sg13g2_fill_8 FILLER_133_328 ();
 sg13g2_fill_8 FILLER_133_368 ();
 sg13g2_fill_4 FILLER_133_376 ();
 sg13g2_fill_8 FILLER_133_415 ();
 sg13g2_fill_4 FILLER_133_423 ();
 sg13g2_fill_1 FILLER_133_427 ();
 sg13g2_fill_2 FILLER_133_464 ();
 sg13g2_fill_1 FILLER_133_466 ();
 sg13g2_fill_2 FILLER_133_474 ();
 sg13g2_fill_1 FILLER_133_476 ();
 sg13g2_fill_8 FILLER_133_495 ();
 sg13g2_fill_8 FILLER_133_503 ();
 sg13g2_fill_2 FILLER_133_511 ();
 sg13g2_fill_1 FILLER_133_513 ();
 sg13g2_fill_8 FILLER_133_524 ();
 sg13g2_fill_4 FILLER_133_532 ();
 sg13g2_fill_2 FILLER_133_536 ();
 sg13g2_fill_1 FILLER_133_538 ();
 sg13g2_fill_2 FILLER_133_544 ();
 sg13g2_fill_8 FILLER_133_550 ();
 sg13g2_fill_8 FILLER_133_558 ();
 sg13g2_fill_8 FILLER_133_576 ();
 sg13g2_fill_8 FILLER_133_584 ();
 sg13g2_fill_4 FILLER_133_592 ();
 sg13g2_fill_8 FILLER_133_601 ();
 sg13g2_fill_4 FILLER_133_609 ();
 sg13g2_fill_4 FILLER_133_621 ();
 sg13g2_fill_4 FILLER_133_635 ();
 sg13g2_fill_2 FILLER_133_639 ();
 sg13g2_fill_1 FILLER_133_641 ();
 sg13g2_fill_2 FILLER_133_663 ();
 sg13g2_fill_1 FILLER_133_685 ();
 sg13g2_fill_2 FILLER_133_696 ();
 sg13g2_fill_1 FILLER_133_698 ();
 sg13g2_fill_1 FILLER_133_725 ();
 sg13g2_fill_8 FILLER_133_752 ();
 sg13g2_fill_8 FILLER_133_760 ();
 sg13g2_fill_2 FILLER_133_768 ();
 sg13g2_fill_1 FILLER_133_770 ();
 sg13g2_fill_8 FILLER_133_801 ();
 sg13g2_fill_8 FILLER_133_809 ();
 sg13g2_fill_8 FILLER_133_817 ();
 sg13g2_fill_2 FILLER_133_825 ();
 sg13g2_fill_1 FILLER_133_827 ();
 sg13g2_fill_4 FILLER_133_838 ();
 sg13g2_fill_4 FILLER_133_845 ();
 sg13g2_fill_1 FILLER_133_849 ();
 sg13g2_fill_2 FILLER_133_855 ();
 sg13g2_fill_1 FILLER_133_857 ();
 sg13g2_fill_2 FILLER_133_868 ();
 sg13g2_fill_8 FILLER_133_875 ();
 sg13g2_fill_2 FILLER_133_883 ();
 sg13g2_fill_1 FILLER_133_885 ();
 sg13g2_fill_8 FILLER_133_895 ();
 sg13g2_fill_8 FILLER_133_903 ();
 sg13g2_fill_8 FILLER_133_911 ();
 sg13g2_fill_8 FILLER_133_919 ();
 sg13g2_fill_1 FILLER_133_927 ();
 sg13g2_fill_8 FILLER_133_949 ();
 sg13g2_fill_4 FILLER_133_957 ();
 sg13g2_fill_8 FILLER_133_969 ();
 sg13g2_fill_1 FILLER_133_977 ();
 sg13g2_fill_4 FILLER_133_994 ();
 sg13g2_fill_1 FILLER_133_998 ();
 sg13g2_fill_8 FILLER_133_1014 ();
 sg13g2_fill_8 FILLER_133_1022 ();
 sg13g2_fill_8 FILLER_133_1055 ();
 sg13g2_fill_4 FILLER_133_1063 ();
 sg13g2_fill_2 FILLER_133_1067 ();
 sg13g2_fill_2 FILLER_133_1074 ();
 sg13g2_fill_1 FILLER_133_1076 ();
 sg13g2_fill_4 FILLER_133_1133 ();
 sg13g2_fill_4 FILLER_133_1141 ();
 sg13g2_fill_1 FILLER_133_1145 ();
 sg13g2_fill_4 FILLER_133_1179 ();
 sg13g2_fill_1 FILLER_133_1183 ();
 sg13g2_fill_2 FILLER_133_1194 ();
 sg13g2_fill_1 FILLER_133_1202 ();
 sg13g2_fill_4 FILLER_133_1206 ();
 sg13g2_fill_2 FILLER_133_1210 ();
 sg13g2_fill_4 FILLER_133_1217 ();
 sg13g2_fill_2 FILLER_133_1221 ();
 sg13g2_fill_1 FILLER_133_1223 ();
 sg13g2_fill_2 FILLER_133_1241 ();
 sg13g2_fill_8 FILLER_133_1257 ();
 sg13g2_fill_4 FILLER_133_1265 ();
 sg13g2_fill_1 FILLER_133_1269 ();
 sg13g2_fill_8 FILLER_133_1273 ();
 sg13g2_fill_8 FILLER_133_1281 ();
 sg13g2_fill_2 FILLER_133_1289 ();
 sg13g2_fill_2 FILLER_133_1296 ();
 sg13g2_fill_4 FILLER_133_1310 ();
 sg13g2_fill_1 FILLER_133_1328 ();
 sg13g2_fill_4 FILLER_133_1337 ();
 sg13g2_fill_2 FILLER_133_1341 ();
 sg13g2_fill_1 FILLER_133_1343 ();
 sg13g2_fill_1 FILLER_133_1353 ();
 sg13g2_fill_2 FILLER_133_1377 ();
 sg13g2_fill_4 FILLER_133_1395 ();
 sg13g2_fill_2 FILLER_133_1399 ();
 sg13g2_fill_1 FILLER_133_1405 ();
 sg13g2_fill_8 FILLER_133_1419 ();
 sg13g2_fill_2 FILLER_133_1427 ();
 sg13g2_fill_1 FILLER_133_1429 ();
 sg13g2_fill_2 FILLER_133_1434 ();
 sg13g2_fill_8 FILLER_133_1462 ();
 sg13g2_fill_2 FILLER_133_1470 ();
 sg13g2_fill_8 FILLER_133_1481 ();
 sg13g2_fill_4 FILLER_133_1489 ();
 sg13g2_fill_1 FILLER_133_1493 ();
 sg13g2_fill_2 FILLER_133_1498 ();
 sg13g2_fill_2 FILLER_133_1506 ();
 sg13g2_fill_2 FILLER_133_1534 ();
 sg13g2_fill_1 FILLER_133_1536 ();
 sg13g2_fill_4 FILLER_133_1548 ();
 sg13g2_fill_1 FILLER_133_1552 ();
 sg13g2_fill_2 FILLER_134_32 ();
 sg13g2_fill_1 FILLER_134_45 ();
 sg13g2_fill_4 FILLER_134_51 ();
 sg13g2_fill_2 FILLER_134_55 ();
 sg13g2_fill_8 FILLER_134_72 ();
 sg13g2_fill_8 FILLER_134_80 ();
 sg13g2_fill_4 FILLER_134_94 ();
 sg13g2_fill_8 FILLER_134_107 ();
 sg13g2_fill_8 FILLER_134_115 ();
 sg13g2_fill_8 FILLER_134_123 ();
 sg13g2_fill_4 FILLER_134_131 ();
 sg13g2_fill_2 FILLER_134_135 ();
 sg13g2_fill_8 FILLER_134_147 ();
 sg13g2_fill_2 FILLER_134_155 ();
 sg13g2_fill_4 FILLER_134_162 ();
 sg13g2_fill_2 FILLER_134_166 ();
 sg13g2_fill_8 FILLER_134_194 ();
 sg13g2_fill_2 FILLER_134_202 ();
 sg13g2_fill_2 FILLER_134_217 ();
 sg13g2_fill_8 FILLER_134_227 ();
 sg13g2_fill_4 FILLER_134_235 ();
 sg13g2_fill_4 FILLER_134_285 ();
 sg13g2_fill_2 FILLER_134_289 ();
 sg13g2_fill_4 FILLER_134_327 ();
 sg13g2_fill_2 FILLER_134_331 ();
 sg13g2_fill_4 FILLER_134_358 ();
 sg13g2_fill_1 FILLER_134_362 ();
 sg13g2_fill_8 FILLER_134_403 ();
 sg13g2_fill_2 FILLER_134_411 ();
 sg13g2_fill_1 FILLER_134_413 ();
 sg13g2_fill_8 FILLER_134_422 ();
 sg13g2_fill_8 FILLER_134_430 ();
 sg13g2_fill_8 FILLER_134_438 ();
 sg13g2_fill_8 FILLER_134_446 ();
 sg13g2_fill_8 FILLER_134_454 ();
 sg13g2_fill_2 FILLER_134_462 ();
 sg13g2_fill_1 FILLER_134_464 ();
 sg13g2_fill_1 FILLER_134_471 ();
 sg13g2_fill_4 FILLER_134_480 ();
 sg13g2_fill_4 FILLER_134_572 ();
 sg13g2_fill_2 FILLER_134_586 ();
 sg13g2_fill_4 FILLER_134_593 ();
 sg13g2_fill_2 FILLER_134_597 ();
 sg13g2_fill_1 FILLER_134_599 ();
 sg13g2_fill_8 FILLER_134_608 ();
 sg13g2_fill_8 FILLER_134_616 ();
 sg13g2_fill_4 FILLER_134_624 ();
 sg13g2_fill_8 FILLER_134_638 ();
 sg13g2_fill_8 FILLER_134_646 ();
 sg13g2_fill_8 FILLER_134_654 ();
 sg13g2_fill_8 FILLER_134_662 ();
 sg13g2_fill_8 FILLER_134_670 ();
 sg13g2_fill_8 FILLER_134_686 ();
 sg13g2_fill_8 FILLER_134_694 ();
 sg13g2_fill_8 FILLER_134_702 ();
 sg13g2_fill_1 FILLER_134_710 ();
 sg13g2_fill_8 FILLER_134_729 ();
 sg13g2_fill_8 FILLER_134_737 ();
 sg13g2_fill_8 FILLER_134_745 ();
 sg13g2_fill_4 FILLER_134_783 ();
 sg13g2_fill_2 FILLER_134_787 ();
 sg13g2_fill_1 FILLER_134_789 ();
 sg13g2_fill_4 FILLER_134_800 ();
 sg13g2_fill_2 FILLER_134_804 ();
 sg13g2_fill_1 FILLER_134_832 ();
 sg13g2_fill_1 FILLER_134_859 ();
 sg13g2_fill_1 FILLER_134_890 ();
 sg13g2_fill_8 FILLER_134_901 ();
 sg13g2_fill_8 FILLER_134_909 ();
 sg13g2_fill_2 FILLER_134_917 ();
 sg13g2_fill_2 FILLER_134_977 ();
 sg13g2_fill_1 FILLER_134_979 ();
 sg13g2_fill_8 FILLER_134_986 ();
 sg13g2_fill_8 FILLER_134_994 ();
 sg13g2_fill_4 FILLER_134_1002 ();
 sg13g2_fill_2 FILLER_134_1006 ();
 sg13g2_fill_4 FILLER_134_1031 ();
 sg13g2_fill_8 FILLER_134_1055 ();
 sg13g2_fill_4 FILLER_134_1082 ();
 sg13g2_fill_1 FILLER_134_1086 ();
 sg13g2_fill_8 FILLER_134_1096 ();
 sg13g2_fill_2 FILLER_134_1104 ();
 sg13g2_fill_1 FILLER_134_1106 ();
 sg13g2_fill_2 FILLER_134_1126 ();
 sg13g2_fill_1 FILLER_134_1128 ();
 sg13g2_fill_2 FILLER_134_1168 ();
 sg13g2_fill_1 FILLER_134_1170 ();
 sg13g2_fill_1 FILLER_134_1181 ();
 sg13g2_fill_2 FILLER_134_1194 ();
 sg13g2_fill_4 FILLER_134_1205 ();
 sg13g2_fill_8 FILLER_134_1220 ();
 sg13g2_fill_2 FILLER_134_1228 ();
 sg13g2_fill_1 FILLER_134_1230 ();
 sg13g2_fill_2 FILLER_134_1236 ();
 sg13g2_fill_4 FILLER_134_1242 ();
 sg13g2_fill_1 FILLER_134_1246 ();
 sg13g2_fill_4 FILLER_134_1252 ();
 sg13g2_fill_2 FILLER_134_1256 ();
 sg13g2_fill_1 FILLER_134_1258 ();
 sg13g2_fill_8 FILLER_134_1273 ();
 sg13g2_fill_8 FILLER_134_1281 ();
 sg13g2_fill_4 FILLER_134_1289 ();
 sg13g2_fill_2 FILLER_134_1293 ();
 sg13g2_fill_1 FILLER_134_1295 ();
 sg13g2_fill_2 FILLER_134_1301 ();
 sg13g2_fill_1 FILLER_134_1303 ();
 sg13g2_fill_2 FILLER_134_1313 ();
 sg13g2_fill_1 FILLER_134_1315 ();
 sg13g2_fill_4 FILLER_134_1337 ();
 sg13g2_fill_8 FILLER_134_1344 ();
 sg13g2_fill_1 FILLER_134_1352 ();
 sg13g2_fill_8 FILLER_134_1387 ();
 sg13g2_fill_8 FILLER_134_1395 ();
 sg13g2_fill_2 FILLER_134_1403 ();
 sg13g2_fill_1 FILLER_134_1405 ();
 sg13g2_fill_4 FILLER_134_1415 ();
 sg13g2_fill_2 FILLER_134_1419 ();
 sg13g2_fill_4 FILLER_134_1442 ();
 sg13g2_fill_1 FILLER_134_1446 ();
 sg13g2_fill_8 FILLER_134_1457 ();
 sg13g2_fill_1 FILLER_134_1465 ();
 sg13g2_fill_8 FILLER_134_1518 ();
 sg13g2_fill_4 FILLER_134_1526 ();
 sg13g2_fill_2 FILLER_134_1530 ();
 sg13g2_fill_1 FILLER_134_1532 ();
 sg13g2_fill_8 FILLER_134_1584 ();
 sg13g2_fill_8 FILLER_135_0 ();
 sg13g2_fill_8 FILLER_135_8 ();
 sg13g2_fill_4 FILLER_135_16 ();
 sg13g2_fill_2 FILLER_135_33 ();
 sg13g2_fill_4 FILLER_135_38 ();
 sg13g2_fill_8 FILLER_135_57 ();
 sg13g2_fill_2 FILLER_135_65 ();
 sg13g2_fill_8 FILLER_135_83 ();
 sg13g2_fill_1 FILLER_135_91 ();
 sg13g2_fill_4 FILLER_135_97 ();
 sg13g2_fill_2 FILLER_135_101 ();
 sg13g2_fill_4 FILLER_135_211 ();
 sg13g2_fill_2 FILLER_135_215 ();
 sg13g2_fill_1 FILLER_135_243 ();
 sg13g2_fill_2 FILLER_135_264 ();
 sg13g2_fill_1 FILLER_135_266 ();
 sg13g2_fill_1 FILLER_135_361 ();
 sg13g2_fill_4 FILLER_135_368 ();
 sg13g2_fill_2 FILLER_135_372 ();
 sg13g2_fill_2 FILLER_135_384 ();
 sg13g2_fill_4 FILLER_135_396 ();
 sg13g2_fill_2 FILLER_135_400 ();
 sg13g2_fill_1 FILLER_135_402 ();
 sg13g2_fill_2 FILLER_135_411 ();
 sg13g2_fill_1 FILLER_135_413 ();
 sg13g2_fill_8 FILLER_135_440 ();
 sg13g2_fill_4 FILLER_135_448 ();
 sg13g2_fill_4 FILLER_135_462 ();
 sg13g2_fill_1 FILLER_135_466 ();
 sg13g2_fill_8 FILLER_135_477 ();
 sg13g2_fill_4 FILLER_135_485 ();
 sg13g2_fill_4 FILLER_135_499 ();
 sg13g2_fill_1 FILLER_135_503 ();
 sg13g2_fill_2 FILLER_135_543 ();
 sg13g2_fill_1 FILLER_135_545 ();
 sg13g2_fill_4 FILLER_135_572 ();
 sg13g2_fill_1 FILLER_135_576 ();
 sg13g2_fill_2 FILLER_135_651 ();
 sg13g2_fill_8 FILLER_135_689 ();
 sg13g2_fill_8 FILLER_135_697 ();
 sg13g2_fill_4 FILLER_135_705 ();
 sg13g2_fill_2 FILLER_135_709 ();
 sg13g2_fill_8 FILLER_135_719 ();
 sg13g2_fill_8 FILLER_135_727 ();
 sg13g2_fill_4 FILLER_135_735 ();
 sg13g2_fill_2 FILLER_135_739 ();
 sg13g2_fill_1 FILLER_135_741 ();
 sg13g2_fill_8 FILLER_135_758 ();
 sg13g2_fill_8 FILLER_135_766 ();
 sg13g2_fill_4 FILLER_135_774 ();
 sg13g2_fill_2 FILLER_135_778 ();
 sg13g2_fill_4 FILLER_135_816 ();
 sg13g2_fill_2 FILLER_135_820 ();
 sg13g2_fill_8 FILLER_135_838 ();
 sg13g2_fill_8 FILLER_135_846 ();
 sg13g2_fill_8 FILLER_135_854 ();
 sg13g2_fill_8 FILLER_135_862 ();
 sg13g2_fill_2 FILLER_135_870 ();
 sg13g2_fill_1 FILLER_135_872 ();
 sg13g2_fill_4 FILLER_135_878 ();
 sg13g2_fill_1 FILLER_135_882 ();
 sg13g2_fill_2 FILLER_135_923 ();
 sg13g2_fill_1 FILLER_135_953 ();
 sg13g2_fill_2 FILLER_135_964 ();
 sg13g2_fill_8 FILLER_135_981 ();
 sg13g2_fill_4 FILLER_135_989 ();
 sg13g2_fill_2 FILLER_135_993 ();
 sg13g2_fill_1 FILLER_135_995 ();
 sg13g2_fill_1 FILLER_135_1001 ();
 sg13g2_fill_4 FILLER_135_1010 ();
 sg13g2_fill_8 FILLER_135_1025 ();
 sg13g2_fill_2 FILLER_135_1033 ();
 sg13g2_fill_1 FILLER_135_1035 ();
 sg13g2_fill_4 FILLER_135_1043 ();
 sg13g2_fill_1 FILLER_135_1047 ();
 sg13g2_fill_4 FILLER_135_1083 ();
 sg13g2_fill_1 FILLER_135_1107 ();
 sg13g2_fill_8 FILLER_135_1134 ();
 sg13g2_fill_4 FILLER_135_1142 ();
 sg13g2_fill_1 FILLER_135_1146 ();
 sg13g2_fill_2 FILLER_135_1200 ();
 sg13g2_fill_2 FILLER_135_1206 ();
 sg13g2_fill_2 FILLER_135_1251 ();
 sg13g2_fill_1 FILLER_135_1253 ();
 sg13g2_fill_4 FILLER_135_1299 ();
 sg13g2_fill_2 FILLER_135_1321 ();
 sg13g2_fill_1 FILLER_135_1323 ();
 sg13g2_fill_4 FILLER_135_1328 ();
 sg13g2_fill_1 FILLER_135_1345 ();
 sg13g2_fill_8 FILLER_135_1351 ();
 sg13g2_fill_1 FILLER_135_1359 ();
 sg13g2_fill_1 FILLER_135_1371 ();
 sg13g2_fill_1 FILLER_135_1381 ();
 sg13g2_fill_4 FILLER_135_1387 ();
 sg13g2_fill_1 FILLER_135_1391 ();
 sg13g2_fill_4 FILLER_135_1437 ();
 sg13g2_fill_2 FILLER_135_1441 ();
 sg13g2_fill_2 FILLER_135_1452 ();
 sg13g2_fill_1 FILLER_135_1454 ();
 sg13g2_fill_4 FILLER_135_1481 ();
 sg13g2_fill_1 FILLER_135_1485 ();
 sg13g2_fill_4 FILLER_135_1535 ();
 sg13g2_fill_4 FILLER_135_1549 ();
 sg13g2_fill_2 FILLER_135_1553 ();
 sg13g2_fill_1 FILLER_135_1555 ();
 sg13g2_fill_8 FILLER_136_0 ();
 sg13g2_fill_8 FILLER_136_8 ();
 sg13g2_fill_1 FILLER_136_19 ();
 sg13g2_fill_2 FILLER_136_26 ();
 sg13g2_fill_1 FILLER_136_28 ();
 sg13g2_fill_2 FILLER_136_41 ();
 sg13g2_fill_1 FILLER_136_43 ();
 sg13g2_fill_8 FILLER_136_49 ();
 sg13g2_fill_2 FILLER_136_57 ();
 sg13g2_fill_1 FILLER_136_59 ();
 sg13g2_fill_8 FILLER_136_66 ();
 sg13g2_fill_4 FILLER_136_74 ();
 sg13g2_fill_1 FILLER_136_78 ();
 sg13g2_fill_4 FILLER_136_130 ();
 sg13g2_fill_2 FILLER_136_134 ();
 sg13g2_fill_1 FILLER_136_136 ();
 sg13g2_fill_8 FILLER_136_182 ();
 sg13g2_fill_8 FILLER_136_190 ();
 sg13g2_fill_8 FILLER_136_198 ();
 sg13g2_fill_4 FILLER_136_206 ();
 sg13g2_fill_2 FILLER_136_210 ();
 sg13g2_fill_8 FILLER_136_222 ();
 sg13g2_fill_8 FILLER_136_230 ();
 sg13g2_fill_8 FILLER_136_238 ();
 sg13g2_fill_8 FILLER_136_246 ();
 sg13g2_fill_8 FILLER_136_254 ();
 sg13g2_fill_8 FILLER_136_262 ();
 sg13g2_fill_2 FILLER_136_270 ();
 sg13g2_fill_1 FILLER_136_272 ();
 sg13g2_fill_8 FILLER_136_283 ();
 sg13g2_fill_8 FILLER_136_291 ();
 sg13g2_fill_4 FILLER_136_299 ();
 sg13g2_fill_2 FILLER_136_303 ();
 sg13g2_fill_1 FILLER_136_305 ();
 sg13g2_fill_8 FILLER_136_331 ();
 sg13g2_fill_4 FILLER_136_339 ();
 sg13g2_fill_8 FILLER_136_353 ();
 sg13g2_fill_8 FILLER_136_361 ();
 sg13g2_fill_8 FILLER_136_369 ();
 sg13g2_fill_8 FILLER_136_377 ();
 sg13g2_fill_8 FILLER_136_385 ();
 sg13g2_fill_2 FILLER_136_393 ();
 sg13g2_fill_1 FILLER_136_395 ();
 sg13g2_fill_4 FILLER_136_404 ();
 sg13g2_fill_4 FILLER_136_416 ();
 sg13g2_fill_2 FILLER_136_420 ();
 sg13g2_fill_1 FILLER_136_422 ();
 sg13g2_fill_2 FILLER_136_459 ();
 sg13g2_fill_4 FILLER_136_503 ();
 sg13g2_fill_2 FILLER_136_507 ();
 sg13g2_fill_1 FILLER_136_509 ();
 sg13g2_fill_4 FILLER_136_536 ();
 sg13g2_fill_1 FILLER_136_540 ();
 sg13g2_fill_8 FILLER_136_551 ();
 sg13g2_fill_8 FILLER_136_559 ();
 sg13g2_fill_1 FILLER_136_567 ();
 sg13g2_fill_8 FILLER_136_593 ();
 sg13g2_fill_2 FILLER_136_601 ();
 sg13g2_fill_8 FILLER_136_656 ();
 sg13g2_fill_8 FILLER_136_664 ();
 sg13g2_fill_8 FILLER_136_672 ();
 sg13g2_fill_2 FILLER_136_680 ();
 sg13g2_fill_4 FILLER_136_692 ();
 sg13g2_fill_1 FILLER_136_696 ();
 sg13g2_fill_4 FILLER_136_741 ();
 sg13g2_fill_2 FILLER_136_745 ();
 sg13g2_fill_8 FILLER_136_773 ();
 sg13g2_fill_4 FILLER_136_781 ();
 sg13g2_fill_2 FILLER_136_795 ();
 sg13g2_fill_1 FILLER_136_797 ();
 sg13g2_fill_4 FILLER_136_824 ();
 sg13g2_fill_1 FILLER_136_828 ();
 sg13g2_fill_2 FILLER_136_888 ();
 sg13g2_fill_8 FILLER_136_900 ();
 sg13g2_fill_8 FILLER_136_908 ();
 sg13g2_fill_2 FILLER_136_916 ();
 sg13g2_fill_1 FILLER_136_918 ();
 sg13g2_fill_2 FILLER_136_947 ();
 sg13g2_fill_1 FILLER_136_949 ();
 sg13g2_fill_4 FILLER_136_954 ();
 sg13g2_fill_2 FILLER_136_958 ();
 sg13g2_fill_1 FILLER_136_960 ();
 sg13g2_fill_8 FILLER_136_970 ();
 sg13g2_fill_4 FILLER_136_978 ();
 sg13g2_fill_1 FILLER_136_982 ();
 sg13g2_fill_1 FILLER_136_988 ();
 sg13g2_fill_4 FILLER_136_994 ();
 sg13g2_fill_2 FILLER_136_998 ();
 sg13g2_fill_1 FILLER_136_1000 ();
 sg13g2_fill_2 FILLER_136_1009 ();
 sg13g2_fill_4 FILLER_136_1020 ();
 sg13g2_fill_8 FILLER_136_1029 ();
 sg13g2_fill_8 FILLER_136_1037 ();
 sg13g2_fill_8 FILLER_136_1045 ();
 sg13g2_fill_8 FILLER_136_1053 ();
 sg13g2_fill_8 FILLER_136_1061 ();
 sg13g2_fill_8 FILLER_136_1073 ();
 sg13g2_fill_8 FILLER_136_1081 ();
 sg13g2_fill_2 FILLER_136_1089 ();
 sg13g2_fill_1 FILLER_136_1091 ();
 sg13g2_fill_1 FILLER_136_1100 ();
 sg13g2_fill_4 FILLER_136_1105 ();
 sg13g2_fill_2 FILLER_136_1109 ();
 sg13g2_fill_1 FILLER_136_1111 ();
 sg13g2_fill_4 FILLER_136_1142 ();
 sg13g2_fill_2 FILLER_136_1156 ();
 sg13g2_fill_2 FILLER_136_1174 ();
 sg13g2_fill_1 FILLER_136_1176 ();
 sg13g2_fill_4 FILLER_136_1190 ();
 sg13g2_fill_2 FILLER_136_1194 ();
 sg13g2_fill_1 FILLER_136_1196 ();
 sg13g2_fill_2 FILLER_136_1210 ();
 sg13g2_fill_8 FILLER_136_1223 ();
 sg13g2_fill_8 FILLER_136_1231 ();
 sg13g2_fill_2 FILLER_136_1239 ();
 sg13g2_fill_1 FILLER_136_1241 ();
 sg13g2_fill_4 FILLER_136_1257 ();
 sg13g2_fill_1 FILLER_136_1266 ();
 sg13g2_fill_8 FILLER_136_1280 ();
 sg13g2_fill_4 FILLER_136_1288 ();
 sg13g2_fill_4 FILLER_136_1298 ();
 sg13g2_fill_2 FILLER_136_1302 ();
 sg13g2_fill_1 FILLER_136_1304 ();
 sg13g2_fill_2 FILLER_136_1314 ();
 sg13g2_fill_8 FILLER_136_1321 ();
 sg13g2_fill_4 FILLER_136_1329 ();
 sg13g2_fill_2 FILLER_136_1354 ();
 sg13g2_fill_1 FILLER_136_1356 ();
 sg13g2_fill_1 FILLER_136_1370 ();
 sg13g2_fill_2 FILLER_136_1379 ();
 sg13g2_fill_1 FILLER_136_1381 ();
 sg13g2_fill_8 FILLER_136_1407 ();
 sg13g2_fill_8 FILLER_136_1415 ();
 sg13g2_fill_8 FILLER_136_1423 ();
 sg13g2_fill_8 FILLER_136_1436 ();
 sg13g2_fill_4 FILLER_136_1444 ();
 sg13g2_fill_2 FILLER_136_1448 ();
 sg13g2_fill_1 FILLER_136_1450 ();
 sg13g2_fill_4 FILLER_136_1461 ();
 sg13g2_fill_1 FILLER_136_1465 ();
 sg13g2_fill_8 FILLER_136_1531 ();
 sg13g2_fill_8 FILLER_136_1539 ();
 sg13g2_fill_8 FILLER_136_1547 ();
 sg13g2_fill_4 FILLER_136_1555 ();
 sg13g2_fill_8 FILLER_136_1571 ();
 sg13g2_fill_8 FILLER_136_1579 ();
 sg13g2_fill_4 FILLER_136_1587 ();
 sg13g2_fill_1 FILLER_136_1591 ();
 sg13g2_fill_4 FILLER_137_0 ();
 sg13g2_fill_4 FILLER_137_14 ();
 sg13g2_fill_2 FILLER_137_18 ();
 sg13g2_fill_1 FILLER_137_20 ();
 sg13g2_fill_1 FILLER_137_27 ();
 sg13g2_fill_2 FILLER_137_46 ();
 sg13g2_fill_1 FILLER_137_48 ();
 sg13g2_fill_2 FILLER_137_54 ();
 sg13g2_fill_2 FILLER_137_64 ();
 sg13g2_fill_8 FILLER_137_80 ();
 sg13g2_fill_8 FILLER_137_88 ();
 sg13g2_fill_8 FILLER_137_96 ();
 sg13g2_fill_8 FILLER_137_104 ();
 sg13g2_fill_2 FILLER_137_143 ();
 sg13g2_fill_4 FILLER_137_171 ();
 sg13g2_fill_8 FILLER_137_183 ();
 sg13g2_fill_8 FILLER_137_191 ();
 sg13g2_fill_8 FILLER_137_199 ();
 sg13g2_fill_8 FILLER_137_207 ();
 sg13g2_fill_1 FILLER_137_215 ();
 sg13g2_fill_1 FILLER_137_242 ();
 sg13g2_fill_8 FILLER_137_255 ();
 sg13g2_fill_2 FILLER_137_279 ();
 sg13g2_fill_2 FILLER_137_286 ();
 sg13g2_fill_8 FILLER_137_294 ();
 sg13g2_fill_2 FILLER_137_302 ();
 sg13g2_fill_1 FILLER_137_304 ();
 sg13g2_fill_1 FILLER_137_318 ();
 sg13g2_fill_8 FILLER_137_329 ();
 sg13g2_fill_8 FILLER_137_337 ();
 sg13g2_fill_4 FILLER_137_345 ();
 sg13g2_fill_1 FILLER_137_349 ();
 sg13g2_fill_8 FILLER_137_360 ();
 sg13g2_fill_1 FILLER_137_368 ();
 sg13g2_fill_8 FILLER_137_413 ();
 sg13g2_fill_4 FILLER_137_421 ();
 sg13g2_fill_2 FILLER_137_425 ();
 sg13g2_fill_8 FILLER_137_437 ();
 sg13g2_fill_4 FILLER_137_445 ();
 sg13g2_fill_2 FILLER_137_449 ();
 sg13g2_fill_1 FILLER_137_461 ();
 sg13g2_fill_4 FILLER_137_468 ();
 sg13g2_fill_2 FILLER_137_472 ();
 sg13g2_fill_8 FILLER_137_482 ();
 sg13g2_fill_4 FILLER_137_490 ();
 sg13g2_fill_1 FILLER_137_494 ();
 sg13g2_fill_8 FILLER_137_505 ();
 sg13g2_fill_8 FILLER_137_513 ();
 sg13g2_fill_1 FILLER_137_521 ();
 sg13g2_fill_8 FILLER_137_530 ();
 sg13g2_fill_8 FILLER_137_538 ();
 sg13g2_fill_8 FILLER_137_546 ();
 sg13g2_fill_8 FILLER_137_554 ();
 sg13g2_fill_4 FILLER_137_562 ();
 sg13g2_fill_2 FILLER_137_566 ();
 sg13g2_fill_4 FILLER_137_590 ();
 sg13g2_fill_8 FILLER_137_599 ();
 sg13g2_fill_4 FILLER_137_607 ();
 sg13g2_fill_4 FILLER_137_636 ();
 sg13g2_fill_1 FILLER_137_686 ();
 sg13g2_fill_2 FILLER_137_713 ();
 sg13g2_fill_1 FILLER_137_715 ();
 sg13g2_fill_8 FILLER_137_724 ();
 sg13g2_fill_4 FILLER_137_732 ();
 sg13g2_fill_8 FILLER_137_744 ();
 sg13g2_fill_8 FILLER_137_752 ();
 sg13g2_fill_8 FILLER_137_760 ();
 sg13g2_fill_8 FILLER_137_773 ();
 sg13g2_fill_4 FILLER_137_781 ();
 sg13g2_fill_8 FILLER_137_795 ();
 sg13g2_fill_8 FILLER_137_803 ();
 sg13g2_fill_8 FILLER_137_811 ();
 sg13g2_fill_1 FILLER_137_843 ();
 sg13g2_fill_2 FILLER_137_849 ();
 sg13g2_fill_1 FILLER_137_851 ();
 sg13g2_fill_8 FILLER_137_858 ();
 sg13g2_fill_8 FILLER_137_866 ();
 sg13g2_fill_2 FILLER_137_874 ();
 sg13g2_fill_1 FILLER_137_881 ();
 sg13g2_fill_4 FILLER_137_892 ();
 sg13g2_fill_2 FILLER_137_896 ();
 sg13g2_fill_1 FILLER_137_898 ();
 sg13g2_fill_8 FILLER_137_934 ();
 sg13g2_fill_4 FILLER_137_942 ();
 sg13g2_fill_8 FILLER_137_951 ();
 sg13g2_fill_4 FILLER_137_959 ();
 sg13g2_fill_1 FILLER_137_963 ();
 sg13g2_fill_2 FILLER_137_976 ();
 sg13g2_fill_8 FILLER_137_995 ();
 sg13g2_fill_2 FILLER_137_1008 ();
 sg13g2_fill_1 FILLER_137_1010 ();
 sg13g2_fill_4 FILLER_137_1023 ();
 sg13g2_fill_1 FILLER_137_1027 ();
 sg13g2_fill_8 FILLER_137_1034 ();
 sg13g2_fill_4 FILLER_137_1042 ();
 sg13g2_fill_1 FILLER_137_1046 ();
 sg13g2_fill_2 FILLER_137_1065 ();
 sg13g2_fill_4 FILLER_137_1080 ();
 sg13g2_fill_8 FILLER_137_1119 ();
 sg13g2_fill_2 FILLER_137_1127 ();
 sg13g2_fill_8 FILLER_137_1134 ();
 sg13g2_fill_8 FILLER_137_1142 ();
 sg13g2_fill_4 FILLER_137_1150 ();
 sg13g2_fill_2 FILLER_137_1154 ();
 sg13g2_fill_2 FILLER_137_1161 ();
 sg13g2_fill_1 FILLER_137_1168 ();
 sg13g2_fill_2 FILLER_137_1177 ();
 sg13g2_fill_8 FILLER_137_1187 ();
 sg13g2_fill_2 FILLER_137_1195 ();
 sg13g2_fill_1 FILLER_137_1202 ();
 sg13g2_fill_8 FILLER_137_1216 ();
 sg13g2_fill_1 FILLER_137_1224 ();
 sg13g2_fill_4 FILLER_137_1229 ();
 sg13g2_fill_8 FILLER_137_1238 ();
 sg13g2_fill_4 FILLER_137_1246 ();
 sg13g2_fill_1 FILLER_137_1250 ();
 sg13g2_fill_8 FILLER_137_1256 ();
 sg13g2_fill_4 FILLER_137_1264 ();
 sg13g2_fill_1 FILLER_137_1268 ();
 sg13g2_fill_2 FILLER_137_1274 ();
 sg13g2_fill_1 FILLER_137_1276 ();
 sg13g2_fill_4 FILLER_137_1282 ();
 sg13g2_fill_2 FILLER_137_1300 ();
 sg13g2_fill_1 FILLER_137_1302 ();
 sg13g2_fill_2 FILLER_137_1307 ();
 sg13g2_fill_2 FILLER_137_1334 ();
 sg13g2_fill_8 FILLER_137_1347 ();
 sg13g2_fill_2 FILLER_137_1374 ();
 sg13g2_fill_1 FILLER_137_1376 ();
 sg13g2_fill_8 FILLER_137_1392 ();
 sg13g2_fill_8 FILLER_137_1400 ();
 sg13g2_fill_1 FILLER_137_1425 ();
 sg13g2_fill_4 FILLER_137_1430 ();
 sg13g2_fill_8 FILLER_137_1438 ();
 sg13g2_fill_2 FILLER_137_1446 ();
 sg13g2_fill_1 FILLER_137_1457 ();
 sg13g2_fill_8 FILLER_137_1484 ();
 sg13g2_fill_2 FILLER_137_1492 ();
 sg13g2_fill_1 FILLER_137_1494 ();
 sg13g2_fill_2 FILLER_137_1540 ();
 sg13g2_fill_8 FILLER_137_1546 ();
 sg13g2_fill_4 FILLER_137_1554 ();
 sg13g2_fill_2 FILLER_137_1558 ();
 sg13g2_fill_1 FILLER_137_1560 ();
 sg13g2_fill_8 FILLER_137_1582 ();
 sg13g2_fill_2 FILLER_137_1590 ();
 sg13g2_fill_8 FILLER_138_26 ();
 sg13g2_fill_4 FILLER_138_34 ();
 sg13g2_fill_8 FILLER_138_48 ();
 sg13g2_fill_2 FILLER_138_56 ();
 sg13g2_fill_1 FILLER_138_58 ();
 sg13g2_fill_2 FILLER_138_68 ();
 sg13g2_fill_4 FILLER_138_100 ();
 sg13g2_fill_2 FILLER_138_104 ();
 sg13g2_fill_2 FILLER_138_126 ();
 sg13g2_fill_1 FILLER_138_128 ();
 sg13g2_fill_4 FILLER_138_156 ();
 sg13g2_fill_2 FILLER_138_160 ();
 sg13g2_fill_4 FILLER_138_168 ();
 sg13g2_fill_2 FILLER_138_172 ();
 sg13g2_fill_8 FILLER_138_192 ();
 sg13g2_fill_2 FILLER_138_200 ();
 sg13g2_fill_1 FILLER_138_225 ();
 sg13g2_fill_2 FILLER_138_271 ();
 sg13g2_fill_1 FILLER_138_304 ();
 sg13g2_fill_2 FILLER_138_313 ();
 sg13g2_fill_4 FILLER_138_351 ();
 sg13g2_fill_8 FILLER_138_386 ();
 sg13g2_fill_8 FILLER_138_402 ();
 sg13g2_fill_4 FILLER_138_410 ();
 sg13g2_fill_2 FILLER_138_414 ();
 sg13g2_fill_2 FILLER_138_429 ();
 sg13g2_fill_1 FILLER_138_431 ();
 sg13g2_fill_8 FILLER_138_442 ();
 sg13g2_fill_4 FILLER_138_450 ();
 sg13g2_fill_1 FILLER_138_454 ();
 sg13g2_fill_4 FILLER_138_465 ();
 sg13g2_fill_8 FILLER_138_479 ();
 sg13g2_fill_1 FILLER_138_533 ();
 sg13g2_fill_8 FILLER_138_554 ();
 sg13g2_fill_4 FILLER_138_562 ();
 sg13g2_fill_2 FILLER_138_587 ();
 sg13g2_fill_1 FILLER_138_589 ();
 sg13g2_fill_1 FILLER_138_634 ();
 sg13g2_fill_4 FILLER_138_641 ();
 sg13g2_fill_2 FILLER_138_645 ();
 sg13g2_fill_1 FILLER_138_647 ();
 sg13g2_fill_8 FILLER_138_660 ();
 sg13g2_fill_8 FILLER_138_668 ();
 sg13g2_fill_8 FILLER_138_676 ();
 sg13g2_fill_2 FILLER_138_684 ();
 sg13g2_fill_1 FILLER_138_726 ();
 sg13g2_fill_4 FILLER_138_735 ();
 sg13g2_fill_1 FILLER_138_739 ();
 sg13g2_fill_2 FILLER_138_750 ();
 sg13g2_fill_8 FILLER_138_781 ();
 sg13g2_fill_2 FILLER_138_799 ();
 sg13g2_fill_1 FILLER_138_801 ();
 sg13g2_fill_8 FILLER_138_865 ();
 sg13g2_fill_8 FILLER_138_873 ();
 sg13g2_fill_4 FILLER_138_881 ();
 sg13g2_fill_8 FILLER_138_920 ();
 sg13g2_fill_1 FILLER_138_928 ();
 sg13g2_fill_4 FILLER_138_935 ();
 sg13g2_fill_8 FILLER_138_972 ();
 sg13g2_fill_1 FILLER_138_980 ();
 sg13g2_fill_2 FILLER_138_992 ();
 sg13g2_fill_4 FILLER_138_1016 ();
 sg13g2_fill_1 FILLER_138_1020 ();
 sg13g2_fill_8 FILLER_138_1031 ();
 sg13g2_fill_2 FILLER_138_1039 ();
 sg13g2_fill_8 FILLER_138_1075 ();
 sg13g2_fill_2 FILLER_138_1083 ();
 sg13g2_fill_1 FILLER_138_1085 ();
 sg13g2_fill_2 FILLER_138_1101 ();
 sg13g2_fill_1 FILLER_138_1103 ();
 sg13g2_fill_1 FILLER_138_1139 ();
 sg13g2_fill_2 FILLER_138_1144 ();
 sg13g2_fill_1 FILLER_138_1146 ();
 sg13g2_fill_2 FILLER_138_1182 ();
 sg13g2_fill_1 FILLER_138_1203 ();
 sg13g2_fill_2 FILLER_138_1219 ();
 sg13g2_fill_1 FILLER_138_1221 ();
 sg13g2_fill_8 FILLER_138_1248 ();
 sg13g2_fill_2 FILLER_138_1256 ();
 sg13g2_fill_1 FILLER_138_1258 ();
 sg13g2_fill_8 FILLER_138_1262 ();
 sg13g2_fill_2 FILLER_138_1270 ();
 sg13g2_fill_1 FILLER_138_1272 ();
 sg13g2_fill_4 FILLER_138_1277 ();
 sg13g2_fill_1 FILLER_138_1281 ();
 sg13g2_fill_2 FILLER_138_1287 ();
 sg13g2_fill_8 FILLER_138_1297 ();
 sg13g2_fill_8 FILLER_138_1305 ();
 sg13g2_fill_2 FILLER_138_1313 ();
 sg13g2_fill_2 FILLER_138_1334 ();
 sg13g2_fill_1 FILLER_138_1346 ();
 sg13g2_fill_8 FILLER_138_1356 ();
 sg13g2_fill_2 FILLER_138_1364 ();
 sg13g2_fill_1 FILLER_138_1366 ();
 sg13g2_fill_8 FILLER_138_1377 ();
 sg13g2_fill_8 FILLER_138_1385 ();
 sg13g2_fill_4 FILLER_138_1393 ();
 sg13g2_fill_1 FILLER_138_1397 ();
 sg13g2_fill_4 FILLER_138_1416 ();
 sg13g2_fill_2 FILLER_138_1420 ();
 sg13g2_fill_1 FILLER_138_1422 ();
 sg13g2_fill_8 FILLER_138_1428 ();
 sg13g2_fill_2 FILLER_138_1436 ();
 sg13g2_fill_2 FILLER_138_1442 ();
 sg13g2_fill_4 FILLER_138_1454 ();
 sg13g2_fill_2 FILLER_138_1515 ();
 sg13g2_fill_4 FILLER_138_1523 ();
 sg13g2_fill_2 FILLER_138_1527 ();
 sg13g2_fill_1 FILLER_138_1529 ();
 sg13g2_fill_2 FILLER_138_1564 ();
 sg13g2_fill_8 FILLER_139_30 ();
 sg13g2_fill_8 FILLER_139_38 ();
 sg13g2_fill_4 FILLER_139_56 ();
 sg13g2_fill_1 FILLER_139_60 ();
 sg13g2_fill_4 FILLER_139_106 ();
 sg13g2_fill_2 FILLER_139_110 ();
 sg13g2_fill_1 FILLER_139_122 ();
 sg13g2_fill_4 FILLER_139_129 ();
 sg13g2_fill_1 FILLER_139_138 ();
 sg13g2_fill_8 FILLER_139_149 ();
 sg13g2_fill_2 FILLER_139_157 ();
 sg13g2_fill_1 FILLER_139_159 ();
 sg13g2_fill_4 FILLER_139_170 ();
 sg13g2_fill_2 FILLER_139_174 ();
 sg13g2_fill_8 FILLER_139_202 ();
 sg13g2_fill_8 FILLER_139_210 ();
 sg13g2_fill_8 FILLER_139_218 ();
 sg13g2_fill_2 FILLER_139_226 ();
 sg13g2_fill_1 FILLER_139_228 ();
 sg13g2_fill_2 FILLER_139_251 ();
 sg13g2_fill_8 FILLER_139_279 ();
 sg13g2_fill_1 FILLER_139_287 ();
 sg13g2_fill_8 FILLER_139_298 ();
 sg13g2_fill_1 FILLER_139_306 ();
 sg13g2_fill_4 FILLER_139_312 ();
 sg13g2_fill_2 FILLER_139_316 ();
 sg13g2_fill_1 FILLER_139_318 ();
 sg13g2_fill_8 FILLER_139_329 ();
 sg13g2_fill_8 FILLER_139_337 ();
 sg13g2_fill_4 FILLER_139_345 ();
 sg13g2_fill_2 FILLER_139_349 ();
 sg13g2_fill_1 FILLER_139_351 ();
 sg13g2_fill_8 FILLER_139_362 ();
 sg13g2_fill_2 FILLER_139_370 ();
 sg13g2_fill_1 FILLER_139_372 ();
 sg13g2_fill_2 FILLER_139_386 ();
 sg13g2_fill_1 FILLER_139_388 ();
 sg13g2_fill_2 FILLER_139_415 ();
 sg13g2_fill_1 FILLER_139_417 ();
 sg13g2_fill_2 FILLER_139_431 ();
 sg13g2_fill_1 FILLER_139_433 ();
 sg13g2_fill_4 FILLER_139_464 ();
 sg13g2_fill_2 FILLER_139_506 ();
 sg13g2_fill_1 FILLER_139_508 ();
 sg13g2_fill_8 FILLER_139_516 ();
 sg13g2_fill_4 FILLER_139_524 ();
 sg13g2_fill_1 FILLER_139_528 ();
 sg13g2_fill_4 FILLER_139_587 ();
 sg13g2_fill_1 FILLER_139_591 ();
 sg13g2_fill_4 FILLER_139_643 ();
 sg13g2_fill_1 FILLER_139_647 ();
 sg13g2_fill_8 FILLER_139_664 ();
 sg13g2_fill_4 FILLER_139_672 ();
 sg13g2_fill_1 FILLER_139_676 ();
 sg13g2_fill_2 FILLER_139_687 ();
 sg13g2_fill_1 FILLER_139_689 ();
 sg13g2_fill_8 FILLER_139_729 ();
 sg13g2_fill_1 FILLER_139_737 ();
 sg13g2_fill_8 FILLER_139_780 ();
 sg13g2_fill_1 FILLER_139_788 ();
 sg13g2_fill_4 FILLER_139_819 ();
 sg13g2_fill_8 FILLER_139_849 ();
 sg13g2_fill_1 FILLER_139_857 ();
 sg13g2_fill_8 FILLER_139_934 ();
 sg13g2_fill_8 FILLER_139_942 ();
 sg13g2_fill_8 FILLER_139_958 ();
 sg13g2_fill_2 FILLER_139_966 ();
 sg13g2_fill_4 FILLER_139_977 ();
 sg13g2_fill_1 FILLER_139_981 ();
 sg13g2_fill_4 FILLER_139_1013 ();
 sg13g2_fill_1 FILLER_139_1022 ();
 sg13g2_fill_8 FILLER_139_1029 ();
 sg13g2_fill_8 FILLER_139_1037 ();
 sg13g2_fill_2 FILLER_139_1045 ();
 sg13g2_fill_1 FILLER_139_1055 ();
 sg13g2_fill_2 FILLER_139_1108 ();
 sg13g2_fill_1 FILLER_139_1110 ();
 sg13g2_fill_8 FILLER_139_1121 ();
 sg13g2_fill_8 FILLER_139_1129 ();
 sg13g2_fill_2 FILLER_139_1137 ();
 sg13g2_fill_1 FILLER_139_1139 ();
 sg13g2_fill_1 FILLER_139_1150 ();
 sg13g2_fill_1 FILLER_139_1195 ();
 sg13g2_fill_2 FILLER_139_1209 ();
 sg13g2_fill_1 FILLER_139_1242 ();
 sg13g2_fill_1 FILLER_139_1278 ();
 sg13g2_fill_4 FILLER_139_1284 ();
 sg13g2_fill_8 FILLER_139_1294 ();
 sg13g2_fill_4 FILLER_139_1302 ();
 sg13g2_fill_2 FILLER_139_1306 ();
 sg13g2_fill_2 FILLER_139_1337 ();
 sg13g2_fill_2 FILLER_139_1372 ();
 sg13g2_fill_1 FILLER_139_1383 ();
 sg13g2_fill_1 FILLER_139_1404 ();
 sg13g2_fill_2 FILLER_139_1410 ();
 sg13g2_fill_1 FILLER_139_1412 ();
 sg13g2_fill_2 FILLER_139_1418 ();
 sg13g2_fill_8 FILLER_139_1435 ();
 sg13g2_fill_2 FILLER_139_1443 ();
 sg13g2_fill_1 FILLER_139_1449 ();
 sg13g2_fill_2 FILLER_139_1464 ();
 sg13g2_fill_2 FILLER_139_1470 ();
 sg13g2_fill_8 FILLER_139_1487 ();
 sg13g2_fill_2 FILLER_139_1495 ();
 sg13g2_fill_1 FILLER_139_1497 ();
 sg13g2_fill_4 FILLER_139_1502 ();
 sg13g2_fill_1 FILLER_139_1506 ();
 sg13g2_fill_4 FILLER_139_1512 ();
 sg13g2_fill_2 FILLER_139_1516 ();
 sg13g2_fill_4 FILLER_139_1527 ();
 sg13g2_fill_2 FILLER_139_1531 ();
 sg13g2_fill_1 FILLER_139_1533 ();
 sg13g2_fill_2 FILLER_139_1548 ();
 sg13g2_fill_1 FILLER_139_1550 ();
 sg13g2_fill_8 FILLER_139_1581 ();
 sg13g2_fill_2 FILLER_139_1589 ();
 sg13g2_fill_1 FILLER_139_1591 ();
 sg13g2_fill_4 FILLER_140_0 ();
 sg13g2_fill_2 FILLER_140_4 ();
 sg13g2_fill_2 FILLER_140_16 ();
 sg13g2_fill_1 FILLER_140_18 ();
 sg13g2_fill_8 FILLER_140_59 ();
 sg13g2_fill_2 FILLER_140_67 ();
 sg13g2_fill_8 FILLER_140_121 ();
 sg13g2_fill_4 FILLER_140_129 ();
 sg13g2_fill_1 FILLER_140_133 ();
 sg13g2_fill_8 FILLER_140_170 ();
 sg13g2_fill_8 FILLER_140_178 ();
 sg13g2_fill_2 FILLER_140_186 ();
 sg13g2_fill_1 FILLER_140_188 ();
 sg13g2_fill_8 FILLER_140_194 ();
 sg13g2_fill_1 FILLER_140_202 ();
 sg13g2_fill_8 FILLER_140_229 ();
 sg13g2_fill_2 FILLER_140_237 ();
 sg13g2_fill_1 FILLER_140_239 ();
 sg13g2_fill_8 FILLER_140_248 ();
 sg13g2_fill_8 FILLER_140_256 ();
 sg13g2_fill_8 FILLER_140_264 ();
 sg13g2_fill_8 FILLER_140_272 ();
 sg13g2_fill_2 FILLER_140_280 ();
 sg13g2_fill_4 FILLER_140_292 ();
 sg13g2_fill_1 FILLER_140_296 ();
 sg13g2_fill_1 FILLER_140_349 ();
 sg13g2_fill_2 FILLER_140_372 ();
 sg13g2_fill_1 FILLER_140_374 ();
 sg13g2_fill_8 FILLER_140_388 ();
 sg13g2_fill_4 FILLER_140_396 ();
 sg13g2_fill_2 FILLER_140_400 ();
 sg13g2_fill_8 FILLER_140_410 ();
 sg13g2_fill_2 FILLER_140_418 ();
 sg13g2_fill_2 FILLER_140_428 ();
 sg13g2_fill_1 FILLER_140_430 ();
 sg13g2_fill_8 FILLER_140_481 ();
 sg13g2_fill_8 FILLER_140_489 ();
 sg13g2_fill_8 FILLER_140_497 ();
 sg13g2_fill_8 FILLER_140_505 ();
 sg13g2_fill_8 FILLER_140_513 ();
 sg13g2_fill_4 FILLER_140_526 ();
 sg13g2_fill_1 FILLER_140_530 ();
 sg13g2_fill_8 FILLER_140_560 ();
 sg13g2_fill_2 FILLER_140_573 ();
 sg13g2_fill_8 FILLER_140_601 ();
 sg13g2_fill_8 FILLER_140_609 ();
 sg13g2_fill_8 FILLER_140_617 ();
 sg13g2_fill_2 FILLER_140_625 ();
 sg13g2_fill_4 FILLER_140_637 ();
 sg13g2_fill_1 FILLER_140_641 ();
 sg13g2_fill_8 FILLER_140_662 ();
 sg13g2_fill_4 FILLER_140_670 ();
 sg13g2_fill_1 FILLER_140_674 ();
 sg13g2_fill_8 FILLER_140_711 ();
 sg13g2_fill_8 FILLER_140_719 ();
 sg13g2_fill_8 FILLER_140_791 ();
 sg13g2_fill_4 FILLER_140_799 ();
 sg13g2_fill_1 FILLER_140_803 ();
 sg13g2_fill_8 FILLER_140_834 ();
 sg13g2_fill_8 FILLER_140_842 ();
 sg13g2_fill_8 FILLER_140_876 ();
 sg13g2_fill_8 FILLER_140_884 ();
 sg13g2_fill_4 FILLER_140_892 ();
 sg13g2_fill_2 FILLER_140_896 ();
 sg13g2_fill_1 FILLER_140_898 ();
 sg13g2_fill_2 FILLER_140_905 ();
 sg13g2_fill_8 FILLER_140_919 ();
 sg13g2_fill_8 FILLER_140_927 ();
 sg13g2_fill_8 FILLER_140_935 ();
 sg13g2_fill_8 FILLER_140_948 ();
 sg13g2_fill_2 FILLER_140_956 ();
 sg13g2_fill_1 FILLER_140_958 ();
 sg13g2_fill_4 FILLER_140_969 ();
 sg13g2_fill_2 FILLER_140_973 ();
 sg13g2_fill_1 FILLER_140_975 ();
 sg13g2_fill_4 FILLER_140_981 ();
 sg13g2_fill_1 FILLER_140_985 ();
 sg13g2_fill_4 FILLER_140_989 ();
 sg13g2_fill_1 FILLER_140_993 ();
 sg13g2_fill_8 FILLER_140_998 ();
 sg13g2_fill_2 FILLER_140_1006 ();
 sg13g2_fill_1 FILLER_140_1008 ();
 sg13g2_fill_8 FILLER_140_1030 ();
 sg13g2_fill_8 FILLER_140_1038 ();
 sg13g2_fill_8 FILLER_140_1046 ();
 sg13g2_fill_4 FILLER_140_1054 ();
 sg13g2_fill_2 FILLER_140_1058 ();
 sg13g2_fill_1 FILLER_140_1060 ();
 sg13g2_fill_4 FILLER_140_1066 ();
 sg13g2_fill_2 FILLER_140_1079 ();
 sg13g2_fill_4 FILLER_140_1090 ();
 sg13g2_fill_8 FILLER_140_1099 ();
 sg13g2_fill_8 FILLER_140_1107 ();
 sg13g2_fill_8 FILLER_140_1115 ();
 sg13g2_fill_8 FILLER_140_1123 ();
 sg13g2_fill_8 FILLER_140_1131 ();
 sg13g2_fill_1 FILLER_140_1139 ();
 sg13g2_fill_8 FILLER_140_1148 ();
 sg13g2_fill_8 FILLER_140_1156 ();
 sg13g2_fill_4 FILLER_140_1164 ();
 sg13g2_fill_1 FILLER_140_1168 ();
 sg13g2_fill_8 FILLER_140_1172 ();
 sg13g2_fill_2 FILLER_140_1184 ();
 sg13g2_fill_2 FILLER_140_1219 ();
 sg13g2_fill_1 FILLER_140_1221 ();
 sg13g2_fill_2 FILLER_140_1228 ();
 sg13g2_fill_1 FILLER_140_1230 ();
 sg13g2_fill_4 FILLER_140_1237 ();
 sg13g2_fill_2 FILLER_140_1241 ();
 sg13g2_fill_4 FILLER_140_1247 ();
 sg13g2_fill_2 FILLER_140_1251 ();
 sg13g2_fill_1 FILLER_140_1253 ();
 sg13g2_fill_2 FILLER_140_1259 ();
 sg13g2_fill_8 FILLER_140_1265 ();
 sg13g2_fill_8 FILLER_140_1273 ();
 sg13g2_fill_1 FILLER_140_1305 ();
 sg13g2_fill_8 FILLER_140_1309 ();
 sg13g2_fill_8 FILLER_140_1317 ();
 sg13g2_fill_2 FILLER_140_1325 ();
 sg13g2_fill_1 FILLER_140_1336 ();
 sg13g2_fill_8 FILLER_140_1345 ();
 sg13g2_fill_8 FILLER_140_1353 ();
 sg13g2_fill_4 FILLER_140_1361 ();
 sg13g2_fill_2 FILLER_140_1365 ();
 sg13g2_fill_1 FILLER_140_1367 ();
 sg13g2_fill_8 FILLER_140_1373 ();
 sg13g2_fill_4 FILLER_140_1381 ();
 sg13g2_fill_1 FILLER_140_1385 ();
 sg13g2_fill_1 FILLER_140_1401 ();
 sg13g2_fill_8 FILLER_140_1407 ();
 sg13g2_fill_8 FILLER_140_1415 ();
 sg13g2_fill_2 FILLER_140_1423 ();
 sg13g2_fill_1 FILLER_140_1425 ();
 sg13g2_fill_4 FILLER_140_1439 ();
 sg13g2_fill_2 FILLER_140_1469 ();
 sg13g2_fill_1 FILLER_140_1471 ();
 sg13g2_fill_8 FILLER_140_1476 ();
 sg13g2_fill_4 FILLER_140_1484 ();
 sg13g2_fill_1 FILLER_140_1488 ();
 sg13g2_fill_2 FILLER_140_1496 ();
 sg13g2_fill_4 FILLER_140_1503 ();
 sg13g2_fill_2 FILLER_140_1507 ();
 sg13g2_fill_1 FILLER_140_1509 ();
 sg13g2_fill_8 FILLER_140_1535 ();
 sg13g2_fill_2 FILLER_140_1543 ();
 sg13g2_fill_4 FILLER_141_0 ();
 sg13g2_fill_1 FILLER_141_4 ();
 sg13g2_fill_8 FILLER_141_13 ();
 sg13g2_fill_8 FILLER_141_21 ();
 sg13g2_fill_8 FILLER_141_29 ();
 sg13g2_fill_8 FILLER_141_37 ();
 sg13g2_fill_2 FILLER_141_45 ();
 sg13g2_fill_1 FILLER_141_47 ();
 sg13g2_fill_4 FILLER_141_74 ();
 sg13g2_fill_1 FILLER_141_78 ();
 sg13g2_fill_8 FILLER_141_89 ();
 sg13g2_fill_8 FILLER_141_97 ();
 sg13g2_fill_2 FILLER_141_105 ();
 sg13g2_fill_1 FILLER_141_107 ();
 sg13g2_fill_4 FILLER_141_118 ();
 sg13g2_fill_2 FILLER_141_122 ();
 sg13g2_fill_1 FILLER_141_124 ();
 sg13g2_fill_8 FILLER_141_135 ();
 sg13g2_fill_8 FILLER_141_143 ();
 sg13g2_fill_2 FILLER_141_151 ();
 sg13g2_fill_1 FILLER_141_153 ();
 sg13g2_fill_8 FILLER_141_162 ();
 sg13g2_fill_1 FILLER_141_175 ();
 sg13g2_fill_8 FILLER_141_186 ();
 sg13g2_fill_4 FILLER_141_194 ();
 sg13g2_fill_2 FILLER_141_198 ();
 sg13g2_fill_1 FILLER_141_200 ();
 sg13g2_fill_8 FILLER_141_211 ();
 sg13g2_fill_2 FILLER_141_219 ();
 sg13g2_fill_1 FILLER_141_221 ();
 sg13g2_fill_4 FILLER_141_232 ();
 sg13g2_fill_4 FILLER_141_252 ();
 sg13g2_fill_8 FILLER_141_302 ();
 sg13g2_fill_8 FILLER_141_310 ();
 sg13g2_fill_4 FILLER_141_318 ();
 sg13g2_fill_8 FILLER_141_330 ();
 sg13g2_fill_8 FILLER_141_338 ();
 sg13g2_fill_1 FILLER_141_372 ();
 sg13g2_fill_4 FILLER_141_394 ();
 sg13g2_fill_2 FILLER_141_398 ();
 sg13g2_fill_1 FILLER_141_400 ();
 sg13g2_fill_8 FILLER_141_411 ();
 sg13g2_fill_2 FILLER_141_419 ();
 sg13g2_fill_4 FILLER_141_431 ();
 sg13g2_fill_1 FILLER_141_435 ();
 sg13g2_fill_2 FILLER_141_462 ();
 sg13g2_fill_1 FILLER_141_464 ();
 sg13g2_fill_8 FILLER_141_475 ();
 sg13g2_fill_4 FILLER_141_483 ();
 sg13g2_fill_2 FILLER_141_487 ();
 sg13g2_fill_2 FILLER_141_521 ();
 sg13g2_fill_1 FILLER_141_561 ();
 sg13g2_fill_2 FILLER_141_572 ();
 sg13g2_fill_1 FILLER_141_574 ();
 sg13g2_fill_8 FILLER_141_585 ();
 sg13g2_fill_8 FILLER_141_593 ();
 sg13g2_fill_8 FILLER_141_601 ();
 sg13g2_fill_8 FILLER_141_609 ();
 sg13g2_fill_4 FILLER_141_617 ();
 sg13g2_fill_1 FILLER_141_621 ();
 sg13g2_fill_4 FILLER_141_630 ();
 sg13g2_fill_1 FILLER_141_634 ();
 sg13g2_fill_4 FILLER_141_641 ();
 sg13g2_fill_8 FILLER_141_651 ();
 sg13g2_fill_8 FILLER_141_685 ();
 sg13g2_fill_8 FILLER_141_693 ();
 sg13g2_fill_8 FILLER_141_701 ();
 sg13g2_fill_8 FILLER_141_709 ();
 sg13g2_fill_1 FILLER_141_717 ();
 sg13g2_fill_2 FILLER_141_755 ();
 sg13g2_fill_1 FILLER_141_757 ();
 sg13g2_fill_4 FILLER_141_765 ();
 sg13g2_fill_8 FILLER_141_782 ();
 sg13g2_fill_2 FILLER_141_790 ();
 sg13g2_fill_1 FILLER_141_792 ();
 sg13g2_fill_8 FILLER_141_855 ();
 sg13g2_fill_4 FILLER_141_863 ();
 sg13g2_fill_1 FILLER_141_867 ();
 sg13g2_fill_4 FILLER_141_1005 ();
 sg13g2_fill_2 FILLER_141_1009 ();
 sg13g2_fill_1 FILLER_141_1011 ();
 sg13g2_fill_2 FILLER_141_1032 ();
 sg13g2_fill_4 FILLER_141_1057 ();
 sg13g2_fill_1 FILLER_141_1061 ();
 sg13g2_fill_1 FILLER_141_1070 ();
 sg13g2_fill_2 FILLER_141_1084 ();
 sg13g2_fill_1 FILLER_141_1112 ();
 sg13g2_fill_2 FILLER_141_1148 ();
 sg13g2_fill_1 FILLER_141_1150 ();
 sg13g2_fill_8 FILLER_141_1192 ();
 sg13g2_fill_4 FILLER_141_1200 ();
 sg13g2_fill_4 FILLER_141_1207 ();
 sg13g2_fill_2 FILLER_141_1211 ();
 sg13g2_fill_1 FILLER_141_1213 ();
 sg13g2_fill_4 FILLER_141_1278 ();
 sg13g2_fill_4 FILLER_141_1287 ();
 sg13g2_fill_1 FILLER_141_1291 ();
 sg13g2_fill_1 FILLER_141_1300 ();
 sg13g2_fill_4 FILLER_141_1314 ();
 sg13g2_fill_2 FILLER_141_1318 ();
 sg13g2_fill_4 FILLER_141_1325 ();
 sg13g2_fill_1 FILLER_141_1329 ();
 sg13g2_fill_4 FILLER_141_1339 ();
 sg13g2_fill_2 FILLER_141_1343 ();
 sg13g2_fill_1 FILLER_141_1345 ();
 sg13g2_fill_4 FILLER_141_1359 ();
 sg13g2_fill_1 FILLER_141_1363 ();
 sg13g2_fill_2 FILLER_141_1379 ();
 sg13g2_fill_2 FILLER_141_1389 ();
 sg13g2_fill_2 FILLER_141_1417 ();
 sg13g2_fill_1 FILLER_141_1419 ();
 sg13g2_fill_8 FILLER_141_1446 ();
 sg13g2_fill_8 FILLER_141_1454 ();
 sg13g2_fill_8 FILLER_141_1462 ();
 sg13g2_fill_8 FILLER_141_1470 ();
 sg13g2_fill_2 FILLER_141_1478 ();
 sg13g2_fill_1 FILLER_141_1480 ();
 sg13g2_fill_2 FILLER_141_1499 ();
 sg13g2_fill_4 FILLER_141_1543 ();
 sg13g2_fill_1 FILLER_141_1547 ();
 sg13g2_fill_8 FILLER_141_1568 ();
 sg13g2_fill_8 FILLER_141_1576 ();
 sg13g2_fill_8 FILLER_141_1584 ();
 sg13g2_fill_4 FILLER_142_0 ();
 sg13g2_fill_2 FILLER_142_4 ();
 sg13g2_fill_1 FILLER_142_6 ();
 sg13g2_fill_8 FILLER_142_43 ();
 sg13g2_fill_4 FILLER_142_51 ();
 sg13g2_fill_2 FILLER_142_55 ();
 sg13g2_fill_1 FILLER_142_57 ();
 sg13g2_fill_4 FILLER_142_84 ();
 sg13g2_fill_2 FILLER_142_88 ();
 sg13g2_fill_8 FILLER_142_100 ();
 sg13g2_fill_1 FILLER_142_108 ();
 sg13g2_fill_2 FILLER_142_171 ();
 sg13g2_fill_1 FILLER_142_173 ();
 sg13g2_fill_8 FILLER_142_252 ();
 sg13g2_fill_8 FILLER_142_260 ();
 sg13g2_fill_8 FILLER_142_268 ();
 sg13g2_fill_8 FILLER_142_276 ();
 sg13g2_fill_8 FILLER_142_284 ();
 sg13g2_fill_1 FILLER_142_292 ();
 sg13g2_fill_4 FILLER_142_301 ();
 sg13g2_fill_1 FILLER_142_305 ();
 sg13g2_fill_8 FILLER_142_319 ();
 sg13g2_fill_1 FILLER_142_327 ();
 sg13g2_fill_8 FILLER_142_336 ();
 sg13g2_fill_1 FILLER_142_344 ();
 sg13g2_fill_8 FILLER_142_376 ();
 sg13g2_fill_8 FILLER_142_436 ();
 sg13g2_fill_8 FILLER_142_444 ();
 sg13g2_fill_8 FILLER_142_452 ();
 sg13g2_fill_4 FILLER_142_460 ();
 sg13g2_fill_2 FILLER_142_464 ();
 sg13g2_fill_1 FILLER_142_466 ();
 sg13g2_fill_2 FILLER_142_503 ();
 sg13g2_fill_2 FILLER_142_515 ();
 sg13g2_fill_1 FILLER_142_543 ();
 sg13g2_fill_4 FILLER_142_552 ();
 sg13g2_fill_2 FILLER_142_592 ();
 sg13g2_fill_1 FILLER_142_594 ();
 sg13g2_fill_8 FILLER_142_654 ();
 sg13g2_fill_4 FILLER_142_662 ();
 sg13g2_fill_1 FILLER_142_666 ();
 sg13g2_fill_8 FILLER_142_677 ();
 sg13g2_fill_4 FILLER_142_685 ();
 sg13g2_fill_2 FILLER_142_689 ();
 sg13g2_fill_1 FILLER_142_691 ();
 sg13g2_fill_8 FILLER_142_702 ();
 sg13g2_fill_4 FILLER_142_710 ();
 sg13g2_fill_1 FILLER_142_714 ();
 sg13g2_fill_8 FILLER_142_725 ();
 sg13g2_fill_8 FILLER_142_733 ();
 sg13g2_fill_8 FILLER_142_741 ();
 sg13g2_fill_2 FILLER_142_749 ();
 sg13g2_fill_1 FILLER_142_751 ();
 sg13g2_fill_4 FILLER_142_756 ();
 sg13g2_fill_1 FILLER_142_760 ();
 sg13g2_fill_8 FILLER_142_776 ();
 sg13g2_fill_4 FILLER_142_784 ();
 sg13g2_fill_2 FILLER_142_788 ();
 sg13g2_fill_2 FILLER_142_816 ();
 sg13g2_fill_1 FILLER_142_818 ();
 sg13g2_fill_8 FILLER_142_829 ();
 sg13g2_fill_8 FILLER_142_837 ();
 sg13g2_fill_8 FILLER_142_845 ();
 sg13g2_fill_8 FILLER_142_853 ();
 sg13g2_fill_8 FILLER_142_861 ();
 sg13g2_fill_2 FILLER_142_869 ();
 sg13g2_fill_1 FILLER_142_871 ();
 sg13g2_fill_2 FILLER_142_902 ();
 sg13g2_fill_4 FILLER_142_912 ();
 sg13g2_fill_2 FILLER_142_916 ();
 sg13g2_fill_8 FILLER_142_938 ();
 sg13g2_fill_8 FILLER_142_946 ();
 sg13g2_fill_4 FILLER_142_954 ();
 sg13g2_fill_1 FILLER_142_958 ();
 sg13g2_fill_4 FILLER_142_965 ();
 sg13g2_fill_1 FILLER_142_969 ();
 sg13g2_fill_2 FILLER_142_1010 ();
 sg13g2_fill_1 FILLER_142_1012 ();
 sg13g2_fill_8 FILLER_142_1023 ();
 sg13g2_fill_8 FILLER_142_1031 ();
 sg13g2_fill_2 FILLER_142_1079 ();
 sg13g2_fill_2 FILLER_142_1095 ();
 sg13g2_fill_1 FILLER_142_1097 ();
 sg13g2_fill_8 FILLER_142_1103 ();
 sg13g2_fill_2 FILLER_142_1141 ();
 sg13g2_fill_4 FILLER_142_1173 ();
 sg13g2_fill_2 FILLER_142_1229 ();
 sg13g2_fill_1 FILLER_142_1264 ();
 sg13g2_fill_4 FILLER_142_1275 ();
 sg13g2_fill_1 FILLER_142_1283 ();
 sg13g2_fill_1 FILLER_142_1318 ();
 sg13g2_fill_4 FILLER_142_1324 ();
 sg13g2_fill_1 FILLER_142_1328 ();
 sg13g2_fill_4 FILLER_142_1334 ();
 sg13g2_fill_2 FILLER_142_1356 ();
 sg13g2_fill_1 FILLER_142_1358 ();
 sg13g2_fill_1 FILLER_142_1377 ();
 sg13g2_fill_2 FILLER_142_1426 ();
 sg13g2_fill_2 FILLER_142_1442 ();
 sg13g2_fill_8 FILLER_142_1452 ();
 sg13g2_fill_2 FILLER_142_1486 ();
 sg13g2_fill_8 FILLER_142_1501 ();
 sg13g2_fill_8 FILLER_142_1509 ();
 sg13g2_fill_8 FILLER_142_1517 ();
 sg13g2_fill_8 FILLER_142_1525 ();
 sg13g2_fill_1 FILLER_142_1533 ();
 sg13g2_fill_4 FILLER_142_1544 ();
 sg13g2_fill_2 FILLER_142_1563 ();
 sg13g2_fill_1 FILLER_142_1591 ();
 sg13g2_fill_8 FILLER_143_0 ();
 sg13g2_fill_8 FILLER_143_18 ();
 sg13g2_fill_2 FILLER_143_26 ();
 sg13g2_fill_1 FILLER_143_28 ();
 sg13g2_fill_8 FILLER_143_39 ();
 sg13g2_fill_8 FILLER_143_47 ();
 sg13g2_fill_2 FILLER_143_55 ();
 sg13g2_fill_1 FILLER_143_57 ();
 sg13g2_fill_8 FILLER_143_84 ();
 sg13g2_fill_1 FILLER_143_92 ();
 sg13g2_fill_2 FILLER_143_119 ();
 sg13g2_fill_1 FILLER_143_121 ();
 sg13g2_fill_8 FILLER_143_144 ();
 sg13g2_fill_2 FILLER_143_152 ();
 sg13g2_fill_1 FILLER_143_154 ();
 sg13g2_fill_8 FILLER_143_160 ();
 sg13g2_fill_8 FILLER_143_168 ();
 sg13g2_fill_4 FILLER_143_176 ();
 sg13g2_fill_2 FILLER_143_201 ();
 sg13g2_fill_8 FILLER_143_213 ();
 sg13g2_fill_8 FILLER_143_221 ();
 sg13g2_fill_8 FILLER_143_229 ();
 sg13g2_fill_4 FILLER_143_237 ();
 sg13g2_fill_1 FILLER_143_249 ();
 sg13g2_fill_2 FILLER_143_276 ();
 sg13g2_fill_4 FILLER_143_304 ();
 sg13g2_fill_8 FILLER_143_313 ();
 sg13g2_fill_2 FILLER_143_321 ();
 sg13g2_fill_8 FILLER_143_366 ();
 sg13g2_fill_8 FILLER_143_374 ();
 sg13g2_fill_8 FILLER_143_382 ();
 sg13g2_fill_8 FILLER_143_390 ();
 sg13g2_fill_8 FILLER_143_398 ();
 sg13g2_fill_8 FILLER_143_406 ();
 sg13g2_fill_8 FILLER_143_414 ();
 sg13g2_fill_8 FILLER_143_422 ();
 sg13g2_fill_4 FILLER_143_430 ();
 sg13g2_fill_8 FILLER_143_439 ();
 sg13g2_fill_2 FILLER_143_460 ();
 sg13g2_fill_1 FILLER_143_462 ();
 sg13g2_fill_8 FILLER_143_489 ();
 sg13g2_fill_2 FILLER_143_497 ();
 sg13g2_fill_1 FILLER_143_499 ();
 sg13g2_fill_8 FILLER_143_517 ();
 sg13g2_fill_4 FILLER_143_525 ();
 sg13g2_fill_1 FILLER_143_529 ();
 sg13g2_fill_8 FILLER_143_556 ();
 sg13g2_fill_1 FILLER_143_564 ();
 sg13g2_fill_8 FILLER_143_579 ();
 sg13g2_fill_8 FILLER_143_587 ();
 sg13g2_fill_4 FILLER_143_595 ();
 sg13g2_fill_2 FILLER_143_599 ();
 sg13g2_fill_1 FILLER_143_601 ();
 sg13g2_fill_8 FILLER_143_608 ();
 sg13g2_fill_8 FILLER_143_616 ();
 sg13g2_fill_8 FILLER_143_624 ();
 sg13g2_fill_4 FILLER_143_632 ();
 sg13g2_fill_2 FILLER_143_636 ();
 sg13g2_fill_2 FILLER_143_649 ();
 sg13g2_fill_1 FILLER_143_662 ();
 sg13g2_fill_2 FILLER_143_725 ();
 sg13g2_fill_4 FILLER_143_750 ();
 sg13g2_fill_2 FILLER_143_800 ();
 sg13g2_fill_1 FILLER_143_802 ();
 sg13g2_fill_8 FILLER_143_808 ();
 sg13g2_fill_1 FILLER_143_841 ();
 sg13g2_fill_2 FILLER_143_847 ();
 sg13g2_fill_4 FILLER_143_854 ();
 sg13g2_fill_2 FILLER_143_858 ();
 sg13g2_fill_1 FILLER_143_860 ();
 sg13g2_fill_8 FILLER_143_881 ();
 sg13g2_fill_8 FILLER_143_889 ();
 sg13g2_fill_8 FILLER_143_897 ();
 sg13g2_fill_8 FILLER_143_905 ();
 sg13g2_fill_2 FILLER_143_913 ();
 sg13g2_fill_1 FILLER_143_915 ();
 sg13g2_fill_8 FILLER_143_941 ();
 sg13g2_fill_8 FILLER_143_949 ();
 sg13g2_fill_1 FILLER_143_957 ();
 sg13g2_fill_2 FILLER_143_961 ();
 sg13g2_fill_8 FILLER_143_976 ();
 sg13g2_fill_8 FILLER_143_984 ();
 sg13g2_fill_2 FILLER_143_1005 ();
 sg13g2_fill_1 FILLER_143_1007 ();
 sg13g2_fill_1 FILLER_143_1013 ();
 sg13g2_fill_8 FILLER_143_1032 ();
 sg13g2_fill_8 FILLER_143_1040 ();
 sg13g2_fill_4 FILLER_143_1048 ();
 sg13g2_fill_2 FILLER_143_1087 ();
 sg13g2_fill_8 FILLER_143_1108 ();
 sg13g2_fill_8 FILLER_143_1116 ();
 sg13g2_fill_2 FILLER_143_1124 ();
 sg13g2_fill_8 FILLER_143_1129 ();
 sg13g2_fill_8 FILLER_143_1166 ();
 sg13g2_fill_2 FILLER_143_1174 ();
 sg13g2_fill_1 FILLER_143_1176 ();
 sg13g2_fill_4 FILLER_143_1189 ();
 sg13g2_fill_1 FILLER_143_1193 ();
 sg13g2_fill_8 FILLER_143_1198 ();
 sg13g2_fill_8 FILLER_143_1206 ();
 sg13g2_fill_8 FILLER_143_1214 ();
 sg13g2_fill_8 FILLER_143_1222 ();
 sg13g2_fill_2 FILLER_143_1230 ();
 sg13g2_fill_1 FILLER_143_1232 ();
 sg13g2_fill_8 FILLER_143_1238 ();
 sg13g2_fill_4 FILLER_143_1246 ();
 sg13g2_fill_2 FILLER_143_1250 ();
 sg13g2_fill_1 FILLER_143_1252 ();
 sg13g2_fill_4 FILLER_143_1256 ();
 sg13g2_fill_1 FILLER_143_1260 ();
 sg13g2_fill_1 FILLER_143_1269 ();
 sg13g2_fill_2 FILLER_143_1273 ();
 sg13g2_fill_4 FILLER_143_1285 ();
 sg13g2_fill_2 FILLER_143_1289 ();
 sg13g2_fill_1 FILLER_143_1291 ();
 sg13g2_fill_2 FILLER_143_1303 ();
 sg13g2_fill_1 FILLER_143_1305 ();
 sg13g2_fill_4 FILLER_143_1316 ();
 sg13g2_fill_1 FILLER_143_1320 ();
 sg13g2_fill_8 FILLER_143_1325 ();
 sg13g2_fill_4 FILLER_143_1333 ();
 sg13g2_fill_2 FILLER_143_1337 ();
 sg13g2_fill_1 FILLER_143_1339 ();
 sg13g2_fill_4 FILLER_143_1345 ();
 sg13g2_fill_2 FILLER_143_1349 ();
 sg13g2_fill_2 FILLER_143_1364 ();
 sg13g2_fill_1 FILLER_143_1377 ();
 sg13g2_fill_2 FILLER_143_1399 ();
 sg13g2_fill_8 FILLER_143_1419 ();
 sg13g2_fill_1 FILLER_143_1427 ();
 sg13g2_fill_8 FILLER_143_1433 ();
 sg13g2_fill_8 FILLER_143_1451 ();
 sg13g2_fill_8 FILLER_143_1459 ();
 sg13g2_fill_8 FILLER_143_1467 ();
 sg13g2_fill_2 FILLER_143_1475 ();
 sg13g2_fill_1 FILLER_143_1477 ();
 sg13g2_fill_4 FILLER_143_1483 ();
 sg13g2_fill_2 FILLER_143_1498 ();
 sg13g2_fill_1 FILLER_143_1500 ();
 sg13g2_fill_2 FILLER_143_1513 ();
 sg13g2_fill_1 FILLER_143_1515 ();
 sg13g2_fill_8 FILLER_143_1542 ();
 sg13g2_fill_4 FILLER_143_1550 ();
 sg13g2_fill_2 FILLER_143_1554 ();
 sg13g2_fill_8 FILLER_144_0 ();
 sg13g2_fill_8 FILLER_144_8 ();
 sg13g2_fill_8 FILLER_144_16 ();
 sg13g2_fill_8 FILLER_144_24 ();
 sg13g2_fill_1 FILLER_144_32 ();
 sg13g2_fill_8 FILLER_144_59 ();
 sg13g2_fill_8 FILLER_144_67 ();
 sg13g2_fill_4 FILLER_144_75 ();
 sg13g2_fill_1 FILLER_144_79 ();
 sg13g2_fill_8 FILLER_144_90 ();
 sg13g2_fill_8 FILLER_144_98 ();
 sg13g2_fill_2 FILLER_144_106 ();
 sg13g2_fill_1 FILLER_144_108 ();
 sg13g2_fill_8 FILLER_144_119 ();
 sg13g2_fill_8 FILLER_144_137 ();
 sg13g2_fill_8 FILLER_144_145 ();
 sg13g2_fill_8 FILLER_144_153 ();
 sg13g2_fill_8 FILLER_144_161 ();
 sg13g2_fill_2 FILLER_144_169 ();
 sg13g2_fill_8 FILLER_144_205 ();
 sg13g2_fill_4 FILLER_144_213 ();
 sg13g2_fill_1 FILLER_144_217 ();
 sg13g2_fill_4 FILLER_144_247 ();
 sg13g2_fill_8 FILLER_144_261 ();
 sg13g2_fill_2 FILLER_144_269 ();
 sg13g2_fill_1 FILLER_144_271 ();
 sg13g2_fill_8 FILLER_144_282 ();
 sg13g2_fill_8 FILLER_144_290 ();
 sg13g2_fill_4 FILLER_144_298 ();
 sg13g2_fill_2 FILLER_144_302 ();
 sg13g2_fill_4 FILLER_144_354 ();
 sg13g2_fill_2 FILLER_144_358 ();
 sg13g2_fill_4 FILLER_144_396 ();
 sg13g2_fill_1 FILLER_144_410 ();
 sg13g2_fill_4 FILLER_144_421 ();
 sg13g2_fill_8 FILLER_144_435 ();
 sg13g2_fill_4 FILLER_144_443 ();
 sg13g2_fill_4 FILLER_144_455 ();
 sg13g2_fill_2 FILLER_144_459 ();
 sg13g2_fill_8 FILLER_144_471 ();
 sg13g2_fill_8 FILLER_144_479 ();
 sg13g2_fill_8 FILLER_144_487 ();
 sg13g2_fill_8 FILLER_144_495 ();
 sg13g2_fill_8 FILLER_144_503 ();
 sg13g2_fill_4 FILLER_144_511 ();
 sg13g2_fill_1 FILLER_144_515 ();
 sg13g2_fill_8 FILLER_144_524 ();
 sg13g2_fill_8 FILLER_144_532 ();
 sg13g2_fill_4 FILLER_144_540 ();
 sg13g2_fill_2 FILLER_144_544 ();
 sg13g2_fill_8 FILLER_144_556 ();
 sg13g2_fill_8 FILLER_144_568 ();
 sg13g2_fill_4 FILLER_144_610 ();
 sg13g2_fill_2 FILLER_144_614 ();
 sg13g2_fill_1 FILLER_144_616 ();
 sg13g2_fill_8 FILLER_144_621 ();
 sg13g2_fill_8 FILLER_144_629 ();
 sg13g2_fill_2 FILLER_144_637 ();
 sg13g2_fill_1 FILLER_144_639 ();
 sg13g2_fill_8 FILLER_144_681 ();
 sg13g2_fill_1 FILLER_144_689 ();
 sg13g2_fill_8 FILLER_144_698 ();
 sg13g2_fill_4 FILLER_144_706 ();
 sg13g2_fill_2 FILLER_144_710 ();
 sg13g2_fill_2 FILLER_144_720 ();
 sg13g2_fill_4 FILLER_144_732 ();
 sg13g2_fill_1 FILLER_144_749 ();
 sg13g2_fill_2 FILLER_144_755 ();
 sg13g2_fill_1 FILLER_144_757 ();
 sg13g2_fill_8 FILLER_144_791 ();
 sg13g2_fill_8 FILLER_144_799 ();
 sg13g2_fill_8 FILLER_144_807 ();
 sg13g2_fill_4 FILLER_144_815 ();
 sg13g2_fill_2 FILLER_144_824 ();
 sg13g2_fill_1 FILLER_144_826 ();
 sg13g2_fill_2 FILLER_144_844 ();
 sg13g2_fill_8 FILLER_144_863 ();
 sg13g2_fill_8 FILLER_144_871 ();
 sg13g2_fill_8 FILLER_144_879 ();
 sg13g2_fill_8 FILLER_144_887 ();
 sg13g2_fill_8 FILLER_144_895 ();
 sg13g2_fill_8 FILLER_144_937 ();
 sg13g2_fill_8 FILLER_144_945 ();
 sg13g2_fill_8 FILLER_144_962 ();
 sg13g2_fill_8 FILLER_144_970 ();
 sg13g2_fill_2 FILLER_144_978 ();
 sg13g2_fill_8 FILLER_144_989 ();
 sg13g2_fill_8 FILLER_144_997 ();
 sg13g2_fill_1 FILLER_144_1005 ();
 sg13g2_fill_1 FILLER_144_1011 ();
 sg13g2_fill_4 FILLER_144_1023 ();
 sg13g2_fill_1 FILLER_144_1027 ();
 sg13g2_fill_1 FILLER_144_1038 ();
 sg13g2_fill_2 FILLER_144_1079 ();
 sg13g2_fill_8 FILLER_144_1115 ();
 sg13g2_fill_8 FILLER_144_1139 ();
 sg13g2_fill_1 FILLER_144_1147 ();
 sg13g2_fill_1 FILLER_144_1153 ();
 sg13g2_fill_2 FILLER_144_1159 ();
 sg13g2_fill_1 FILLER_144_1161 ();
 sg13g2_fill_4 FILLER_144_1172 ();
 sg13g2_fill_1 FILLER_144_1176 ();
 sg13g2_fill_8 FILLER_144_1188 ();
 sg13g2_fill_8 FILLER_144_1196 ();
 sg13g2_fill_2 FILLER_144_1204 ();
 sg13g2_fill_1 FILLER_144_1209 ();
 sg13g2_fill_4 FILLER_144_1225 ();
 sg13g2_fill_1 FILLER_144_1229 ();
 sg13g2_fill_2 FILLER_144_1235 ();
 sg13g2_fill_1 FILLER_144_1237 ();
 sg13g2_fill_4 FILLER_144_1249 ();
 sg13g2_fill_1 FILLER_144_1264 ();
 sg13g2_fill_2 FILLER_144_1273 ();
 sg13g2_fill_2 FILLER_144_1289 ();
 sg13g2_fill_1 FILLER_144_1291 ();
 sg13g2_fill_1 FILLER_144_1295 ();
 sg13g2_fill_8 FILLER_144_1303 ();
 sg13g2_fill_8 FILLER_144_1311 ();
 sg13g2_fill_4 FILLER_144_1319 ();
 sg13g2_fill_1 FILLER_144_1323 ();
 sg13g2_fill_8 FILLER_144_1334 ();
 sg13g2_fill_8 FILLER_144_1342 ();
 sg13g2_fill_8 FILLER_144_1350 ();
 sg13g2_fill_2 FILLER_144_1409 ();
 sg13g2_fill_2 FILLER_144_1419 ();
 sg13g2_fill_8 FILLER_144_1428 ();
 sg13g2_fill_8 FILLER_144_1441 ();
 sg13g2_fill_4 FILLER_144_1449 ();
 sg13g2_fill_1 FILLER_144_1453 ();
 sg13g2_fill_2 FILLER_144_1496 ();
 sg13g2_fill_4 FILLER_144_1507 ();
 sg13g2_fill_8 FILLER_144_1530 ();
 sg13g2_fill_4 FILLER_144_1550 ();
 sg13g2_fill_8 FILLER_144_1565 ();
 sg13g2_fill_8 FILLER_144_1573 ();
 sg13g2_fill_8 FILLER_144_1581 ();
 sg13g2_fill_2 FILLER_144_1589 ();
 sg13g2_fill_1 FILLER_144_1591 ();
 sg13g2_fill_8 FILLER_145_0 ();
 sg13g2_fill_4 FILLER_145_8 ();
 sg13g2_fill_1 FILLER_145_12 ();
 sg13g2_fill_4 FILLER_145_68 ();
 sg13g2_fill_2 FILLER_145_72 ();
 sg13g2_fill_1 FILLER_145_74 ();
 sg13g2_fill_4 FILLER_145_85 ();
 sg13g2_fill_8 FILLER_145_99 ();
 sg13g2_fill_4 FILLER_145_107 ();
 sg13g2_fill_2 FILLER_145_111 ();
 sg13g2_fill_1 FILLER_145_113 ();
 sg13g2_fill_4 FILLER_145_124 ();
 sg13g2_fill_2 FILLER_145_128 ();
 sg13g2_fill_1 FILLER_145_130 ();
 sg13g2_fill_2 FILLER_145_142 ();
 sg13g2_fill_2 FILLER_145_149 ();
 sg13g2_fill_1 FILLER_145_151 ();
 sg13g2_fill_8 FILLER_145_213 ();
 sg13g2_fill_4 FILLER_145_221 ();
 sg13g2_fill_2 FILLER_145_225 ();
 sg13g2_fill_1 FILLER_145_227 ();
 sg13g2_fill_8 FILLER_145_263 ();
 sg13g2_fill_8 FILLER_145_271 ();
 sg13g2_fill_2 FILLER_145_279 ();
 sg13g2_fill_1 FILLER_145_281 ();
 sg13g2_fill_1 FILLER_145_326 ();
 sg13g2_fill_8 FILLER_145_337 ();
 sg13g2_fill_4 FILLER_145_345 ();
 sg13g2_fill_1 FILLER_145_349 ();
 sg13g2_fill_8 FILLER_145_371 ();
 sg13g2_fill_8 FILLER_145_379 ();
 sg13g2_fill_2 FILLER_145_387 ();
 sg13g2_fill_4 FILLER_145_415 ();
 sg13g2_fill_2 FILLER_145_419 ();
 sg13g2_fill_1 FILLER_145_475 ();
 sg13g2_fill_2 FILLER_145_515 ();
 sg13g2_fill_1 FILLER_145_517 ();
 sg13g2_fill_2 FILLER_145_526 ();
 sg13g2_fill_1 FILLER_145_528 ();
 sg13g2_fill_2 FILLER_145_636 ();
 sg13g2_fill_4 FILLER_145_659 ();
 sg13g2_fill_2 FILLER_145_663 ();
 sg13g2_fill_1 FILLER_145_675 ();
 sg13g2_fill_8 FILLER_145_702 ();
 sg13g2_fill_8 FILLER_145_710 ();
 sg13g2_fill_4 FILLER_145_718 ();
 sg13g2_fill_8 FILLER_145_726 ();
 sg13g2_fill_2 FILLER_145_734 ();
 sg13g2_fill_1 FILLER_145_736 ();
 sg13g2_fill_2 FILLER_145_754 ();
 sg13g2_fill_1 FILLER_145_756 ();
 sg13g2_fill_1 FILLER_145_765 ();
 sg13g2_fill_8 FILLER_145_786 ();
 sg13g2_fill_2 FILLER_145_794 ();
 sg13g2_fill_1 FILLER_145_796 ();
 sg13g2_fill_4 FILLER_145_802 ();
 sg13g2_fill_1 FILLER_145_806 ();
 sg13g2_fill_1 FILLER_145_811 ();
 sg13g2_fill_1 FILLER_145_817 ();
 sg13g2_fill_8 FILLER_145_827 ();
 sg13g2_fill_8 FILLER_145_835 ();
 sg13g2_fill_2 FILLER_145_848 ();
 sg13g2_fill_1 FILLER_145_860 ();
 sg13g2_fill_2 FILLER_145_870 ();
 sg13g2_fill_4 FILLER_145_886 ();
 sg13g2_fill_1 FILLER_145_890 ();
 sg13g2_fill_1 FILLER_145_957 ();
 sg13g2_fill_1 FILLER_145_966 ();
 sg13g2_fill_2 FILLER_145_983 ();
 sg13g2_fill_8 FILLER_145_996 ();
 sg13g2_fill_4 FILLER_145_1004 ();
 sg13g2_fill_2 FILLER_145_1008 ();
 sg13g2_fill_2 FILLER_145_1015 ();
 sg13g2_fill_1 FILLER_145_1017 ();
 sg13g2_fill_4 FILLER_145_1023 ();
 sg13g2_fill_2 FILLER_145_1027 ();
 sg13g2_fill_2 FILLER_145_1034 ();
 sg13g2_fill_2 FILLER_145_1064 ();
 sg13g2_fill_1 FILLER_145_1066 ();
 sg13g2_fill_8 FILLER_145_1071 ();
 sg13g2_fill_4 FILLER_145_1079 ();
 sg13g2_fill_8 FILLER_145_1087 ();
 sg13g2_fill_2 FILLER_145_1095 ();
 sg13g2_fill_4 FILLER_145_1102 ();
 sg13g2_fill_4 FILLER_145_1110 ();
 sg13g2_fill_2 FILLER_145_1114 ();
 sg13g2_fill_1 FILLER_145_1131 ();
 sg13g2_fill_8 FILLER_145_1167 ();
 sg13g2_fill_2 FILLER_145_1175 ();
 sg13g2_fill_8 FILLER_145_1186 ();
 sg13g2_fill_8 FILLER_145_1194 ();
 sg13g2_fill_1 FILLER_145_1202 ();
 sg13g2_fill_8 FILLER_145_1210 ();
 sg13g2_fill_2 FILLER_145_1218 ();
 sg13g2_fill_2 FILLER_145_1229 ();
 sg13g2_fill_2 FILLER_145_1236 ();
 sg13g2_fill_1 FILLER_145_1238 ();
 sg13g2_fill_2 FILLER_145_1245 ();
 sg13g2_fill_1 FILLER_145_1247 ();
 sg13g2_fill_2 FILLER_145_1269 ();
 sg13g2_fill_8 FILLER_145_1275 ();
 sg13g2_fill_4 FILLER_145_1283 ();
 sg13g2_fill_2 FILLER_145_1287 ();
 sg13g2_fill_2 FILLER_145_1299 ();
 sg13g2_fill_1 FILLER_145_1301 ();
 sg13g2_fill_8 FILLER_145_1308 ();
 sg13g2_fill_1 FILLER_145_1316 ();
 sg13g2_fill_4 FILLER_145_1342 ();
 sg13g2_fill_1 FILLER_145_1346 ();
 sg13g2_fill_1 FILLER_145_1360 ();
 sg13g2_fill_1 FILLER_145_1399 ();
 sg13g2_fill_4 FILLER_145_1417 ();
 sg13g2_fill_1 FILLER_145_1430 ();
 sg13g2_fill_8 FILLER_145_1450 ();
 sg13g2_fill_8 FILLER_145_1458 ();
 sg13g2_fill_8 FILLER_145_1466 ();
 sg13g2_fill_4 FILLER_145_1474 ();
 sg13g2_fill_2 FILLER_145_1541 ();
 sg13g2_fill_2 FILLER_145_1553 ();
 sg13g2_fill_1 FILLER_145_1555 ();
 sg13g2_fill_8 FILLER_146_0 ();
 sg13g2_fill_8 FILLER_146_8 ();
 sg13g2_fill_8 FILLER_146_16 ();
 sg13g2_fill_4 FILLER_146_24 ();
 sg13g2_fill_4 FILLER_146_54 ();
 sg13g2_fill_8 FILLER_146_84 ();
 sg13g2_fill_8 FILLER_146_118 ();
 sg13g2_fill_1 FILLER_146_126 ();
 sg13g2_fill_8 FILLER_146_155 ();
 sg13g2_fill_8 FILLER_146_163 ();
 sg13g2_fill_1 FILLER_146_171 ();
 sg13g2_fill_4 FILLER_146_198 ();
 sg13g2_fill_2 FILLER_146_249 ();
 sg13g2_fill_4 FILLER_146_298 ();
 sg13g2_fill_4 FILLER_146_323 ();
 sg13g2_fill_1 FILLER_146_327 ();
 sg13g2_fill_8 FILLER_146_364 ();
 sg13g2_fill_8 FILLER_146_372 ();
 sg13g2_fill_8 FILLER_146_380 ();
 sg13g2_fill_8 FILLER_146_388 ();
 sg13g2_fill_8 FILLER_146_396 ();
 sg13g2_fill_2 FILLER_146_404 ();
 sg13g2_fill_1 FILLER_146_406 ();
 sg13g2_fill_8 FILLER_146_417 ();
 sg13g2_fill_2 FILLER_146_425 ();
 sg13g2_fill_8 FILLER_146_439 ();
 sg13g2_fill_8 FILLER_146_447 ();
 sg13g2_fill_8 FILLER_146_455 ();
 sg13g2_fill_4 FILLER_146_463 ();
 sg13g2_fill_1 FILLER_146_467 ();
 sg13g2_fill_2 FILLER_146_542 ();
 sg13g2_fill_1 FILLER_146_544 ();
 sg13g2_fill_8 FILLER_146_549 ();
 sg13g2_fill_8 FILLER_146_557 ();
 sg13g2_fill_4 FILLER_146_591 ();
 sg13g2_fill_2 FILLER_146_595 ();
 sg13g2_fill_2 FILLER_146_608 ();
 sg13g2_fill_8 FILLER_146_636 ();
 sg13g2_fill_1 FILLER_146_644 ();
 sg13g2_fill_8 FILLER_146_691 ();
 sg13g2_fill_4 FILLER_146_699 ();
 sg13g2_fill_8 FILLER_146_713 ();
 sg13g2_fill_4 FILLER_146_721 ();
 sg13g2_fill_2 FILLER_146_725 ();
 sg13g2_fill_8 FILLER_146_737 ();
 sg13g2_fill_8 FILLER_146_745 ();
 sg13g2_fill_1 FILLER_146_753 ();
 sg13g2_fill_4 FILLER_146_765 ();
 sg13g2_fill_2 FILLER_146_769 ();
 sg13g2_fill_8 FILLER_146_776 ();
 sg13g2_fill_1 FILLER_146_784 ();
 sg13g2_fill_1 FILLER_146_795 ();
 sg13g2_fill_1 FILLER_146_801 ();
 sg13g2_fill_4 FILLER_146_825 ();
 sg13g2_fill_2 FILLER_146_829 ();
 sg13g2_fill_1 FILLER_146_831 ();
 sg13g2_fill_8 FILLER_146_837 ();
 sg13g2_fill_8 FILLER_146_845 ();
 sg13g2_fill_8 FILLER_146_858 ();
 sg13g2_fill_1 FILLER_146_866 ();
 sg13g2_fill_4 FILLER_146_893 ();
 sg13g2_fill_4 FILLER_146_905 ();
 sg13g2_fill_4 FILLER_146_922 ();
 sg13g2_fill_1 FILLER_146_926 ();
 sg13g2_fill_8 FILLER_146_958 ();
 sg13g2_fill_8 FILLER_146_966 ();
 sg13g2_fill_4 FILLER_146_974 ();
 sg13g2_fill_1 FILLER_146_978 ();
 sg13g2_fill_4 FILLER_146_1014 ();
 sg13g2_fill_1 FILLER_146_1018 ();
 sg13g2_fill_4 FILLER_146_1024 ();
 sg13g2_fill_2 FILLER_146_1028 ();
 sg13g2_fill_4 FILLER_146_1053 ();
 sg13g2_fill_1 FILLER_146_1057 ();
 sg13g2_fill_2 FILLER_146_1071 ();
 sg13g2_fill_2 FILLER_146_1086 ();
 sg13g2_fill_1 FILLER_146_1088 ();
 sg13g2_fill_1 FILLER_146_1103 ();
 sg13g2_fill_4 FILLER_146_1134 ();
 sg13g2_fill_2 FILLER_146_1138 ();
 sg13g2_fill_1 FILLER_146_1140 ();
 sg13g2_fill_8 FILLER_146_1160 ();
 sg13g2_fill_1 FILLER_146_1168 ();
 sg13g2_fill_4 FILLER_146_1173 ();
 sg13g2_fill_2 FILLER_146_1206 ();
 sg13g2_fill_4 FILLER_146_1234 ();
 sg13g2_fill_2 FILLER_146_1250 ();
 sg13g2_fill_1 FILLER_146_1252 ();
 sg13g2_fill_2 FILLER_146_1277 ();
 sg13g2_fill_1 FILLER_146_1279 ();
 sg13g2_fill_1 FILLER_146_1285 ();
 sg13g2_fill_4 FILLER_146_1290 ();
 sg13g2_fill_1 FILLER_146_1298 ();
 sg13g2_fill_4 FILLER_146_1320 ();
 sg13g2_fill_2 FILLER_146_1324 ();
 sg13g2_fill_1 FILLER_146_1326 ();
 sg13g2_fill_2 FILLER_146_1342 ();
 sg13g2_fill_2 FILLER_146_1364 ();
 sg13g2_fill_2 FILLER_146_1397 ();
 sg13g2_fill_1 FILLER_146_1399 ();
 sg13g2_fill_2 FILLER_146_1424 ();
 sg13g2_fill_2 FILLER_146_1454 ();
 sg13g2_fill_4 FILLER_146_1494 ();
 sg13g2_fill_2 FILLER_146_1524 ();
 sg13g2_fill_1 FILLER_146_1526 ();
 sg13g2_fill_4 FILLER_146_1553 ();
 sg13g2_fill_1 FILLER_146_1557 ();
 sg13g2_fill_4 FILLER_146_1562 ();
 sg13g2_fill_1 FILLER_146_1591 ();
 sg13g2_fill_8 FILLER_147_0 ();
 sg13g2_fill_8 FILLER_147_8 ();
 sg13g2_fill_8 FILLER_147_16 ();
 sg13g2_fill_4 FILLER_147_24 ();
 sg13g2_fill_8 FILLER_147_64 ();
 sg13g2_fill_8 FILLER_147_72 ();
 sg13g2_fill_2 FILLER_147_80 ();
 sg13g2_fill_1 FILLER_147_82 ();
 sg13g2_fill_8 FILLER_147_89 ();
 sg13g2_fill_1 FILLER_147_97 ();
 sg13g2_fill_2 FILLER_147_133 ();
 sg13g2_fill_2 FILLER_147_160 ();
 sg13g2_fill_1 FILLER_147_162 ();
 sg13g2_fill_8 FILLER_147_188 ();
 sg13g2_fill_4 FILLER_147_196 ();
 sg13g2_fill_4 FILLER_147_223 ();
 sg13g2_fill_1 FILLER_147_227 ();
 sg13g2_fill_4 FILLER_147_231 ();
 sg13g2_fill_2 FILLER_147_243 ();
 sg13g2_fill_1 FILLER_147_245 ();
 sg13g2_fill_8 FILLER_147_251 ();
 sg13g2_fill_8 FILLER_147_259 ();
 sg13g2_fill_8 FILLER_147_267 ();
 sg13g2_fill_1 FILLER_147_296 ();
 sg13g2_fill_2 FILLER_147_327 ();
 sg13g2_fill_4 FILLER_147_354 ();
 sg13g2_fill_2 FILLER_147_358 ();
 sg13g2_fill_1 FILLER_147_360 ();
 sg13g2_fill_8 FILLER_147_387 ();
 sg13g2_fill_2 FILLER_147_395 ();
 sg13g2_fill_2 FILLER_147_407 ();
 sg13g2_fill_4 FILLER_147_439 ();
 sg13g2_fill_8 FILLER_147_453 ();
 sg13g2_fill_8 FILLER_147_461 ();
 sg13g2_fill_1 FILLER_147_469 ();
 sg13g2_fill_8 FILLER_147_521 ();
 sg13g2_fill_8 FILLER_147_529 ();
 sg13g2_fill_8 FILLER_147_537 ();
 sg13g2_fill_4 FILLER_147_545 ();
 sg13g2_fill_8 FILLER_147_553 ();
 sg13g2_fill_8 FILLER_147_575 ();
 sg13g2_fill_8 FILLER_147_583 ();
 sg13g2_fill_8 FILLER_147_591 ();
 sg13g2_fill_4 FILLER_147_599 ();
 sg13g2_fill_8 FILLER_147_607 ();
 sg13g2_fill_8 FILLER_147_615 ();
 sg13g2_fill_2 FILLER_147_623 ();
 sg13g2_fill_8 FILLER_147_651 ();
 sg13g2_fill_8 FILLER_147_659 ();
 sg13g2_fill_8 FILLER_147_667 ();
 sg13g2_fill_1 FILLER_147_675 ();
 sg13g2_fill_4 FILLER_147_684 ();
 sg13g2_fill_2 FILLER_147_688 ();
 sg13g2_fill_8 FILLER_147_752 ();
 sg13g2_fill_4 FILLER_147_760 ();
 sg13g2_fill_8 FILLER_147_768 ();
 sg13g2_fill_4 FILLER_147_776 ();
 sg13g2_fill_1 FILLER_147_780 ();
 sg13g2_fill_4 FILLER_147_805 ();
 sg13g2_fill_2 FILLER_147_809 ();
 sg13g2_fill_8 FILLER_147_820 ();
 sg13g2_fill_1 FILLER_147_828 ();
 sg13g2_fill_2 FILLER_147_840 ();
 sg13g2_fill_4 FILLER_147_848 ();
 sg13g2_fill_4 FILLER_147_870 ();
 sg13g2_fill_2 FILLER_147_874 ();
 sg13g2_fill_8 FILLER_147_886 ();
 sg13g2_fill_4 FILLER_147_894 ();
 sg13g2_fill_2 FILLER_147_898 ();
 sg13g2_fill_1 FILLER_147_900 ();
 sg13g2_fill_4 FILLER_147_939 ();
 sg13g2_fill_4 FILLER_147_957 ();
 sg13g2_fill_8 FILLER_147_973 ();
 sg13g2_fill_4 FILLER_147_981 ();
 sg13g2_fill_2 FILLER_147_985 ();
 sg13g2_fill_1 FILLER_147_987 ();
 sg13g2_fill_2 FILLER_147_993 ();
 sg13g2_fill_2 FILLER_147_1005 ();
 sg13g2_fill_1 FILLER_147_1007 ();
 sg13g2_fill_2 FILLER_147_1034 ();
 sg13g2_fill_8 FILLER_147_1042 ();
 sg13g2_fill_8 FILLER_147_1050 ();
 sg13g2_fill_4 FILLER_147_1058 ();
 sg13g2_fill_8 FILLER_147_1068 ();
 sg13g2_fill_8 FILLER_147_1076 ();
 sg13g2_fill_8 FILLER_147_1084 ();
 sg13g2_fill_2 FILLER_147_1092 ();
 sg13g2_fill_8 FILLER_147_1098 ();
 sg13g2_fill_8 FILLER_147_1106 ();
 sg13g2_fill_8 FILLER_147_1114 ();
 sg13g2_fill_4 FILLER_147_1122 ();
 sg13g2_fill_8 FILLER_147_1135 ();
 sg13g2_fill_2 FILLER_147_1143 ();
 sg13g2_fill_1 FILLER_147_1145 ();
 sg13g2_fill_8 FILLER_147_1154 ();
 sg13g2_fill_4 FILLER_147_1162 ();
 sg13g2_fill_1 FILLER_147_1166 ();
 sg13g2_fill_8 FILLER_147_1218 ();
 sg13g2_fill_8 FILLER_147_1226 ();
 sg13g2_fill_2 FILLER_147_1234 ();
 sg13g2_fill_1 FILLER_147_1236 ();
 sg13g2_fill_8 FILLER_147_1242 ();
 sg13g2_fill_8 FILLER_147_1250 ();
 sg13g2_fill_2 FILLER_147_1258 ();
 sg13g2_fill_1 FILLER_147_1260 ();
 sg13g2_fill_8 FILLER_147_1291 ();
 sg13g2_fill_1 FILLER_147_1299 ();
 sg13g2_fill_1 FILLER_147_1312 ();
 sg13g2_fill_8 FILLER_147_1332 ();
 sg13g2_fill_8 FILLER_147_1340 ();
 sg13g2_fill_8 FILLER_147_1348 ();
 sg13g2_fill_1 FILLER_147_1363 ();
 sg13g2_fill_2 FILLER_147_1374 ();
 sg13g2_fill_2 FILLER_147_1389 ();
 sg13g2_fill_8 FILLER_147_1416 ();
 sg13g2_fill_4 FILLER_147_1432 ();
 sg13g2_fill_1 FILLER_147_1436 ();
 sg13g2_fill_8 FILLER_147_1445 ();
 sg13g2_fill_8 FILLER_147_1453 ();
 sg13g2_fill_8 FILLER_147_1461 ();
 sg13g2_fill_1 FILLER_147_1485 ();
 sg13g2_fill_2 FILLER_147_1496 ();
 sg13g2_fill_1 FILLER_147_1498 ();
 sg13g2_fill_4 FILLER_147_1503 ();
 sg13g2_fill_1 FILLER_147_1507 ();
 sg13g2_fill_4 FILLER_147_1514 ();
 sg13g2_fill_2 FILLER_147_1518 ();
 sg13g2_fill_8 FILLER_147_1524 ();
 sg13g2_fill_8 FILLER_147_1532 ();
 sg13g2_fill_8 FILLER_147_1540 ();
 sg13g2_fill_2 FILLER_147_1548 ();
 sg13g2_fill_1 FILLER_147_1550 ();
 sg13g2_fill_8 FILLER_148_0 ();
 sg13g2_fill_8 FILLER_148_8 ();
 sg13g2_fill_8 FILLER_148_16 ();
 sg13g2_fill_8 FILLER_148_24 ();
 sg13g2_fill_8 FILLER_148_32 ();
 sg13g2_fill_8 FILLER_148_40 ();
 sg13g2_fill_2 FILLER_148_48 ();
 sg13g2_fill_1 FILLER_148_50 ();
 sg13g2_fill_8 FILLER_148_61 ();
 sg13g2_fill_2 FILLER_148_69 ();
 sg13g2_fill_1 FILLER_148_71 ();
 sg13g2_fill_2 FILLER_148_82 ();
 sg13g2_fill_4 FILLER_148_120 ();
 sg13g2_fill_2 FILLER_148_124 ();
 sg13g2_fill_1 FILLER_148_126 ();
 sg13g2_fill_2 FILLER_148_171 ();
 sg13g2_fill_1 FILLER_148_173 ();
 sg13g2_fill_8 FILLER_148_200 ();
 sg13g2_fill_4 FILLER_148_234 ();
 sg13g2_fill_1 FILLER_148_238 ();
 sg13g2_fill_8 FILLER_148_275 ();
 sg13g2_fill_4 FILLER_148_283 ();
 sg13g2_fill_2 FILLER_148_287 ();
 sg13g2_fill_2 FILLER_148_297 ();
 sg13g2_fill_1 FILLER_148_299 ();
 sg13g2_fill_1 FILLER_148_379 ();
 sg13g2_fill_2 FILLER_148_406 ();
 sg13g2_fill_1 FILLER_148_408 ();
 sg13g2_fill_2 FILLER_148_441 ();
 sg13g2_fill_8 FILLER_148_469 ();
 sg13g2_fill_8 FILLER_148_477 ();
 sg13g2_fill_4 FILLER_148_485 ();
 sg13g2_fill_2 FILLER_148_489 ();
 sg13g2_fill_4 FILLER_148_501 ();
 sg13g2_fill_2 FILLER_148_505 ();
 sg13g2_fill_8 FILLER_148_525 ();
 sg13g2_fill_2 FILLER_148_533 ();
 sg13g2_fill_1 FILLER_148_535 ();
 sg13g2_fill_4 FILLER_148_560 ();
 sg13g2_fill_2 FILLER_148_564 ();
 sg13g2_fill_1 FILLER_148_566 ();
 sg13g2_fill_2 FILLER_148_607 ();
 sg13g2_fill_1 FILLER_148_609 ();
 sg13g2_fill_4 FILLER_148_620 ();
 sg13g2_fill_2 FILLER_148_640 ();
 sg13g2_fill_1 FILLER_148_642 ();
 sg13g2_fill_4 FILLER_148_689 ();
 sg13g2_fill_2 FILLER_148_693 ();
 sg13g2_fill_1 FILLER_148_720 ();
 sg13g2_fill_8 FILLER_148_731 ();
 sg13g2_fill_8 FILLER_148_739 ();
 sg13g2_fill_1 FILLER_148_752 ();
 sg13g2_fill_8 FILLER_148_782 ();
 sg13g2_fill_8 FILLER_148_799 ();
 sg13g2_fill_4 FILLER_148_807 ();
 sg13g2_fill_1 FILLER_148_826 ();
 sg13g2_fill_1 FILLER_148_839 ();
 sg13g2_fill_4 FILLER_148_852 ();
 sg13g2_fill_2 FILLER_148_856 ();
 sg13g2_fill_8 FILLER_148_864 ();
 sg13g2_fill_2 FILLER_148_872 ();
 sg13g2_fill_1 FILLER_148_874 ();
 sg13g2_fill_2 FILLER_148_880 ();
 sg13g2_fill_4 FILLER_148_892 ();
 sg13g2_fill_2 FILLER_148_896 ();
 sg13g2_fill_2 FILLER_148_909 ();
 sg13g2_fill_1 FILLER_148_911 ();
 sg13g2_fill_1 FILLER_148_918 ();
 sg13g2_fill_2 FILLER_148_927 ();
 sg13g2_fill_1 FILLER_148_929 ();
 sg13g2_fill_1 FILLER_148_940 ();
 sg13g2_fill_8 FILLER_148_990 ();
 sg13g2_fill_8 FILLER_148_998 ();
 sg13g2_fill_4 FILLER_148_1010 ();
 sg13g2_fill_2 FILLER_148_1014 ();
 sg13g2_fill_1 FILLER_148_1016 ();
 sg13g2_fill_8 FILLER_148_1027 ();
 sg13g2_fill_4 FILLER_148_1035 ();
 sg13g2_fill_2 FILLER_148_1039 ();
 sg13g2_fill_4 FILLER_148_1054 ();
 sg13g2_fill_2 FILLER_148_1058 ();
 sg13g2_fill_1 FILLER_148_1060 ();
 sg13g2_fill_4 FILLER_148_1075 ();
 sg13g2_fill_4 FILLER_148_1099 ();
 sg13g2_fill_2 FILLER_148_1110 ();
 sg13g2_fill_1 FILLER_148_1120 ();
 sg13g2_fill_4 FILLER_148_1137 ();
 sg13g2_fill_1 FILLER_148_1141 ();
 sg13g2_fill_1 FILLER_148_1147 ();
 sg13g2_fill_1 FILLER_148_1188 ();
 sg13g2_fill_1 FILLER_148_1218 ();
 sg13g2_fill_1 FILLER_148_1226 ();
 sg13g2_fill_1 FILLER_148_1247 ();
 sg13g2_fill_4 FILLER_148_1252 ();
 sg13g2_fill_2 FILLER_148_1256 ();
 sg13g2_fill_1 FILLER_148_1258 ();
 sg13g2_fill_8 FILLER_148_1271 ();
 sg13g2_fill_4 FILLER_148_1279 ();
 sg13g2_fill_8 FILLER_148_1288 ();
 sg13g2_fill_4 FILLER_148_1296 ();
 sg13g2_fill_2 FILLER_148_1304 ();
 sg13g2_fill_1 FILLER_148_1306 ();
 sg13g2_fill_2 FILLER_148_1327 ();
 sg13g2_fill_1 FILLER_148_1329 ();
 sg13g2_fill_4 FILLER_148_1340 ();
 sg13g2_fill_2 FILLER_148_1344 ();
 sg13g2_fill_1 FILLER_148_1346 ();
 sg13g2_fill_4 FILLER_148_1358 ();
 sg13g2_fill_2 FILLER_148_1362 ();
 sg13g2_fill_2 FILLER_148_1378 ();
 sg13g2_fill_1 FILLER_148_1380 ();
 sg13g2_fill_1 FILLER_148_1403 ();
 sg13g2_fill_2 FILLER_148_1411 ();
 sg13g2_fill_1 FILLER_148_1413 ();
 sg13g2_fill_2 FILLER_148_1423 ();
 sg13g2_fill_1 FILLER_148_1425 ();
 sg13g2_fill_8 FILLER_148_1436 ();
 sg13g2_fill_8 FILLER_148_1444 ();
 sg13g2_fill_8 FILLER_148_1452 ();
 sg13g2_fill_2 FILLER_148_1460 ();
 sg13g2_fill_4 FILLER_148_1492 ();
 sg13g2_fill_2 FILLER_148_1522 ();
 sg13g2_fill_8 FILLER_148_1532 ();
 sg13g2_fill_4 FILLER_148_1540 ();
 sg13g2_fill_4 FILLER_148_1560 ();
 sg13g2_fill_2 FILLER_148_1564 ();
 sg13g2_fill_8 FILLER_149_0 ();
 sg13g2_fill_8 FILLER_149_8 ();
 sg13g2_fill_8 FILLER_149_16 ();
 sg13g2_fill_8 FILLER_149_24 ();
 sg13g2_fill_1 FILLER_149_32 ();
 sg13g2_fill_8 FILLER_149_59 ();
 sg13g2_fill_4 FILLER_149_67 ();
 sg13g2_fill_2 FILLER_149_71 ();
 sg13g2_fill_1 FILLER_149_73 ();
 sg13g2_fill_8 FILLER_149_90 ();
 sg13g2_fill_2 FILLER_149_98 ();
 sg13g2_fill_8 FILLER_149_116 ();
 sg13g2_fill_4 FILLER_149_124 ();
 sg13g2_fill_1 FILLER_149_128 ();
 sg13g2_fill_4 FILLER_149_160 ();
 sg13g2_fill_2 FILLER_149_164 ();
 sg13g2_fill_4 FILLER_149_176 ();
 sg13g2_fill_2 FILLER_149_180 ();
 sg13g2_fill_8 FILLER_149_192 ();
 sg13g2_fill_8 FILLER_149_200 ();
 sg13g2_fill_8 FILLER_149_208 ();
 sg13g2_fill_8 FILLER_149_216 ();
 sg13g2_fill_8 FILLER_149_224 ();
 sg13g2_fill_2 FILLER_149_232 ();
 sg13g2_fill_1 FILLER_149_234 ();
 sg13g2_fill_8 FILLER_149_243 ();
 sg13g2_fill_8 FILLER_149_251 ();
 sg13g2_fill_8 FILLER_149_259 ();
 sg13g2_fill_2 FILLER_149_267 ();
 sg13g2_fill_4 FILLER_149_298 ();
 sg13g2_fill_1 FILLER_149_302 ();
 sg13g2_fill_8 FILLER_149_313 ();
 sg13g2_fill_8 FILLER_149_321 ();
 sg13g2_fill_4 FILLER_149_329 ();
 sg13g2_fill_2 FILLER_149_333 ();
 sg13g2_fill_1 FILLER_149_335 ();
 sg13g2_fill_4 FILLER_149_357 ();
 sg13g2_fill_8 FILLER_149_387 ();
 sg13g2_fill_8 FILLER_149_395 ();
 sg13g2_fill_4 FILLER_149_403 ();
 sg13g2_fill_2 FILLER_149_407 ();
 sg13g2_fill_2 FILLER_149_419 ();
 sg13g2_fill_2 FILLER_149_433 ();
 sg13g2_fill_8 FILLER_149_460 ();
 sg13g2_fill_8 FILLER_149_546 ();
 sg13g2_fill_1 FILLER_149_554 ();
 sg13g2_fill_8 FILLER_149_573 ();
 sg13g2_fill_8 FILLER_149_591 ();
 sg13g2_fill_4 FILLER_149_599 ();
 sg13g2_fill_2 FILLER_149_603 ();
 sg13g2_fill_8 FILLER_149_631 ();
 sg13g2_fill_4 FILLER_149_639 ();
 sg13g2_fill_2 FILLER_149_643 ();
 sg13g2_fill_1 FILLER_149_645 ();
 sg13g2_fill_8 FILLER_149_656 ();
 sg13g2_fill_8 FILLER_149_664 ();
 sg13g2_fill_8 FILLER_149_672 ();
 sg13g2_fill_8 FILLER_149_680 ();
 sg13g2_fill_1 FILLER_149_714 ();
 sg13g2_fill_8 FILLER_149_725 ();
 sg13g2_fill_4 FILLER_149_733 ();
 sg13g2_fill_1 FILLER_149_737 ();
 sg13g2_fill_1 FILLER_149_760 ();
 sg13g2_fill_8 FILLER_149_765 ();
 sg13g2_fill_8 FILLER_149_773 ();
 sg13g2_fill_2 FILLER_149_781 ();
 sg13g2_fill_8 FILLER_149_802 ();
 sg13g2_fill_4 FILLER_149_810 ();
 sg13g2_fill_2 FILLER_149_814 ();
 sg13g2_fill_8 FILLER_149_826 ();
 sg13g2_fill_4 FILLER_149_834 ();
 sg13g2_fill_1 FILLER_149_838 ();
 sg13g2_fill_1 FILLER_149_849 ();
 sg13g2_fill_2 FILLER_149_880 ();
 sg13g2_fill_1 FILLER_149_882 ();
 sg13g2_fill_8 FILLER_149_903 ();
 sg13g2_fill_8 FILLER_149_911 ();
 sg13g2_fill_2 FILLER_149_919 ();
 sg13g2_fill_8 FILLER_149_971 ();
 sg13g2_fill_8 FILLER_149_979 ();
 sg13g2_fill_4 FILLER_149_987 ();
 sg13g2_fill_2 FILLER_149_991 ();
 sg13g2_fill_1 FILLER_149_993 ();
 sg13g2_fill_8 FILLER_149_1009 ();
 sg13g2_fill_8 FILLER_149_1017 ();
 sg13g2_fill_2 FILLER_149_1038 ();
 sg13g2_fill_1 FILLER_149_1040 ();
 sg13g2_fill_2 FILLER_149_1057 ();
 sg13g2_fill_1 FILLER_149_1059 ();
 sg13g2_fill_1 FILLER_149_1081 ();
 sg13g2_fill_8 FILLER_149_1101 ();
 sg13g2_fill_8 FILLER_149_1109 ();
 sg13g2_fill_4 FILLER_149_1117 ();
 sg13g2_fill_2 FILLER_149_1121 ();
 sg13g2_fill_2 FILLER_149_1135 ();
 sg13g2_fill_4 FILLER_149_1152 ();
 sg13g2_fill_1 FILLER_149_1156 ();
 sg13g2_fill_2 FILLER_149_1166 ();
 sg13g2_fill_4 FILLER_149_1184 ();
 sg13g2_fill_2 FILLER_149_1188 ();
 sg13g2_fill_1 FILLER_149_1224 ();
 sg13g2_fill_1 FILLER_149_1237 ();
 sg13g2_fill_8 FILLER_149_1298 ();
 sg13g2_fill_2 FILLER_149_1306 ();
 sg13g2_fill_1 FILLER_149_1308 ();
 sg13g2_fill_4 FILLER_149_1368 ();
 sg13g2_fill_2 FILLER_149_1372 ();
 sg13g2_fill_1 FILLER_149_1374 ();
 sg13g2_fill_2 FILLER_149_1384 ();
 sg13g2_fill_1 FILLER_149_1386 ();
 sg13g2_fill_1 FILLER_149_1390 ();
 sg13g2_fill_1 FILLER_149_1395 ();
 sg13g2_fill_2 FILLER_149_1405 ();
 sg13g2_fill_1 FILLER_149_1407 ();
 sg13g2_fill_2 FILLER_149_1439 ();
 sg13g2_fill_1 FILLER_149_1441 ();
 sg13g2_fill_4 FILLER_149_1468 ();
 sg13g2_fill_2 FILLER_149_1472 ();
 sg13g2_fill_4 FILLER_149_1503 ();
 sg13g2_fill_2 FILLER_149_1507 ();
 sg13g2_fill_1 FILLER_149_1509 ();
 sg13g2_fill_4 FILLER_149_1518 ();
 sg13g2_fill_1 FILLER_149_1551 ();
 sg13g2_fill_1 FILLER_149_1556 ();
 sg13g2_fill_8 FILLER_149_1567 ();
 sg13g2_fill_8 FILLER_149_1575 ();
 sg13g2_fill_8 FILLER_149_1583 ();
 sg13g2_fill_1 FILLER_149_1591 ();
 sg13g2_fill_8 FILLER_150_0 ();
 sg13g2_fill_8 FILLER_150_8 ();
 sg13g2_fill_8 FILLER_150_16 ();
 sg13g2_fill_8 FILLER_150_24 ();
 sg13g2_fill_2 FILLER_150_32 ();
 sg13g2_fill_1 FILLER_150_34 ();
 sg13g2_fill_8 FILLER_150_91 ();
 sg13g2_fill_4 FILLER_150_99 ();
 sg13g2_fill_2 FILLER_150_103 ();
 sg13g2_fill_1 FILLER_150_131 ();
 sg13g2_fill_2 FILLER_150_176 ();
 sg13g2_fill_8 FILLER_150_199 ();
 sg13g2_fill_2 FILLER_150_207 ();
 sg13g2_fill_1 FILLER_150_209 ();
 sg13g2_fill_2 FILLER_150_236 ();
 sg13g2_fill_4 FILLER_150_246 ();
 sg13g2_fill_1 FILLER_150_250 ();
 sg13g2_fill_4 FILLER_150_298 ();
 sg13g2_fill_2 FILLER_150_302 ();
 sg13g2_fill_4 FILLER_150_330 ();
 sg13g2_fill_1 FILLER_150_334 ();
 sg13g2_fill_2 FILLER_150_361 ();
 sg13g2_fill_2 FILLER_150_381 ();
 sg13g2_fill_8 FILLER_150_419 ();
 sg13g2_fill_8 FILLER_150_427 ();
 sg13g2_fill_1 FILLER_150_435 ();
 sg13g2_fill_4 FILLER_150_451 ();
 sg13g2_fill_2 FILLER_150_455 ();
 sg13g2_fill_1 FILLER_150_457 ();
 sg13g2_fill_2 FILLER_150_468 ();
 sg13g2_fill_1 FILLER_150_480 ();
 sg13g2_fill_8 FILLER_150_505 ();
 sg13g2_fill_8 FILLER_150_513 ();
 sg13g2_fill_8 FILLER_150_521 ();
 sg13g2_fill_8 FILLER_150_529 ();
 sg13g2_fill_8 FILLER_150_537 ();
 sg13g2_fill_8 FILLER_150_545 ();
 sg13g2_fill_8 FILLER_150_558 ();
 sg13g2_fill_8 FILLER_150_566 ();
 sg13g2_fill_2 FILLER_150_574 ();
 sg13g2_fill_1 FILLER_150_602 ();
 sg13g2_fill_8 FILLER_150_613 ();
 sg13g2_fill_4 FILLER_150_621 ();
 sg13g2_fill_4 FILLER_150_635 ();
 sg13g2_fill_2 FILLER_150_639 ();
 sg13g2_fill_1 FILLER_150_641 ();
 sg13g2_fill_4 FILLER_150_678 ();
 sg13g2_fill_2 FILLER_150_682 ();
 sg13g2_fill_4 FILLER_150_719 ();
 sg13g2_fill_1 FILLER_150_749 ();
 sg13g2_fill_8 FILLER_150_754 ();
 sg13g2_fill_8 FILLER_150_775 ();
 sg13g2_fill_1 FILLER_150_783 ();
 sg13g2_fill_8 FILLER_150_826 ();
 sg13g2_fill_8 FILLER_150_834 ();
 sg13g2_fill_2 FILLER_150_842 ();
 sg13g2_fill_1 FILLER_150_844 ();
 sg13g2_fill_8 FILLER_150_849 ();
 sg13g2_fill_4 FILLER_150_875 ();
 sg13g2_fill_2 FILLER_150_879 ();
 sg13g2_fill_2 FILLER_150_902 ();
 sg13g2_fill_2 FILLER_150_929 ();
 sg13g2_fill_1 FILLER_150_934 ();
 sg13g2_fill_8 FILLER_150_938 ();
 sg13g2_fill_8 FILLER_150_946 ();
 sg13g2_fill_2 FILLER_150_954 ();
 sg13g2_fill_1 FILLER_150_956 ();
 sg13g2_fill_4 FILLER_150_963 ();
 sg13g2_fill_2 FILLER_150_967 ();
 sg13g2_fill_1 FILLER_150_969 ();
 sg13g2_fill_8 FILLER_150_974 ();
 sg13g2_fill_4 FILLER_150_982 ();
 sg13g2_fill_1 FILLER_150_986 ();
 sg13g2_fill_2 FILLER_150_1002 ();
 sg13g2_fill_8 FILLER_150_1010 ();
 sg13g2_fill_4 FILLER_150_1018 ();
 sg13g2_fill_4 FILLER_150_1039 ();
 sg13g2_fill_2 FILLER_150_1043 ();
 sg13g2_fill_8 FILLER_150_1050 ();
 sg13g2_fill_4 FILLER_150_1058 ();
 sg13g2_fill_2 FILLER_150_1062 ();
 sg13g2_fill_1 FILLER_150_1064 ();
 sg13g2_fill_8 FILLER_150_1075 ();
 sg13g2_fill_8 FILLER_150_1083 ();
 sg13g2_fill_2 FILLER_150_1091 ();
 sg13g2_fill_1 FILLER_150_1093 ();
 sg13g2_fill_1 FILLER_150_1110 ();
 sg13g2_fill_8 FILLER_150_1127 ();
 sg13g2_fill_4 FILLER_150_1135 ();
 sg13g2_fill_2 FILLER_150_1139 ();
 sg13g2_fill_1 FILLER_150_1141 ();
 sg13g2_fill_8 FILLER_150_1145 ();
 sg13g2_fill_8 FILLER_150_1153 ();
 sg13g2_fill_8 FILLER_150_1161 ();
 sg13g2_fill_8 FILLER_150_1169 ();
 sg13g2_fill_4 FILLER_150_1177 ();
 sg13g2_fill_8 FILLER_150_1191 ();
 sg13g2_fill_2 FILLER_150_1205 ();
 sg13g2_fill_1 FILLER_150_1207 ();
 sg13g2_fill_4 FILLER_150_1213 ();
 sg13g2_fill_2 FILLER_150_1217 ();
 sg13g2_fill_8 FILLER_150_1233 ();
 sg13g2_fill_8 FILLER_150_1241 ();
 sg13g2_fill_8 FILLER_150_1249 ();
 sg13g2_fill_8 FILLER_150_1257 ();
 sg13g2_fill_8 FILLER_150_1265 ();
 sg13g2_fill_4 FILLER_150_1273 ();
 sg13g2_fill_2 FILLER_150_1277 ();
 sg13g2_fill_2 FILLER_150_1309 ();
 sg13g2_fill_1 FILLER_150_1311 ();
 sg13g2_fill_4 FILLER_150_1340 ();
 sg13g2_fill_2 FILLER_150_1344 ();
 sg13g2_fill_2 FILLER_150_1352 ();
 sg13g2_fill_1 FILLER_150_1354 ();
 sg13g2_fill_8 FILLER_150_1363 ();
 sg13g2_fill_8 FILLER_150_1371 ();
 sg13g2_fill_2 FILLER_150_1379 ();
 sg13g2_fill_8 FILLER_150_1389 ();
 sg13g2_fill_8 FILLER_150_1397 ();
 sg13g2_fill_8 FILLER_150_1405 ();
 sg13g2_fill_2 FILLER_150_1413 ();
 sg13g2_fill_1 FILLER_150_1415 ();
 sg13g2_fill_2 FILLER_150_1423 ();
 sg13g2_fill_1 FILLER_150_1425 ();
 sg13g2_fill_2 FILLER_150_1437 ();
 sg13g2_fill_1 FILLER_150_1439 ();
 sg13g2_fill_2 FILLER_150_1448 ();
 sg13g2_fill_1 FILLER_150_1450 ();
 sg13g2_fill_8 FILLER_150_1481 ();
 sg13g2_fill_8 FILLER_150_1489 ();
 sg13g2_fill_4 FILLER_150_1497 ();
 sg13g2_fill_2 FILLER_150_1501 ();
 sg13g2_fill_1 FILLER_150_1503 ();
 sg13g2_fill_8 FILLER_150_1508 ();
 sg13g2_fill_8 FILLER_150_1516 ();
 sg13g2_fill_4 FILLER_150_1524 ();
 sg13g2_fill_8 FILLER_150_1531 ();
 sg13g2_fill_4 FILLER_150_1539 ();
 sg13g2_fill_1 FILLER_150_1543 ();
 sg13g2_fill_2 FILLER_150_1552 ();
 sg13g2_fill_8 FILLER_150_1564 ();
 sg13g2_fill_8 FILLER_150_1572 ();
 sg13g2_fill_8 FILLER_150_1580 ();
 sg13g2_fill_4 FILLER_150_1588 ();
 sg13g2_fill_8 FILLER_151_0 ();
 sg13g2_fill_8 FILLER_151_8 ();
 sg13g2_fill_8 FILLER_151_16 ();
 sg13g2_fill_8 FILLER_151_24 ();
 sg13g2_fill_8 FILLER_151_32 ();
 sg13g2_fill_8 FILLER_151_40 ();
 sg13g2_fill_4 FILLER_151_48 ();
 sg13g2_fill_2 FILLER_151_52 ();
 sg13g2_fill_1 FILLER_151_54 ();
 sg13g2_fill_8 FILLER_151_65 ();
 sg13g2_fill_8 FILLER_151_73 ();
 sg13g2_fill_8 FILLER_151_81 ();
 sg13g2_fill_8 FILLER_151_89 ();
 sg13g2_fill_4 FILLER_151_97 ();
 sg13g2_fill_1 FILLER_151_101 ();
 sg13g2_fill_8 FILLER_151_110 ();
 sg13g2_fill_4 FILLER_151_118 ();
 sg13g2_fill_2 FILLER_151_122 ();
 sg13g2_fill_8 FILLER_151_134 ();
 sg13g2_fill_2 FILLER_151_142 ();
 sg13g2_fill_8 FILLER_151_152 ();
 sg13g2_fill_8 FILLER_151_160 ();
 sg13g2_fill_8 FILLER_151_168 ();
 sg13g2_fill_1 FILLER_151_176 ();
 sg13g2_fill_4 FILLER_151_245 ();
 sg13g2_fill_8 FILLER_151_269 ();
 sg13g2_fill_8 FILLER_151_277 ();
 sg13g2_fill_8 FILLER_151_285 ();
 sg13g2_fill_4 FILLER_151_293 ();
 sg13g2_fill_1 FILLER_151_297 ();
 sg13g2_fill_8 FILLER_151_306 ();
 sg13g2_fill_8 FILLER_151_314 ();
 sg13g2_fill_1 FILLER_151_322 ();
 sg13g2_fill_8 FILLER_151_333 ();
 sg13g2_fill_8 FILLER_151_341 ();
 sg13g2_fill_1 FILLER_151_349 ();
 sg13g2_fill_1 FILLER_151_358 ();
 sg13g2_fill_8 FILLER_151_389 ();
 sg13g2_fill_8 FILLER_151_397 ();
 sg13g2_fill_8 FILLER_151_405 ();
 sg13g2_fill_2 FILLER_151_413 ();
 sg13g2_fill_1 FILLER_151_415 ();
 sg13g2_fill_8 FILLER_151_426 ();
 sg13g2_fill_2 FILLER_151_434 ();
 sg13g2_fill_1 FILLER_151_472 ();
 sg13g2_fill_8 FILLER_151_479 ();
 sg13g2_fill_2 FILLER_151_487 ();
 sg13g2_fill_1 FILLER_151_489 ();
 sg13g2_fill_1 FILLER_151_496 ();
 sg13g2_fill_8 FILLER_151_503 ();
 sg13g2_fill_1 FILLER_151_511 ();
 sg13g2_fill_4 FILLER_151_517 ();
 sg13g2_fill_2 FILLER_151_521 ();
 sg13g2_fill_2 FILLER_151_533 ();
 sg13g2_fill_1 FILLER_151_535 ();
 sg13g2_fill_4 FILLER_151_546 ();
 sg13g2_fill_8 FILLER_151_576 ();
 sg13g2_fill_8 FILLER_151_584 ();
 sg13g2_fill_2 FILLER_151_592 ();
 sg13g2_fill_1 FILLER_151_594 ();
 sg13g2_fill_4 FILLER_151_620 ();
 sg13g2_fill_2 FILLER_151_624 ();
 sg13g2_fill_1 FILLER_151_626 ();
 sg13g2_fill_4 FILLER_151_637 ();
 sg13g2_fill_8 FILLER_151_651 ();
 sg13g2_fill_8 FILLER_151_659 ();
 sg13g2_fill_4 FILLER_151_667 ();
 sg13g2_fill_2 FILLER_151_671 ();
 sg13g2_fill_1 FILLER_151_673 ();
 sg13g2_fill_4 FILLER_151_682 ();
 sg13g2_fill_2 FILLER_151_686 ();
 sg13g2_fill_1 FILLER_151_688 ();
 sg13g2_fill_1 FILLER_151_704 ();
 sg13g2_fill_8 FILLER_151_723 ();
 sg13g2_fill_8 FILLER_151_731 ();
 sg13g2_fill_4 FILLER_151_739 ();
 sg13g2_fill_2 FILLER_151_743 ();
 sg13g2_fill_4 FILLER_151_758 ();
 sg13g2_fill_1 FILLER_151_762 ();
 sg13g2_fill_2 FILLER_151_771 ();
 sg13g2_fill_1 FILLER_151_773 ();
 sg13g2_fill_8 FILLER_151_779 ();
 sg13g2_fill_4 FILLER_151_787 ();
 sg13g2_fill_1 FILLER_151_791 ();
 sg13g2_fill_2 FILLER_151_802 ();
 sg13g2_fill_1 FILLER_151_804 ();
 sg13g2_fill_8 FILLER_151_810 ();
 sg13g2_fill_1 FILLER_151_824 ();
 sg13g2_fill_4 FILLER_151_829 ();
 sg13g2_fill_2 FILLER_151_833 ();
 sg13g2_fill_1 FILLER_151_835 ();
 sg13g2_fill_1 FILLER_151_851 ();
 sg13g2_fill_8 FILLER_151_857 ();
 sg13g2_fill_8 FILLER_151_865 ();
 sg13g2_fill_8 FILLER_151_873 ();
 sg13g2_fill_8 FILLER_151_881 ();
 sg13g2_fill_8 FILLER_151_889 ();
 sg13g2_fill_8 FILLER_151_897 ();
 sg13g2_fill_1 FILLER_151_905 ();
 sg13g2_fill_1 FILLER_151_934 ();
 sg13g2_fill_1 FILLER_151_946 ();
 sg13g2_fill_8 FILLER_151_1000 ();
 sg13g2_fill_8 FILLER_151_1021 ();
 sg13g2_fill_4 FILLER_151_1033 ();
 sg13g2_fill_4 FILLER_151_1042 ();
 sg13g2_fill_2 FILLER_151_1046 ();
 sg13g2_fill_2 FILLER_151_1060 ();
 sg13g2_fill_1 FILLER_151_1062 ();
 sg13g2_fill_4 FILLER_151_1070 ();
 sg13g2_fill_2 FILLER_151_1074 ();
 sg13g2_fill_2 FILLER_151_1080 ();
 sg13g2_fill_4 FILLER_151_1086 ();
 sg13g2_fill_2 FILLER_151_1105 ();
 sg13g2_fill_1 FILLER_151_1107 ();
 sg13g2_fill_4 FILLER_151_1119 ();
 sg13g2_fill_1 FILLER_151_1133 ();
 sg13g2_fill_8 FILLER_151_1151 ();
 sg13g2_fill_1 FILLER_151_1159 ();
 sg13g2_fill_1 FILLER_151_1169 ();
 sg13g2_fill_1 FILLER_151_1176 ();
 sg13g2_fill_8 FILLER_151_1182 ();
 sg13g2_fill_2 FILLER_151_1190 ();
 sg13g2_fill_4 FILLER_151_1242 ();
 sg13g2_fill_2 FILLER_151_1254 ();
 sg13g2_fill_8 FILLER_151_1274 ();
 sg13g2_fill_8 FILLER_151_1282 ();
 sg13g2_fill_2 FILLER_151_1290 ();
 sg13g2_fill_1 FILLER_151_1292 ();
 sg13g2_fill_8 FILLER_151_1299 ();
 sg13g2_fill_2 FILLER_151_1307 ();
 sg13g2_fill_1 FILLER_151_1309 ();
 sg13g2_fill_8 FILLER_151_1326 ();
 sg13g2_fill_8 FILLER_151_1334 ();
 sg13g2_fill_4 FILLER_151_1342 ();
 sg13g2_fill_1 FILLER_151_1352 ();
 sg13g2_fill_2 FILLER_151_1364 ();
 sg13g2_fill_1 FILLER_151_1366 ();
 sg13g2_fill_4 FILLER_151_1378 ();
 sg13g2_fill_1 FILLER_151_1382 ();
 sg13g2_fill_8 FILLER_151_1399 ();
 sg13g2_fill_8 FILLER_151_1407 ();
 sg13g2_fill_8 FILLER_151_1415 ();
 sg13g2_fill_8 FILLER_151_1423 ();
 sg13g2_fill_4 FILLER_151_1431 ();
 sg13g2_fill_2 FILLER_151_1435 ();
 sg13g2_fill_1 FILLER_151_1437 ();
 sg13g2_fill_4 FILLER_151_1443 ();
 sg13g2_fill_4 FILLER_151_1457 ();
 sg13g2_fill_2 FILLER_151_1461 ();
 sg13g2_fill_1 FILLER_151_1463 ();
 sg13g2_fill_2 FILLER_151_1490 ();
 sg13g2_fill_1 FILLER_151_1492 ();
 sg13g2_fill_8 FILLER_151_1519 ();
 sg13g2_fill_4 FILLER_151_1535 ();
 sg13g2_fill_1 FILLER_151_1539 ();
 sg13g2_fill_8 FILLER_151_1545 ();
 sg13g2_fill_2 FILLER_151_1553 ();
 sg13g2_fill_1 FILLER_151_1563 ();
 sg13g2_fill_2 FILLER_151_1590 ();
 sg13g2_fill_8 FILLER_152_0 ();
 sg13g2_fill_8 FILLER_152_8 ();
 sg13g2_fill_8 FILLER_152_16 ();
 sg13g2_fill_8 FILLER_152_24 ();
 sg13g2_fill_8 FILLER_152_32 ();
 sg13g2_fill_8 FILLER_152_40 ();
 sg13g2_fill_8 FILLER_152_48 ();
 sg13g2_fill_4 FILLER_152_56 ();
 sg13g2_fill_1 FILLER_152_60 ();
 sg13g2_fill_4 FILLER_152_64 ();
 sg13g2_fill_1 FILLER_152_68 ();
 sg13g2_fill_4 FILLER_152_105 ();
 sg13g2_fill_1 FILLER_152_109 ();
 sg13g2_fill_4 FILLER_152_120 ();
 sg13g2_fill_2 FILLER_152_124 ();
 sg13g2_fill_1 FILLER_152_126 ();
 sg13g2_fill_8 FILLER_152_142 ();
 sg13g2_fill_2 FILLER_152_150 ();
 sg13g2_fill_1 FILLER_152_152 ();
 sg13g2_fill_8 FILLER_152_161 ();
 sg13g2_fill_8 FILLER_152_169 ();
 sg13g2_fill_8 FILLER_152_177 ();
 sg13g2_fill_4 FILLER_152_218 ();
 sg13g2_fill_4 FILLER_152_243 ();
 sg13g2_fill_2 FILLER_152_247 ();
 sg13g2_fill_1 FILLER_152_249 ();
 sg13g2_fill_4 FILLER_152_285 ();
 sg13g2_fill_2 FILLER_152_289 ();
 sg13g2_fill_1 FILLER_152_299 ();
 sg13g2_fill_4 FILLER_152_310 ();
 sg13g2_fill_2 FILLER_152_413 ();
 sg13g2_fill_1 FILLER_152_415 ();
 sg13g2_fill_8 FILLER_152_449 ();
 sg13g2_fill_8 FILLER_152_457 ();
 sg13g2_fill_2 FILLER_152_465 ();
 sg13g2_fill_8 FILLER_152_477 ();
 sg13g2_fill_1 FILLER_152_485 ();
 sg13g2_fill_1 FILLER_152_496 ();
 sg13g2_fill_8 FILLER_152_523 ();
 sg13g2_fill_1 FILLER_152_531 ();
 sg13g2_fill_1 FILLER_152_547 ();
 sg13g2_fill_2 FILLER_152_574 ();
 sg13g2_fill_1 FILLER_152_576 ();
 sg13g2_fill_8 FILLER_152_639 ();
 sg13g2_fill_8 FILLER_152_647 ();
 sg13g2_fill_8 FILLER_152_655 ();
 sg13g2_fill_1 FILLER_152_663 ();
 sg13g2_fill_4 FILLER_152_674 ();
 sg13g2_fill_8 FILLER_152_719 ();
 sg13g2_fill_4 FILLER_152_727 ();
 sg13g2_fill_4 FILLER_152_737 ();
 sg13g2_fill_8 FILLER_152_751 ();
 sg13g2_fill_4 FILLER_152_759 ();
 sg13g2_fill_2 FILLER_152_763 ();
 sg13g2_fill_1 FILLER_152_765 ();
 sg13g2_fill_8 FILLER_152_771 ();
 sg13g2_fill_4 FILLER_152_779 ();
 sg13g2_fill_1 FILLER_152_783 ();
 sg13g2_fill_4 FILLER_152_789 ();
 sg13g2_fill_2 FILLER_152_793 ();
 sg13g2_fill_1 FILLER_152_795 ();
 sg13g2_fill_2 FILLER_152_816 ();
 sg13g2_fill_1 FILLER_152_832 ();
 sg13g2_fill_2 FILLER_152_854 ();
 sg13g2_fill_2 FILLER_152_870 ();
 sg13g2_fill_4 FILLER_152_877 ();
 sg13g2_fill_2 FILLER_152_886 ();
 sg13g2_fill_4 FILLER_152_897 ();
 sg13g2_fill_2 FILLER_152_901 ();
 sg13g2_fill_1 FILLER_152_903 ();
 sg13g2_fill_8 FILLER_152_909 ();
 sg13g2_fill_8 FILLER_152_917 ();
 sg13g2_fill_4 FILLER_152_925 ();
 sg13g2_fill_2 FILLER_152_929 ();
 sg13g2_fill_1 FILLER_152_952 ();
 sg13g2_fill_2 FILLER_152_969 ();
 sg13g2_fill_2 FILLER_152_997 ();
 sg13g2_fill_4 FILLER_152_1028 ();
 sg13g2_fill_4 FILLER_152_1060 ();
 sg13g2_fill_2 FILLER_152_1064 ();
 sg13g2_fill_1 FILLER_152_1070 ();
 sg13g2_fill_8 FILLER_152_1075 ();
 sg13g2_fill_2 FILLER_152_1083 ();
 sg13g2_fill_4 FILLER_152_1089 ();
 sg13g2_fill_4 FILLER_152_1101 ();
 sg13g2_fill_4 FILLER_152_1114 ();
 sg13g2_fill_1 FILLER_152_1118 ();
 sg13g2_fill_4 FILLER_152_1127 ();
 sg13g2_fill_1 FILLER_152_1131 ();
 sg13g2_fill_1 FILLER_152_1145 ();
 sg13g2_fill_1 FILLER_152_1158 ();
 sg13g2_fill_4 FILLER_152_1209 ();
 sg13g2_fill_2 FILLER_152_1213 ();
 sg13g2_fill_1 FILLER_152_1223 ();
 sg13g2_fill_4 FILLER_152_1234 ();
 sg13g2_fill_2 FILLER_152_1238 ();
 sg13g2_fill_8 FILLER_152_1261 ();
 sg13g2_fill_1 FILLER_152_1269 ();
 sg13g2_fill_8 FILLER_152_1276 ();
 sg13g2_fill_4 FILLER_152_1284 ();
 sg13g2_fill_4 FILLER_152_1292 ();
 sg13g2_fill_1 FILLER_152_1296 ();
 sg13g2_fill_1 FILLER_152_1362 ();
 sg13g2_fill_8 FILLER_152_1385 ();
 sg13g2_fill_2 FILLER_152_1393 ();
 sg13g2_fill_8 FILLER_152_1412 ();
 sg13g2_fill_1 FILLER_152_1420 ();
 sg13g2_fill_8 FILLER_152_1429 ();
 sg13g2_fill_8 FILLER_152_1445 ();
 sg13g2_fill_8 FILLER_152_1453 ();
 sg13g2_fill_2 FILLER_152_1461 ();
 sg13g2_fill_2 FILLER_152_1489 ();
 sg13g2_fill_4 FILLER_152_1512 ();
 sg13g2_fill_2 FILLER_152_1516 ();
 sg13g2_fill_1 FILLER_152_1518 ();
 sg13g2_fill_8 FILLER_152_1530 ();
 sg13g2_fill_4 FILLER_152_1538 ();
 sg13g2_fill_1 FILLER_152_1542 ();
 sg13g2_fill_1 FILLER_152_1555 ();
 sg13g2_fill_8 FILLER_153_0 ();
 sg13g2_fill_8 FILLER_153_8 ();
 sg13g2_fill_8 FILLER_153_16 ();
 sg13g2_fill_8 FILLER_153_24 ();
 sg13g2_fill_8 FILLER_153_32 ();
 sg13g2_fill_8 FILLER_153_40 ();
 sg13g2_fill_4 FILLER_153_48 ();
 sg13g2_fill_2 FILLER_153_52 ();
 sg13g2_fill_1 FILLER_153_54 ();
 sg13g2_fill_4 FILLER_153_81 ();
 sg13g2_fill_2 FILLER_153_85 ();
 sg13g2_fill_2 FILLER_153_123 ();
 sg13g2_fill_1 FILLER_153_125 ();
 sg13g2_fill_1 FILLER_153_147 ();
 sg13g2_fill_8 FILLER_153_202 ();
 sg13g2_fill_8 FILLER_153_210 ();
 sg13g2_fill_8 FILLER_153_218 ();
 sg13g2_fill_8 FILLER_153_226 ();
 sg13g2_fill_4 FILLER_153_234 ();
 sg13g2_fill_2 FILLER_153_238 ();
 sg13g2_fill_4 FILLER_153_326 ();
 sg13g2_fill_2 FILLER_153_330 ();
 sg13g2_fill_1 FILLER_153_332 ();
 sg13g2_fill_8 FILLER_153_354 ();
 sg13g2_fill_2 FILLER_153_362 ();
 sg13g2_fill_1 FILLER_153_364 ();
 sg13g2_fill_8 FILLER_153_370 ();
 sg13g2_fill_8 FILLER_153_378 ();
 sg13g2_fill_8 FILLER_153_386 ();
 sg13g2_fill_8 FILLER_153_394 ();
 sg13g2_fill_1 FILLER_153_402 ();
 sg13g2_fill_8 FILLER_153_413 ();
 sg13g2_fill_2 FILLER_153_421 ();
 sg13g2_fill_8 FILLER_153_431 ();
 sg13g2_fill_4 FILLER_153_439 ();
 sg13g2_fill_2 FILLER_153_479 ();
 sg13g2_fill_1 FILLER_153_481 ();
 sg13g2_fill_8 FILLER_153_502 ();
 sg13g2_fill_2 FILLER_153_510 ();
 sg13g2_fill_1 FILLER_153_512 ();
 sg13g2_fill_4 FILLER_153_549 ();
 sg13g2_fill_1 FILLER_153_553 ();
 sg13g2_fill_8 FILLER_153_579 ();
 sg13g2_fill_1 FILLER_153_587 ();
 sg13g2_fill_8 FILLER_153_592 ();
 sg13g2_fill_8 FILLER_153_600 ();
 sg13g2_fill_8 FILLER_153_608 ();
 sg13g2_fill_8 FILLER_153_616 ();
 sg13g2_fill_4 FILLER_153_624 ();
 sg13g2_fill_1 FILLER_153_628 ();
 sg13g2_fill_8 FILLER_153_691 ();
 sg13g2_fill_8 FILLER_153_699 ();
 sg13g2_fill_8 FILLER_153_707 ();
 sg13g2_fill_8 FILLER_153_715 ();
 sg13g2_fill_2 FILLER_153_723 ();
 sg13g2_fill_1 FILLER_153_725 ();
 sg13g2_fill_2 FILLER_153_752 ();
 sg13g2_fill_1 FILLER_153_754 ();
 sg13g2_fill_2 FILLER_153_783 ();
 sg13g2_fill_1 FILLER_153_785 ();
 sg13g2_fill_1 FILLER_153_795 ();
 sg13g2_fill_8 FILLER_153_802 ();
 sg13g2_fill_4 FILLER_153_810 ();
 sg13g2_fill_2 FILLER_153_820 ();
 sg13g2_fill_2 FILLER_153_832 ();
 sg13g2_fill_1 FILLER_153_834 ();
 sg13g2_fill_8 FILLER_153_841 ();
 sg13g2_fill_2 FILLER_153_849 ();
 sg13g2_fill_4 FILLER_153_869 ();
 sg13g2_fill_2 FILLER_153_873 ();
 sg13g2_fill_1 FILLER_153_875 ();
 sg13g2_fill_2 FILLER_153_896 ();
 sg13g2_fill_8 FILLER_153_922 ();
 sg13g2_fill_2 FILLER_153_969 ();
 sg13g2_fill_2 FILLER_153_1007 ();
 sg13g2_fill_4 FILLER_153_1027 ();
 sg13g2_fill_1 FILLER_153_1031 ();
 sg13g2_fill_1 FILLER_153_1048 ();
 sg13g2_fill_2 FILLER_153_1057 ();
 sg13g2_fill_1 FILLER_153_1059 ();
 sg13g2_fill_1 FILLER_153_1079 ();
 sg13g2_fill_1 FILLER_153_1088 ();
 sg13g2_fill_1 FILLER_153_1099 ();
 sg13g2_fill_8 FILLER_153_1106 ();
 sg13g2_fill_8 FILLER_153_1114 ();
 sg13g2_fill_2 FILLER_153_1122 ();
 sg13g2_fill_1 FILLER_153_1128 ();
 sg13g2_fill_8 FILLER_153_1134 ();
 sg13g2_fill_8 FILLER_153_1142 ();
 sg13g2_fill_2 FILLER_153_1150 ();
 sg13g2_fill_1 FILLER_153_1152 ();
 sg13g2_fill_8 FILLER_153_1165 ();
 sg13g2_fill_8 FILLER_153_1173 ();
 sg13g2_fill_8 FILLER_153_1181 ();
 sg13g2_fill_1 FILLER_153_1189 ();
 sg13g2_fill_8 FILLER_153_1195 ();
 sg13g2_fill_8 FILLER_153_1203 ();
 sg13g2_fill_1 FILLER_153_1211 ();
 sg13g2_fill_8 FILLER_153_1215 ();
 sg13g2_fill_8 FILLER_153_1223 ();
 sg13g2_fill_8 FILLER_153_1231 ();
 sg13g2_fill_8 FILLER_153_1239 ();
 sg13g2_fill_2 FILLER_153_1247 ();
 sg13g2_fill_1 FILLER_153_1249 ();
 sg13g2_fill_1 FILLER_153_1261 ();
 sg13g2_fill_2 FILLER_153_1270 ();
 sg13g2_fill_8 FILLER_153_1279 ();
 sg13g2_fill_4 FILLER_153_1287 ();
 sg13g2_fill_1 FILLER_153_1295 ();
 sg13g2_fill_8 FILLER_153_1300 ();
 sg13g2_fill_8 FILLER_153_1308 ();
 sg13g2_fill_4 FILLER_153_1316 ();
 sg13g2_fill_2 FILLER_153_1320 ();
 sg13g2_fill_8 FILLER_153_1332 ();
 sg13g2_fill_2 FILLER_153_1340 ();
 sg13g2_fill_1 FILLER_153_1342 ();
 sg13g2_fill_4 FILLER_153_1348 ();
 sg13g2_fill_2 FILLER_153_1352 ();
 sg13g2_fill_1 FILLER_153_1354 ();
 sg13g2_fill_1 FILLER_153_1366 ();
 sg13g2_fill_4 FILLER_153_1373 ();
 sg13g2_fill_1 FILLER_153_1377 ();
 sg13g2_fill_2 FILLER_153_1386 ();
 sg13g2_fill_2 FILLER_153_1411 ();
 sg13g2_fill_1 FILLER_153_1429 ();
 sg13g2_fill_4 FILLER_153_1435 ();
 sg13g2_fill_1 FILLER_153_1439 ();
 sg13g2_fill_8 FILLER_153_1455 ();
 sg13g2_fill_8 FILLER_153_1463 ();
 sg13g2_fill_8 FILLER_153_1471 ();
 sg13g2_fill_8 FILLER_153_1479 ();
 sg13g2_fill_8 FILLER_153_1487 ();
 sg13g2_fill_8 FILLER_153_1495 ();
 sg13g2_fill_8 FILLER_153_1503 ();
 sg13g2_fill_4 FILLER_153_1511 ();
 sg13g2_fill_1 FILLER_153_1515 ();
 sg13g2_fill_4 FILLER_153_1550 ();
 sg13g2_fill_1 FILLER_153_1554 ();
 sg13g2_fill_2 FILLER_153_1569 ();
 sg13g2_fill_1 FILLER_153_1571 ();
 sg13g2_fill_8 FILLER_153_1580 ();
 sg13g2_fill_4 FILLER_153_1588 ();
 sg13g2_fill_8 FILLER_154_0 ();
 sg13g2_fill_8 FILLER_154_8 ();
 sg13g2_fill_8 FILLER_154_16 ();
 sg13g2_fill_8 FILLER_154_24 ();
 sg13g2_fill_4 FILLER_154_32 ();
 sg13g2_fill_8 FILLER_154_97 ();
 sg13g2_fill_8 FILLER_154_105 ();
 sg13g2_fill_8 FILLER_154_113 ();
 sg13g2_fill_8 FILLER_154_121 ();
 sg13g2_fill_2 FILLER_154_129 ();
 sg13g2_fill_8 FILLER_154_137 ();
 sg13g2_fill_8 FILLER_154_145 ();
 sg13g2_fill_4 FILLER_154_153 ();
 sg13g2_fill_2 FILLER_154_157 ();
 sg13g2_fill_8 FILLER_154_194 ();
 sg13g2_fill_8 FILLER_154_228 ();
 sg13g2_fill_4 FILLER_154_236 ();
 sg13g2_fill_1 FILLER_154_248 ();
 sg13g2_fill_8 FILLER_154_254 ();
 sg13g2_fill_8 FILLER_154_262 ();
 sg13g2_fill_8 FILLER_154_270 ();
 sg13g2_fill_8 FILLER_154_278 ();
 sg13g2_fill_8 FILLER_154_286 ();
 sg13g2_fill_8 FILLER_154_294 ();
 sg13g2_fill_2 FILLER_154_302 ();
 sg13g2_fill_1 FILLER_154_304 ();
 sg13g2_fill_8 FILLER_154_313 ();
 sg13g2_fill_8 FILLER_154_321 ();
 sg13g2_fill_8 FILLER_154_329 ();
 sg13g2_fill_8 FILLER_154_337 ();
 sg13g2_fill_8 FILLER_154_345 ();
 sg13g2_fill_8 FILLER_154_353 ();
 sg13g2_fill_2 FILLER_154_361 ();
 sg13g2_fill_4 FILLER_154_389 ();
 sg13g2_fill_2 FILLER_154_393 ();
 sg13g2_fill_1 FILLER_154_395 ();
 sg13g2_fill_2 FILLER_154_422 ();
 sg13g2_fill_8 FILLER_154_460 ();
 sg13g2_fill_8 FILLER_154_494 ();
 sg13g2_fill_8 FILLER_154_502 ();
 sg13g2_fill_8 FILLER_154_510 ();
 sg13g2_fill_1 FILLER_154_518 ();
 sg13g2_fill_8 FILLER_154_529 ();
 sg13g2_fill_2 FILLER_154_537 ();
 sg13g2_fill_4 FILLER_154_549 ();
 sg13g2_fill_8 FILLER_154_579 ();
 sg13g2_fill_8 FILLER_154_587 ();
 sg13g2_fill_8 FILLER_154_595 ();
 sg13g2_fill_2 FILLER_154_603 ();
 sg13g2_fill_1 FILLER_154_605 ();
 sg13g2_fill_4 FILLER_154_632 ();
 sg13g2_fill_1 FILLER_154_636 ();
 sg13g2_fill_8 FILLER_154_668 ();
 sg13g2_fill_2 FILLER_154_676 ();
 sg13g2_fill_1 FILLER_154_678 ();
 sg13g2_fill_8 FILLER_154_687 ();
 sg13g2_fill_4 FILLER_154_741 ();
 sg13g2_fill_2 FILLER_154_745 ();
 sg13g2_fill_1 FILLER_154_747 ();
 sg13g2_fill_2 FILLER_154_758 ();
 sg13g2_fill_1 FILLER_154_760 ();
 sg13g2_fill_2 FILLER_154_765 ();
 sg13g2_fill_1 FILLER_154_767 ();
 sg13g2_fill_4 FILLER_154_773 ();
 sg13g2_fill_2 FILLER_154_782 ();
 sg13g2_fill_1 FILLER_154_808 ();
 sg13g2_fill_8 FILLER_154_814 ();
 sg13g2_fill_1 FILLER_154_822 ();
 sg13g2_fill_8 FILLER_154_828 ();
 sg13g2_fill_8 FILLER_154_836 ();
 sg13g2_fill_4 FILLER_154_844 ();
 sg13g2_fill_8 FILLER_154_854 ();
 sg13g2_fill_8 FILLER_154_862 ();
 sg13g2_fill_4 FILLER_154_874 ();
 sg13g2_fill_2 FILLER_154_878 ();
 sg13g2_fill_1 FILLER_154_880 ();
 sg13g2_fill_1 FILLER_154_890 ();
 sg13g2_fill_1 FILLER_154_895 ();
 sg13g2_fill_4 FILLER_154_899 ();
 sg13g2_fill_2 FILLER_154_903 ();
 sg13g2_fill_4 FILLER_154_910 ();
 sg13g2_fill_8 FILLER_154_922 ();
 sg13g2_fill_8 FILLER_154_930 ();
 sg13g2_fill_2 FILLER_154_938 ();
 sg13g2_fill_8 FILLER_154_946 ();
 sg13g2_fill_1 FILLER_154_965 ();
 sg13g2_fill_2 FILLER_154_974 ();
 sg13g2_fill_4 FILLER_154_992 ();
 sg13g2_fill_1 FILLER_154_1000 ();
 sg13g2_fill_8 FILLER_154_1009 ();
 sg13g2_fill_8 FILLER_154_1017 ();
 sg13g2_fill_8 FILLER_154_1025 ();
 sg13g2_fill_2 FILLER_154_1033 ();
 sg13g2_fill_4 FILLER_154_1040 ();
 sg13g2_fill_2 FILLER_154_1044 ();
 sg13g2_fill_1 FILLER_154_1046 ();
 sg13g2_fill_4 FILLER_154_1051 ();
 sg13g2_fill_2 FILLER_154_1055 ();
 sg13g2_fill_4 FILLER_154_1067 ();
 sg13g2_fill_2 FILLER_154_1085 ();
 sg13g2_fill_8 FILLER_154_1118 ();
 sg13g2_fill_1 FILLER_154_1126 ();
 sg13g2_fill_8 FILLER_154_1135 ();
 sg13g2_fill_8 FILLER_154_1143 ();
 sg13g2_fill_8 FILLER_154_1156 ();
 sg13g2_fill_8 FILLER_154_1164 ();
 sg13g2_fill_8 FILLER_154_1172 ();
 sg13g2_fill_2 FILLER_154_1184 ();
 sg13g2_fill_4 FILLER_154_1190 ();
 sg13g2_fill_1 FILLER_154_1194 ();
 sg13g2_fill_2 FILLER_154_1203 ();
 sg13g2_fill_1 FILLER_154_1215 ();
 sg13g2_fill_2 FILLER_154_1225 ();
 sg13g2_fill_1 FILLER_154_1227 ();
 sg13g2_fill_4 FILLER_154_1237 ();
 sg13g2_fill_2 FILLER_154_1241 ();
 sg13g2_fill_2 FILLER_154_1269 ();
 sg13g2_fill_2 FILLER_154_1287 ();
 sg13g2_fill_1 FILLER_154_1289 ();
 sg13g2_fill_8 FILLER_154_1305 ();
 sg13g2_fill_8 FILLER_154_1313 ();
 sg13g2_fill_8 FILLER_154_1321 ();
 sg13g2_fill_8 FILLER_154_1329 ();
 sg13g2_fill_8 FILLER_154_1337 ();
 sg13g2_fill_8 FILLER_154_1345 ();
 sg13g2_fill_8 FILLER_154_1353 ();
 sg13g2_fill_8 FILLER_154_1361 ();
 sg13g2_fill_8 FILLER_154_1369 ();
 sg13g2_fill_1 FILLER_154_1377 ();
 sg13g2_fill_4 FILLER_154_1381 ();
 sg13g2_fill_1 FILLER_154_1385 ();
 sg13g2_fill_4 FILLER_154_1415 ();
 sg13g2_fill_2 FILLER_154_1432 ();
 sg13g2_fill_1 FILLER_154_1442 ();
 sg13g2_fill_8 FILLER_154_1453 ();
 sg13g2_fill_8 FILLER_154_1461 ();
 sg13g2_fill_8 FILLER_154_1469 ();
 sg13g2_fill_8 FILLER_154_1477 ();
 sg13g2_fill_8 FILLER_154_1485 ();
 sg13g2_fill_4 FILLER_154_1493 ();
 sg13g2_fill_1 FILLER_154_1518 ();
 sg13g2_fill_4 FILLER_154_1529 ();
 sg13g2_fill_8 FILLER_154_1551 ();
 sg13g2_fill_4 FILLER_154_1559 ();
 sg13g2_fill_2 FILLER_154_1563 ();
 sg13g2_fill_1 FILLER_154_1565 ();
 sg13g2_fill_8 FILLER_155_0 ();
 sg13g2_fill_8 FILLER_155_8 ();
 sg13g2_fill_8 FILLER_155_16 ();
 sg13g2_fill_8 FILLER_155_24 ();
 sg13g2_fill_8 FILLER_155_32 ();
 sg13g2_fill_2 FILLER_155_40 ();
 sg13g2_fill_2 FILLER_155_82 ();
 sg13g2_fill_8 FILLER_155_90 ();
 sg13g2_fill_8 FILLER_155_98 ();
 sg13g2_fill_1 FILLER_155_106 ();
 sg13g2_fill_8 FILLER_155_143 ();
 sg13g2_fill_2 FILLER_155_151 ();
 sg13g2_fill_1 FILLER_155_163 ();
 sg13g2_fill_2 FILLER_155_190 ();
 sg13g2_fill_8 FILLER_155_197 ();
 sg13g2_fill_1 FILLER_155_205 ();
 sg13g2_fill_8 FILLER_155_250 ();
 sg13g2_fill_8 FILLER_155_258 ();
 sg13g2_fill_4 FILLER_155_266 ();
 sg13g2_fill_4 FILLER_155_291 ();
 sg13g2_fill_2 FILLER_155_295 ();
 sg13g2_fill_8 FILLER_155_305 ();
 sg13g2_fill_4 FILLER_155_313 ();
 sg13g2_fill_4 FILLER_155_358 ();
 sg13g2_fill_1 FILLER_155_398 ();
 sg13g2_fill_1 FILLER_155_404 ();
 sg13g2_fill_8 FILLER_155_410 ();
 sg13g2_fill_1 FILLER_155_418 ();
 sg13g2_fill_8 FILLER_155_462 ();
 sg13g2_fill_1 FILLER_155_470 ();
 sg13g2_fill_8 FILLER_155_477 ();
 sg13g2_fill_8 FILLER_155_485 ();
 sg13g2_fill_8 FILLER_155_493 ();
 sg13g2_fill_8 FILLER_155_501 ();
 sg13g2_fill_8 FILLER_155_509 ();
 sg13g2_fill_4 FILLER_155_517 ();
 sg13g2_fill_2 FILLER_155_521 ();
 sg13g2_fill_8 FILLER_155_539 ();
 sg13g2_fill_4 FILLER_155_557 ();
 sg13g2_fill_2 FILLER_155_606 ();
 sg13g2_fill_4 FILLER_155_613 ();
 sg13g2_fill_4 FILLER_155_625 ();
 sg13g2_fill_2 FILLER_155_629 ();
 sg13g2_fill_1 FILLER_155_631 ();
 sg13g2_fill_8 FILLER_155_657 ();
 sg13g2_fill_8 FILLER_155_665 ();
 sg13g2_fill_8 FILLER_155_673 ();
 sg13g2_fill_8 FILLER_155_717 ();
 sg13g2_fill_8 FILLER_155_725 ();
 sg13g2_fill_8 FILLER_155_733 ();
 sg13g2_fill_8 FILLER_155_741 ();
 sg13g2_fill_2 FILLER_155_749 ();
 sg13g2_fill_8 FILLER_155_765 ();
 sg13g2_fill_8 FILLER_155_773 ();
 sg13g2_fill_4 FILLER_155_781 ();
 sg13g2_fill_2 FILLER_155_785 ();
 sg13g2_fill_1 FILLER_155_787 ();
 sg13g2_fill_4 FILLER_155_797 ();
 sg13g2_fill_2 FILLER_155_801 ();
 sg13g2_fill_1 FILLER_155_803 ();
 sg13g2_fill_8 FILLER_155_809 ();
 sg13g2_fill_4 FILLER_155_817 ();
 sg13g2_fill_2 FILLER_155_821 ();
 sg13g2_fill_1 FILLER_155_842 ();
 sg13g2_fill_2 FILLER_155_859 ();
 sg13g2_fill_1 FILLER_155_871 ();
 sg13g2_fill_8 FILLER_155_885 ();
 sg13g2_fill_4 FILLER_155_893 ();
 sg13g2_fill_2 FILLER_155_903 ();
 sg13g2_fill_1 FILLER_155_905 ();
 sg13g2_fill_8 FILLER_155_926 ();
 sg13g2_fill_2 FILLER_155_934 ();
 sg13g2_fill_1 FILLER_155_936 ();
 sg13g2_fill_8 FILLER_155_957 ();
 sg13g2_fill_1 FILLER_155_965 ();
 sg13g2_fill_2 FILLER_155_969 ();
 sg13g2_fill_1 FILLER_155_971 ();
 sg13g2_fill_8 FILLER_155_988 ();
 sg13g2_fill_1 FILLER_155_996 ();
 sg13g2_fill_2 FILLER_155_1006 ();
 sg13g2_fill_2 FILLER_155_1013 ();
 sg13g2_fill_1 FILLER_155_1015 ();
 sg13g2_fill_4 FILLER_155_1024 ();
 sg13g2_fill_2 FILLER_155_1028 ();
 sg13g2_fill_8 FILLER_155_1038 ();
 sg13g2_fill_8 FILLER_155_1046 ();
 sg13g2_fill_8 FILLER_155_1054 ();
 sg13g2_fill_8 FILLER_155_1062 ();
 sg13g2_fill_4 FILLER_155_1090 ();
 sg13g2_fill_2 FILLER_155_1094 ();
 sg13g2_fill_1 FILLER_155_1096 ();
 sg13g2_fill_1 FILLER_155_1100 ();
 sg13g2_fill_2 FILLER_155_1113 ();
 sg13g2_fill_2 FILLER_155_1130 ();
 sg13g2_fill_4 FILLER_155_1175 ();
 sg13g2_fill_2 FILLER_155_1179 ();
 sg13g2_fill_1 FILLER_155_1181 ();
 sg13g2_fill_2 FILLER_155_1199 ();
 sg13g2_fill_1 FILLER_155_1201 ();
 sg13g2_fill_1 FILLER_155_1221 ();
 sg13g2_fill_4 FILLER_155_1246 ();
 sg13g2_fill_2 FILLER_155_1250 ();
 sg13g2_fill_2 FILLER_155_1256 ();
 sg13g2_fill_1 FILLER_155_1258 ();
 sg13g2_fill_4 FILLER_155_1267 ();
 sg13g2_fill_2 FILLER_155_1271 ();
 sg13g2_fill_1 FILLER_155_1286 ();
 sg13g2_fill_2 FILLER_155_1292 ();
 sg13g2_fill_8 FILLER_155_1307 ();
 sg13g2_fill_1 FILLER_155_1315 ();
 sg13g2_fill_8 FILLER_155_1334 ();
 sg13g2_fill_2 FILLER_155_1342 ();
 sg13g2_fill_1 FILLER_155_1344 ();
 sg13g2_fill_8 FILLER_155_1361 ();
 sg13g2_fill_1 FILLER_155_1369 ();
 sg13g2_fill_2 FILLER_155_1382 ();
 sg13g2_fill_4 FILLER_155_1398 ();
 sg13g2_fill_8 FILLER_155_1407 ();
 sg13g2_fill_8 FILLER_155_1415 ();
 sg13g2_fill_1 FILLER_155_1423 ();
 sg13g2_fill_4 FILLER_155_1432 ();
 sg13g2_fill_2 FILLER_155_1436 ();
 sg13g2_fill_1 FILLER_155_1438 ();
 sg13g2_fill_8 FILLER_155_1446 ();
 sg13g2_fill_8 FILLER_155_1454 ();
 sg13g2_fill_8 FILLER_155_1462 ();
 sg13g2_fill_8 FILLER_155_1470 ();
 sg13g2_fill_2 FILLER_155_1478 ();
 sg13g2_fill_1 FILLER_155_1480 ();
 sg13g2_fill_8 FILLER_155_1507 ();
 sg13g2_fill_8 FILLER_155_1515 ();
 sg13g2_fill_8 FILLER_155_1523 ();
 sg13g2_fill_2 FILLER_155_1531 ();
 sg13g2_fill_1 FILLER_155_1533 ();
 sg13g2_fill_4 FILLER_155_1545 ();
 sg13g2_fill_1 FILLER_155_1549 ();
 sg13g2_fill_8 FILLER_155_1571 ();
 sg13g2_fill_8 FILLER_155_1579 ();
 sg13g2_fill_4 FILLER_155_1587 ();
 sg13g2_fill_1 FILLER_155_1591 ();
 sg13g2_fill_8 FILLER_156_0 ();
 sg13g2_fill_8 FILLER_156_8 ();
 sg13g2_fill_8 FILLER_156_16 ();
 sg13g2_fill_8 FILLER_156_24 ();
 sg13g2_fill_8 FILLER_156_32 ();
 sg13g2_fill_4 FILLER_156_40 ();
 sg13g2_fill_2 FILLER_156_44 ();
 sg13g2_fill_1 FILLER_156_46 ();
 sg13g2_fill_1 FILLER_156_83 ();
 sg13g2_fill_1 FILLER_156_90 ();
 sg13g2_fill_8 FILLER_156_101 ();
 sg13g2_fill_8 FILLER_156_109 ();
 sg13g2_fill_8 FILLER_156_117 ();
 sg13g2_fill_4 FILLER_156_125 ();
 sg13g2_fill_1 FILLER_156_129 ();
 sg13g2_fill_2 FILLER_156_166 ();
 sg13g2_fill_1 FILLER_156_168 ();
 sg13g2_fill_8 FILLER_156_182 ();
 sg13g2_fill_8 FILLER_156_190 ();
 sg13g2_fill_8 FILLER_156_198 ();
 sg13g2_fill_8 FILLER_156_206 ();
 sg13g2_fill_8 FILLER_156_214 ();
 sg13g2_fill_8 FILLER_156_222 ();
 sg13g2_fill_8 FILLER_156_230 ();
 sg13g2_fill_8 FILLER_156_238 ();
 sg13g2_fill_4 FILLER_156_246 ();
 sg13g2_fill_1 FILLER_156_250 ();
 sg13g2_fill_8 FILLER_156_277 ();
 sg13g2_fill_8 FILLER_156_321 ();
 sg13g2_fill_8 FILLER_156_329 ();
 sg13g2_fill_4 FILLER_156_337 ();
 sg13g2_fill_8 FILLER_156_380 ();
 sg13g2_fill_8 FILLER_156_388 ();
 sg13g2_fill_4 FILLER_156_396 ();
 sg13g2_fill_2 FILLER_156_400 ();
 sg13g2_fill_1 FILLER_156_410 ();
 sg13g2_fill_8 FILLER_156_457 ();
 sg13g2_fill_4 FILLER_156_465 ();
 sg13g2_fill_4 FILLER_156_479 ();
 sg13g2_fill_2 FILLER_156_527 ();
 sg13g2_fill_4 FILLER_156_539 ();
 sg13g2_fill_4 FILLER_156_548 ();
 sg13g2_fill_8 FILLER_156_562 ();
 sg13g2_fill_4 FILLER_156_570 ();
 sg13g2_fill_1 FILLER_156_574 ();
 sg13g2_fill_4 FILLER_156_585 ();
 sg13g2_fill_1 FILLER_156_589 ();
 sg13g2_fill_4 FILLER_156_608 ();
 sg13g2_fill_2 FILLER_156_612 ();
 sg13g2_fill_8 FILLER_156_620 ();
 sg13g2_fill_4 FILLER_156_628 ();
 sg13g2_fill_1 FILLER_156_632 ();
 sg13g2_fill_8 FILLER_156_643 ();
 sg13g2_fill_8 FILLER_156_651 ();
 sg13g2_fill_8 FILLER_156_659 ();
 sg13g2_fill_4 FILLER_156_667 ();
 sg13g2_fill_4 FILLER_156_689 ();
 sg13g2_fill_2 FILLER_156_693 ();
 sg13g2_fill_4 FILLER_156_705 ();
 sg13g2_fill_2 FILLER_156_735 ();
 sg13g2_fill_1 FILLER_156_737 ();
 sg13g2_fill_2 FILLER_156_748 ();
 sg13g2_fill_1 FILLER_156_750 ();
 sg13g2_fill_8 FILLER_156_761 ();
 sg13g2_fill_4 FILLER_156_769 ();
 sg13g2_fill_2 FILLER_156_773 ();
 sg13g2_fill_1 FILLER_156_775 ();
 sg13g2_fill_8 FILLER_156_798 ();
 sg13g2_fill_2 FILLER_156_806 ();
 sg13g2_fill_2 FILLER_156_818 ();
 sg13g2_fill_8 FILLER_156_838 ();
 sg13g2_fill_8 FILLER_156_846 ();
 sg13g2_fill_1 FILLER_156_859 ();
 sg13g2_fill_8 FILLER_156_894 ();
 sg13g2_fill_4 FILLER_156_906 ();
 sg13g2_fill_8 FILLER_156_922 ();
 sg13g2_fill_8 FILLER_156_960 ();
 sg13g2_fill_1 FILLER_156_968 ();
 sg13g2_fill_2 FILLER_156_994 ();
 sg13g2_fill_2 FILLER_156_1001 ();
 sg13g2_fill_2 FILLER_156_1008 ();
 sg13g2_fill_8 FILLER_156_1018 ();
 sg13g2_fill_4 FILLER_156_1026 ();
 sg13g2_fill_1 FILLER_156_1030 ();
 sg13g2_fill_4 FILLER_156_1039 ();
 sg13g2_fill_4 FILLER_156_1051 ();
 sg13g2_fill_1 FILLER_156_1063 ();
 sg13g2_fill_4 FILLER_156_1072 ();
 sg13g2_fill_2 FILLER_156_1082 ();
 sg13g2_fill_4 FILLER_156_1103 ();
 sg13g2_fill_2 FILLER_156_1107 ();
 sg13g2_fill_1 FILLER_156_1109 ();
 sg13g2_fill_8 FILLER_156_1120 ();
 sg13g2_fill_8 FILLER_156_1136 ();
 sg13g2_fill_1 FILLER_156_1144 ();
 sg13g2_fill_8 FILLER_156_1154 ();
 sg13g2_fill_1 FILLER_156_1162 ();
 sg13g2_fill_4 FILLER_156_1167 ();
 sg13g2_fill_2 FILLER_156_1196 ();
 sg13g2_fill_1 FILLER_156_1198 ();
 sg13g2_fill_4 FILLER_156_1203 ();
 sg13g2_fill_2 FILLER_156_1207 ();
 sg13g2_fill_1 FILLER_156_1209 ();
 sg13g2_fill_2 FILLER_156_1244 ();
 sg13g2_fill_4 FILLER_156_1257 ();
 sg13g2_fill_2 FILLER_156_1261 ();
 sg13g2_fill_2 FILLER_156_1274 ();
 sg13g2_fill_2 FILLER_156_1292 ();
 sg13g2_fill_2 FILLER_156_1306 ();
 sg13g2_fill_2 FILLER_156_1335 ();
 sg13g2_fill_2 FILLER_156_1386 ();
 sg13g2_fill_1 FILLER_156_1388 ();
 sg13g2_fill_8 FILLER_156_1409 ();
 sg13g2_fill_4 FILLER_156_1417 ();
 sg13g2_fill_2 FILLER_156_1425 ();
 sg13g2_fill_8 FILLER_156_1431 ();
 sg13g2_fill_1 FILLER_156_1439 ();
 sg13g2_fill_8 FILLER_156_1448 ();
 sg13g2_fill_8 FILLER_156_1456 ();
 sg13g2_fill_8 FILLER_156_1464 ();
 sg13g2_fill_8 FILLER_156_1472 ();
 sg13g2_fill_8 FILLER_156_1480 ();
 sg13g2_fill_8 FILLER_156_1488 ();
 sg13g2_fill_2 FILLER_156_1496 ();
 sg13g2_fill_1 FILLER_156_1498 ();
 sg13g2_fill_8 FILLER_156_1528 ();
 sg13g2_fill_1 FILLER_156_1536 ();
 sg13g2_fill_4 FILLER_156_1562 ();
 sg13g2_fill_8 FILLER_157_0 ();
 sg13g2_fill_8 FILLER_157_8 ();
 sg13g2_fill_8 FILLER_157_16 ();
 sg13g2_fill_8 FILLER_157_24 ();
 sg13g2_fill_8 FILLER_157_32 ();
 sg13g2_fill_8 FILLER_157_40 ();
 sg13g2_fill_8 FILLER_157_48 ();
 sg13g2_fill_8 FILLER_157_56 ();
 sg13g2_fill_8 FILLER_157_64 ();
 sg13g2_fill_8 FILLER_157_72 ();
 sg13g2_fill_8 FILLER_157_80 ();
 sg13g2_fill_2 FILLER_157_88 ();
 sg13g2_fill_4 FILLER_157_116 ();
 sg13g2_fill_2 FILLER_157_140 ();
 sg13g2_fill_4 FILLER_157_148 ();
 sg13g2_fill_1 FILLER_157_152 ();
 sg13g2_fill_8 FILLER_157_158 ();
 sg13g2_fill_4 FILLER_157_166 ();
 sg13g2_fill_2 FILLER_157_170 ();
 sg13g2_fill_1 FILLER_157_172 ();
 sg13g2_fill_8 FILLER_157_199 ();
 sg13g2_fill_8 FILLER_157_207 ();
 sg13g2_fill_2 FILLER_157_215 ();
 sg13g2_fill_8 FILLER_157_258 ();
 sg13g2_fill_2 FILLER_157_266 ();
 sg13g2_fill_1 FILLER_157_268 ();
 sg13g2_fill_8 FILLER_157_298 ();
 sg13g2_fill_4 FILLER_157_306 ();
 sg13g2_fill_2 FILLER_157_310 ();
 sg13g2_fill_1 FILLER_157_312 ();
 sg13g2_fill_4 FILLER_157_339 ();
 sg13g2_fill_2 FILLER_157_343 ();
 sg13g2_fill_1 FILLER_157_345 ();
 sg13g2_fill_8 FILLER_157_355 ();
 sg13g2_fill_2 FILLER_157_363 ();
 sg13g2_fill_1 FILLER_157_365 ();
 sg13g2_fill_8 FILLER_157_391 ();
 sg13g2_fill_2 FILLER_157_407 ();
 sg13g2_fill_8 FILLER_157_414 ();
 sg13g2_fill_4 FILLER_157_422 ();
 sg13g2_fill_2 FILLER_157_426 ();
 sg13g2_fill_8 FILLER_157_433 ();
 sg13g2_fill_8 FILLER_157_441 ();
 sg13g2_fill_2 FILLER_157_449 ();
 sg13g2_fill_1 FILLER_157_487 ();
 sg13g2_fill_8 FILLER_157_501 ();
 sg13g2_fill_4 FILLER_157_509 ();
 sg13g2_fill_8 FILLER_157_523 ();
 sg13g2_fill_8 FILLER_157_531 ();
 sg13g2_fill_1 FILLER_157_539 ();
 sg13g2_fill_8 FILLER_157_553 ();
 sg13g2_fill_4 FILLER_157_561 ();
 sg13g2_fill_2 FILLER_157_593 ();
 sg13g2_fill_2 FILLER_157_600 ();
 sg13g2_fill_1 FILLER_157_602 ();
 sg13g2_fill_2 FILLER_157_677 ();
 sg13g2_fill_1 FILLER_157_679 ();
 sg13g2_fill_8 FILLER_157_690 ();
 sg13g2_fill_4 FILLER_157_698 ();
 sg13g2_fill_2 FILLER_157_702 ();
 sg13g2_fill_1 FILLER_157_704 ();
 sg13g2_fill_4 FILLER_157_715 ();
 sg13g2_fill_1 FILLER_157_719 ();
 sg13g2_fill_1 FILLER_157_752 ();
 sg13g2_fill_1 FILLER_157_766 ();
 sg13g2_fill_2 FILLER_157_777 ();
 sg13g2_fill_2 FILLER_157_795 ();
 sg13g2_fill_1 FILLER_157_803 ();
 sg13g2_fill_2 FILLER_157_818 ();
 sg13g2_fill_1 FILLER_157_820 ();
 sg13g2_fill_2 FILLER_157_830 ();
 sg13g2_fill_8 FILLER_157_847 ();
 sg13g2_fill_8 FILLER_157_855 ();
 sg13g2_fill_4 FILLER_157_863 ();
 sg13g2_fill_1 FILLER_157_867 ();
 sg13g2_fill_8 FILLER_157_873 ();
 sg13g2_fill_4 FILLER_157_881 ();
 sg13g2_fill_4 FILLER_157_890 ();
 sg13g2_fill_2 FILLER_157_894 ();
 sg13g2_fill_8 FILLER_157_917 ();
 sg13g2_fill_8 FILLER_157_925 ();
 sg13g2_fill_8 FILLER_157_933 ();
 sg13g2_fill_8 FILLER_157_941 ();
 sg13g2_fill_8 FILLER_157_949 ();
 sg13g2_fill_8 FILLER_157_957 ();
 sg13g2_fill_8 FILLER_157_965 ();
 sg13g2_fill_1 FILLER_157_973 ();
 sg13g2_fill_4 FILLER_157_989 ();
 sg13g2_fill_2 FILLER_157_993 ();
 sg13g2_fill_1 FILLER_157_1003 ();
 sg13g2_fill_1 FILLER_157_1019 ();
 sg13g2_fill_4 FILLER_157_1027 ();
 sg13g2_fill_2 FILLER_157_1031 ();
 sg13g2_fill_1 FILLER_157_1038 ();
 sg13g2_fill_1 FILLER_157_1080 ();
 sg13g2_fill_2 FILLER_157_1087 ();
 sg13g2_fill_2 FILLER_157_1113 ();
 sg13g2_fill_2 FILLER_157_1131 ();
 sg13g2_fill_2 FILLER_157_1146 ();
 sg13g2_fill_4 FILLER_157_1152 ();
 sg13g2_fill_8 FILLER_157_1161 ();
 sg13g2_fill_4 FILLER_157_1169 ();
 sg13g2_fill_2 FILLER_157_1178 ();
 sg13g2_fill_4 FILLER_157_1184 ();
 sg13g2_fill_2 FILLER_157_1188 ();
 sg13g2_fill_8 FILLER_157_1194 ();
 sg13g2_fill_8 FILLER_157_1202 ();
 sg13g2_fill_2 FILLER_157_1210 ();
 sg13g2_fill_1 FILLER_157_1212 ();
 sg13g2_fill_4 FILLER_157_1217 ();
 sg13g2_fill_2 FILLER_157_1221 ();
 sg13g2_fill_1 FILLER_157_1223 ();
 sg13g2_fill_1 FILLER_157_1270 ();
 sg13g2_fill_2 FILLER_157_1278 ();
 sg13g2_fill_1 FILLER_157_1290 ();
 sg13g2_fill_8 FILLER_157_1305 ();
 sg13g2_fill_2 FILLER_157_1313 ();
 sg13g2_fill_8 FILLER_157_1324 ();
 sg13g2_fill_4 FILLER_157_1332 ();
 sg13g2_fill_1 FILLER_157_1336 ();
 sg13g2_fill_2 FILLER_157_1350 ();
 sg13g2_fill_1 FILLER_157_1352 ();
 sg13g2_fill_8 FILLER_157_1363 ();
 sg13g2_fill_2 FILLER_157_1371 ();
 sg13g2_fill_1 FILLER_157_1373 ();
 sg13g2_fill_4 FILLER_157_1387 ();
 sg13g2_fill_1 FILLER_157_1391 ();
 sg13g2_fill_2 FILLER_157_1411 ();
 sg13g2_fill_1 FILLER_157_1413 ();
 sg13g2_fill_2 FILLER_157_1435 ();
 sg13g2_fill_1 FILLER_157_1437 ();
 sg13g2_fill_8 FILLER_157_1459 ();
 sg13g2_fill_8 FILLER_157_1467 ();
 sg13g2_fill_8 FILLER_157_1475 ();
 sg13g2_fill_4 FILLER_157_1483 ();
 sg13g2_fill_4 FILLER_157_1513 ();
 sg13g2_fill_2 FILLER_157_1517 ();
 sg13g2_fill_8 FILLER_157_1582 ();
 sg13g2_fill_2 FILLER_157_1590 ();
 sg13g2_fill_8 FILLER_158_0 ();
 sg13g2_fill_8 FILLER_158_8 ();
 sg13g2_fill_8 FILLER_158_16 ();
 sg13g2_fill_8 FILLER_158_24 ();
 sg13g2_fill_8 FILLER_158_32 ();
 sg13g2_fill_8 FILLER_158_40 ();
 sg13g2_fill_4 FILLER_158_48 ();
 sg13g2_fill_2 FILLER_158_52 ();
 sg13g2_fill_1 FILLER_158_54 ();
 sg13g2_fill_1 FILLER_158_81 ();
 sg13g2_fill_2 FILLER_158_92 ();
 sg13g2_fill_4 FILLER_158_120 ();
 sg13g2_fill_2 FILLER_158_124 ();
 sg13g2_fill_1 FILLER_158_126 ();
 sg13g2_fill_4 FILLER_158_137 ();
 sg13g2_fill_2 FILLER_158_162 ();
 sg13g2_fill_8 FILLER_158_210 ();
 sg13g2_fill_4 FILLER_158_239 ();
 sg13g2_fill_4 FILLER_158_279 ();
 sg13g2_fill_2 FILLER_158_283 ();
 sg13g2_fill_8 FILLER_158_293 ();
 sg13g2_fill_4 FILLER_158_301 ();
 sg13g2_fill_2 FILLER_158_305 ();
 sg13g2_fill_1 FILLER_158_307 ();
 sg13g2_fill_8 FILLER_158_344 ();
 sg13g2_fill_2 FILLER_158_352 ();
 sg13g2_fill_2 FILLER_158_411 ();
 sg13g2_fill_8 FILLER_158_418 ();
 sg13g2_fill_8 FILLER_158_426 ();
 sg13g2_fill_8 FILLER_158_434 ();
 sg13g2_fill_8 FILLER_158_442 ();
 sg13g2_fill_1 FILLER_158_450 ();
 sg13g2_fill_1 FILLER_158_461 ();
 sg13g2_fill_2 FILLER_158_482 ();
 sg13g2_fill_2 FILLER_158_537 ();
 sg13g2_fill_2 FILLER_158_552 ();
 sg13g2_fill_1 FILLER_158_554 ();
 sg13g2_fill_2 FILLER_158_597 ();
 sg13g2_fill_1 FILLER_158_599 ();
 sg13g2_fill_8 FILLER_158_635 ();
 sg13g2_fill_8 FILLER_158_643 ();
 sg13g2_fill_8 FILLER_158_651 ();
 sg13g2_fill_4 FILLER_158_659 ();
 sg13g2_fill_1 FILLER_158_663 ();
 sg13g2_fill_8 FILLER_158_674 ();
 sg13g2_fill_4 FILLER_158_708 ();
 sg13g2_fill_2 FILLER_158_712 ();
 sg13g2_fill_8 FILLER_158_754 ();
 sg13g2_fill_2 FILLER_158_762 ();
 sg13g2_fill_8 FILLER_158_771 ();
 sg13g2_fill_8 FILLER_158_779 ();
 sg13g2_fill_2 FILLER_158_787 ();
 sg13g2_fill_4 FILLER_158_794 ();
 sg13g2_fill_1 FILLER_158_798 ();
 sg13g2_fill_8 FILLER_158_809 ();
 sg13g2_fill_8 FILLER_158_817 ();
 sg13g2_fill_8 FILLER_158_825 ();
 sg13g2_fill_2 FILLER_158_833 ();
 sg13g2_fill_4 FILLER_158_865 ();
 sg13g2_fill_4 FILLER_158_878 ();
 sg13g2_fill_2 FILLER_158_882 ();
 sg13g2_fill_1 FILLER_158_884 ();
 sg13g2_fill_1 FILLER_158_906 ();
 sg13g2_fill_8 FILLER_158_925 ();
 sg13g2_fill_8 FILLER_158_933 ();
 sg13g2_fill_8 FILLER_158_941 ();
 sg13g2_fill_8 FILLER_158_949 ();
 sg13g2_fill_8 FILLER_158_957 ();
 sg13g2_fill_8 FILLER_158_965 ();
 sg13g2_fill_8 FILLER_158_973 ();
 sg13g2_fill_2 FILLER_158_981 ();
 sg13g2_fill_4 FILLER_158_991 ();
 sg13g2_fill_4 FILLER_158_1009 ();
 sg13g2_fill_2 FILLER_158_1013 ();
 sg13g2_fill_4 FILLER_158_1020 ();
 sg13g2_fill_1 FILLER_158_1024 ();
 sg13g2_fill_2 FILLER_158_1030 ();
 sg13g2_fill_2 FILLER_158_1054 ();
 sg13g2_fill_2 FILLER_158_1061 ();
 sg13g2_fill_1 FILLER_158_1072 ();
 sg13g2_fill_2 FILLER_158_1078 ();
 sg13g2_fill_1 FILLER_158_1095 ();
 sg13g2_fill_8 FILLER_158_1101 ();
 sg13g2_fill_4 FILLER_158_1109 ();
 sg13g2_fill_2 FILLER_158_1113 ();
 sg13g2_fill_1 FILLER_158_1115 ();
 sg13g2_fill_2 FILLER_158_1128 ();
 sg13g2_fill_1 FILLER_158_1130 ();
 sg13g2_fill_4 FILLER_158_1136 ();
 sg13g2_fill_1 FILLER_158_1140 ();
 sg13g2_fill_2 FILLER_158_1146 ();
 sg13g2_fill_2 FILLER_158_1166 ();
 sg13g2_fill_1 FILLER_158_1168 ();
 sg13g2_fill_1 FILLER_158_1218 ();
 sg13g2_fill_2 FILLER_158_1222 ();
 sg13g2_fill_1 FILLER_158_1237 ();
 sg13g2_fill_2 FILLER_158_1249 ();
 sg13g2_fill_1 FILLER_158_1272 ();
 sg13g2_fill_1 FILLER_158_1290 ();
 sg13g2_fill_4 FILLER_158_1306 ();
 sg13g2_fill_8 FILLER_158_1318 ();
 sg13g2_fill_8 FILLER_158_1334 ();
 sg13g2_fill_2 FILLER_158_1342 ();
 sg13g2_fill_1 FILLER_158_1344 ();
 sg13g2_fill_8 FILLER_158_1350 ();
 sg13g2_fill_8 FILLER_158_1358 ();
 sg13g2_fill_8 FILLER_158_1366 ();
 sg13g2_fill_8 FILLER_158_1374 ();
 sg13g2_fill_8 FILLER_158_1382 ();
 sg13g2_fill_4 FILLER_158_1390 ();
 sg13g2_fill_2 FILLER_158_1394 ();
 sg13g2_fill_1 FILLER_158_1396 ();
 sg13g2_fill_8 FILLER_158_1402 ();
 sg13g2_fill_8 FILLER_158_1410 ();
 sg13g2_fill_2 FILLER_158_1418 ();
 sg13g2_fill_1 FILLER_158_1420 ();
 sg13g2_fill_4 FILLER_158_1434 ();
 sg13g2_fill_2 FILLER_158_1438 ();
 sg13g2_fill_8 FILLER_158_1459 ();
 sg13g2_fill_8 FILLER_158_1467 ();
 sg13g2_fill_8 FILLER_158_1475 ();
 sg13g2_fill_8 FILLER_158_1483 ();
 sg13g2_fill_8 FILLER_158_1491 ();
 sg13g2_fill_8 FILLER_158_1499 ();
 sg13g2_fill_8 FILLER_158_1507 ();
 sg13g2_fill_8 FILLER_158_1515 ();
 sg13g2_fill_8 FILLER_158_1523 ();
 sg13g2_fill_8 FILLER_158_1531 ();
 sg13g2_fill_4 FILLER_158_1539 ();
 sg13g2_fill_2 FILLER_158_1543 ();
 sg13g2_fill_1 FILLER_158_1545 ();
 sg13g2_fill_8 FILLER_158_1556 ();
 sg13g2_fill_8 FILLER_158_1564 ();
 sg13g2_fill_8 FILLER_158_1572 ();
 sg13g2_fill_8 FILLER_158_1580 ();
 sg13g2_fill_4 FILLER_158_1588 ();
 sg13g2_fill_8 FILLER_159_0 ();
 sg13g2_fill_2 FILLER_159_8 ();
 sg13g2_fill_8 FILLER_159_18 ();
 sg13g2_fill_8 FILLER_159_26 ();
 sg13g2_fill_8 FILLER_159_34 ();
 sg13g2_fill_4 FILLER_159_42 ();
 sg13g2_fill_8 FILLER_159_82 ();
 sg13g2_fill_1 FILLER_159_90 ();
 sg13g2_fill_2 FILLER_159_101 ();
 sg13g2_fill_1 FILLER_159_103 ();
 sg13g2_fill_2 FILLER_159_149 ();
 sg13g2_fill_1 FILLER_159_151 ();
 sg13g2_fill_4 FILLER_159_168 ();
 sg13g2_fill_1 FILLER_159_172 ();
 sg13g2_fill_8 FILLER_159_183 ();
 sg13g2_fill_8 FILLER_159_191 ();
 sg13g2_fill_2 FILLER_159_199 ();
 sg13g2_fill_8 FILLER_159_253 ();
 sg13g2_fill_8 FILLER_159_261 ();
 sg13g2_fill_4 FILLER_159_269 ();
 sg13g2_fill_1 FILLER_159_273 ();
 sg13g2_fill_4 FILLER_159_300 ();
 sg13g2_fill_4 FILLER_159_360 ();
 sg13g2_fill_2 FILLER_159_364 ();
 sg13g2_fill_8 FILLER_159_370 ();
 sg13g2_fill_8 FILLER_159_378 ();
 sg13g2_fill_8 FILLER_159_386 ();
 sg13g2_fill_4 FILLER_159_394 ();
 sg13g2_fill_2 FILLER_159_398 ();
 sg13g2_fill_2 FILLER_159_405 ();
 sg13g2_fill_2 FILLER_159_449 ();
 sg13g2_fill_1 FILLER_159_451 ();
 sg13g2_fill_8 FILLER_159_462 ();
 sg13g2_fill_8 FILLER_159_470 ();
 sg13g2_fill_8 FILLER_159_478 ();
 sg13g2_fill_8 FILLER_159_486 ();
 sg13g2_fill_8 FILLER_159_494 ();
 sg13g2_fill_1 FILLER_159_502 ();
 sg13g2_fill_8 FILLER_159_508 ();
 sg13g2_fill_8 FILLER_159_516 ();
 sg13g2_fill_2 FILLER_159_524 ();
 sg13g2_fill_4 FILLER_159_542 ();
 sg13g2_fill_4 FILLER_159_605 ();
 sg13g2_fill_2 FILLER_159_609 ();
 sg13g2_fill_4 FILLER_159_660 ();
 sg13g2_fill_8 FILLER_159_674 ();
 sg13g2_fill_8 FILLER_159_682 ();
 sg13g2_fill_1 FILLER_159_690 ();
 sg13g2_fill_4 FILLER_159_726 ();
 sg13g2_fill_8 FILLER_159_766 ();
 sg13g2_fill_4 FILLER_159_774 ();
 sg13g2_fill_1 FILLER_159_778 ();
 sg13g2_fill_1 FILLER_159_784 ();
 sg13g2_fill_2 FILLER_159_791 ();
 sg13g2_fill_1 FILLER_159_793 ();
 sg13g2_fill_1 FILLER_159_804 ();
 sg13g2_fill_2 FILLER_159_831 ();
 sg13g2_fill_1 FILLER_159_833 ();
 sg13g2_fill_8 FILLER_159_844 ();
 sg13g2_fill_2 FILLER_159_852 ();
 sg13g2_fill_1 FILLER_159_854 ();
 sg13g2_fill_2 FILLER_159_876 ();
 sg13g2_fill_1 FILLER_159_878 ();
 sg13g2_fill_2 FILLER_159_893 ();
 sg13g2_fill_8 FILLER_159_899 ();
 sg13g2_fill_1 FILLER_159_907 ();
 sg13g2_fill_8 FILLER_159_913 ();
 sg13g2_fill_8 FILLER_159_921 ();
 sg13g2_fill_8 FILLER_159_929 ();
 sg13g2_fill_8 FILLER_159_937 ();
 sg13g2_fill_8 FILLER_159_945 ();
 sg13g2_fill_2 FILLER_159_953 ();
 sg13g2_fill_1 FILLER_159_955 ();
 sg13g2_fill_8 FILLER_159_980 ();
 sg13g2_fill_4 FILLER_159_988 ();
 sg13g2_fill_8 FILLER_159_1002 ();
 sg13g2_fill_8 FILLER_159_1010 ();
 sg13g2_fill_1 FILLER_159_1018 ();
 sg13g2_fill_4 FILLER_159_1027 ();
 sg13g2_fill_1 FILLER_159_1031 ();
 sg13g2_fill_4 FILLER_159_1035 ();
 sg13g2_fill_8 FILLER_159_1043 ();
 sg13g2_fill_2 FILLER_159_1051 ();
 sg13g2_fill_1 FILLER_159_1053 ();
 sg13g2_fill_1 FILLER_159_1069 ();
 sg13g2_fill_2 FILLER_159_1082 ();
 sg13g2_fill_4 FILLER_159_1096 ();
 sg13g2_fill_2 FILLER_159_1100 ();
 sg13g2_fill_8 FILLER_159_1109 ();
 sg13g2_fill_8 FILLER_159_1117 ();
 sg13g2_fill_4 FILLER_159_1125 ();
 sg13g2_fill_2 FILLER_159_1129 ();
 sg13g2_fill_1 FILLER_159_1131 ();
 sg13g2_fill_4 FILLER_159_1144 ();
 sg13g2_fill_8 FILLER_159_1159 ();
 sg13g2_fill_2 FILLER_159_1170 ();
 sg13g2_fill_1 FILLER_159_1172 ();
 sg13g2_fill_1 FILLER_159_1178 ();
 sg13g2_fill_8 FILLER_159_1184 ();
 sg13g2_fill_1 FILLER_159_1192 ();
 sg13g2_fill_1 FILLER_159_1203 ();
 sg13g2_fill_1 FILLER_159_1215 ();
 sg13g2_fill_2 FILLER_159_1235 ();
 sg13g2_fill_1 FILLER_159_1237 ();
 sg13g2_fill_2 FILLER_159_1241 ();
 sg13g2_fill_8 FILLER_159_1297 ();
 sg13g2_fill_8 FILLER_159_1305 ();
 sg13g2_fill_4 FILLER_159_1313 ();
 sg13g2_fill_2 FILLER_159_1317 ();
 sg13g2_fill_1 FILLER_159_1319 ();
 sg13g2_fill_4 FILLER_159_1350 ();
 sg13g2_fill_8 FILLER_159_1362 ();
 sg13g2_fill_8 FILLER_159_1378 ();
 sg13g2_fill_4 FILLER_159_1386 ();
 sg13g2_fill_2 FILLER_159_1390 ();
 sg13g2_fill_1 FILLER_159_1392 ();
 sg13g2_fill_8 FILLER_159_1409 ();
 sg13g2_fill_1 FILLER_159_1417 ();
 sg13g2_fill_1 FILLER_159_1421 ();
 sg13g2_fill_4 FILLER_159_1431 ();
 sg13g2_fill_2 FILLER_159_1435 ();
 sg13g2_fill_2 FILLER_159_1445 ();
 sg13g2_fill_1 FILLER_159_1447 ();
 sg13g2_fill_8 FILLER_159_1453 ();
 sg13g2_fill_8 FILLER_159_1461 ();
 sg13g2_fill_8 FILLER_159_1469 ();
 sg13g2_fill_8 FILLER_159_1477 ();
 sg13g2_fill_8 FILLER_159_1485 ();
 sg13g2_fill_8 FILLER_159_1493 ();
 sg13g2_fill_8 FILLER_159_1501 ();
 sg13g2_fill_8 FILLER_159_1509 ();
 sg13g2_fill_8 FILLER_159_1517 ();
 sg13g2_fill_8 FILLER_159_1525 ();
 sg13g2_fill_8 FILLER_159_1533 ();
 sg13g2_fill_8 FILLER_159_1541 ();
 sg13g2_fill_8 FILLER_159_1549 ();
 sg13g2_fill_8 FILLER_159_1557 ();
 sg13g2_fill_8 FILLER_159_1565 ();
 sg13g2_fill_8 FILLER_159_1573 ();
 sg13g2_fill_8 FILLER_159_1581 ();
 sg13g2_fill_2 FILLER_159_1589 ();
 sg13g2_fill_1 FILLER_159_1591 ();
 sg13g2_fill_8 FILLER_160_0 ();
 sg13g2_fill_8 FILLER_160_8 ();
 sg13g2_fill_8 FILLER_160_16 ();
 sg13g2_fill_8 FILLER_160_24 ();
 sg13g2_fill_8 FILLER_160_32 ();
 sg13g2_fill_8 FILLER_160_40 ();
 sg13g2_fill_4 FILLER_160_48 ();
 sg13g2_fill_2 FILLER_160_52 ();
 sg13g2_fill_4 FILLER_160_64 ();
 sg13g2_fill_2 FILLER_160_68 ();
 sg13g2_fill_2 FILLER_160_137 ();
 sg13g2_fill_1 FILLER_160_139 ();
 sg13g2_fill_2 FILLER_160_156 ();
 sg13g2_fill_8 FILLER_160_184 ();
 sg13g2_fill_8 FILLER_160_192 ();
 sg13g2_fill_2 FILLER_160_200 ();
 sg13g2_fill_1 FILLER_160_202 ();
 sg13g2_fill_1 FILLER_160_228 ();
 sg13g2_fill_8 FILLER_160_244 ();
 sg13g2_fill_8 FILLER_160_252 ();
 sg13g2_fill_8 FILLER_160_260 ();
 sg13g2_fill_2 FILLER_160_268 ();
 sg13g2_fill_8 FILLER_160_280 ();
 sg13g2_fill_8 FILLER_160_288 ();
 sg13g2_fill_2 FILLER_160_296 ();
 sg13g2_fill_2 FILLER_160_308 ();
 sg13g2_fill_4 FILLER_160_360 ();
 sg13g2_fill_2 FILLER_160_364 ();
 sg13g2_fill_1 FILLER_160_366 ();
 sg13g2_fill_4 FILLER_160_403 ();
 sg13g2_fill_2 FILLER_160_443 ();
 sg13g2_fill_4 FILLER_160_477 ();
 sg13g2_fill_4 FILLER_160_540 ();
 sg13g2_fill_2 FILLER_160_544 ();
 sg13g2_fill_1 FILLER_160_546 ();
 sg13g2_fill_8 FILLER_160_557 ();
 sg13g2_fill_8 FILLER_160_565 ();
 sg13g2_fill_8 FILLER_160_573 ();
 sg13g2_fill_4 FILLER_160_581 ();
 sg13g2_fill_8 FILLER_160_592 ();
 sg13g2_fill_8 FILLER_160_600 ();
 sg13g2_fill_1 FILLER_160_608 ();
 sg13g2_fill_8 FILLER_160_619 ();
 sg13g2_fill_8 FILLER_160_627 ();
 sg13g2_fill_8 FILLER_160_635 ();
 sg13g2_fill_8 FILLER_160_643 ();
 sg13g2_fill_1 FILLER_160_651 ();
 sg13g2_fill_8 FILLER_160_678 ();
 sg13g2_fill_8 FILLER_160_686 ();
 sg13g2_fill_8 FILLER_160_694 ();
 sg13g2_fill_4 FILLER_160_702 ();
 sg13g2_fill_2 FILLER_160_706 ();
 sg13g2_fill_4 FILLER_160_734 ();
 sg13g2_fill_2 FILLER_160_738 ();
 sg13g2_fill_2 FILLER_160_775 ();
 sg13g2_fill_1 FILLER_160_777 ();
 sg13g2_fill_1 FILLER_160_783 ();
 sg13g2_fill_2 FILLER_160_799 ();
 sg13g2_fill_8 FILLER_160_821 ();
 sg13g2_fill_2 FILLER_160_845 ();
 sg13g2_fill_8 FILLER_160_852 ();
 sg13g2_fill_8 FILLER_160_860 ();
 sg13g2_fill_2 FILLER_160_868 ();
 sg13g2_fill_8 FILLER_160_875 ();
 sg13g2_fill_8 FILLER_160_883 ();
 sg13g2_fill_8 FILLER_160_891 ();
 sg13g2_fill_2 FILLER_160_899 ();
 sg13g2_fill_1 FILLER_160_910 ();
 sg13g2_fill_8 FILLER_160_920 ();
 sg13g2_fill_8 FILLER_160_928 ();
 sg13g2_fill_8 FILLER_160_936 ();
 sg13g2_fill_8 FILLER_160_944 ();
 sg13g2_fill_8 FILLER_160_952 ();
 sg13g2_fill_1 FILLER_160_984 ();
 sg13g2_fill_8 FILLER_160_1004 ();
 sg13g2_fill_8 FILLER_160_1012 ();
 sg13g2_fill_2 FILLER_160_1020 ();
 sg13g2_fill_8 FILLER_160_1027 ();
 sg13g2_fill_8 FILLER_160_1035 ();
 sg13g2_fill_8 FILLER_160_1043 ();
 sg13g2_fill_1 FILLER_160_1051 ();
 sg13g2_fill_1 FILLER_160_1060 ();
 sg13g2_fill_8 FILLER_160_1080 ();
 sg13g2_fill_8 FILLER_160_1088 ();
 sg13g2_fill_8 FILLER_160_1116 ();
 sg13g2_fill_4 FILLER_160_1124 ();
 sg13g2_fill_8 FILLER_160_1155 ();
 sg13g2_fill_1 FILLER_160_1163 ();
 sg13g2_fill_8 FILLER_160_1171 ();
 sg13g2_fill_8 FILLER_160_1187 ();
 sg13g2_fill_8 FILLER_160_1195 ();
 sg13g2_fill_1 FILLER_160_1203 ();
 sg13g2_fill_2 FILLER_160_1209 ();
 sg13g2_fill_4 FILLER_160_1214 ();
 sg13g2_fill_2 FILLER_160_1218 ();
 sg13g2_fill_1 FILLER_160_1220 ();
 sg13g2_fill_1 FILLER_160_1227 ();
 sg13g2_fill_1 FILLER_160_1233 ();
 sg13g2_fill_8 FILLER_160_1251 ();
 sg13g2_fill_4 FILLER_160_1259 ();
 sg13g2_fill_1 FILLER_160_1282 ();
 sg13g2_fill_4 FILLER_160_1300 ();
 sg13g2_fill_1 FILLER_160_1304 ();
 sg13g2_fill_1 FILLER_160_1324 ();
 sg13g2_fill_8 FILLER_160_1333 ();
 sg13g2_fill_8 FILLER_160_1341 ();
 sg13g2_fill_8 FILLER_160_1349 ();
 sg13g2_fill_4 FILLER_160_1357 ();
 sg13g2_fill_4 FILLER_160_1385 ();
 sg13g2_fill_2 FILLER_160_1389 ();
 sg13g2_fill_2 FILLER_160_1406 ();
 sg13g2_fill_1 FILLER_160_1408 ();
 sg13g2_fill_4 FILLER_160_1428 ();
 sg13g2_fill_2 FILLER_160_1432 ();
 sg13g2_fill_8 FILLER_160_1461 ();
 sg13g2_fill_8 FILLER_160_1469 ();
 sg13g2_fill_8 FILLER_160_1477 ();
 sg13g2_fill_8 FILLER_160_1485 ();
 sg13g2_fill_8 FILLER_160_1493 ();
 sg13g2_fill_8 FILLER_160_1501 ();
 sg13g2_fill_8 FILLER_160_1509 ();
 sg13g2_fill_8 FILLER_160_1517 ();
 sg13g2_fill_8 FILLER_160_1525 ();
 sg13g2_fill_8 FILLER_160_1533 ();
 sg13g2_fill_8 FILLER_160_1541 ();
 sg13g2_fill_8 FILLER_160_1549 ();
 sg13g2_fill_8 FILLER_160_1557 ();
 sg13g2_fill_8 FILLER_160_1565 ();
 sg13g2_fill_8 FILLER_160_1573 ();
 sg13g2_fill_8 FILLER_160_1581 ();
 sg13g2_fill_2 FILLER_160_1589 ();
 sg13g2_fill_1 FILLER_160_1591 ();
 sg13g2_fill_8 FILLER_161_0 ();
 sg13g2_fill_8 FILLER_161_8 ();
 sg13g2_fill_8 FILLER_161_16 ();
 sg13g2_fill_8 FILLER_161_24 ();
 sg13g2_fill_8 FILLER_161_32 ();
 sg13g2_fill_8 FILLER_161_40 ();
 sg13g2_fill_8 FILLER_161_48 ();
 sg13g2_fill_8 FILLER_161_56 ();
 sg13g2_fill_8 FILLER_161_64 ();
 sg13g2_fill_8 FILLER_161_72 ();
 sg13g2_fill_4 FILLER_161_83 ();
 sg13g2_fill_8 FILLER_161_121 ();
 sg13g2_fill_8 FILLER_161_129 ();
 sg13g2_fill_4 FILLER_161_142 ();
 sg13g2_fill_8 FILLER_161_166 ();
 sg13g2_fill_2 FILLER_161_174 ();
 sg13g2_fill_2 FILLER_161_202 ();
 sg13g2_fill_1 FILLER_161_204 ();
 sg13g2_fill_8 FILLER_161_267 ();
 sg13g2_fill_8 FILLER_161_275 ();
 sg13g2_fill_4 FILLER_161_283 ();
 sg13g2_fill_2 FILLER_161_287 ();
 sg13g2_fill_1 FILLER_161_289 ();
 sg13g2_fill_2 FILLER_161_298 ();
 sg13g2_fill_8 FILLER_161_326 ();
 sg13g2_fill_1 FILLER_161_334 ();
 sg13g2_fill_4 FILLER_161_364 ();
 sg13g2_fill_2 FILLER_161_368 ();
 sg13g2_fill_1 FILLER_161_370 ();
 sg13g2_fill_8 FILLER_161_379 ();
 sg13g2_fill_8 FILLER_161_387 ();
 sg13g2_fill_8 FILLER_161_395 ();
 sg13g2_fill_8 FILLER_161_403 ();
 sg13g2_fill_8 FILLER_161_421 ();
 sg13g2_fill_4 FILLER_161_429 ();
 sg13g2_fill_2 FILLER_161_433 ();
 sg13g2_fill_1 FILLER_161_435 ();
 sg13g2_fill_8 FILLER_161_446 ();
 sg13g2_fill_4 FILLER_161_454 ();
 sg13g2_fill_1 FILLER_161_458 ();
 sg13g2_fill_2 FILLER_161_464 ();
 sg13g2_fill_8 FILLER_161_547 ();
 sg13g2_fill_8 FILLER_161_555 ();
 sg13g2_fill_8 FILLER_161_563 ();
 sg13g2_fill_8 FILLER_161_571 ();
 sg13g2_fill_4 FILLER_161_589 ();
 sg13g2_fill_1 FILLER_161_593 ();
 sg13g2_fill_8 FILLER_161_640 ();
 sg13g2_fill_2 FILLER_161_648 ();
 sg13g2_fill_1 FILLER_161_650 ();
 sg13g2_fill_8 FILLER_161_656 ();
 sg13g2_fill_4 FILLER_161_664 ();
 sg13g2_fill_4 FILLER_161_714 ();
 sg13g2_fill_8 FILLER_161_726 ();
 sg13g2_fill_8 FILLER_161_734 ();
 sg13g2_fill_2 FILLER_161_742 ();
 sg13g2_fill_1 FILLER_161_744 ();
 sg13g2_fill_2 FILLER_161_754 ();
 sg13g2_fill_1 FILLER_161_761 ();
 sg13g2_fill_8 FILLER_161_766 ();
 sg13g2_fill_8 FILLER_161_774 ();
 sg13g2_fill_4 FILLER_161_786 ();
 sg13g2_fill_2 FILLER_161_790 ();
 sg13g2_fill_8 FILLER_161_805 ();
 sg13g2_fill_8 FILLER_161_813 ();
 sg13g2_fill_8 FILLER_161_821 ();
 sg13g2_fill_4 FILLER_161_834 ();
 sg13g2_fill_2 FILLER_161_843 ();
 sg13g2_fill_4 FILLER_161_851 ();
 sg13g2_fill_2 FILLER_161_860 ();
 sg13g2_fill_1 FILLER_161_862 ();
 sg13g2_fill_4 FILLER_161_867 ();
 sg13g2_fill_2 FILLER_161_871 ();
 sg13g2_fill_8 FILLER_161_878 ();
 sg13g2_fill_4 FILLER_161_895 ();
 sg13g2_fill_1 FILLER_161_899 ();
 sg13g2_fill_8 FILLER_161_924 ();
 sg13g2_fill_8 FILLER_161_932 ();
 sg13g2_fill_8 FILLER_161_940 ();
 sg13g2_fill_4 FILLER_161_948 ();
 sg13g2_fill_1 FILLER_161_952 ();
 sg13g2_fill_1 FILLER_161_966 ();
 sg13g2_fill_8 FILLER_161_972 ();
 sg13g2_fill_2 FILLER_161_990 ();
 sg13g2_fill_2 FILLER_161_997 ();
 sg13g2_fill_1 FILLER_161_999 ();
 sg13g2_fill_8 FILLER_161_1015 ();
 sg13g2_fill_1 FILLER_161_1023 ();
 sg13g2_fill_2 FILLER_161_1038 ();
 sg13g2_fill_8 FILLER_161_1049 ();
 sg13g2_fill_2 FILLER_161_1057 ();
 sg13g2_fill_1 FILLER_161_1059 ();
 sg13g2_fill_2 FILLER_161_1073 ();
 sg13g2_fill_1 FILLER_161_1075 ();
 sg13g2_fill_2 FILLER_161_1095 ();
 sg13g2_fill_1 FILLER_161_1112 ();
 sg13g2_fill_1 FILLER_161_1125 ();
 sg13g2_fill_1 FILLER_161_1131 ();
 sg13g2_fill_4 FILLER_161_1137 ();
 sg13g2_fill_1 FILLER_161_1141 ();
 sg13g2_fill_2 FILLER_161_1155 ();
 sg13g2_fill_2 FILLER_161_1164 ();
 sg13g2_fill_1 FILLER_161_1166 ();
 sg13g2_fill_4 FILLER_161_1170 ();
 sg13g2_fill_4 FILLER_161_1207 ();
 sg13g2_fill_8 FILLER_161_1229 ();
 sg13g2_fill_4 FILLER_161_1237 ();
 sg13g2_fill_2 FILLER_161_1241 ();
 sg13g2_fill_4 FILLER_161_1261 ();
 sg13g2_fill_1 FILLER_161_1265 ();
 sg13g2_fill_2 FILLER_161_1293 ();
 sg13g2_fill_8 FILLER_161_1319 ();
 sg13g2_fill_8 FILLER_161_1327 ();
 sg13g2_fill_8 FILLER_161_1335 ();
 sg13g2_fill_4 FILLER_161_1343 ();
 sg13g2_fill_2 FILLER_161_1347 ();
 sg13g2_fill_8 FILLER_161_1354 ();
 sg13g2_fill_4 FILLER_161_1362 ();
 sg13g2_fill_2 FILLER_161_1366 ();
 sg13g2_fill_1 FILLER_161_1368 ();
 sg13g2_fill_8 FILLER_161_1377 ();
 sg13g2_fill_4 FILLER_161_1385 ();
 sg13g2_fill_8 FILLER_161_1401 ();
 sg13g2_fill_8 FILLER_161_1409 ();
 sg13g2_fill_8 FILLER_161_1417 ();
 sg13g2_fill_8 FILLER_161_1425 ();
 sg13g2_fill_8 FILLER_161_1458 ();
 sg13g2_fill_8 FILLER_161_1466 ();
 sg13g2_fill_8 FILLER_161_1474 ();
 sg13g2_fill_8 FILLER_161_1482 ();
 sg13g2_fill_8 FILLER_161_1490 ();
 sg13g2_fill_8 FILLER_161_1498 ();
 sg13g2_fill_8 FILLER_161_1506 ();
 sg13g2_fill_8 FILLER_161_1514 ();
 sg13g2_fill_8 FILLER_161_1522 ();
 sg13g2_fill_8 FILLER_161_1530 ();
 sg13g2_fill_8 FILLER_161_1538 ();
 sg13g2_fill_8 FILLER_161_1546 ();
 sg13g2_fill_8 FILLER_161_1554 ();
 sg13g2_fill_8 FILLER_161_1562 ();
 sg13g2_fill_8 FILLER_161_1570 ();
 sg13g2_fill_8 FILLER_161_1578 ();
 sg13g2_fill_4 FILLER_161_1586 ();
 sg13g2_fill_2 FILLER_161_1590 ();
 sg13g2_fill_8 FILLER_162_0 ();
 sg13g2_fill_8 FILLER_162_8 ();
 sg13g2_fill_8 FILLER_162_16 ();
 sg13g2_fill_8 FILLER_162_24 ();
 sg13g2_fill_8 FILLER_162_32 ();
 sg13g2_fill_8 FILLER_162_40 ();
 sg13g2_fill_8 FILLER_162_48 ();
 sg13g2_fill_1 FILLER_162_56 ();
 sg13g2_fill_8 FILLER_162_83 ();
 sg13g2_fill_8 FILLER_162_117 ();
 sg13g2_fill_4 FILLER_162_125 ();
 sg13g2_fill_2 FILLER_162_129 ();
 sg13g2_fill_8 FILLER_162_141 ();
 sg13g2_fill_8 FILLER_162_149 ();
 sg13g2_fill_8 FILLER_162_157 ();
 sg13g2_fill_8 FILLER_162_165 ();
 sg13g2_fill_8 FILLER_162_173 ();
 sg13g2_fill_8 FILLER_162_181 ();
 sg13g2_fill_8 FILLER_162_189 ();
 sg13g2_fill_4 FILLER_162_244 ();
 sg13g2_fill_2 FILLER_162_284 ();
 sg13g2_fill_8 FILLER_162_291 ();
 sg13g2_fill_1 FILLER_162_299 ();
 sg13g2_fill_8 FILLER_162_310 ();
 sg13g2_fill_8 FILLER_162_318 ();
 sg13g2_fill_1 FILLER_162_336 ();
 sg13g2_fill_8 FILLER_162_363 ();
 sg13g2_fill_4 FILLER_162_376 ();
 sg13g2_fill_2 FILLER_162_380 ();
 sg13g2_fill_2 FILLER_162_413 ();
 sg13g2_fill_4 FILLER_162_425 ();
 sg13g2_fill_8 FILLER_162_434 ();
 sg13g2_fill_8 FILLER_162_442 ();
 sg13g2_fill_8 FILLER_162_475 ();
 sg13g2_fill_8 FILLER_162_483 ();
 sg13g2_fill_8 FILLER_162_491 ();
 sg13g2_fill_2 FILLER_162_499 ();
 sg13g2_fill_8 FILLER_162_506 ();
 sg13g2_fill_4 FILLER_162_514 ();
 sg13g2_fill_8 FILLER_162_528 ();
 sg13g2_fill_4 FILLER_162_536 ();
 sg13g2_fill_2 FILLER_162_540 ();
 sg13g2_fill_2 FILLER_162_558 ();
 sg13g2_fill_1 FILLER_162_560 ();
 sg13g2_fill_2 FILLER_162_586 ();
 sg13g2_fill_1 FILLER_162_588 ();
 sg13g2_fill_8 FILLER_162_615 ();
 sg13g2_fill_8 FILLER_162_623 ();
 sg13g2_fill_8 FILLER_162_631 ();
 sg13g2_fill_4 FILLER_162_669 ();
 sg13g2_fill_1 FILLER_162_673 ();
 sg13g2_fill_8 FILLER_162_682 ();
 sg13g2_fill_4 FILLER_162_690 ();
 sg13g2_fill_1 FILLER_162_694 ();
 sg13g2_fill_8 FILLER_162_705 ();
 sg13g2_fill_8 FILLER_162_713 ();
 sg13g2_fill_1 FILLER_162_721 ();
 sg13g2_fill_8 FILLER_162_732 ();
 sg13g2_fill_8 FILLER_162_740 ();
 sg13g2_fill_8 FILLER_162_748 ();
 sg13g2_fill_4 FILLER_162_756 ();
 sg13g2_fill_2 FILLER_162_760 ();
 sg13g2_fill_2 FILLER_162_766 ();
 sg13g2_fill_1 FILLER_162_768 ();
 sg13g2_fill_8 FILLER_162_774 ();
 sg13g2_fill_8 FILLER_162_782 ();
 sg13g2_fill_2 FILLER_162_790 ();
 sg13g2_fill_1 FILLER_162_792 ();
 sg13g2_fill_1 FILLER_162_801 ();
 sg13g2_fill_4 FILLER_162_806 ();
 sg13g2_fill_2 FILLER_162_820 ();
 sg13g2_fill_2 FILLER_162_833 ();
 sg13g2_fill_1 FILLER_162_835 ();
 sg13g2_fill_8 FILLER_162_841 ();
 sg13g2_fill_1 FILLER_162_849 ();
 sg13g2_fill_1 FILLER_162_865 ();
 sg13g2_fill_2 FILLER_162_880 ();
 sg13g2_fill_1 FILLER_162_882 ();
 sg13g2_fill_2 FILLER_162_904 ();
 sg13g2_fill_2 FILLER_162_910 ();
 sg13g2_fill_1 FILLER_162_912 ();
 sg13g2_fill_8 FILLER_162_918 ();
 sg13g2_fill_8 FILLER_162_926 ();
 sg13g2_fill_8 FILLER_162_934 ();
 sg13g2_fill_4 FILLER_162_942 ();
 sg13g2_fill_2 FILLER_162_946 ();
 sg13g2_fill_1 FILLER_162_948 ();
 sg13g2_fill_4 FILLER_162_974 ();
 sg13g2_fill_1 FILLER_162_978 ();
 sg13g2_fill_4 FILLER_162_1014 ();
 sg13g2_fill_1 FILLER_162_1018 ();
 sg13g2_fill_8 FILLER_162_1056 ();
 sg13g2_fill_8 FILLER_162_1064 ();
 sg13g2_fill_8 FILLER_162_1072 ();
 sg13g2_fill_1 FILLER_162_1080 ();
 sg13g2_fill_4 FILLER_162_1086 ();
 sg13g2_fill_1 FILLER_162_1090 ();
 sg13g2_fill_4 FILLER_162_1096 ();
 sg13g2_fill_1 FILLER_162_1100 ();
 sg13g2_fill_2 FILLER_162_1109 ();
 sg13g2_fill_8 FILLER_162_1116 ();
 sg13g2_fill_4 FILLER_162_1124 ();
 sg13g2_fill_2 FILLER_162_1128 ();
 sg13g2_fill_8 FILLER_162_1135 ();
 sg13g2_fill_8 FILLER_162_1143 ();
 sg13g2_fill_4 FILLER_162_1151 ();
 sg13g2_fill_2 FILLER_162_1155 ();
 sg13g2_fill_1 FILLER_162_1157 ();
 sg13g2_fill_1 FILLER_162_1163 ();
 sg13g2_fill_8 FILLER_162_1174 ();
 sg13g2_fill_8 FILLER_162_1182 ();
 sg13g2_fill_2 FILLER_162_1190 ();
 sg13g2_fill_1 FILLER_162_1192 ();
 sg13g2_fill_8 FILLER_162_1199 ();
 sg13g2_fill_2 FILLER_162_1207 ();
 sg13g2_fill_1 FILLER_162_1209 ();
 sg13g2_fill_1 FILLER_162_1217 ();
 sg13g2_fill_4 FILLER_162_1225 ();
 sg13g2_fill_1 FILLER_162_1237 ();
 sg13g2_fill_8 FILLER_162_1258 ();
 sg13g2_fill_2 FILLER_162_1266 ();
 sg13g2_fill_1 FILLER_162_1268 ();
 sg13g2_fill_1 FILLER_162_1272 ();
 sg13g2_fill_1 FILLER_162_1301 ();
 sg13g2_fill_1 FILLER_162_1306 ();
 sg13g2_fill_1 FILLER_162_1328 ();
 sg13g2_fill_8 FILLER_162_1371 ();
 sg13g2_fill_8 FILLER_162_1379 ();
 sg13g2_fill_2 FILLER_162_1387 ();
 sg13g2_fill_4 FILLER_162_1401 ();
 sg13g2_fill_8 FILLER_162_1417 ();
 sg13g2_fill_8 FILLER_162_1425 ();
 sg13g2_fill_4 FILLER_162_1433 ();
 sg13g2_fill_2 FILLER_162_1437 ();
 sg13g2_fill_1 FILLER_162_1439 ();
 sg13g2_fill_8 FILLER_162_1444 ();
 sg13g2_fill_8 FILLER_162_1452 ();
 sg13g2_fill_8 FILLER_162_1460 ();
 sg13g2_fill_8 FILLER_162_1468 ();
 sg13g2_fill_8 FILLER_162_1476 ();
 sg13g2_fill_8 FILLER_162_1484 ();
 sg13g2_fill_8 FILLER_162_1492 ();
 sg13g2_fill_8 FILLER_162_1500 ();
 sg13g2_fill_8 FILLER_162_1508 ();
 sg13g2_fill_8 FILLER_162_1516 ();
 sg13g2_fill_8 FILLER_162_1524 ();
 sg13g2_fill_8 FILLER_162_1532 ();
 sg13g2_fill_8 FILLER_162_1540 ();
 sg13g2_fill_8 FILLER_162_1548 ();
 sg13g2_fill_8 FILLER_162_1556 ();
 sg13g2_fill_8 FILLER_162_1564 ();
 sg13g2_fill_8 FILLER_162_1572 ();
 sg13g2_fill_8 FILLER_162_1580 ();
 sg13g2_fill_4 FILLER_162_1588 ();
 sg13g2_fill_8 FILLER_163_0 ();
 sg13g2_fill_8 FILLER_163_8 ();
 sg13g2_fill_8 FILLER_163_16 ();
 sg13g2_fill_8 FILLER_163_24 ();
 sg13g2_fill_8 FILLER_163_32 ();
 sg13g2_fill_8 FILLER_163_40 ();
 sg13g2_fill_4 FILLER_163_48 ();
 sg13g2_fill_2 FILLER_163_52 ();
 sg13g2_fill_1 FILLER_163_54 ();
 sg13g2_fill_8 FILLER_163_65 ();
 sg13g2_fill_4 FILLER_163_73 ();
 sg13g2_fill_1 FILLER_163_77 ();
 sg13g2_fill_8 FILLER_163_88 ();
 sg13g2_fill_2 FILLER_163_96 ();
 sg13g2_fill_2 FILLER_163_150 ();
 sg13g2_fill_1 FILLER_163_152 ();
 sg13g2_fill_8 FILLER_163_161 ();
 sg13g2_fill_4 FILLER_163_169 ();
 sg13g2_fill_2 FILLER_163_173 ();
 sg13g2_fill_1 FILLER_163_175 ();
 sg13g2_fill_8 FILLER_163_181 ();
 sg13g2_fill_4 FILLER_163_189 ();
 sg13g2_fill_2 FILLER_163_193 ();
 sg13g2_fill_1 FILLER_163_195 ();
 sg13g2_fill_8 FILLER_163_206 ();
 sg13g2_fill_8 FILLER_163_214 ();
 sg13g2_fill_8 FILLER_163_222 ();
 sg13g2_fill_8 FILLER_163_230 ();
 sg13g2_fill_2 FILLER_163_238 ();
 sg13g2_fill_4 FILLER_163_263 ();
 sg13g2_fill_2 FILLER_163_267 ();
 sg13g2_fill_8 FILLER_163_290 ();
 sg13g2_fill_2 FILLER_163_324 ();
 sg13g2_fill_2 FILLER_163_347 ();
 sg13g2_fill_1 FILLER_163_349 ();
 sg13g2_fill_4 FILLER_163_396 ();
 sg13g2_fill_1 FILLER_163_400 ();
 sg13g2_fill_2 FILLER_163_427 ();
 sg13g2_fill_1 FILLER_163_446 ();
 sg13g2_fill_2 FILLER_163_475 ();
 sg13g2_fill_1 FILLER_163_477 ();
 sg13g2_fill_2 FILLER_163_488 ();
 sg13g2_fill_2 FILLER_163_500 ();
 sg13g2_fill_2 FILLER_163_510 ();
 sg13g2_fill_8 FILLER_163_522 ();
 sg13g2_fill_8 FILLER_163_530 ();
 sg13g2_fill_2 FILLER_163_538 ();
 sg13g2_fill_4 FILLER_163_545 ();
 sg13g2_fill_2 FILLER_163_559 ();
 sg13g2_fill_2 FILLER_163_595 ();
 sg13g2_fill_1 FILLER_163_597 ();
 sg13g2_fill_8 FILLER_163_606 ();
 sg13g2_fill_8 FILLER_163_614 ();
 sg13g2_fill_8 FILLER_163_622 ();
 sg13g2_fill_2 FILLER_163_665 ();
 sg13g2_fill_1 FILLER_163_667 ();
 sg13g2_fill_4 FILLER_163_694 ();
 sg13g2_fill_2 FILLER_163_698 ();
 sg13g2_fill_1 FILLER_163_726 ();
 sg13g2_fill_1 FILLER_163_753 ();
 sg13g2_fill_2 FILLER_163_781 ();
 sg13g2_fill_1 FILLER_163_788 ();
 sg13g2_fill_8 FILLER_163_794 ();
 sg13g2_fill_4 FILLER_163_802 ();
 sg13g2_fill_2 FILLER_163_806 ();
 sg13g2_fill_8 FILLER_163_830 ();
 sg13g2_fill_2 FILLER_163_838 ();
 sg13g2_fill_1 FILLER_163_840 ();
 sg13g2_fill_2 FILLER_163_846 ();
 sg13g2_fill_1 FILLER_163_869 ();
 sg13g2_fill_1 FILLER_163_875 ();
 sg13g2_fill_2 FILLER_163_880 ();
 sg13g2_fill_1 FILLER_163_882 ();
 sg13g2_fill_8 FILLER_163_896 ();
 sg13g2_fill_4 FILLER_163_904 ();
 sg13g2_fill_1 FILLER_163_912 ();
 sg13g2_fill_8 FILLER_163_923 ();
 sg13g2_fill_8 FILLER_163_931 ();
 sg13g2_fill_8 FILLER_163_939 ();
 sg13g2_fill_8 FILLER_163_947 ();
 sg13g2_fill_1 FILLER_163_955 ();
 sg13g2_fill_8 FILLER_163_970 ();
 sg13g2_fill_8 FILLER_163_978 ();
 sg13g2_fill_8 FILLER_163_986 ();
 sg13g2_fill_2 FILLER_163_994 ();
 sg13g2_fill_8 FILLER_163_1007 ();
 sg13g2_fill_4 FILLER_163_1015 ();
 sg13g2_fill_2 FILLER_163_1019 ();
 sg13g2_fill_1 FILLER_163_1021 ();
 sg13g2_fill_2 FILLER_163_1038 ();
 sg13g2_fill_1 FILLER_163_1040 ();
 sg13g2_fill_8 FILLER_163_1057 ();
 sg13g2_fill_8 FILLER_163_1065 ();
 sg13g2_fill_8 FILLER_163_1108 ();
 sg13g2_fill_8 FILLER_163_1116 ();
 sg13g2_fill_4 FILLER_163_1144 ();
 sg13g2_fill_1 FILLER_163_1148 ();
 sg13g2_fill_2 FILLER_163_1161 ();
 sg13g2_fill_4 FILLER_163_1173 ();
 sg13g2_fill_2 FILLER_163_1185 ();
 sg13g2_fill_8 FILLER_163_1192 ();
 sg13g2_fill_8 FILLER_163_1200 ();
 sg13g2_fill_4 FILLER_163_1208 ();
 sg13g2_fill_1 FILLER_163_1212 ();
 sg13g2_fill_2 FILLER_163_1218 ();
 sg13g2_fill_1 FILLER_163_1220 ();
 sg13g2_fill_4 FILLER_163_1232 ();
 sg13g2_fill_2 FILLER_163_1236 ();
 sg13g2_fill_8 FILLER_163_1246 ();
 sg13g2_fill_2 FILLER_163_1254 ();
 sg13g2_fill_1 FILLER_163_1256 ();
 sg13g2_fill_8 FILLER_163_1280 ();
 sg13g2_fill_8 FILLER_163_1288 ();
 sg13g2_fill_2 FILLER_163_1296 ();
 sg13g2_fill_1 FILLER_163_1298 ();
 sg13g2_fill_8 FILLER_163_1307 ();
 sg13g2_fill_8 FILLER_163_1320 ();
 sg13g2_fill_4 FILLER_163_1328 ();
 sg13g2_fill_2 FILLER_163_1332 ();
 sg13g2_fill_2 FILLER_163_1346 ();
 sg13g2_fill_1 FILLER_163_1348 ();
 sg13g2_fill_1 FILLER_163_1379 ();
 sg13g2_fill_2 FILLER_163_1396 ();
 sg13g2_fill_4 FILLER_163_1435 ();
 sg13g2_fill_2 FILLER_163_1439 ();
 sg13g2_fill_8 FILLER_163_1453 ();
 sg13g2_fill_8 FILLER_163_1461 ();
 sg13g2_fill_8 FILLER_163_1469 ();
 sg13g2_fill_8 FILLER_163_1477 ();
 sg13g2_fill_8 FILLER_163_1485 ();
 sg13g2_fill_8 FILLER_163_1493 ();
 sg13g2_fill_8 FILLER_163_1501 ();
 sg13g2_fill_8 FILLER_163_1509 ();
 sg13g2_fill_8 FILLER_163_1517 ();
 sg13g2_fill_8 FILLER_163_1525 ();
 sg13g2_fill_8 FILLER_163_1533 ();
 sg13g2_fill_8 FILLER_163_1541 ();
 sg13g2_fill_8 FILLER_163_1549 ();
 sg13g2_fill_8 FILLER_163_1557 ();
 sg13g2_fill_8 FILLER_163_1565 ();
 sg13g2_fill_8 FILLER_163_1573 ();
 sg13g2_fill_8 FILLER_163_1581 ();
 sg13g2_fill_2 FILLER_163_1589 ();
 sg13g2_fill_1 FILLER_163_1591 ();
 sg13g2_fill_8 FILLER_164_0 ();
 sg13g2_fill_8 FILLER_164_8 ();
 sg13g2_fill_8 FILLER_164_16 ();
 sg13g2_fill_8 FILLER_164_24 ();
 sg13g2_fill_8 FILLER_164_32 ();
 sg13g2_fill_8 FILLER_164_40 ();
 sg13g2_fill_2 FILLER_164_48 ();
 sg13g2_fill_1 FILLER_164_50 ();
 sg13g2_fill_1 FILLER_164_77 ();
 sg13g2_fill_8 FILLER_164_100 ();
 sg13g2_fill_8 FILLER_164_108 ();
 sg13g2_fill_4 FILLER_164_116 ();
 sg13g2_fill_2 FILLER_164_120 ();
 sg13g2_fill_1 FILLER_164_122 ();
 sg13g2_fill_2 FILLER_164_133 ();
 sg13g2_fill_4 FILLER_164_151 ();
 sg13g2_fill_8 FILLER_164_210 ();
 sg13g2_fill_1 FILLER_164_218 ();
 sg13g2_fill_8 FILLER_164_229 ();
 sg13g2_fill_4 FILLER_164_237 ();
 sg13g2_fill_2 FILLER_164_241 ();
 sg13g2_fill_1 FILLER_164_243 ();
 sg13g2_fill_1 FILLER_164_270 ();
 sg13g2_fill_2 FILLER_164_292 ();
 sg13g2_fill_1 FILLER_164_294 ();
 sg13g2_fill_8 FILLER_164_360 ();
 sg13g2_fill_4 FILLER_164_368 ();
 sg13g2_fill_1 FILLER_164_372 ();
 sg13g2_fill_8 FILLER_164_378 ();
 sg13g2_fill_8 FILLER_164_386 ();
 sg13g2_fill_8 FILLER_164_394 ();
 sg13g2_fill_8 FILLER_164_402 ();
 sg13g2_fill_8 FILLER_164_410 ();
 sg13g2_fill_8 FILLER_164_418 ();
 sg13g2_fill_4 FILLER_164_426 ();
 sg13g2_fill_1 FILLER_164_440 ();
 sg13g2_fill_2 FILLER_164_454 ();
 sg13g2_fill_1 FILLER_164_456 ();
 sg13g2_fill_2 FILLER_164_489 ();
 sg13g2_fill_1 FILLER_164_491 ();
 sg13g2_fill_8 FILLER_164_551 ();
 sg13g2_fill_8 FILLER_164_559 ();
 sg13g2_fill_4 FILLER_164_567 ();
 sg13g2_fill_1 FILLER_164_571 ();
 sg13g2_fill_8 FILLER_164_588 ();
 sg13g2_fill_8 FILLER_164_596 ();
 sg13g2_fill_8 FILLER_164_604 ();
 sg13g2_fill_8 FILLER_164_612 ();
 sg13g2_fill_1 FILLER_164_620 ();
 sg13g2_fill_2 FILLER_164_655 ();
 sg13g2_fill_1 FILLER_164_657 ();
 sg13g2_fill_8 FILLER_164_668 ();
 sg13g2_fill_8 FILLER_164_676 ();
 sg13g2_fill_4 FILLER_164_684 ();
 sg13g2_fill_1 FILLER_164_698 ();
 sg13g2_fill_8 FILLER_164_724 ();
 sg13g2_fill_8 FILLER_164_752 ();
 sg13g2_fill_2 FILLER_164_760 ();
 sg13g2_fill_8 FILLER_164_767 ();
 sg13g2_fill_2 FILLER_164_775 ();
 sg13g2_fill_4 FILLER_164_810 ();
 sg13g2_fill_2 FILLER_164_814 ();
 sg13g2_fill_8 FILLER_164_821 ();
 sg13g2_fill_4 FILLER_164_829 ();
 sg13g2_fill_2 FILLER_164_839 ();
 sg13g2_fill_1 FILLER_164_841 ();
 sg13g2_fill_8 FILLER_164_861 ();
 sg13g2_fill_8 FILLER_164_869 ();
 sg13g2_fill_1 FILLER_164_877 ();
 sg13g2_fill_8 FILLER_164_888 ();
 sg13g2_fill_4 FILLER_164_896 ();
 sg13g2_fill_2 FILLER_164_900 ();
 sg13g2_fill_8 FILLER_164_915 ();
 sg13g2_fill_8 FILLER_164_923 ();
 sg13g2_fill_8 FILLER_164_931 ();
 sg13g2_fill_8 FILLER_164_939 ();
 sg13g2_fill_8 FILLER_164_947 ();
 sg13g2_fill_2 FILLER_164_955 ();
 sg13g2_fill_4 FILLER_164_973 ();
 sg13g2_fill_1 FILLER_164_977 ();
 sg13g2_fill_8 FILLER_164_981 ();
 sg13g2_fill_1 FILLER_164_989 ();
 sg13g2_fill_8 FILLER_164_1008 ();
 sg13g2_fill_8 FILLER_164_1016 ();
 sg13g2_fill_4 FILLER_164_1024 ();
 sg13g2_fill_2 FILLER_164_1028 ();
 sg13g2_fill_4 FILLER_164_1039 ();
 sg13g2_fill_2 FILLER_164_1043 ();
 sg13g2_fill_4 FILLER_164_1050 ();
 sg13g2_fill_2 FILLER_164_1054 ();
 sg13g2_fill_1 FILLER_164_1056 ();
 sg13g2_fill_4 FILLER_164_1073 ();
 sg13g2_fill_2 FILLER_164_1077 ();
 sg13g2_fill_1 FILLER_164_1087 ();
 sg13g2_fill_1 FILLER_164_1092 ();
 sg13g2_fill_2 FILLER_164_1107 ();
 sg13g2_fill_1 FILLER_164_1109 ();
 sg13g2_fill_1 FILLER_164_1118 ();
 sg13g2_fill_2 FILLER_164_1124 ();
 sg13g2_fill_4 FILLER_164_1139 ();
 sg13g2_fill_2 FILLER_164_1143 ();
 sg13g2_fill_1 FILLER_164_1145 ();
 sg13g2_fill_4 FILLER_164_1189 ();
 sg13g2_fill_1 FILLER_164_1193 ();
 sg13g2_fill_1 FILLER_164_1199 ();
 sg13g2_fill_4 FILLER_164_1204 ();
 sg13g2_fill_2 FILLER_164_1208 ();
 sg13g2_fill_1 FILLER_164_1210 ();
 sg13g2_fill_8 FILLER_164_1220 ();
 sg13g2_fill_8 FILLER_164_1228 ();
 sg13g2_fill_8 FILLER_164_1236 ();
 sg13g2_fill_2 FILLER_164_1244 ();
 sg13g2_fill_1 FILLER_164_1246 ();
 sg13g2_fill_8 FILLER_164_1255 ();
 sg13g2_fill_8 FILLER_164_1263 ();
 sg13g2_fill_8 FILLER_164_1279 ();
 sg13g2_fill_2 FILLER_164_1287 ();
 sg13g2_fill_1 FILLER_164_1289 ();
 sg13g2_fill_2 FILLER_164_1298 ();
 sg13g2_fill_1 FILLER_164_1300 ();
 sg13g2_fill_8 FILLER_164_1305 ();
 sg13g2_fill_2 FILLER_164_1313 ();
 sg13g2_fill_1 FILLER_164_1315 ();
 sg13g2_fill_4 FILLER_164_1331 ();
 sg13g2_fill_2 FILLER_164_1340 ();
 sg13g2_fill_1 FILLER_164_1353 ();
 sg13g2_fill_2 FILLER_164_1375 ();
 sg13g2_fill_8 FILLER_164_1391 ();
 sg13g2_fill_8 FILLER_164_1399 ();
 sg13g2_fill_2 FILLER_164_1407 ();
 sg13g2_fill_1 FILLER_164_1409 ();
 sg13g2_fill_1 FILLER_164_1415 ();
 sg13g2_fill_8 FILLER_164_1456 ();
 sg13g2_fill_8 FILLER_164_1464 ();
 sg13g2_fill_8 FILLER_164_1472 ();
 sg13g2_fill_8 FILLER_164_1480 ();
 sg13g2_fill_8 FILLER_164_1488 ();
 sg13g2_fill_8 FILLER_164_1496 ();
 sg13g2_fill_8 FILLER_164_1504 ();
 sg13g2_fill_8 FILLER_164_1512 ();
 sg13g2_fill_8 FILLER_164_1520 ();
 sg13g2_fill_8 FILLER_164_1528 ();
 sg13g2_fill_8 FILLER_164_1536 ();
 sg13g2_fill_8 FILLER_164_1544 ();
 sg13g2_fill_8 FILLER_164_1552 ();
 sg13g2_fill_8 FILLER_164_1560 ();
 sg13g2_fill_8 FILLER_164_1568 ();
 sg13g2_fill_8 FILLER_164_1576 ();
 sg13g2_fill_8 FILLER_164_1584 ();
 sg13g2_fill_8 FILLER_165_0 ();
 sg13g2_fill_8 FILLER_165_8 ();
 sg13g2_fill_8 FILLER_165_16 ();
 sg13g2_fill_8 FILLER_165_24 ();
 sg13g2_fill_8 FILLER_165_32 ();
 sg13g2_fill_8 FILLER_165_40 ();
 sg13g2_fill_4 FILLER_165_48 ();
 sg13g2_fill_2 FILLER_165_52 ();
 sg13g2_fill_8 FILLER_165_64 ();
 sg13g2_fill_2 FILLER_165_72 ();
 sg13g2_fill_1 FILLER_165_74 ();
 sg13g2_fill_8 FILLER_165_85 ();
 sg13g2_fill_8 FILLER_165_93 ();
 sg13g2_fill_8 FILLER_165_101 ();
 sg13g2_fill_8 FILLER_165_109 ();
 sg13g2_fill_8 FILLER_165_117 ();
 sg13g2_fill_8 FILLER_165_125 ();
 sg13g2_fill_2 FILLER_165_133 ();
 sg13g2_fill_4 FILLER_165_145 ();
 sg13g2_fill_2 FILLER_165_169 ();
 sg13g2_fill_8 FILLER_165_179 ();
 sg13g2_fill_8 FILLER_165_187 ();
 sg13g2_fill_8 FILLER_165_205 ();
 sg13g2_fill_8 FILLER_165_239 ();
 sg13g2_fill_2 FILLER_165_247 ();
 sg13g2_fill_1 FILLER_165_249 ();
 sg13g2_fill_8 FILLER_165_285 ();
 sg13g2_fill_8 FILLER_165_293 ();
 sg13g2_fill_8 FILLER_165_301 ();
 sg13g2_fill_8 FILLER_165_309 ();
 sg13g2_fill_8 FILLER_165_317 ();
 sg13g2_fill_8 FILLER_165_325 ();
 sg13g2_fill_8 FILLER_165_333 ();
 sg13g2_fill_8 FILLER_165_341 ();
 sg13g2_fill_8 FILLER_165_349 ();
 sg13g2_fill_2 FILLER_165_357 ();
 sg13g2_fill_1 FILLER_165_369 ();
 sg13g2_fill_2 FILLER_165_376 ();
 sg13g2_fill_1 FILLER_165_378 ();
 sg13g2_fill_4 FILLER_165_389 ();
 sg13g2_fill_8 FILLER_165_399 ();
 sg13g2_fill_4 FILLER_165_407 ();
 sg13g2_fill_1 FILLER_165_411 ();
 sg13g2_fill_8 FILLER_165_422 ();
 sg13g2_fill_8 FILLER_165_430 ();
 sg13g2_fill_8 FILLER_165_444 ();
 sg13g2_fill_8 FILLER_165_452 ();
 sg13g2_fill_8 FILLER_165_460 ();
 sg13g2_fill_8 FILLER_165_468 ();
 sg13g2_fill_1 FILLER_165_476 ();
 sg13g2_fill_8 FILLER_165_487 ();
 sg13g2_fill_8 FILLER_165_495 ();
 sg13g2_fill_8 FILLER_165_503 ();
 sg13g2_fill_8 FILLER_165_511 ();
 sg13g2_fill_8 FILLER_165_519 ();
 sg13g2_fill_2 FILLER_165_527 ();
 sg13g2_fill_1 FILLER_165_529 ();
 sg13g2_fill_4 FILLER_165_535 ();
 sg13g2_fill_2 FILLER_165_539 ();
 sg13g2_fill_1 FILLER_165_551 ();
 sg13g2_fill_1 FILLER_165_588 ();
 sg13g2_fill_4 FILLER_165_645 ();
 sg13g2_fill_2 FILLER_165_649 ();
 sg13g2_fill_1 FILLER_165_651 ();
 sg13g2_fill_4 FILLER_165_675 ();
 sg13g2_fill_2 FILLER_165_679 ();
 sg13g2_fill_1 FILLER_165_681 ();
 sg13g2_fill_4 FILLER_165_728 ();
 sg13g2_fill_8 FILLER_165_742 ();
 sg13g2_fill_8 FILLER_165_750 ();
 sg13g2_fill_8 FILLER_165_758 ();
 sg13g2_fill_2 FILLER_165_766 ();
 sg13g2_fill_1 FILLER_165_768 ();
 sg13g2_fill_8 FILLER_165_777 ();
 sg13g2_fill_2 FILLER_165_785 ();
 sg13g2_fill_1 FILLER_165_787 ();
 sg13g2_fill_1 FILLER_165_792 ();
 sg13g2_fill_8 FILLER_165_798 ();
 sg13g2_fill_8 FILLER_165_806 ();
 sg13g2_fill_1 FILLER_165_814 ();
 sg13g2_fill_1 FILLER_165_826 ();
 sg13g2_fill_1 FILLER_165_840 ();
 sg13g2_fill_2 FILLER_165_845 ();
 sg13g2_fill_2 FILLER_165_852 ();
 sg13g2_fill_1 FILLER_165_854 ();
 sg13g2_fill_4 FILLER_165_860 ();
 sg13g2_fill_1 FILLER_165_864 ();
 sg13g2_fill_2 FILLER_165_870 ();
 sg13g2_fill_8 FILLER_165_915 ();
 sg13g2_fill_8 FILLER_165_923 ();
 sg13g2_fill_8 FILLER_165_931 ();
 sg13g2_fill_8 FILLER_165_939 ();
 sg13g2_fill_8 FILLER_165_947 ();
 sg13g2_fill_8 FILLER_165_955 ();
 sg13g2_fill_8 FILLER_165_963 ();
 sg13g2_fill_2 FILLER_165_971 ();
 sg13g2_fill_4 FILLER_165_983 ();
 sg13g2_fill_1 FILLER_165_987 ();
 sg13g2_fill_8 FILLER_165_1008 ();
 sg13g2_fill_2 FILLER_165_1016 ();
 sg13g2_fill_1 FILLER_165_1018 ();
 sg13g2_fill_8 FILLER_165_1077 ();
 sg13g2_fill_8 FILLER_165_1085 ();
 sg13g2_fill_8 FILLER_165_1097 ();
 sg13g2_fill_8 FILLER_165_1105 ();
 sg13g2_fill_8 FILLER_165_1113 ();
 sg13g2_fill_8 FILLER_165_1121 ();
 sg13g2_fill_2 FILLER_165_1129 ();
 sg13g2_fill_8 FILLER_165_1136 ();
 sg13g2_fill_1 FILLER_165_1144 ();
 sg13g2_fill_8 FILLER_165_1154 ();
 sg13g2_fill_8 FILLER_165_1162 ();
 sg13g2_fill_4 FILLER_165_1170 ();
 sg13g2_fill_2 FILLER_165_1174 ();
 sg13g2_fill_1 FILLER_165_1176 ();
 sg13g2_fill_2 FILLER_165_1182 ();
 sg13g2_fill_2 FILLER_165_1196 ();
 sg13g2_fill_4 FILLER_165_1215 ();
 sg13g2_fill_8 FILLER_165_1236 ();
 sg13g2_fill_1 FILLER_165_1244 ();
 sg13g2_fill_4 FILLER_165_1266 ();
 sg13g2_fill_1 FILLER_165_1270 ();
 sg13g2_fill_2 FILLER_165_1310 ();
 sg13g2_fill_1 FILLER_165_1317 ();
 sg13g2_fill_4 FILLER_165_1330 ();
 sg13g2_fill_1 FILLER_165_1334 ();
 sg13g2_fill_8 FILLER_165_1346 ();
 sg13g2_fill_4 FILLER_165_1354 ();
 sg13g2_fill_2 FILLER_165_1358 ();
 sg13g2_fill_1 FILLER_165_1360 ();
 sg13g2_fill_2 FILLER_165_1374 ();
 sg13g2_fill_8 FILLER_165_1381 ();
 sg13g2_fill_8 FILLER_165_1389 ();
 sg13g2_fill_8 FILLER_165_1397 ();
 sg13g2_fill_8 FILLER_165_1405 ();
 sg13g2_fill_8 FILLER_165_1431 ();
 sg13g2_fill_8 FILLER_165_1450 ();
 sg13g2_fill_8 FILLER_165_1458 ();
 sg13g2_fill_8 FILLER_165_1466 ();
 sg13g2_fill_8 FILLER_165_1474 ();
 sg13g2_fill_8 FILLER_165_1482 ();
 sg13g2_fill_8 FILLER_165_1490 ();
 sg13g2_fill_8 FILLER_165_1498 ();
 sg13g2_fill_8 FILLER_165_1506 ();
 sg13g2_fill_8 FILLER_165_1514 ();
 sg13g2_fill_8 FILLER_165_1522 ();
 sg13g2_fill_8 FILLER_165_1530 ();
 sg13g2_fill_8 FILLER_165_1538 ();
 sg13g2_fill_8 FILLER_165_1546 ();
 sg13g2_fill_8 FILLER_165_1554 ();
 sg13g2_fill_8 FILLER_165_1562 ();
 sg13g2_fill_8 FILLER_165_1570 ();
 sg13g2_fill_8 FILLER_165_1578 ();
 sg13g2_fill_4 FILLER_165_1586 ();
 sg13g2_fill_2 FILLER_165_1590 ();
 sg13g2_fill_8 FILLER_166_0 ();
 sg13g2_fill_8 FILLER_166_8 ();
 sg13g2_fill_8 FILLER_166_16 ();
 sg13g2_fill_8 FILLER_166_24 ();
 sg13g2_fill_8 FILLER_166_32 ();
 sg13g2_fill_8 FILLER_166_40 ();
 sg13g2_fill_2 FILLER_166_48 ();
 sg13g2_fill_1 FILLER_166_76 ();
 sg13g2_fill_4 FILLER_166_87 ();
 sg13g2_fill_2 FILLER_166_91 ();
 sg13g2_fill_4 FILLER_166_129 ();
 sg13g2_fill_1 FILLER_166_133 ();
 sg13g2_fill_4 FILLER_166_194 ();
 sg13g2_fill_2 FILLER_166_198 ();
 sg13g2_fill_1 FILLER_166_200 ();
 sg13g2_fill_8 FILLER_166_221 ();
 sg13g2_fill_8 FILLER_166_229 ();
 sg13g2_fill_2 FILLER_166_237 ();
 sg13g2_fill_4 FILLER_166_275 ();
 sg13g2_fill_8 FILLER_166_305 ();
 sg13g2_fill_8 FILLER_166_313 ();
 sg13g2_fill_2 FILLER_166_321 ();
 sg13g2_fill_1 FILLER_166_323 ();
 sg13g2_fill_2 FILLER_166_350 ();
 sg13g2_fill_8 FILLER_166_362 ();
 sg13g2_fill_8 FILLER_166_370 ();
 sg13g2_fill_2 FILLER_166_378 ();
 sg13g2_fill_2 FILLER_166_390 ();
 sg13g2_fill_1 FILLER_166_392 ();
 sg13g2_fill_2 FILLER_166_408 ();
 sg13g2_fill_4 FILLER_166_436 ();
 sg13g2_fill_4 FILLER_166_450 ();
 sg13g2_fill_2 FILLER_166_454 ();
 sg13g2_fill_8 FILLER_166_466 ();
 sg13g2_fill_2 FILLER_166_474 ();
 sg13g2_fill_1 FILLER_166_476 ();
 sg13g2_fill_8 FILLER_166_493 ();
 sg13g2_fill_1 FILLER_166_501 ();
 sg13g2_fill_8 FILLER_166_507 ();
 sg13g2_fill_8 FILLER_166_515 ();
 sg13g2_fill_4 FILLER_166_523 ();
 sg13g2_fill_8 FILLER_166_580 ();
 sg13g2_fill_4 FILLER_166_588 ();
 sg13g2_fill_2 FILLER_166_592 ();
 sg13g2_fill_8 FILLER_166_599 ();
 sg13g2_fill_8 FILLER_166_607 ();
 sg13g2_fill_1 FILLER_166_615 ();
 sg13g2_fill_8 FILLER_166_626 ();
 sg13g2_fill_8 FILLER_166_634 ();
 sg13g2_fill_8 FILLER_166_642 ();
 sg13g2_fill_4 FILLER_166_650 ();
 sg13g2_fill_1 FILLER_166_654 ();
 sg13g2_fill_4 FILLER_166_663 ();
 sg13g2_fill_1 FILLER_166_667 ();
 sg13g2_fill_4 FILLER_166_694 ();
 sg13g2_fill_1 FILLER_166_698 ();
 sg13g2_fill_8 FILLER_166_724 ();
 sg13g2_fill_2 FILLER_166_732 ();
 sg13g2_fill_2 FILLER_166_754 ();
 sg13g2_fill_4 FILLER_166_760 ();
 sg13g2_fill_1 FILLER_166_764 ();
 sg13g2_fill_1 FILLER_166_781 ();
 sg13g2_fill_2 FILLER_166_786 ();
 sg13g2_fill_1 FILLER_166_788 ();
 sg13g2_fill_4 FILLER_166_794 ();
 sg13g2_fill_2 FILLER_166_798 ();
 sg13g2_fill_1 FILLER_166_800 ();
 sg13g2_fill_2 FILLER_166_814 ();
 sg13g2_fill_4 FILLER_166_821 ();
 sg13g2_fill_8 FILLER_166_839 ();
 sg13g2_fill_8 FILLER_166_853 ();
 sg13g2_fill_4 FILLER_166_861 ();
 sg13g2_fill_1 FILLER_166_865 ();
 sg13g2_fill_4 FILLER_166_871 ();
 sg13g2_fill_1 FILLER_166_875 ();
 sg13g2_fill_4 FILLER_166_886 ();
 sg13g2_fill_2 FILLER_166_890 ();
 sg13g2_fill_1 FILLER_166_892 ();
 sg13g2_fill_4 FILLER_166_897 ();
 sg13g2_fill_1 FILLER_166_901 ();
 sg13g2_fill_2 FILLER_166_908 ();
 sg13g2_fill_8 FILLER_166_919 ();
 sg13g2_fill_8 FILLER_166_927 ();
 sg13g2_fill_8 FILLER_166_935 ();
 sg13g2_fill_8 FILLER_166_943 ();
 sg13g2_fill_8 FILLER_166_951 ();
 sg13g2_fill_2 FILLER_166_959 ();
 sg13g2_fill_1 FILLER_166_981 ();
 sg13g2_fill_1 FILLER_166_987 ();
 sg13g2_fill_1 FILLER_166_993 ();
 sg13g2_fill_8 FILLER_166_1002 ();
 sg13g2_fill_4 FILLER_166_1010 ();
 sg13g2_fill_1 FILLER_166_1014 ();
 sg13g2_fill_1 FILLER_166_1035 ();
 sg13g2_fill_2 FILLER_166_1043 ();
 sg13g2_fill_8 FILLER_166_1049 ();
 sg13g2_fill_4 FILLER_166_1057 ();
 sg13g2_fill_2 FILLER_166_1061 ();
 sg13g2_fill_1 FILLER_166_1063 ();
 sg13g2_fill_8 FILLER_166_1068 ();
 sg13g2_fill_8 FILLER_166_1076 ();
 sg13g2_fill_4 FILLER_166_1084 ();
 sg13g2_fill_1 FILLER_166_1088 ();
 sg13g2_fill_4 FILLER_166_1094 ();
 sg13g2_fill_1 FILLER_166_1110 ();
 sg13g2_fill_8 FILLER_166_1116 ();
 sg13g2_fill_2 FILLER_166_1136 ();
 sg13g2_fill_1 FILLER_166_1138 ();
 sg13g2_fill_2 FILLER_166_1147 ();
 sg13g2_fill_8 FILLER_166_1168 ();
 sg13g2_fill_2 FILLER_166_1176 ();
 sg13g2_fill_8 FILLER_166_1187 ();
 sg13g2_fill_1 FILLER_166_1195 ();
 sg13g2_fill_2 FILLER_166_1200 ();
 sg13g2_fill_4 FILLER_166_1211 ();
 sg13g2_fill_4 FILLER_166_1271 ();
 sg13g2_fill_2 FILLER_166_1275 ();
 sg13g2_fill_1 FILLER_166_1277 ();
 sg13g2_fill_1 FILLER_166_1295 ();
 sg13g2_fill_2 FILLER_166_1301 ();
 sg13g2_fill_1 FILLER_166_1303 ();
 sg13g2_fill_8 FILLER_166_1335 ();
 sg13g2_fill_4 FILLER_166_1343 ();
 sg13g2_fill_2 FILLER_166_1347 ();
 sg13g2_fill_8 FILLER_166_1354 ();
 sg13g2_fill_8 FILLER_166_1362 ();
 sg13g2_fill_8 FILLER_166_1386 ();
 sg13g2_fill_1 FILLER_166_1394 ();
 sg13g2_fill_8 FILLER_166_1411 ();
 sg13g2_fill_8 FILLER_166_1419 ();
 sg13g2_fill_8 FILLER_166_1431 ();
 sg13g2_fill_8 FILLER_166_1439 ();
 sg13g2_fill_8 FILLER_166_1447 ();
 sg13g2_fill_8 FILLER_166_1455 ();
 sg13g2_fill_8 FILLER_166_1463 ();
 sg13g2_fill_8 FILLER_166_1471 ();
 sg13g2_fill_8 FILLER_166_1479 ();
 sg13g2_fill_8 FILLER_166_1487 ();
 sg13g2_fill_8 FILLER_166_1495 ();
 sg13g2_fill_8 FILLER_166_1503 ();
 sg13g2_fill_8 FILLER_166_1511 ();
 sg13g2_fill_8 FILLER_166_1519 ();
 sg13g2_fill_8 FILLER_166_1527 ();
 sg13g2_fill_8 FILLER_166_1535 ();
 sg13g2_fill_8 FILLER_166_1543 ();
 sg13g2_fill_8 FILLER_166_1551 ();
 sg13g2_fill_8 FILLER_166_1559 ();
 sg13g2_fill_8 FILLER_166_1567 ();
 sg13g2_fill_8 FILLER_166_1575 ();
 sg13g2_fill_8 FILLER_166_1583 ();
 sg13g2_fill_1 FILLER_166_1591 ();
 sg13g2_fill_8 FILLER_167_0 ();
 sg13g2_fill_8 FILLER_167_8 ();
 sg13g2_fill_8 FILLER_167_16 ();
 sg13g2_fill_8 FILLER_167_24 ();
 sg13g2_fill_8 FILLER_167_32 ();
 sg13g2_fill_8 FILLER_167_40 ();
 sg13g2_fill_8 FILLER_167_48 ();
 sg13g2_fill_2 FILLER_167_56 ();
 sg13g2_fill_1 FILLER_167_58 ();
 sg13g2_fill_8 FILLER_167_69 ();
 sg13g2_fill_8 FILLER_167_77 ();
 sg13g2_fill_8 FILLER_167_95 ();
 sg13g2_fill_8 FILLER_167_103 ();
 sg13g2_fill_2 FILLER_167_111 ();
 sg13g2_fill_2 FILLER_167_149 ();
 sg13g2_fill_8 FILLER_167_192 ();
 sg13g2_fill_4 FILLER_167_200 ();
 sg13g2_fill_1 FILLER_167_204 ();
 sg13g2_fill_8 FILLER_167_239 ();
 sg13g2_fill_8 FILLER_167_247 ();
 sg13g2_fill_8 FILLER_167_255 ();
 sg13g2_fill_4 FILLER_167_263 ();
 sg13g2_fill_8 FILLER_167_277 ();
 sg13g2_fill_4 FILLER_167_285 ();
 sg13g2_fill_2 FILLER_167_294 ();
 sg13g2_fill_1 FILLER_167_296 ();
 sg13g2_fill_4 FILLER_167_302 ();
 sg13g2_fill_1 FILLER_167_306 ();
 sg13g2_fill_8 FILLER_167_348 ();
 sg13g2_fill_8 FILLER_167_392 ();
 sg13g2_fill_8 FILLER_167_400 ();
 sg13g2_fill_8 FILLER_167_408 ();
 sg13g2_fill_1 FILLER_167_452 ();
 sg13g2_fill_4 FILLER_167_479 ();
 sg13g2_fill_2 FILLER_167_483 ();
 sg13g2_fill_8 FILLER_167_521 ();
 sg13g2_fill_8 FILLER_167_529 ();
 sg13g2_fill_4 FILLER_167_537 ();
 sg13g2_fill_1 FILLER_167_541 ();
 sg13g2_fill_8 FILLER_167_567 ();
 sg13g2_fill_4 FILLER_167_575 ();
 sg13g2_fill_2 FILLER_167_579 ();
 sg13g2_fill_1 FILLER_167_581 ();
 sg13g2_fill_4 FILLER_167_592 ();
 sg13g2_fill_1 FILLER_167_596 ();
 sg13g2_fill_2 FILLER_167_623 ();
 sg13g2_fill_1 FILLER_167_625 ();
 sg13g2_fill_2 FILLER_167_662 ();
 sg13g2_fill_4 FILLER_167_684 ();
 sg13g2_fill_2 FILLER_167_688 ();
 sg13g2_fill_1 FILLER_167_690 ();
 sg13g2_fill_8 FILLER_167_701 ();
 sg13g2_fill_8 FILLER_167_735 ();
 sg13g2_fill_1 FILLER_167_743 ();
 sg13g2_fill_8 FILLER_167_770 ();
 sg13g2_fill_2 FILLER_167_794 ();
 sg13g2_fill_8 FILLER_167_817 ();
 sg13g2_fill_8 FILLER_167_825 ();
 sg13g2_fill_2 FILLER_167_833 ();
 sg13g2_fill_8 FILLER_167_844 ();
 sg13g2_fill_2 FILLER_167_852 ();
 sg13g2_fill_8 FILLER_167_866 ();
 sg13g2_fill_2 FILLER_167_874 ();
 sg13g2_fill_1 FILLER_167_876 ();
 sg13g2_fill_4 FILLER_167_885 ();
 sg13g2_fill_2 FILLER_167_889 ();
 sg13g2_fill_8 FILLER_167_917 ();
 sg13g2_fill_8 FILLER_167_925 ();
 sg13g2_fill_8 FILLER_167_933 ();
 sg13g2_fill_8 FILLER_167_941 ();
 sg13g2_fill_8 FILLER_167_949 ();
 sg13g2_fill_8 FILLER_167_957 ();
 sg13g2_fill_4 FILLER_167_965 ();
 sg13g2_fill_2 FILLER_167_969 ();
 sg13g2_fill_8 FILLER_167_992 ();
 sg13g2_fill_4 FILLER_167_1000 ();
 sg13g2_fill_2 FILLER_167_1004 ();
 sg13g2_fill_8 FILLER_167_1026 ();
 sg13g2_fill_8 FILLER_167_1034 ();
 sg13g2_fill_8 FILLER_167_1042 ();
 sg13g2_fill_8 FILLER_167_1050 ();
 sg13g2_fill_2 FILLER_167_1058 ();
 sg13g2_fill_1 FILLER_167_1060 ();
 sg13g2_fill_4 FILLER_167_1069 ();
 sg13g2_fill_2 FILLER_167_1073 ();
 sg13g2_fill_1 FILLER_167_1075 ();
 sg13g2_fill_2 FILLER_167_1092 ();
 sg13g2_fill_1 FILLER_167_1094 ();
 sg13g2_fill_8 FILLER_167_1130 ();
 sg13g2_fill_1 FILLER_167_1138 ();
 sg13g2_fill_8 FILLER_167_1148 ();
 sg13g2_fill_8 FILLER_167_1156 ();
 sg13g2_fill_1 FILLER_167_1164 ();
 sg13g2_fill_1 FILLER_167_1201 ();
 sg13g2_fill_1 FILLER_167_1211 ();
 sg13g2_fill_1 FILLER_167_1225 ();
 sg13g2_fill_8 FILLER_167_1230 ();
 sg13g2_fill_8 FILLER_167_1238 ();
 sg13g2_fill_1 FILLER_167_1246 ();
 sg13g2_fill_1 FILLER_167_1252 ();
 sg13g2_fill_8 FILLER_167_1263 ();
 sg13g2_fill_8 FILLER_167_1271 ();
 sg13g2_fill_8 FILLER_167_1279 ();
 sg13g2_fill_8 FILLER_167_1287 ();
 sg13g2_fill_8 FILLER_167_1295 ();
 sg13g2_fill_1 FILLER_167_1303 ();
 sg13g2_fill_4 FILLER_167_1313 ();
 sg13g2_fill_2 FILLER_167_1317 ();
 sg13g2_fill_8 FILLER_167_1324 ();
 sg13g2_fill_8 FILLER_167_1332 ();
 sg13g2_fill_1 FILLER_167_1340 ();
 sg13g2_fill_4 FILLER_167_1362 ();
 sg13g2_fill_8 FILLER_167_1386 ();
 sg13g2_fill_2 FILLER_167_1394 ();
 sg13g2_fill_4 FILLER_167_1404 ();
 sg13g2_fill_8 FILLER_167_1442 ();
 sg13g2_fill_8 FILLER_167_1450 ();
 sg13g2_fill_8 FILLER_167_1458 ();
 sg13g2_fill_8 FILLER_167_1466 ();
 sg13g2_fill_8 FILLER_167_1474 ();
 sg13g2_fill_8 FILLER_167_1482 ();
 sg13g2_fill_8 FILLER_167_1490 ();
 sg13g2_fill_8 FILLER_167_1498 ();
 sg13g2_fill_8 FILLER_167_1506 ();
 sg13g2_fill_8 FILLER_167_1514 ();
 sg13g2_fill_8 FILLER_167_1522 ();
 sg13g2_fill_8 FILLER_167_1530 ();
 sg13g2_fill_8 FILLER_167_1538 ();
 sg13g2_fill_8 FILLER_167_1546 ();
 sg13g2_fill_8 FILLER_167_1554 ();
 sg13g2_fill_8 FILLER_167_1562 ();
 sg13g2_fill_8 FILLER_167_1570 ();
 sg13g2_fill_8 FILLER_167_1578 ();
 sg13g2_fill_4 FILLER_167_1586 ();
 sg13g2_fill_2 FILLER_167_1590 ();
 sg13g2_fill_8 FILLER_168_0 ();
 sg13g2_fill_8 FILLER_168_8 ();
 sg13g2_fill_8 FILLER_168_16 ();
 sg13g2_fill_8 FILLER_168_24 ();
 sg13g2_fill_8 FILLER_168_32 ();
 sg13g2_fill_8 FILLER_168_40 ();
 sg13g2_fill_4 FILLER_168_48 ();
 sg13g2_fill_2 FILLER_168_52 ();
 sg13g2_fill_1 FILLER_168_54 ();
 sg13g2_fill_8 FILLER_168_81 ();
 sg13g2_fill_1 FILLER_168_125 ();
 sg13g2_fill_4 FILLER_168_136 ();
 sg13g2_fill_1 FILLER_168_140 ();
 sg13g2_fill_1 FILLER_168_153 ();
 sg13g2_fill_4 FILLER_168_171 ();
 sg13g2_fill_8 FILLER_168_211 ();
 sg13g2_fill_4 FILLER_168_219 ();
 sg13g2_fill_2 FILLER_168_223 ();
 sg13g2_fill_1 FILLER_168_225 ();
 sg13g2_fill_1 FILLER_168_252 ();
 sg13g2_fill_4 FILLER_168_279 ();
 sg13g2_fill_2 FILLER_168_283 ();
 sg13g2_fill_1 FILLER_168_285 ();
 sg13g2_fill_4 FILLER_168_312 ();
 sg13g2_fill_2 FILLER_168_316 ();
 sg13g2_fill_8 FILLER_168_328 ();
 sg13g2_fill_8 FILLER_168_336 ();
 sg13g2_fill_8 FILLER_168_344 ();
 sg13g2_fill_8 FILLER_168_352 ();
 sg13g2_fill_8 FILLER_168_360 ();
 sg13g2_fill_4 FILLER_168_368 ();
 sg13g2_fill_2 FILLER_168_372 ();
 sg13g2_fill_1 FILLER_168_374 ();
 sg13g2_fill_4 FILLER_168_381 ();
 sg13g2_fill_2 FILLER_168_385 ();
 sg13g2_fill_1 FILLER_168_387 ();
 sg13g2_fill_8 FILLER_168_414 ();
 sg13g2_fill_8 FILLER_168_422 ();
 sg13g2_fill_8 FILLER_168_446 ();
 sg13g2_fill_8 FILLER_168_454 ();
 sg13g2_fill_8 FILLER_168_462 ();
 sg13g2_fill_4 FILLER_168_470 ();
 sg13g2_fill_4 FILLER_168_484 ();
 sg13g2_fill_1 FILLER_168_488 ();
 sg13g2_fill_8 FILLER_168_495 ();
 sg13g2_fill_8 FILLER_168_503 ();
 sg13g2_fill_1 FILLER_168_511 ();
 sg13g2_fill_2 FILLER_168_522 ();
 sg13g2_fill_2 FILLER_168_530 ();
 sg13g2_fill_4 FILLER_168_542 ();
 sg13g2_fill_4 FILLER_168_561 ();
 sg13g2_fill_2 FILLER_168_565 ();
 sg13g2_fill_4 FILLER_168_593 ();
 sg13g2_fill_8 FILLER_168_607 ();
 sg13g2_fill_8 FILLER_168_615 ();
 sg13g2_fill_4 FILLER_168_623 ();
 sg13g2_fill_1 FILLER_168_627 ();
 sg13g2_fill_8 FILLER_168_638 ();
 sg13g2_fill_8 FILLER_168_646 ();
 sg13g2_fill_4 FILLER_168_659 ();
 sg13g2_fill_1 FILLER_168_663 ();
 sg13g2_fill_4 FILLER_168_690 ();
 sg13g2_fill_1 FILLER_168_694 ();
 sg13g2_fill_1 FILLER_168_724 ();
 sg13g2_fill_8 FILLER_168_745 ();
 sg13g2_fill_8 FILLER_168_753 ();
 sg13g2_fill_8 FILLER_168_761 ();
 sg13g2_fill_8 FILLER_168_790 ();
 sg13g2_fill_8 FILLER_168_798 ();
 sg13g2_fill_4 FILLER_168_806 ();
 sg13g2_fill_2 FILLER_168_810 ();
 sg13g2_fill_1 FILLER_168_812 ();
 sg13g2_fill_8 FILLER_168_818 ();
 sg13g2_fill_8 FILLER_168_843 ();
 sg13g2_fill_8 FILLER_168_856 ();
 sg13g2_fill_4 FILLER_168_864 ();
 sg13g2_fill_2 FILLER_168_868 ();
 sg13g2_fill_2 FILLER_168_879 ();
 sg13g2_fill_1 FILLER_168_881 ();
 sg13g2_fill_8 FILLER_168_895 ();
 sg13g2_fill_8 FILLER_168_903 ();
 sg13g2_fill_8 FILLER_168_911 ();
 sg13g2_fill_8 FILLER_168_919 ();
 sg13g2_fill_8 FILLER_168_927 ();
 sg13g2_fill_8 FILLER_168_935 ();
 sg13g2_fill_8 FILLER_168_943 ();
 sg13g2_fill_8 FILLER_168_951 ();
 sg13g2_fill_8 FILLER_168_959 ();
 sg13g2_fill_4 FILLER_168_967 ();
 sg13g2_fill_2 FILLER_168_971 ();
 sg13g2_fill_1 FILLER_168_979 ();
 sg13g2_fill_1 FILLER_168_984 ();
 sg13g2_fill_4 FILLER_168_995 ();
 sg13g2_fill_1 FILLER_168_999 ();
 sg13g2_fill_4 FILLER_168_1033 ();
 sg13g2_fill_2 FILLER_168_1037 ();
 sg13g2_fill_1 FILLER_168_1039 ();
 sg13g2_fill_4 FILLER_168_1048 ();
 sg13g2_fill_2 FILLER_168_1052 ();
 sg13g2_fill_2 FILLER_168_1059 ();
 sg13g2_fill_1 FILLER_168_1061 ();
 sg13g2_fill_2 FILLER_168_1082 ();
 sg13g2_fill_1 FILLER_168_1084 ();
 sg13g2_fill_2 FILLER_168_1089 ();
 sg13g2_fill_4 FILLER_168_1099 ();
 sg13g2_fill_2 FILLER_168_1103 ();
 sg13g2_fill_1 FILLER_168_1105 ();
 sg13g2_fill_8 FILLER_168_1162 ();
 sg13g2_fill_4 FILLER_168_1170 ();
 sg13g2_fill_2 FILLER_168_1174 ();
 sg13g2_fill_1 FILLER_168_1176 ();
 sg13g2_fill_8 FILLER_168_1184 ();
 sg13g2_fill_1 FILLER_168_1192 ();
 sg13g2_fill_8 FILLER_168_1214 ();
 sg13g2_fill_8 FILLER_168_1229 ();
 sg13g2_fill_8 FILLER_168_1237 ();
 sg13g2_fill_8 FILLER_168_1245 ();
 sg13g2_fill_8 FILLER_168_1253 ();
 sg13g2_fill_8 FILLER_168_1261 ();
 sg13g2_fill_2 FILLER_168_1280 ();
 sg13g2_fill_2 FILLER_168_1290 ();
 sg13g2_fill_1 FILLER_168_1292 ();
 sg13g2_fill_8 FILLER_168_1316 ();
 sg13g2_fill_2 FILLER_168_1337 ();
 sg13g2_fill_1 FILLER_168_1339 ();
 sg13g2_fill_4 FILLER_168_1357 ();
 sg13g2_fill_2 FILLER_168_1361 ();
 sg13g2_fill_8 FILLER_168_1389 ();
 sg13g2_fill_8 FILLER_168_1397 ();
 sg13g2_fill_4 FILLER_168_1405 ();
 sg13g2_fill_2 FILLER_168_1419 ();
 sg13g2_fill_1 FILLER_168_1421 ();
 sg13g2_fill_1 FILLER_168_1428 ();
 sg13g2_fill_8 FILLER_168_1434 ();
 sg13g2_fill_8 FILLER_168_1442 ();
 sg13g2_fill_8 FILLER_168_1450 ();
 sg13g2_fill_8 FILLER_168_1458 ();
 sg13g2_fill_8 FILLER_168_1466 ();
 sg13g2_fill_8 FILLER_168_1474 ();
 sg13g2_fill_8 FILLER_168_1482 ();
 sg13g2_fill_8 FILLER_168_1490 ();
 sg13g2_fill_8 FILLER_168_1498 ();
 sg13g2_fill_8 FILLER_168_1506 ();
 sg13g2_fill_8 FILLER_168_1514 ();
 sg13g2_fill_8 FILLER_168_1522 ();
 sg13g2_fill_8 FILLER_168_1530 ();
 sg13g2_fill_8 FILLER_168_1538 ();
 sg13g2_fill_8 FILLER_168_1546 ();
 sg13g2_fill_8 FILLER_168_1554 ();
 sg13g2_fill_8 FILLER_168_1562 ();
 sg13g2_fill_8 FILLER_168_1570 ();
 sg13g2_fill_8 FILLER_168_1578 ();
 sg13g2_fill_4 FILLER_168_1586 ();
 sg13g2_fill_2 FILLER_168_1590 ();
 sg13g2_fill_8 FILLER_169_0 ();
 sg13g2_fill_8 FILLER_169_8 ();
 sg13g2_fill_8 FILLER_169_16 ();
 sg13g2_fill_8 FILLER_169_24 ();
 sg13g2_fill_8 FILLER_169_32 ();
 sg13g2_fill_8 FILLER_169_40 ();
 sg13g2_fill_8 FILLER_169_48 ();
 sg13g2_fill_1 FILLER_169_56 ();
 sg13g2_fill_2 FILLER_169_147 ();
 sg13g2_fill_1 FILLER_169_149 ();
 sg13g2_fill_8 FILLER_169_160 ();
 sg13g2_fill_2 FILLER_169_168 ();
 sg13g2_fill_2 FILLER_169_175 ();
 sg13g2_fill_8 FILLER_169_183 ();
 sg13g2_fill_8 FILLER_169_191 ();
 sg13g2_fill_8 FILLER_169_199 ();
 sg13g2_fill_8 FILLER_169_207 ();
 sg13g2_fill_8 FILLER_169_215 ();
 sg13g2_fill_4 FILLER_169_223 ();
 sg13g2_fill_8 FILLER_169_243 ();
 sg13g2_fill_8 FILLER_169_251 ();
 sg13g2_fill_8 FILLER_169_259 ();
 sg13g2_fill_8 FILLER_169_267 ();
 sg13g2_fill_8 FILLER_169_275 ();
 sg13g2_fill_8 FILLER_169_283 ();
 sg13g2_fill_2 FILLER_169_291 ();
 sg13g2_fill_1 FILLER_169_293 ();
 sg13g2_fill_8 FILLER_169_327 ();
 sg13g2_fill_8 FILLER_169_335 ();
 sg13g2_fill_8 FILLER_169_343 ();
 sg13g2_fill_4 FILLER_169_351 ();
 sg13g2_fill_1 FILLER_169_355 ();
 sg13g2_fill_4 FILLER_169_379 ();
 sg13g2_fill_2 FILLER_169_383 ();
 sg13g2_fill_4 FILLER_169_421 ();
 sg13g2_fill_4 FILLER_169_435 ();
 sg13g2_fill_1 FILLER_169_455 ();
 sg13g2_fill_8 FILLER_169_466 ();
 sg13g2_fill_8 FILLER_169_474 ();
 sg13g2_fill_2 FILLER_169_482 ();
 sg13g2_fill_4 FILLER_169_500 ();
 sg13g2_fill_2 FILLER_169_546 ();
 sg13g2_fill_8 FILLER_169_574 ();
 sg13g2_fill_4 FILLER_169_582 ();
 sg13g2_fill_2 FILLER_169_586 ();
 sg13g2_fill_4 FILLER_169_598 ();
 sg13g2_fill_1 FILLER_169_602 ();
 sg13g2_fill_4 FILLER_169_613 ();
 sg13g2_fill_2 FILLER_169_617 ();
 sg13g2_fill_1 FILLER_169_619 ();
 sg13g2_fill_4 FILLER_169_681 ();
 sg13g2_fill_4 FILLER_169_703 ();
 sg13g2_fill_1 FILLER_169_707 ();
 sg13g2_fill_8 FILLER_169_753 ();
 sg13g2_fill_1 FILLER_169_761 ();
 sg13g2_fill_1 FILLER_169_773 ();
 sg13g2_fill_4 FILLER_169_778 ();
 sg13g2_fill_4 FILLER_169_789 ();
 sg13g2_fill_4 FILLER_169_798 ();
 sg13g2_fill_2 FILLER_169_825 ();
 sg13g2_fill_8 FILLER_169_840 ();
 sg13g2_fill_2 FILLER_169_848 ();
 sg13g2_fill_1 FILLER_169_850 ();
 sg13g2_fill_2 FILLER_169_871 ();
 sg13g2_fill_4 FILLER_169_888 ();
 sg13g2_fill_8 FILLER_169_906 ();
 sg13g2_fill_8 FILLER_169_914 ();
 sg13g2_fill_8 FILLER_169_922 ();
 sg13g2_fill_8 FILLER_169_930 ();
 sg13g2_fill_8 FILLER_169_938 ();
 sg13g2_fill_8 FILLER_169_946 ();
 sg13g2_fill_8 FILLER_169_954 ();
 sg13g2_fill_4 FILLER_169_962 ();
 sg13g2_fill_2 FILLER_169_970 ();
 sg13g2_fill_2 FILLER_169_977 ();
 sg13g2_fill_1 FILLER_169_979 ();
 sg13g2_fill_8 FILLER_169_997 ();
 sg13g2_fill_4 FILLER_169_1005 ();
 sg13g2_fill_2 FILLER_169_1009 ();
 sg13g2_fill_8 FILLER_169_1027 ();
 sg13g2_fill_4 FILLER_169_1035 ();
 sg13g2_fill_2 FILLER_169_1039 ();
 sg13g2_fill_1 FILLER_169_1041 ();
 sg13g2_fill_8 FILLER_169_1083 ();
 sg13g2_fill_8 FILLER_169_1091 ();
 sg13g2_fill_8 FILLER_169_1099 ();
 sg13g2_fill_8 FILLER_169_1107 ();
 sg13g2_fill_8 FILLER_169_1115 ();
 sg13g2_fill_8 FILLER_169_1123 ();
 sg13g2_fill_8 FILLER_169_1131 ();
 sg13g2_fill_1 FILLER_169_1139 ();
 sg13g2_fill_2 FILLER_169_1151 ();
 sg13g2_fill_1 FILLER_169_1153 ();
 sg13g2_fill_2 FILLER_169_1172 ();
 sg13g2_fill_8 FILLER_169_1178 ();
 sg13g2_fill_2 FILLER_169_1186 ();
 sg13g2_fill_1 FILLER_169_1188 ();
 sg13g2_fill_8 FILLER_169_1195 ();
 sg13g2_fill_1 FILLER_169_1203 ();
 sg13g2_fill_2 FILLER_169_1212 ();
 sg13g2_fill_1 FILLER_169_1214 ();
 sg13g2_fill_4 FILLER_169_1233 ();
 sg13g2_fill_1 FILLER_169_1237 ();
 sg13g2_fill_8 FILLER_169_1254 ();
 sg13g2_fill_1 FILLER_169_1262 ();
 sg13g2_fill_2 FILLER_169_1268 ();
 sg13g2_fill_8 FILLER_169_1290 ();
 sg13g2_fill_4 FILLER_169_1298 ();
 sg13g2_fill_8 FILLER_169_1306 ();
 sg13g2_fill_8 FILLER_169_1314 ();
 sg13g2_fill_8 FILLER_169_1322 ();
 sg13g2_fill_4 FILLER_169_1330 ();
 sg13g2_fill_1 FILLER_169_1343 ();
 sg13g2_fill_2 FILLER_169_1360 ();
 sg13g2_fill_1 FILLER_169_1362 ();
 sg13g2_fill_4 FILLER_169_1385 ();
 sg13g2_fill_2 FILLER_169_1389 ();
 sg13g2_fill_1 FILLER_169_1391 ();
 sg13g2_fill_1 FILLER_169_1401 ();
 sg13g2_fill_4 FILLER_169_1407 ();
 sg13g2_fill_2 FILLER_169_1423 ();
 sg13g2_fill_8 FILLER_169_1432 ();
 sg13g2_fill_8 FILLER_169_1440 ();
 sg13g2_fill_8 FILLER_169_1448 ();
 sg13g2_fill_8 FILLER_169_1456 ();
 sg13g2_fill_8 FILLER_169_1464 ();
 sg13g2_fill_8 FILLER_169_1472 ();
 sg13g2_fill_8 FILLER_169_1480 ();
 sg13g2_fill_8 FILLER_169_1488 ();
 sg13g2_fill_8 FILLER_169_1496 ();
 sg13g2_fill_8 FILLER_169_1504 ();
 sg13g2_fill_8 FILLER_169_1512 ();
 sg13g2_fill_8 FILLER_169_1520 ();
 sg13g2_fill_8 FILLER_169_1528 ();
 sg13g2_fill_8 FILLER_169_1536 ();
 sg13g2_fill_8 FILLER_169_1544 ();
 sg13g2_fill_8 FILLER_169_1552 ();
 sg13g2_fill_8 FILLER_169_1560 ();
 sg13g2_fill_8 FILLER_169_1568 ();
 sg13g2_fill_8 FILLER_169_1576 ();
 sg13g2_fill_8 FILLER_169_1584 ();
 sg13g2_fill_8 FILLER_170_0 ();
 sg13g2_fill_8 FILLER_170_8 ();
 sg13g2_fill_8 FILLER_170_16 ();
 sg13g2_fill_8 FILLER_170_24 ();
 sg13g2_fill_8 FILLER_170_32 ();
 sg13g2_fill_8 FILLER_170_40 ();
 sg13g2_fill_8 FILLER_170_48 ();
 sg13g2_fill_8 FILLER_170_56 ();
 sg13g2_fill_2 FILLER_170_64 ();
 sg13g2_fill_1 FILLER_170_66 ();
 sg13g2_fill_8 FILLER_170_73 ();
 sg13g2_fill_1 FILLER_170_133 ();
 sg13g2_fill_2 FILLER_170_154 ();
 sg13g2_fill_1 FILLER_170_156 ();
 sg13g2_fill_8 FILLER_170_177 ();
 sg13g2_fill_4 FILLER_170_185 ();
 sg13g2_fill_2 FILLER_170_189 ();
 sg13g2_fill_1 FILLER_170_191 ();
 sg13g2_fill_4 FILLER_170_200 ();
 sg13g2_fill_2 FILLER_170_204 ();
 sg13g2_fill_1 FILLER_170_206 ();
 sg13g2_fill_2 FILLER_170_248 ();
 sg13g2_fill_1 FILLER_170_250 ();
 sg13g2_fill_8 FILLER_170_277 ();
 sg13g2_fill_8 FILLER_170_285 ();
 sg13g2_fill_4 FILLER_170_293 ();
 sg13g2_fill_1 FILLER_170_297 ();
 sg13g2_fill_4 FILLER_170_304 ();
 sg13g2_fill_2 FILLER_170_308 ();
 sg13g2_fill_1 FILLER_170_310 ();
 sg13g2_fill_4 FILLER_170_321 ();
 sg13g2_fill_2 FILLER_170_325 ();
 sg13g2_fill_4 FILLER_170_348 ();
 sg13g2_fill_8 FILLER_170_360 ();
 sg13g2_fill_8 FILLER_170_368 ();
 sg13g2_fill_1 FILLER_170_376 ();
 sg13g2_fill_4 FILLER_170_408 ();
 sg13g2_fill_2 FILLER_170_412 ();
 sg13g2_fill_1 FILLER_170_414 ();
 sg13g2_fill_2 FILLER_170_425 ();
 sg13g2_fill_2 FILLER_170_452 ();
 sg13g2_fill_4 FILLER_170_480 ();
 sg13g2_fill_8 FILLER_170_494 ();
 sg13g2_fill_8 FILLER_170_502 ();
 sg13g2_fill_8 FILLER_170_510 ();
 sg13g2_fill_8 FILLER_170_518 ();
 sg13g2_fill_8 FILLER_170_526 ();
 sg13g2_fill_8 FILLER_170_534 ();
 sg13g2_fill_2 FILLER_170_542 ();
 sg13g2_fill_1 FILLER_170_544 ();
 sg13g2_fill_8 FILLER_170_560 ();
 sg13g2_fill_8 FILLER_170_568 ();
 sg13g2_fill_2 FILLER_170_576 ();
 sg13g2_fill_2 FILLER_170_596 ();
 sg13g2_fill_8 FILLER_170_634 ();
 sg13g2_fill_4 FILLER_170_642 ();
 sg13g2_fill_1 FILLER_170_646 ();
 sg13g2_fill_8 FILLER_170_655 ();
 sg13g2_fill_1 FILLER_170_663 ();
 sg13g2_fill_2 FILLER_170_699 ();
 sg13g2_fill_1 FILLER_170_701 ();
 sg13g2_fill_1 FILLER_170_728 ();
 sg13g2_fill_1 FILLER_170_785 ();
 sg13g2_fill_8 FILLER_170_798 ();
 sg13g2_fill_4 FILLER_170_806 ();
 sg13g2_fill_4 FILLER_170_820 ();
 sg13g2_fill_4 FILLER_170_829 ();
 sg13g2_fill_1 FILLER_170_833 ();
 sg13g2_fill_2 FILLER_170_848 ();
 sg13g2_fill_1 FILLER_170_850 ();
 sg13g2_fill_1 FILLER_170_864 ();
 sg13g2_fill_8 FILLER_170_892 ();
 sg13g2_fill_8 FILLER_170_900 ();
 sg13g2_fill_8 FILLER_170_908 ();
 sg13g2_fill_8 FILLER_170_916 ();
 sg13g2_fill_8 FILLER_170_924 ();
 sg13g2_fill_8 FILLER_170_932 ();
 sg13g2_fill_8 FILLER_170_940 ();
 sg13g2_fill_8 FILLER_170_948 ();
 sg13g2_fill_1 FILLER_170_956 ();
 sg13g2_fill_8 FILLER_170_983 ();
 sg13g2_fill_8 FILLER_170_991 ();
 sg13g2_fill_8 FILLER_170_999 ();
 sg13g2_fill_8 FILLER_170_1007 ();
 sg13g2_fill_4 FILLER_170_1015 ();
 sg13g2_fill_2 FILLER_170_1019 ();
 sg13g2_fill_8 FILLER_170_1026 ();
 sg13g2_fill_4 FILLER_170_1034 ();
 sg13g2_fill_2 FILLER_170_1038 ();
 sg13g2_fill_8 FILLER_170_1046 ();
 sg13g2_fill_2 FILLER_170_1054 ();
 sg13g2_fill_1 FILLER_170_1056 ();
 sg13g2_fill_8 FILLER_170_1072 ();
 sg13g2_fill_8 FILLER_170_1080 ();
 sg13g2_fill_2 FILLER_170_1088 ();
 sg13g2_fill_1 FILLER_170_1090 ();
 sg13g2_fill_8 FILLER_170_1099 ();
 sg13g2_fill_4 FILLER_170_1107 ();
 sg13g2_fill_8 FILLER_170_1120 ();
 sg13g2_fill_8 FILLER_170_1128 ();
 sg13g2_fill_8 FILLER_170_1136 ();
 sg13g2_fill_4 FILLER_170_1144 ();
 sg13g2_fill_2 FILLER_170_1148 ();
 sg13g2_fill_4 FILLER_170_1159 ();
 sg13g2_fill_2 FILLER_170_1168 ();
 sg13g2_fill_1 FILLER_170_1170 ();
 sg13g2_fill_2 FILLER_170_1180 ();
 sg13g2_fill_4 FILLER_170_1192 ();
 sg13g2_fill_8 FILLER_170_1199 ();
 sg13g2_fill_4 FILLER_170_1207 ();
 sg13g2_fill_2 FILLER_170_1211 ();
 sg13g2_fill_1 FILLER_170_1213 ();
 sg13g2_fill_8 FILLER_170_1223 ();
 sg13g2_fill_8 FILLER_170_1231 ();
 sg13g2_fill_2 FILLER_170_1239 ();
 sg13g2_fill_1 FILLER_170_1241 ();
 sg13g2_fill_1 FILLER_170_1263 ();
 sg13g2_fill_2 FILLER_170_1275 ();
 sg13g2_fill_1 FILLER_170_1277 ();
 sg13g2_fill_4 FILLER_170_1294 ();
 sg13g2_fill_2 FILLER_170_1298 ();
 sg13g2_fill_1 FILLER_170_1300 ();
 sg13g2_fill_4 FILLER_170_1306 ();
 sg13g2_fill_2 FILLER_170_1310 ();
 sg13g2_fill_1 FILLER_170_1328 ();
 sg13g2_fill_2 FILLER_170_1337 ();
 sg13g2_fill_1 FILLER_170_1339 ();
 sg13g2_fill_8 FILLER_170_1352 ();
 sg13g2_fill_8 FILLER_170_1360 ();
 sg13g2_fill_4 FILLER_170_1368 ();
 sg13g2_fill_2 FILLER_170_1372 ();
 sg13g2_fill_1 FILLER_170_1374 ();
 sg13g2_fill_8 FILLER_170_1379 ();
 sg13g2_fill_2 FILLER_170_1387 ();
 sg13g2_fill_2 FILLER_170_1401 ();
 sg13g2_fill_8 FILLER_170_1437 ();
 sg13g2_fill_8 FILLER_170_1445 ();
 sg13g2_fill_8 FILLER_170_1453 ();
 sg13g2_fill_8 FILLER_170_1461 ();
 sg13g2_fill_8 FILLER_170_1469 ();
 sg13g2_fill_8 FILLER_170_1477 ();
 sg13g2_fill_8 FILLER_170_1485 ();
 sg13g2_fill_8 FILLER_170_1493 ();
 sg13g2_fill_8 FILLER_170_1501 ();
 sg13g2_fill_8 FILLER_170_1509 ();
 sg13g2_fill_8 FILLER_170_1517 ();
 sg13g2_fill_8 FILLER_170_1525 ();
 sg13g2_fill_8 FILLER_170_1533 ();
 sg13g2_fill_8 FILLER_170_1541 ();
 sg13g2_fill_8 FILLER_170_1549 ();
 sg13g2_fill_8 FILLER_170_1557 ();
 sg13g2_fill_8 FILLER_170_1565 ();
 sg13g2_fill_8 FILLER_170_1573 ();
 sg13g2_fill_8 FILLER_170_1581 ();
 sg13g2_fill_2 FILLER_170_1589 ();
 sg13g2_fill_1 FILLER_170_1591 ();
 sg13g2_fill_8 FILLER_171_0 ();
 sg13g2_fill_8 FILLER_171_8 ();
 sg13g2_fill_8 FILLER_171_16 ();
 sg13g2_fill_8 FILLER_171_24 ();
 sg13g2_fill_8 FILLER_171_32 ();
 sg13g2_fill_8 FILLER_171_40 ();
 sg13g2_fill_8 FILLER_171_48 ();
 sg13g2_fill_8 FILLER_171_56 ();
 sg13g2_fill_8 FILLER_171_64 ();
 sg13g2_fill_2 FILLER_171_72 ();
 sg13g2_fill_8 FILLER_171_113 ();
 sg13g2_fill_8 FILLER_171_121 ();
 sg13g2_fill_8 FILLER_171_129 ();
 sg13g2_fill_4 FILLER_171_137 ();
 sg13g2_fill_2 FILLER_171_141 ();
 sg13g2_fill_2 FILLER_171_195 ();
 sg13g2_fill_4 FILLER_171_268 ();
 sg13g2_fill_1 FILLER_171_303 ();
 sg13g2_fill_2 FILLER_171_330 ();
 sg13g2_fill_2 FILLER_171_353 ();
 sg13g2_fill_1 FILLER_171_355 ();
 sg13g2_fill_2 FILLER_171_382 ();
 sg13g2_fill_1 FILLER_171_384 ();
 sg13g2_fill_8 FILLER_171_447 ();
 sg13g2_fill_8 FILLER_171_455 ();
 sg13g2_fill_4 FILLER_171_463 ();
 sg13g2_fill_2 FILLER_171_467 ();
 sg13g2_fill_1 FILLER_171_505 ();
 sg13g2_fill_2 FILLER_171_542 ();
 sg13g2_fill_1 FILLER_171_544 ();
 sg13g2_fill_4 FILLER_171_553 ();
 sg13g2_fill_2 FILLER_171_557 ();
 sg13g2_fill_1 FILLER_171_559 ();
 sg13g2_fill_1 FILLER_171_586 ();
 sg13g2_fill_4 FILLER_171_632 ();
 sg13g2_fill_8 FILLER_171_662 ();
 sg13g2_fill_8 FILLER_171_706 ();
 sg13g2_fill_4 FILLER_171_714 ();
 sg13g2_fill_4 FILLER_171_728 ();
 sg13g2_fill_4 FILLER_171_757 ();
 sg13g2_fill_2 FILLER_171_761 ();
 sg13g2_fill_1 FILLER_171_763 ();
 sg13g2_fill_4 FILLER_171_769 ();
 sg13g2_fill_2 FILLER_171_773 ();
 sg13g2_fill_2 FILLER_171_786 ();
 sg13g2_fill_4 FILLER_171_798 ();
 sg13g2_fill_2 FILLER_171_802 ();
 sg13g2_fill_8 FILLER_171_809 ();
 sg13g2_fill_8 FILLER_171_817 ();
 sg13g2_fill_4 FILLER_171_825 ();
 sg13g2_fill_8 FILLER_171_838 ();
 sg13g2_fill_2 FILLER_171_846 ();
 sg13g2_fill_2 FILLER_171_856 ();
 sg13g2_fill_8 FILLER_171_866 ();
 sg13g2_fill_8 FILLER_171_874 ();
 sg13g2_fill_8 FILLER_171_882 ();
 sg13g2_fill_8 FILLER_171_890 ();
 sg13g2_fill_8 FILLER_171_898 ();
 sg13g2_fill_8 FILLER_171_906 ();
 sg13g2_fill_8 FILLER_171_914 ();
 sg13g2_fill_8 FILLER_171_922 ();
 sg13g2_fill_8 FILLER_171_930 ();
 sg13g2_fill_8 FILLER_171_938 ();
 sg13g2_fill_8 FILLER_171_946 ();
 sg13g2_fill_4 FILLER_171_954 ();
 sg13g2_fill_2 FILLER_171_958 ();
 sg13g2_fill_1 FILLER_171_960 ();
 sg13g2_fill_2 FILLER_171_969 ();
 sg13g2_fill_1 FILLER_171_971 ();
 sg13g2_fill_2 FILLER_171_991 ();
 sg13g2_fill_1 FILLER_171_993 ();
 sg13g2_fill_2 FILLER_171_1010 ();
 sg13g2_fill_1 FILLER_171_1012 ();
 sg13g2_fill_1 FILLER_171_1017 ();
 sg13g2_fill_1 FILLER_171_1033 ();
 sg13g2_fill_8 FILLER_171_1044 ();
 sg13g2_fill_8 FILLER_171_1052 ();
 sg13g2_fill_1 FILLER_171_1060 ();
 sg13g2_fill_8 FILLER_171_1069 ();
 sg13g2_fill_1 FILLER_171_1077 ();
 sg13g2_fill_2 FILLER_171_1103 ();
 sg13g2_fill_1 FILLER_171_1105 ();
 sg13g2_fill_8 FILLER_171_1132 ();
 sg13g2_fill_2 FILLER_171_1140 ();
 sg13g2_fill_1 FILLER_171_1142 ();
 sg13g2_fill_2 FILLER_171_1151 ();
 sg13g2_fill_1 FILLER_171_1164 ();
 sg13g2_fill_2 FILLER_171_1186 ();
 sg13g2_fill_4 FILLER_171_1218 ();
 sg13g2_fill_2 FILLER_171_1232 ();
 sg13g2_fill_1 FILLER_171_1234 ();
 sg13g2_fill_4 FILLER_171_1238 ();
 sg13g2_fill_1 FILLER_171_1245 ();
 sg13g2_fill_4 FILLER_171_1252 ();
 sg13g2_fill_4 FILLER_171_1269 ();
 sg13g2_fill_4 FILLER_171_1290 ();
 sg13g2_fill_1 FILLER_171_1294 ();
 sg13g2_fill_8 FILLER_171_1326 ();
 sg13g2_fill_2 FILLER_171_1334 ();
 sg13g2_fill_1 FILLER_171_1336 ();
 sg13g2_fill_8 FILLER_171_1346 ();
 sg13g2_fill_8 FILLER_171_1354 ();
 sg13g2_fill_4 FILLER_171_1362 ();
 sg13g2_fill_8 FILLER_171_1382 ();
 sg13g2_fill_4 FILLER_171_1390 ();
 sg13g2_fill_1 FILLER_171_1394 ();
 sg13g2_fill_8 FILLER_171_1414 ();
 sg13g2_fill_4 FILLER_171_1431 ();
 sg13g2_fill_2 FILLER_171_1440 ();
 sg13g2_fill_1 FILLER_171_1442 ();
 sg13g2_fill_8 FILLER_171_1446 ();
 sg13g2_fill_8 FILLER_171_1454 ();
 sg13g2_fill_8 FILLER_171_1462 ();
 sg13g2_fill_8 FILLER_171_1470 ();
 sg13g2_fill_8 FILLER_171_1478 ();
 sg13g2_fill_8 FILLER_171_1486 ();
 sg13g2_fill_8 FILLER_171_1494 ();
 sg13g2_fill_8 FILLER_171_1502 ();
 sg13g2_fill_8 FILLER_171_1510 ();
 sg13g2_fill_8 FILLER_171_1518 ();
 sg13g2_fill_8 FILLER_171_1526 ();
 sg13g2_fill_8 FILLER_171_1534 ();
 sg13g2_fill_8 FILLER_171_1542 ();
 sg13g2_fill_8 FILLER_171_1550 ();
 sg13g2_fill_8 FILLER_171_1558 ();
 sg13g2_fill_8 FILLER_171_1566 ();
 sg13g2_fill_8 FILLER_171_1574 ();
 sg13g2_fill_8 FILLER_171_1582 ();
 sg13g2_fill_2 FILLER_171_1590 ();
 sg13g2_fill_8 FILLER_172_0 ();
 sg13g2_fill_8 FILLER_172_8 ();
 sg13g2_fill_8 FILLER_172_16 ();
 sg13g2_fill_8 FILLER_172_24 ();
 sg13g2_fill_8 FILLER_172_32 ();
 sg13g2_fill_8 FILLER_172_40 ();
 sg13g2_fill_8 FILLER_172_48 ();
 sg13g2_fill_8 FILLER_172_56 ();
 sg13g2_fill_8 FILLER_172_64 ();
 sg13g2_fill_8 FILLER_172_72 ();
 sg13g2_fill_8 FILLER_172_80 ();
 sg13g2_fill_8 FILLER_172_88 ();
 sg13g2_fill_8 FILLER_172_96 ();
 sg13g2_fill_8 FILLER_172_104 ();
 sg13g2_fill_8 FILLER_172_112 ();
 sg13g2_fill_8 FILLER_172_120 ();
 sg13g2_fill_1 FILLER_172_128 ();
 sg13g2_fill_8 FILLER_172_135 ();
 sg13g2_fill_8 FILLER_172_143 ();
 sg13g2_fill_8 FILLER_172_151 ();
 sg13g2_fill_4 FILLER_172_159 ();
 sg13g2_fill_1 FILLER_172_163 ();
 sg13g2_fill_8 FILLER_172_174 ();
 sg13g2_fill_4 FILLER_172_182 ();
 sg13g2_fill_2 FILLER_172_202 ();
 sg13g2_fill_1 FILLER_172_204 ();
 sg13g2_fill_8 FILLER_172_215 ();
 sg13g2_fill_2 FILLER_172_223 ();
 sg13g2_fill_8 FILLER_172_229 ();
 sg13g2_fill_1 FILLER_172_294 ();
 sg13g2_fill_8 FILLER_172_305 ();
 sg13g2_fill_4 FILLER_172_313 ();
 sg13g2_fill_1 FILLER_172_317 ();
 sg13g2_fill_8 FILLER_172_326 ();
 sg13g2_fill_2 FILLER_172_334 ();
 sg13g2_fill_4 FILLER_172_367 ();
 sg13g2_fill_1 FILLER_172_371 ();
 sg13g2_fill_8 FILLER_172_398 ();
 sg13g2_fill_8 FILLER_172_406 ();
 sg13g2_fill_8 FILLER_172_414 ();
 sg13g2_fill_4 FILLER_172_422 ();
 sg13g2_fill_1 FILLER_172_426 ();
 sg13g2_fill_8 FILLER_172_440 ();
 sg13g2_fill_1 FILLER_172_448 ();
 sg13g2_fill_4 FILLER_172_510 ();
 sg13g2_fill_2 FILLER_172_514 ();
 sg13g2_fill_1 FILLER_172_516 ();
 sg13g2_fill_8 FILLER_172_527 ();
 sg13g2_fill_4 FILLER_172_535 ();
 sg13g2_fill_1 FILLER_172_539 ();
 sg13g2_fill_8 FILLER_172_557 ();
 sg13g2_fill_8 FILLER_172_565 ();
 sg13g2_fill_4 FILLER_172_573 ();
 sg13g2_fill_2 FILLER_172_577 ();
 sg13g2_fill_8 FILLER_172_584 ();
 sg13g2_fill_8 FILLER_172_592 ();
 sg13g2_fill_1 FILLER_172_600 ();
 sg13g2_fill_4 FILLER_172_627 ();
 sg13g2_fill_8 FILLER_172_649 ();
 sg13g2_fill_8 FILLER_172_657 ();
 sg13g2_fill_1 FILLER_172_665 ();
 sg13g2_fill_8 FILLER_172_701 ();
 sg13g2_fill_8 FILLER_172_709 ();
 sg13g2_fill_2 FILLER_172_717 ();
 sg13g2_fill_4 FILLER_172_752 ();
 sg13g2_fill_2 FILLER_172_756 ();
 sg13g2_fill_1 FILLER_172_758 ();
 sg13g2_fill_8 FILLER_172_769 ();
 sg13g2_fill_4 FILLER_172_788 ();
 sg13g2_fill_8 FILLER_172_813 ();
 sg13g2_fill_8 FILLER_172_821 ();
 sg13g2_fill_8 FILLER_172_829 ();
 sg13g2_fill_8 FILLER_172_837 ();
 sg13g2_fill_2 FILLER_172_845 ();
 sg13g2_fill_1 FILLER_172_847 ();
 sg13g2_fill_8 FILLER_172_860 ();
 sg13g2_fill_8 FILLER_172_868 ();
 sg13g2_fill_8 FILLER_172_876 ();
 sg13g2_fill_8 FILLER_172_884 ();
 sg13g2_fill_8 FILLER_172_892 ();
 sg13g2_fill_8 FILLER_172_900 ();
 sg13g2_fill_8 FILLER_172_908 ();
 sg13g2_fill_8 FILLER_172_916 ();
 sg13g2_fill_8 FILLER_172_924 ();
 sg13g2_fill_8 FILLER_172_932 ();
 sg13g2_fill_8 FILLER_172_940 ();
 sg13g2_fill_8 FILLER_172_948 ();
 sg13g2_fill_8 FILLER_172_956 ();
 sg13g2_fill_8 FILLER_172_983 ();
 sg13g2_fill_8 FILLER_172_991 ();
 sg13g2_fill_2 FILLER_172_999 ();
 sg13g2_fill_2 FILLER_172_1009 ();
 sg13g2_fill_1 FILLER_172_1011 ();
 sg13g2_fill_2 FILLER_172_1017 ();
 sg13g2_fill_2 FILLER_172_1052 ();
 sg13g2_fill_1 FILLER_172_1054 ();
 sg13g2_fill_8 FILLER_172_1075 ();
 sg13g2_fill_1 FILLER_172_1083 ();
 sg13g2_fill_2 FILLER_172_1092 ();
 sg13g2_fill_1 FILLER_172_1126 ();
 sg13g2_fill_2 FILLER_172_1141 ();
 sg13g2_fill_1 FILLER_172_1143 ();
 sg13g2_fill_4 FILLER_172_1152 ();
 sg13g2_fill_2 FILLER_172_1156 ();
 sg13g2_fill_1 FILLER_172_1158 ();
 sg13g2_fill_8 FILLER_172_1167 ();
 sg13g2_fill_4 FILLER_172_1184 ();
 sg13g2_fill_1 FILLER_172_1188 ();
 sg13g2_fill_8 FILLER_172_1204 ();
 sg13g2_fill_8 FILLER_172_1212 ();
 sg13g2_fill_4 FILLER_172_1220 ();
 sg13g2_fill_2 FILLER_172_1224 ();
 sg13g2_fill_1 FILLER_172_1226 ();
 sg13g2_fill_8 FILLER_172_1243 ();
 sg13g2_fill_8 FILLER_172_1251 ();
 sg13g2_fill_8 FILLER_172_1259 ();
 sg13g2_fill_2 FILLER_172_1267 ();
 sg13g2_fill_2 FILLER_172_1274 ();
 sg13g2_fill_1 FILLER_172_1276 ();
 sg13g2_fill_8 FILLER_172_1284 ();
 sg13g2_fill_1 FILLER_172_1292 ();
 sg13g2_fill_8 FILLER_172_1306 ();
 sg13g2_fill_8 FILLER_172_1314 ();
 sg13g2_fill_8 FILLER_172_1322 ();
 sg13g2_fill_4 FILLER_172_1330 ();
 sg13g2_fill_2 FILLER_172_1334 ();
 sg13g2_fill_1 FILLER_172_1336 ();
 sg13g2_fill_4 FILLER_172_1348 ();
 sg13g2_fill_2 FILLER_172_1363 ();
 sg13g2_fill_4 FILLER_172_1389 ();
 sg13g2_fill_1 FILLER_172_1393 ();
 sg13g2_fill_8 FILLER_172_1402 ();
 sg13g2_fill_8 FILLER_172_1410 ();
 sg13g2_fill_8 FILLER_172_1418 ();
 sg13g2_fill_8 FILLER_172_1426 ();
 sg13g2_fill_1 FILLER_172_1434 ();
 sg13g2_fill_8 FILLER_172_1442 ();
 sg13g2_fill_8 FILLER_172_1450 ();
 sg13g2_fill_8 FILLER_172_1458 ();
 sg13g2_fill_8 FILLER_172_1466 ();
 sg13g2_fill_8 FILLER_172_1474 ();
 sg13g2_fill_8 FILLER_172_1482 ();
 sg13g2_fill_8 FILLER_172_1490 ();
 sg13g2_fill_8 FILLER_172_1498 ();
 sg13g2_fill_8 FILLER_172_1506 ();
 sg13g2_fill_8 FILLER_172_1514 ();
 sg13g2_fill_8 FILLER_172_1522 ();
 sg13g2_fill_8 FILLER_172_1530 ();
 sg13g2_fill_8 FILLER_172_1538 ();
 sg13g2_fill_8 FILLER_172_1546 ();
 sg13g2_fill_8 FILLER_172_1554 ();
 sg13g2_fill_8 FILLER_172_1562 ();
 sg13g2_fill_8 FILLER_172_1570 ();
 sg13g2_fill_8 FILLER_172_1578 ();
 sg13g2_fill_4 FILLER_172_1586 ();
 sg13g2_fill_2 FILLER_172_1590 ();
 sg13g2_fill_8 FILLER_173_0 ();
 sg13g2_fill_8 FILLER_173_8 ();
 sg13g2_fill_8 FILLER_173_16 ();
 sg13g2_fill_8 FILLER_173_24 ();
 sg13g2_fill_8 FILLER_173_32 ();
 sg13g2_fill_8 FILLER_173_40 ();
 sg13g2_fill_8 FILLER_173_48 ();
 sg13g2_fill_8 FILLER_173_56 ();
 sg13g2_fill_8 FILLER_173_64 ();
 sg13g2_fill_4 FILLER_173_72 ();
 sg13g2_fill_2 FILLER_173_76 ();
 sg13g2_fill_8 FILLER_173_88 ();
 sg13g2_fill_8 FILLER_173_96 ();
 sg13g2_fill_4 FILLER_173_104 ();
 sg13g2_fill_4 FILLER_173_118 ();
 sg13g2_fill_2 FILLER_173_122 ();
 sg13g2_fill_1 FILLER_173_124 ();
 sg13g2_fill_2 FILLER_173_141 ();
 sg13g2_fill_1 FILLER_173_143 ();
 sg13g2_fill_1 FILLER_173_154 ();
 sg13g2_fill_8 FILLER_173_169 ();
 sg13g2_fill_1 FILLER_173_177 ();
 sg13g2_fill_8 FILLER_173_184 ();
 sg13g2_fill_4 FILLER_173_192 ();
 sg13g2_fill_2 FILLER_173_196 ();
 sg13g2_fill_8 FILLER_173_204 ();
 sg13g2_fill_8 FILLER_173_212 ();
 sg13g2_fill_4 FILLER_173_220 ();
 sg13g2_fill_2 FILLER_173_224 ();
 sg13g2_fill_1 FILLER_173_226 ();
 sg13g2_fill_4 FILLER_173_233 ();
 sg13g2_fill_2 FILLER_173_237 ();
 sg13g2_fill_4 FILLER_173_255 ();
 sg13g2_fill_2 FILLER_173_259 ();
 sg13g2_fill_2 FILLER_173_271 ();
 sg13g2_fill_8 FILLER_173_309 ();
 sg13g2_fill_8 FILLER_173_317 ();
 sg13g2_fill_8 FILLER_173_325 ();
 sg13g2_fill_8 FILLER_173_333 ();
 sg13g2_fill_1 FILLER_173_341 ();
 sg13g2_fill_8 FILLER_173_398 ();
 sg13g2_fill_1 FILLER_173_406 ();
 sg13g2_fill_8 FILLER_173_415 ();
 sg13g2_fill_1 FILLER_173_423 ();
 sg13g2_fill_8 FILLER_173_460 ();
 sg13g2_fill_8 FILLER_173_468 ();
 sg13g2_fill_4 FILLER_173_476 ();
 sg13g2_fill_4 FILLER_173_539 ();
 sg13g2_fill_1 FILLER_173_543 ();
 sg13g2_fill_8 FILLER_173_580 ();
 sg13g2_fill_8 FILLER_173_588 ();
 sg13g2_fill_2 FILLER_173_596 ();
 sg13g2_fill_8 FILLER_173_608 ();
 sg13g2_fill_8 FILLER_173_616 ();
 sg13g2_fill_8 FILLER_173_624 ();
 sg13g2_fill_4 FILLER_173_632 ();
 sg13g2_fill_1 FILLER_173_636 ();
 sg13g2_fill_8 FILLER_173_642 ();
 sg13g2_fill_2 FILLER_173_650 ();
 sg13g2_fill_2 FILLER_173_687 ();
 sg13g2_fill_1 FILLER_173_689 ();
 sg13g2_fill_2 FILLER_173_721 ();
 sg13g2_fill_4 FILLER_173_753 ();
 sg13g2_fill_1 FILLER_173_757 ();
 sg13g2_fill_8 FILLER_173_779 ();
 sg13g2_fill_8 FILLER_173_787 ();
 sg13g2_fill_4 FILLER_173_795 ();
 sg13g2_fill_8 FILLER_173_835 ();
 sg13g2_fill_8 FILLER_173_843 ();
 sg13g2_fill_8 FILLER_173_851 ();
 sg13g2_fill_8 FILLER_173_859 ();
 sg13g2_fill_8 FILLER_173_867 ();
 sg13g2_fill_8 FILLER_173_875 ();
 sg13g2_fill_8 FILLER_173_883 ();
 sg13g2_fill_8 FILLER_173_891 ();
 sg13g2_fill_8 FILLER_173_899 ();
 sg13g2_fill_8 FILLER_173_907 ();
 sg13g2_fill_8 FILLER_173_915 ();
 sg13g2_fill_8 FILLER_173_923 ();
 sg13g2_fill_8 FILLER_173_931 ();
 sg13g2_fill_8 FILLER_173_939 ();
 sg13g2_fill_8 FILLER_173_947 ();
 sg13g2_fill_8 FILLER_173_955 ();
 sg13g2_fill_4 FILLER_173_963 ();
 sg13g2_fill_4 FILLER_173_971 ();
 sg13g2_fill_2 FILLER_173_983 ();
 sg13g2_fill_8 FILLER_173_990 ();
 sg13g2_fill_2 FILLER_173_998 ();
 sg13g2_fill_1 FILLER_173_1000 ();
 sg13g2_fill_2 FILLER_173_1030 ();
 sg13g2_fill_1 FILLER_173_1032 ();
 sg13g2_fill_2 FILLER_173_1052 ();
 sg13g2_fill_2 FILLER_173_1083 ();
 sg13g2_fill_1 FILLER_173_1085 ();
 sg13g2_fill_4 FILLER_173_1098 ();
 sg13g2_fill_2 FILLER_173_1102 ();
 sg13g2_fill_4 FILLER_173_1119 ();
 sg13g2_fill_2 FILLER_173_1123 ();
 sg13g2_fill_1 FILLER_173_1125 ();
 sg13g2_fill_4 FILLER_173_1136 ();
 sg13g2_fill_4 FILLER_173_1153 ();
 sg13g2_fill_1 FILLER_173_1157 ();
 sg13g2_fill_4 FILLER_173_1187 ();
 sg13g2_fill_2 FILLER_173_1191 ();
 sg13g2_fill_1 FILLER_173_1193 ();
 sg13g2_fill_8 FILLER_173_1199 ();
 sg13g2_fill_8 FILLER_173_1207 ();
 sg13g2_fill_8 FILLER_173_1215 ();
 sg13g2_fill_4 FILLER_173_1239 ();
 sg13g2_fill_2 FILLER_173_1243 ();
 sg13g2_fill_1 FILLER_173_1245 ();
 sg13g2_fill_8 FILLER_173_1262 ();
 sg13g2_fill_8 FILLER_173_1270 ();
 sg13g2_fill_2 FILLER_173_1278 ();
 sg13g2_fill_1 FILLER_173_1280 ();
 sg13g2_fill_4 FILLER_173_1287 ();
 sg13g2_fill_8 FILLER_173_1298 ();
 sg13g2_fill_8 FILLER_173_1306 ();
 sg13g2_fill_2 FILLER_173_1314 ();
 sg13g2_fill_2 FILLER_173_1324 ();
 sg13g2_fill_1 FILLER_173_1326 ();
 sg13g2_fill_4 FILLER_173_1348 ();
 sg13g2_fill_1 FILLER_173_1352 ();
 sg13g2_fill_4 FILLER_173_1357 ();
 sg13g2_fill_8 FILLER_173_1386 ();
 sg13g2_fill_4 FILLER_173_1394 ();
 sg13g2_fill_2 FILLER_173_1405 ();
 sg13g2_fill_1 FILLER_173_1407 ();
 sg13g2_fill_8 FILLER_173_1417 ();
 sg13g2_fill_4 FILLER_173_1425 ();
 sg13g2_fill_2 FILLER_173_1429 ();
 sg13g2_fill_8 FILLER_173_1452 ();
 sg13g2_fill_8 FILLER_173_1460 ();
 sg13g2_fill_8 FILLER_173_1468 ();
 sg13g2_fill_8 FILLER_173_1476 ();
 sg13g2_fill_8 FILLER_173_1484 ();
 sg13g2_fill_8 FILLER_173_1492 ();
 sg13g2_fill_8 FILLER_173_1500 ();
 sg13g2_fill_8 FILLER_173_1508 ();
 sg13g2_fill_8 FILLER_173_1516 ();
 sg13g2_fill_8 FILLER_173_1524 ();
 sg13g2_fill_8 FILLER_173_1532 ();
 sg13g2_fill_8 FILLER_173_1540 ();
 sg13g2_fill_8 FILLER_173_1548 ();
 sg13g2_fill_8 FILLER_173_1556 ();
 sg13g2_fill_8 FILLER_173_1564 ();
 sg13g2_fill_8 FILLER_173_1572 ();
 sg13g2_fill_8 FILLER_173_1580 ();
 sg13g2_fill_4 FILLER_173_1588 ();
 sg13g2_fill_8 FILLER_174_0 ();
 sg13g2_fill_8 FILLER_174_8 ();
 sg13g2_fill_8 FILLER_174_16 ();
 sg13g2_fill_8 FILLER_174_24 ();
 sg13g2_fill_8 FILLER_174_32 ();
 sg13g2_fill_8 FILLER_174_40 ();
 sg13g2_fill_8 FILLER_174_48 ();
 sg13g2_fill_8 FILLER_174_56 ();
 sg13g2_fill_8 FILLER_174_64 ();
 sg13g2_fill_8 FILLER_174_72 ();
 sg13g2_fill_1 FILLER_174_106 ();
 sg13g2_fill_2 FILLER_174_143 ();
 sg13g2_fill_4 FILLER_174_163 ();
 sg13g2_fill_4 FILLER_174_177 ();
 sg13g2_fill_1 FILLER_174_181 ();
 sg13g2_fill_2 FILLER_174_188 ();
 sg13g2_fill_1 FILLER_174_237 ();
 sg13g2_fill_2 FILLER_174_254 ();
 sg13g2_fill_2 FILLER_174_282 ();
 sg13g2_fill_1 FILLER_174_284 ();
 sg13g2_fill_2 FILLER_174_311 ();
 sg13g2_fill_1 FILLER_174_321 ();
 sg13g2_fill_4 FILLER_174_383 ();
 sg13g2_fill_2 FILLER_174_387 ();
 sg13g2_fill_2 FILLER_174_415 ();
 sg13g2_fill_8 FILLER_174_427 ();
 sg13g2_fill_4 FILLER_174_435 ();
 sg13g2_fill_2 FILLER_174_449 ();
 sg13g2_fill_8 FILLER_174_455 ();
 sg13g2_fill_8 FILLER_174_489 ();
 sg13g2_fill_8 FILLER_174_507 ();
 sg13g2_fill_8 FILLER_174_515 ();
 sg13g2_fill_4 FILLER_174_523 ();
 sg13g2_fill_1 FILLER_174_527 ();
 sg13g2_fill_4 FILLER_174_574 ();
 sg13g2_fill_2 FILLER_174_578 ();
 sg13g2_fill_8 FILLER_174_600 ();
 sg13g2_fill_8 FILLER_174_608 ();
 sg13g2_fill_8 FILLER_174_626 ();
 sg13g2_fill_8 FILLER_174_634 ();
 sg13g2_fill_1 FILLER_174_642 ();
 sg13g2_fill_4 FILLER_174_669 ();
 sg13g2_fill_2 FILLER_174_709 ();
 sg13g2_fill_1 FILLER_174_711 ();
 sg13g2_fill_4 FILLER_174_722 ();
 sg13g2_fill_1 FILLER_174_726 ();
 sg13g2_fill_8 FILLER_174_753 ();
 sg13g2_fill_8 FILLER_174_761 ();
 sg13g2_fill_8 FILLER_174_769 ();
 sg13g2_fill_8 FILLER_174_777 ();
 sg13g2_fill_8 FILLER_174_785 ();
 sg13g2_fill_8 FILLER_174_793 ();
 sg13g2_fill_8 FILLER_174_801 ();
 sg13g2_fill_8 FILLER_174_809 ();
 sg13g2_fill_8 FILLER_174_817 ();
 sg13g2_fill_8 FILLER_174_825 ();
 sg13g2_fill_8 FILLER_174_833 ();
 sg13g2_fill_8 FILLER_174_841 ();
 sg13g2_fill_8 FILLER_174_849 ();
 sg13g2_fill_8 FILLER_174_857 ();
 sg13g2_fill_8 FILLER_174_865 ();
 sg13g2_fill_8 FILLER_174_873 ();
 sg13g2_fill_8 FILLER_174_881 ();
 sg13g2_fill_8 FILLER_174_889 ();
 sg13g2_fill_8 FILLER_174_897 ();
 sg13g2_fill_8 FILLER_174_905 ();
 sg13g2_fill_8 FILLER_174_913 ();
 sg13g2_fill_8 FILLER_174_921 ();
 sg13g2_fill_8 FILLER_174_929 ();
 sg13g2_fill_8 FILLER_174_937 ();
 sg13g2_fill_8 FILLER_174_945 ();
 sg13g2_fill_8 FILLER_174_953 ();
 sg13g2_fill_8 FILLER_174_961 ();
 sg13g2_fill_1 FILLER_174_969 ();
 sg13g2_fill_2 FILLER_174_976 ();
 sg13g2_fill_1 FILLER_174_978 ();
 sg13g2_fill_4 FILLER_174_1000 ();
 sg13g2_fill_2 FILLER_174_1004 ();
 sg13g2_fill_8 FILLER_174_1023 ();
 sg13g2_fill_8 FILLER_174_1031 ();
 sg13g2_fill_8 FILLER_174_1039 ();
 sg13g2_fill_8 FILLER_174_1047 ();
 sg13g2_fill_8 FILLER_174_1055 ();
 sg13g2_fill_2 FILLER_174_1063 ();
 sg13g2_fill_1 FILLER_174_1065 ();
 sg13g2_fill_2 FILLER_174_1074 ();
 sg13g2_fill_1 FILLER_174_1076 ();
 sg13g2_fill_8 FILLER_174_1090 ();
 sg13g2_fill_8 FILLER_174_1106 ();
 sg13g2_fill_4 FILLER_174_1114 ();
 sg13g2_fill_4 FILLER_174_1126 ();
 sg13g2_fill_2 FILLER_174_1135 ();
 sg13g2_fill_1 FILLER_174_1137 ();
 sg13g2_fill_8 FILLER_174_1143 ();
 sg13g2_fill_8 FILLER_174_1151 ();
 sg13g2_fill_8 FILLER_174_1159 ();
 sg13g2_fill_8 FILLER_174_1167 ();
 sg13g2_fill_8 FILLER_174_1175 ();
 sg13g2_fill_8 FILLER_174_1183 ();
 sg13g2_fill_2 FILLER_174_1222 ();
 sg13g2_fill_1 FILLER_174_1224 ();
 sg13g2_fill_2 FILLER_174_1233 ();
 sg13g2_fill_1 FILLER_174_1235 ();
 sg13g2_fill_2 FILLER_174_1270 ();
 sg13g2_fill_2 FILLER_174_1277 ();
 sg13g2_fill_1 FILLER_174_1279 ();
 sg13g2_fill_4 FILLER_174_1305 ();
 sg13g2_fill_1 FILLER_174_1309 ();
 sg13g2_fill_2 FILLER_174_1337 ();
 sg13g2_fill_1 FILLER_174_1351 ();
 sg13g2_fill_2 FILLER_174_1363 ();
 sg13g2_fill_1 FILLER_174_1374 ();
 sg13g2_fill_8 FILLER_174_1380 ();
 sg13g2_fill_8 FILLER_174_1388 ();
 sg13g2_fill_2 FILLER_174_1396 ();
 sg13g2_fill_1 FILLER_174_1398 ();
 sg13g2_fill_4 FILLER_174_1429 ();
 sg13g2_fill_1 FILLER_174_1433 ();
 sg13g2_fill_4 FILLER_174_1437 ();
 sg13g2_fill_8 FILLER_174_1447 ();
 sg13g2_fill_8 FILLER_174_1455 ();
 sg13g2_fill_8 FILLER_174_1463 ();
 sg13g2_fill_8 FILLER_174_1471 ();
 sg13g2_fill_8 FILLER_174_1479 ();
 sg13g2_fill_8 FILLER_174_1487 ();
 sg13g2_fill_8 FILLER_174_1495 ();
 sg13g2_fill_8 FILLER_174_1503 ();
 sg13g2_fill_8 FILLER_174_1511 ();
 sg13g2_fill_8 FILLER_174_1519 ();
 sg13g2_fill_8 FILLER_174_1527 ();
 sg13g2_fill_8 FILLER_174_1535 ();
 sg13g2_fill_8 FILLER_174_1543 ();
 sg13g2_fill_8 FILLER_174_1551 ();
 sg13g2_fill_8 FILLER_174_1559 ();
 sg13g2_fill_8 FILLER_174_1567 ();
 sg13g2_fill_8 FILLER_174_1575 ();
 sg13g2_fill_8 FILLER_174_1583 ();
 sg13g2_fill_1 FILLER_174_1591 ();
 sg13g2_fill_8 FILLER_175_0 ();
 sg13g2_fill_8 FILLER_175_8 ();
 sg13g2_fill_8 FILLER_175_16 ();
 sg13g2_fill_8 FILLER_175_24 ();
 sg13g2_fill_8 FILLER_175_32 ();
 sg13g2_fill_8 FILLER_175_40 ();
 sg13g2_fill_8 FILLER_175_48 ();
 sg13g2_fill_8 FILLER_175_56 ();
 sg13g2_fill_4 FILLER_175_64 ();
 sg13g2_fill_2 FILLER_175_68 ();
 sg13g2_fill_1 FILLER_175_70 ();
 sg13g2_fill_8 FILLER_175_117 ();
 sg13g2_fill_1 FILLER_175_125 ();
 sg13g2_fill_8 FILLER_175_136 ();
 sg13g2_fill_4 FILLER_175_144 ();
 sg13g2_fill_2 FILLER_175_189 ();
 sg13g2_fill_1 FILLER_175_191 ();
 sg13g2_fill_4 FILLER_175_207 ();
 sg13g2_fill_8 FILLER_175_231 ();
 sg13g2_fill_4 FILLER_175_239 ();
 sg13g2_fill_1 FILLER_175_243 ();
 sg13g2_fill_8 FILLER_175_254 ();
 sg13g2_fill_8 FILLER_175_262 ();
 sg13g2_fill_4 FILLER_175_270 ();
 sg13g2_fill_2 FILLER_175_274 ();
 sg13g2_fill_1 FILLER_175_276 ();
 sg13g2_fill_8 FILLER_175_287 ();
 sg13g2_fill_8 FILLER_175_295 ();
 sg13g2_fill_4 FILLER_175_303 ();
 sg13g2_fill_2 FILLER_175_307 ();
 sg13g2_fill_1 FILLER_175_309 ();
 sg13g2_fill_4 FILLER_175_346 ();
 sg13g2_fill_2 FILLER_175_350 ();
 sg13g2_fill_1 FILLER_175_352 ();
 sg13g2_fill_8 FILLER_175_396 ();
 sg13g2_fill_8 FILLER_175_404 ();
 sg13g2_fill_2 FILLER_175_412 ();
 sg13g2_fill_4 FILLER_175_450 ();
 sg13g2_fill_2 FILLER_175_454 ();
 sg13g2_fill_1 FILLER_175_456 ();
 sg13g2_fill_4 FILLER_175_493 ();
 sg13g2_fill_4 FILLER_175_523 ();
 sg13g2_fill_1 FILLER_175_527 ();
 sg13g2_fill_4 FILLER_175_553 ();
 sg13g2_fill_2 FILLER_175_567 ();
 sg13g2_fill_2 FILLER_175_595 ();
 sg13g2_fill_1 FILLER_175_597 ();
 sg13g2_fill_1 FILLER_175_650 ();
 sg13g2_fill_4 FILLER_175_671 ();
 sg13g2_fill_8 FILLER_175_710 ();
 sg13g2_fill_4 FILLER_175_718 ();
 sg13g2_fill_8 FILLER_175_732 ();
 sg13g2_fill_2 FILLER_175_740 ();
 sg13g2_fill_4 FILLER_175_752 ();
 sg13g2_fill_2 FILLER_175_756 ();
 sg13g2_fill_1 FILLER_175_758 ();
 sg13g2_fill_4 FILLER_175_769 ();
 sg13g2_fill_4 FILLER_175_799 ();
 sg13g2_fill_2 FILLER_175_803 ();
 sg13g2_fill_8 FILLER_175_815 ();
 sg13g2_fill_8 FILLER_175_823 ();
 sg13g2_fill_8 FILLER_175_831 ();
 sg13g2_fill_8 FILLER_175_839 ();
 sg13g2_fill_8 FILLER_175_847 ();
 sg13g2_fill_8 FILLER_175_855 ();
 sg13g2_fill_8 FILLER_175_863 ();
 sg13g2_fill_8 FILLER_175_871 ();
 sg13g2_fill_8 FILLER_175_879 ();
 sg13g2_fill_8 FILLER_175_887 ();
 sg13g2_fill_8 FILLER_175_895 ();
 sg13g2_fill_8 FILLER_175_903 ();
 sg13g2_fill_8 FILLER_175_911 ();
 sg13g2_fill_8 FILLER_175_919 ();
 sg13g2_fill_8 FILLER_175_927 ();
 sg13g2_fill_8 FILLER_175_935 ();
 sg13g2_fill_8 FILLER_175_943 ();
 sg13g2_fill_8 FILLER_175_951 ();
 sg13g2_fill_8 FILLER_175_959 ();
 sg13g2_fill_8 FILLER_175_967 ();
 sg13g2_fill_4 FILLER_175_975 ();
 sg13g2_fill_2 FILLER_175_979 ();
 sg13g2_fill_1 FILLER_175_981 ();
 sg13g2_fill_8 FILLER_175_993 ();
 sg13g2_fill_8 FILLER_175_1001 ();
 sg13g2_fill_8 FILLER_175_1009 ();
 sg13g2_fill_4 FILLER_175_1017 ();
 sg13g2_fill_1 FILLER_175_1021 ();
 sg13g2_fill_8 FILLER_175_1025 ();
 sg13g2_fill_8 FILLER_175_1033 ();
 sg13g2_fill_8 FILLER_175_1041 ();
 sg13g2_fill_8 FILLER_175_1049 ();
 sg13g2_fill_4 FILLER_175_1057 ();
 sg13g2_fill_2 FILLER_175_1061 ();
 sg13g2_fill_2 FILLER_175_1071 ();
 sg13g2_fill_8 FILLER_175_1076 ();
 sg13g2_fill_8 FILLER_175_1084 ();
 sg13g2_fill_1 FILLER_175_1092 ();
 sg13g2_fill_2 FILLER_175_1099 ();
 sg13g2_fill_4 FILLER_175_1106 ();
 sg13g2_fill_2 FILLER_175_1110 ();
 sg13g2_fill_4 FILLER_175_1117 ();
 sg13g2_fill_2 FILLER_175_1121 ();
 sg13g2_fill_2 FILLER_175_1134 ();
 sg13g2_fill_8 FILLER_175_1144 ();
 sg13g2_fill_4 FILLER_175_1152 ();
 sg13g2_fill_1 FILLER_175_1165 ();
 sg13g2_fill_4 FILLER_175_1174 ();
 sg13g2_fill_1 FILLER_175_1178 ();
 sg13g2_fill_8 FILLER_175_1187 ();
 sg13g2_fill_4 FILLER_175_1195 ();
 sg13g2_fill_2 FILLER_175_1199 ();
 sg13g2_fill_2 FILLER_175_1225 ();
 sg13g2_fill_8 FILLER_175_1232 ();
 sg13g2_fill_8 FILLER_175_1240 ();
 sg13g2_fill_2 FILLER_175_1248 ();
 sg13g2_fill_4 FILLER_175_1258 ();
 sg13g2_fill_1 FILLER_175_1262 ();
 sg13g2_fill_4 FILLER_175_1287 ();
 sg13g2_fill_8 FILLER_175_1296 ();
 sg13g2_fill_8 FILLER_175_1316 ();
 sg13g2_fill_8 FILLER_175_1324 ();
 sg13g2_fill_8 FILLER_175_1332 ();
 sg13g2_fill_4 FILLER_175_1340 ();
 sg13g2_fill_8 FILLER_175_1348 ();
 sg13g2_fill_8 FILLER_175_1356 ();
 sg13g2_fill_2 FILLER_175_1364 ();
 sg13g2_fill_1 FILLER_175_1366 ();
 sg13g2_fill_8 FILLER_175_1372 ();
 sg13g2_fill_1 FILLER_175_1387 ();
 sg13g2_fill_1 FILLER_175_1397 ();
 sg13g2_fill_4 FILLER_175_1417 ();
 sg13g2_fill_2 FILLER_175_1421 ();
 sg13g2_fill_1 FILLER_175_1423 ();
 sg13g2_fill_1 FILLER_175_1428 ();
 sg13g2_fill_8 FILLER_175_1447 ();
 sg13g2_fill_8 FILLER_175_1455 ();
 sg13g2_fill_8 FILLER_175_1463 ();
 sg13g2_fill_8 FILLER_175_1471 ();
 sg13g2_fill_8 FILLER_175_1479 ();
 sg13g2_fill_8 FILLER_175_1487 ();
 sg13g2_fill_8 FILLER_175_1495 ();
 sg13g2_fill_8 FILLER_175_1503 ();
 sg13g2_fill_8 FILLER_175_1511 ();
 sg13g2_fill_8 FILLER_175_1519 ();
 sg13g2_fill_8 FILLER_175_1527 ();
 sg13g2_fill_8 FILLER_175_1535 ();
 sg13g2_fill_8 FILLER_175_1543 ();
 sg13g2_fill_8 FILLER_175_1551 ();
 sg13g2_fill_8 FILLER_175_1559 ();
 sg13g2_fill_8 FILLER_175_1567 ();
 sg13g2_fill_8 FILLER_175_1575 ();
 sg13g2_fill_8 FILLER_175_1583 ();
 sg13g2_fill_1 FILLER_175_1591 ();
 sg13g2_fill_8 FILLER_176_0 ();
 sg13g2_fill_8 FILLER_176_8 ();
 sg13g2_fill_8 FILLER_176_24 ();
 sg13g2_fill_8 FILLER_176_32 ();
 sg13g2_fill_8 FILLER_176_40 ();
 sg13g2_fill_8 FILLER_176_48 ();
 sg13g2_fill_8 FILLER_176_56 ();
 sg13g2_fill_8 FILLER_176_64 ();
 sg13g2_fill_8 FILLER_176_72 ();
 sg13g2_fill_8 FILLER_176_80 ();
 sg13g2_fill_8 FILLER_176_88 ();
 sg13g2_fill_8 FILLER_176_96 ();
 sg13g2_fill_8 FILLER_176_104 ();
 sg13g2_fill_8 FILLER_176_112 ();
 sg13g2_fill_8 FILLER_176_120 ();
 sg13g2_fill_8 FILLER_176_128 ();
 sg13g2_fill_1 FILLER_176_136 ();
 sg13g2_fill_4 FILLER_176_147 ();
 sg13g2_fill_2 FILLER_176_151 ();
 sg13g2_fill_1 FILLER_176_153 ();
 sg13g2_fill_1 FILLER_176_160 ();
 sg13g2_fill_2 FILLER_176_166 ();
 sg13g2_fill_2 FILLER_176_178 ();
 sg13g2_fill_8 FILLER_176_215 ();
 sg13g2_fill_8 FILLER_176_223 ();
 sg13g2_fill_8 FILLER_176_231 ();
 sg13g2_fill_8 FILLER_176_239 ();
 sg13g2_fill_8 FILLER_176_247 ();
 sg13g2_fill_8 FILLER_176_255 ();
 sg13g2_fill_8 FILLER_176_263 ();
 sg13g2_fill_8 FILLER_176_271 ();
 sg13g2_fill_8 FILLER_176_279 ();
 sg13g2_fill_8 FILLER_176_287 ();
 sg13g2_fill_8 FILLER_176_305 ();
 sg13g2_fill_2 FILLER_176_313 ();
 sg13g2_fill_2 FILLER_176_320 ();
 sg13g2_fill_8 FILLER_176_330 ();
 sg13g2_fill_8 FILLER_176_338 ();
 sg13g2_fill_1 FILLER_176_346 ();
 sg13g2_fill_8 FILLER_176_394 ();
 sg13g2_fill_8 FILLER_176_402 ();
 sg13g2_fill_4 FILLER_176_410 ();
 sg13g2_fill_1 FILLER_176_414 ();
 sg13g2_fill_8 FILLER_176_425 ();
 sg13g2_fill_8 FILLER_176_433 ();
 sg13g2_fill_8 FILLER_176_441 ();
 sg13g2_fill_4 FILLER_176_449 ();
 sg13g2_fill_2 FILLER_176_453 ();
 sg13g2_fill_8 FILLER_176_500 ();
 sg13g2_fill_4 FILLER_176_508 ();
 sg13g2_fill_1 FILLER_176_512 ();
 sg13g2_fill_4 FILLER_176_549 ();
 sg13g2_fill_8 FILLER_176_578 ();
 sg13g2_fill_8 FILLER_176_586 ();
 sg13g2_fill_4 FILLER_176_604 ();
 sg13g2_fill_2 FILLER_176_608 ();
 sg13g2_fill_4 FILLER_176_630 ();
 sg13g2_fill_1 FILLER_176_634 ();
 sg13g2_fill_4 FILLER_176_660 ();
 sg13g2_fill_4 FILLER_176_725 ();
 sg13g2_fill_2 FILLER_176_729 ();
 sg13g2_fill_2 FILLER_176_741 ();
 sg13g2_fill_2 FILLER_176_766 ();
 sg13g2_fill_2 FILLER_176_790 ();
 sg13g2_fill_1 FILLER_176_792 ();
 sg13g2_fill_8 FILLER_176_839 ();
 sg13g2_fill_8 FILLER_176_847 ();
 sg13g2_fill_8 FILLER_176_855 ();
 sg13g2_fill_8 FILLER_176_863 ();
 sg13g2_fill_8 FILLER_176_871 ();
 sg13g2_fill_8 FILLER_176_879 ();
 sg13g2_fill_8 FILLER_176_887 ();
 sg13g2_fill_8 FILLER_176_895 ();
 sg13g2_fill_8 FILLER_176_903 ();
 sg13g2_fill_8 FILLER_176_911 ();
 sg13g2_fill_8 FILLER_176_919 ();
 sg13g2_fill_8 FILLER_176_927 ();
 sg13g2_fill_8 FILLER_176_935 ();
 sg13g2_fill_8 FILLER_176_943 ();
 sg13g2_fill_8 FILLER_176_951 ();
 sg13g2_fill_8 FILLER_176_959 ();
 sg13g2_fill_4 FILLER_176_967 ();
 sg13g2_fill_2 FILLER_176_971 ();
 sg13g2_fill_8 FILLER_176_981 ();
 sg13g2_fill_2 FILLER_176_989 ();
 sg13g2_fill_2 FILLER_176_999 ();
 sg13g2_fill_1 FILLER_176_1001 ();
 sg13g2_fill_1 FILLER_176_1016 ();
 sg13g2_fill_1 FILLER_176_1030 ();
 sg13g2_fill_1 FILLER_176_1045 ();
 sg13g2_fill_2 FILLER_176_1059 ();
 sg13g2_fill_1 FILLER_176_1093 ();
 sg13g2_fill_2 FILLER_176_1100 ();
 sg13g2_fill_1 FILLER_176_1102 ();
 sg13g2_fill_8 FILLER_176_1109 ();
 sg13g2_fill_1 FILLER_176_1117 ();
 sg13g2_fill_8 FILLER_176_1126 ();
 sg13g2_fill_8 FILLER_176_1134 ();
 sg13g2_fill_2 FILLER_176_1142 ();
 sg13g2_fill_1 FILLER_176_1144 ();
 sg13g2_fill_2 FILLER_176_1171 ();
 sg13g2_fill_8 FILLER_176_1196 ();
 sg13g2_fill_2 FILLER_176_1204 ();
 sg13g2_fill_1 FILLER_176_1206 ();
 sg13g2_fill_2 FILLER_176_1212 ();
 sg13g2_fill_1 FILLER_176_1214 ();
 sg13g2_fill_2 FILLER_176_1220 ();
 sg13g2_fill_4 FILLER_176_1226 ();
 sg13g2_fill_2 FILLER_176_1230 ();
 sg13g2_fill_8 FILLER_176_1237 ();
 sg13g2_fill_4 FILLER_176_1245 ();
 sg13g2_fill_1 FILLER_176_1249 ();
 sg13g2_fill_8 FILLER_176_1261 ();
 sg13g2_fill_8 FILLER_176_1274 ();
 sg13g2_fill_8 FILLER_176_1282 ();
 sg13g2_fill_8 FILLER_176_1290 ();
 sg13g2_fill_8 FILLER_176_1303 ();
 sg13g2_fill_4 FILLER_176_1311 ();
 sg13g2_fill_1 FILLER_176_1315 ();
 sg13g2_fill_4 FILLER_176_1324 ();
 sg13g2_fill_2 FILLER_176_1340 ();
 sg13g2_fill_8 FILLER_176_1347 ();
 sg13g2_fill_4 FILLER_176_1355 ();
 sg13g2_fill_2 FILLER_176_1371 ();
 sg13g2_fill_1 FILLER_176_1412 ();
 sg13g2_fill_8 FILLER_176_1454 ();
 sg13g2_fill_8 FILLER_176_1462 ();
 sg13g2_fill_8 FILLER_176_1470 ();
 sg13g2_fill_8 FILLER_176_1478 ();
 sg13g2_fill_8 FILLER_176_1486 ();
 sg13g2_fill_8 FILLER_176_1494 ();
 sg13g2_fill_8 FILLER_176_1502 ();
 sg13g2_fill_8 FILLER_176_1510 ();
 sg13g2_fill_8 FILLER_176_1518 ();
 sg13g2_fill_8 FILLER_176_1526 ();
 sg13g2_fill_8 FILLER_176_1534 ();
 sg13g2_fill_8 FILLER_176_1542 ();
 sg13g2_fill_8 FILLER_176_1550 ();
 sg13g2_fill_8 FILLER_176_1558 ();
 sg13g2_fill_8 FILLER_176_1566 ();
 sg13g2_fill_8 FILLER_176_1574 ();
 sg13g2_fill_8 FILLER_176_1582 ();
 sg13g2_fill_2 FILLER_176_1590 ();
 sg13g2_fill_8 FILLER_177_0 ();
 sg13g2_fill_8 FILLER_177_8 ();
 sg13g2_fill_8 FILLER_177_16 ();
 sg13g2_fill_8 FILLER_177_24 ();
 sg13g2_fill_8 FILLER_177_32 ();
 sg13g2_fill_8 FILLER_177_40 ();
 sg13g2_fill_8 FILLER_177_48 ();
 sg13g2_fill_8 FILLER_177_56 ();
 sg13g2_fill_4 FILLER_177_64 ();
 sg13g2_fill_2 FILLER_177_68 ();
 sg13g2_fill_8 FILLER_177_75 ();
 sg13g2_fill_2 FILLER_177_83 ();
 sg13g2_fill_1 FILLER_177_85 ();
 sg13g2_fill_4 FILLER_177_96 ();
 sg13g2_fill_2 FILLER_177_100 ();
 sg13g2_fill_4 FILLER_177_112 ();
 sg13g2_fill_8 FILLER_177_121 ();
 sg13g2_fill_1 FILLER_177_165 ();
 sg13g2_fill_4 FILLER_177_176 ();
 sg13g2_fill_2 FILLER_177_231 ();
 sg13g2_fill_1 FILLER_177_233 ();
 sg13g2_fill_2 FILLER_177_252 ();
 sg13g2_fill_1 FILLER_177_280 ();
 sg13g2_fill_4 FILLER_177_291 ();
 sg13g2_fill_1 FILLER_177_295 ();
 sg13g2_fill_4 FILLER_177_306 ();
 sg13g2_fill_2 FILLER_177_310 ();
 sg13g2_fill_1 FILLER_177_312 ();
 sg13g2_fill_2 FILLER_177_318 ();
 sg13g2_fill_8 FILLER_177_332 ();
 sg13g2_fill_8 FILLER_177_340 ();
 sg13g2_fill_4 FILLER_177_348 ();
 sg13g2_fill_2 FILLER_177_352 ();
 sg13g2_fill_4 FILLER_177_416 ();
 sg13g2_fill_8 FILLER_177_446 ();
 sg13g2_fill_8 FILLER_177_454 ();
 sg13g2_fill_2 FILLER_177_462 ();
 sg13g2_fill_1 FILLER_177_464 ();
 sg13g2_fill_8 FILLER_177_471 ();
 sg13g2_fill_8 FILLER_177_479 ();
 sg13g2_fill_8 FILLER_177_487 ();
 sg13g2_fill_4 FILLER_177_495 ();
 sg13g2_fill_2 FILLER_177_499 ();
 sg13g2_fill_1 FILLER_177_501 ();
 sg13g2_fill_4 FILLER_177_512 ();
 sg13g2_fill_2 FILLER_177_516 ();
 sg13g2_fill_2 FILLER_177_553 ();
 sg13g2_fill_1 FILLER_177_555 ();
 sg13g2_fill_2 FILLER_177_576 ();
 sg13g2_fill_8 FILLER_177_614 ();
 sg13g2_fill_2 FILLER_177_622 ();
 sg13g2_fill_1 FILLER_177_624 ();
 sg13g2_fill_2 FILLER_177_673 ();
 sg13g2_fill_1 FILLER_177_675 ();
 sg13g2_fill_4 FILLER_177_712 ();
 sg13g2_fill_2 FILLER_177_777 ();
 sg13g2_fill_8 FILLER_177_789 ();
 sg13g2_fill_4 FILLER_177_797 ();
 sg13g2_fill_8 FILLER_177_811 ();
 sg13g2_fill_8 FILLER_177_819 ();
 sg13g2_fill_8 FILLER_177_827 ();
 sg13g2_fill_8 FILLER_177_835 ();
 sg13g2_fill_8 FILLER_177_843 ();
 sg13g2_fill_8 FILLER_177_851 ();
 sg13g2_fill_8 FILLER_177_859 ();
 sg13g2_fill_8 FILLER_177_867 ();
 sg13g2_fill_8 FILLER_177_875 ();
 sg13g2_fill_8 FILLER_177_883 ();
 sg13g2_fill_8 FILLER_177_891 ();
 sg13g2_fill_8 FILLER_177_899 ();
 sg13g2_fill_8 FILLER_177_907 ();
 sg13g2_fill_8 FILLER_177_915 ();
 sg13g2_fill_8 FILLER_177_923 ();
 sg13g2_fill_8 FILLER_177_931 ();
 sg13g2_fill_8 FILLER_177_939 ();
 sg13g2_fill_8 FILLER_177_947 ();
 sg13g2_fill_8 FILLER_177_955 ();
 sg13g2_fill_4 FILLER_177_963 ();
 sg13g2_fill_2 FILLER_177_967 ();
 sg13g2_fill_8 FILLER_177_985 ();
 sg13g2_fill_4 FILLER_177_993 ();
 sg13g2_fill_1 FILLER_177_997 ();
 sg13g2_fill_2 FILLER_177_1016 ();
 sg13g2_fill_2 FILLER_177_1037 ();
 sg13g2_fill_4 FILLER_177_1060 ();
 sg13g2_fill_2 FILLER_177_1064 ();
 sg13g2_fill_1 FILLER_177_1066 ();
 sg13g2_fill_8 FILLER_177_1072 ();
 sg13g2_fill_4 FILLER_177_1096 ();
 sg13g2_fill_1 FILLER_177_1100 ();
 sg13g2_fill_2 FILLER_177_1119 ();
 sg13g2_fill_4 FILLER_177_1133 ();
 sg13g2_fill_8 FILLER_177_1145 ();
 sg13g2_fill_1 FILLER_177_1153 ();
 sg13g2_fill_8 FILLER_177_1163 ();
 sg13g2_fill_2 FILLER_177_1171 ();
 sg13g2_fill_1 FILLER_177_1173 ();
 sg13g2_fill_4 FILLER_177_1191 ();
 sg13g2_fill_4 FILLER_177_1222 ();
 sg13g2_fill_4 FILLER_177_1236 ();
 sg13g2_fill_1 FILLER_177_1240 ();
 sg13g2_fill_8 FILLER_177_1262 ();
 sg13g2_fill_1 FILLER_177_1270 ();
 sg13g2_fill_8 FILLER_177_1277 ();
 sg13g2_fill_2 FILLER_177_1285 ();
 sg13g2_fill_1 FILLER_177_1287 ();
 sg13g2_fill_4 FILLER_177_1294 ();
 sg13g2_fill_2 FILLER_177_1309 ();
 sg13g2_fill_2 FILLER_177_1339 ();
 sg13g2_fill_8 FILLER_177_1357 ();
 sg13g2_fill_1 FILLER_177_1365 ();
 sg13g2_fill_4 FILLER_177_1375 ();
 sg13g2_fill_2 FILLER_177_1379 ();
 sg13g2_fill_8 FILLER_177_1393 ();
 sg13g2_fill_8 FILLER_177_1408 ();
 sg13g2_fill_8 FILLER_177_1416 ();
 sg13g2_fill_2 FILLER_177_1424 ();
 sg13g2_fill_1 FILLER_177_1436 ();
 sg13g2_fill_8 FILLER_177_1447 ();
 sg13g2_fill_8 FILLER_177_1455 ();
 sg13g2_fill_8 FILLER_177_1463 ();
 sg13g2_fill_8 FILLER_177_1471 ();
 sg13g2_fill_8 FILLER_177_1479 ();
 sg13g2_fill_8 FILLER_177_1487 ();
 sg13g2_fill_8 FILLER_177_1495 ();
 sg13g2_fill_8 FILLER_177_1503 ();
 sg13g2_fill_8 FILLER_177_1511 ();
 sg13g2_fill_8 FILLER_177_1519 ();
 sg13g2_fill_8 FILLER_177_1527 ();
 sg13g2_fill_8 FILLER_177_1535 ();
 sg13g2_fill_8 FILLER_177_1543 ();
 sg13g2_fill_8 FILLER_177_1551 ();
 sg13g2_fill_8 FILLER_177_1559 ();
 sg13g2_fill_8 FILLER_177_1567 ();
 sg13g2_fill_8 FILLER_177_1575 ();
 sg13g2_fill_8 FILLER_177_1583 ();
 sg13g2_fill_1 FILLER_177_1591 ();
 sg13g2_fill_8 FILLER_178_0 ();
 sg13g2_fill_8 FILLER_178_8 ();
 sg13g2_fill_8 FILLER_178_16 ();
 sg13g2_fill_8 FILLER_178_24 ();
 sg13g2_fill_8 FILLER_178_32 ();
 sg13g2_fill_8 FILLER_178_40 ();
 sg13g2_fill_8 FILLER_178_48 ();
 sg13g2_fill_8 FILLER_178_56 ();
 sg13g2_fill_8 FILLER_178_64 ();
 sg13g2_fill_8 FILLER_178_72 ();
 sg13g2_fill_8 FILLER_178_142 ();
 sg13g2_fill_8 FILLER_178_150 ();
 sg13g2_fill_8 FILLER_178_158 ();
 sg13g2_fill_2 FILLER_178_192 ();
 sg13g2_fill_1 FILLER_178_194 ();
 sg13g2_fill_4 FILLER_178_205 ();
 sg13g2_fill_2 FILLER_178_209 ();
 sg13g2_fill_2 FILLER_178_221 ();
 sg13g2_fill_2 FILLER_178_259 ();
 sg13g2_fill_8 FILLER_178_313 ();
 sg13g2_fill_2 FILLER_178_321 ();
 sg13g2_fill_8 FILLER_178_359 ();
 sg13g2_fill_8 FILLER_178_367 ();
 sg13g2_fill_8 FILLER_178_375 ();
 sg13g2_fill_8 FILLER_178_383 ();
 sg13g2_fill_8 FILLER_178_391 ();
 sg13g2_fill_8 FILLER_178_399 ();
 sg13g2_fill_1 FILLER_178_407 ();
 sg13g2_fill_8 FILLER_178_416 ();
 sg13g2_fill_8 FILLER_178_424 ();
 sg13g2_fill_8 FILLER_178_432 ();
 sg13g2_fill_8 FILLER_178_440 ();
 sg13g2_fill_8 FILLER_178_448 ();
 sg13g2_fill_8 FILLER_178_456 ();
 sg13g2_fill_8 FILLER_178_464 ();
 sg13g2_fill_8 FILLER_178_472 ();
 sg13g2_fill_8 FILLER_178_480 ();
 sg13g2_fill_4 FILLER_178_488 ();
 sg13g2_fill_2 FILLER_178_518 ();
 sg13g2_fill_1 FILLER_178_520 ();
 sg13g2_fill_2 FILLER_178_547 ();
 sg13g2_fill_1 FILLER_178_549 ();
 sg13g2_fill_8 FILLER_178_589 ();
 sg13g2_fill_8 FILLER_178_597 ();
 sg13g2_fill_8 FILLER_178_605 ();
 sg13g2_fill_4 FILLER_178_613 ();
 sg13g2_fill_8 FILLER_178_635 ();
 sg13g2_fill_4 FILLER_178_669 ();
 sg13g2_fill_2 FILLER_178_673 ();
 sg13g2_fill_8 FILLER_178_710 ();
 sg13g2_fill_8 FILLER_178_718 ();
 sg13g2_fill_8 FILLER_178_726 ();
 sg13g2_fill_8 FILLER_178_734 ();
 sg13g2_fill_4 FILLER_178_762 ();
 sg13g2_fill_2 FILLER_178_766 ();
 sg13g2_fill_1 FILLER_178_768 ();
 sg13g2_fill_4 FILLER_178_784 ();
 sg13g2_fill_2 FILLER_178_788 ();
 sg13g2_fill_1 FILLER_178_790 ();
 sg13g2_fill_2 FILLER_178_811 ();
 sg13g2_fill_8 FILLER_178_839 ();
 sg13g2_fill_8 FILLER_178_847 ();
 sg13g2_fill_8 FILLER_178_855 ();
 sg13g2_fill_8 FILLER_178_863 ();
 sg13g2_fill_8 FILLER_178_871 ();
 sg13g2_fill_8 FILLER_178_879 ();
 sg13g2_fill_8 FILLER_178_887 ();
 sg13g2_fill_8 FILLER_178_895 ();
 sg13g2_fill_8 FILLER_178_903 ();
 sg13g2_fill_8 FILLER_178_911 ();
 sg13g2_fill_8 FILLER_178_919 ();
 sg13g2_fill_8 FILLER_178_927 ();
 sg13g2_fill_8 FILLER_178_935 ();
 sg13g2_fill_8 FILLER_178_943 ();
 sg13g2_fill_8 FILLER_178_951 ();
 sg13g2_fill_8 FILLER_178_959 ();
 sg13g2_fill_4 FILLER_178_967 ();
 sg13g2_fill_2 FILLER_178_971 ();
 sg13g2_fill_1 FILLER_178_973 ();
 sg13g2_fill_4 FILLER_178_984 ();
 sg13g2_fill_1 FILLER_178_988 ();
 sg13g2_fill_2 FILLER_178_999 ();
 sg13g2_fill_1 FILLER_178_1001 ();
 sg13g2_fill_8 FILLER_178_1008 ();
 sg13g2_fill_4 FILLER_178_1016 ();
 sg13g2_fill_1 FILLER_178_1020 ();
 sg13g2_fill_4 FILLER_178_1039 ();
 sg13g2_fill_2 FILLER_178_1043 ();
 sg13g2_fill_8 FILLER_178_1053 ();
 sg13g2_fill_8 FILLER_178_1061 ();
 sg13g2_fill_4 FILLER_178_1069 ();
 sg13g2_fill_2 FILLER_178_1073 ();
 sg13g2_fill_8 FILLER_178_1083 ();
 sg13g2_fill_1 FILLER_178_1091 ();
 sg13g2_fill_8 FILLER_178_1104 ();
 sg13g2_fill_4 FILLER_178_1112 ();
 sg13g2_fill_2 FILLER_178_1116 ();
 sg13g2_fill_1 FILLER_178_1118 ();
 sg13g2_fill_8 FILLER_178_1140 ();
 sg13g2_fill_2 FILLER_178_1148 ();
 sg13g2_fill_4 FILLER_178_1161 ();
 sg13g2_fill_2 FILLER_178_1165 ();
 sg13g2_fill_1 FILLER_178_1167 ();
 sg13g2_fill_8 FILLER_178_1173 ();
 sg13g2_fill_1 FILLER_178_1181 ();
 sg13g2_fill_8 FILLER_178_1187 ();
 sg13g2_fill_8 FILLER_178_1195 ();
 sg13g2_fill_4 FILLER_178_1203 ();
 sg13g2_fill_8 FILLER_178_1228 ();
 sg13g2_fill_4 FILLER_178_1236 ();
 sg13g2_fill_2 FILLER_178_1240 ();
 sg13g2_fill_1 FILLER_178_1242 ();
 sg13g2_fill_4 FILLER_178_1259 ();
 sg13g2_fill_1 FILLER_178_1263 ();
 sg13g2_fill_4 FILLER_178_1286 ();
 sg13g2_fill_2 FILLER_178_1290 ();
 sg13g2_fill_1 FILLER_178_1292 ();
 sg13g2_fill_8 FILLER_178_1306 ();
 sg13g2_fill_1 FILLER_178_1314 ();
 sg13g2_fill_8 FILLER_178_1323 ();
 sg13g2_fill_2 FILLER_178_1331 ();
 sg13g2_fill_8 FILLER_178_1361 ();
 sg13g2_fill_8 FILLER_178_1369 ();
 sg13g2_fill_8 FILLER_178_1377 ();
 sg13g2_fill_8 FILLER_178_1385 ();
 sg13g2_fill_8 FILLER_178_1393 ();
 sg13g2_fill_4 FILLER_178_1401 ();
 sg13g2_fill_2 FILLER_178_1405 ();
 sg13g2_fill_1 FILLER_178_1412 ();
 sg13g2_fill_4 FILLER_178_1418 ();
 sg13g2_fill_2 FILLER_178_1422 ();
 sg13g2_fill_1 FILLER_178_1424 ();
 sg13g2_fill_1 FILLER_178_1430 ();
 sg13g2_fill_8 FILLER_178_1440 ();
 sg13g2_fill_8 FILLER_178_1448 ();
 sg13g2_fill_8 FILLER_178_1456 ();
 sg13g2_fill_8 FILLER_178_1464 ();
 sg13g2_fill_8 FILLER_178_1472 ();
 sg13g2_fill_8 FILLER_178_1480 ();
 sg13g2_fill_8 FILLER_178_1488 ();
 sg13g2_fill_8 FILLER_178_1496 ();
 sg13g2_fill_8 FILLER_178_1504 ();
 sg13g2_fill_8 FILLER_178_1512 ();
 sg13g2_fill_8 FILLER_178_1520 ();
 sg13g2_fill_8 FILLER_178_1528 ();
 sg13g2_fill_8 FILLER_178_1536 ();
 sg13g2_fill_8 FILLER_178_1544 ();
 sg13g2_fill_8 FILLER_178_1552 ();
 sg13g2_fill_8 FILLER_178_1560 ();
 sg13g2_fill_8 FILLER_178_1568 ();
 sg13g2_fill_8 FILLER_178_1576 ();
 sg13g2_fill_8 FILLER_178_1584 ();
 sg13g2_fill_8 FILLER_179_0 ();
 sg13g2_fill_8 FILLER_179_8 ();
 sg13g2_fill_8 FILLER_179_16 ();
 sg13g2_fill_8 FILLER_179_24 ();
 sg13g2_fill_8 FILLER_179_32 ();
 sg13g2_fill_8 FILLER_179_40 ();
 sg13g2_fill_8 FILLER_179_48 ();
 sg13g2_fill_8 FILLER_179_56 ();
 sg13g2_fill_8 FILLER_179_64 ();
 sg13g2_fill_8 FILLER_179_72 ();
 sg13g2_fill_8 FILLER_179_80 ();
 sg13g2_fill_8 FILLER_179_88 ();
 sg13g2_fill_8 FILLER_179_96 ();
 sg13g2_fill_8 FILLER_179_104 ();
 sg13g2_fill_4 FILLER_179_112 ();
 sg13g2_fill_8 FILLER_179_122 ();
 sg13g2_fill_2 FILLER_179_130 ();
 sg13g2_fill_1 FILLER_179_186 ();
 sg13g2_fill_2 FILLER_179_195 ();
 sg13g2_fill_1 FILLER_179_197 ();
 sg13g2_fill_8 FILLER_179_216 ();
 sg13g2_fill_4 FILLER_179_224 ();
 sg13g2_fill_1 FILLER_179_228 ();
 sg13g2_fill_8 FILLER_179_234 ();
 sg13g2_fill_8 FILLER_179_252 ();
 sg13g2_fill_8 FILLER_179_260 ();
 sg13g2_fill_8 FILLER_179_268 ();
 sg13g2_fill_8 FILLER_179_276 ();
 sg13g2_fill_8 FILLER_179_284 ();
 sg13g2_fill_8 FILLER_179_292 ();
 sg13g2_fill_4 FILLER_179_300 ();
 sg13g2_fill_2 FILLER_179_325 ();
 sg13g2_fill_1 FILLER_179_327 ();
 sg13g2_fill_8 FILLER_179_349 ();
 sg13g2_fill_4 FILLER_179_357 ();
 sg13g2_fill_2 FILLER_179_382 ();
 sg13g2_fill_8 FILLER_179_405 ();
 sg13g2_fill_8 FILLER_179_413 ();
 sg13g2_fill_8 FILLER_179_421 ();
 sg13g2_fill_8 FILLER_179_429 ();
 sg13g2_fill_8 FILLER_179_437 ();
 sg13g2_fill_8 FILLER_179_445 ();
 sg13g2_fill_8 FILLER_179_453 ();
 sg13g2_fill_8 FILLER_179_461 ();
 sg13g2_fill_8 FILLER_179_469 ();
 sg13g2_fill_8 FILLER_179_477 ();
 sg13g2_fill_8 FILLER_179_485 ();
 sg13g2_fill_8 FILLER_179_493 ();
 sg13g2_fill_8 FILLER_179_501 ();
 sg13g2_fill_2 FILLER_179_509 ();
 sg13g2_fill_8 FILLER_179_521 ();
 sg13g2_fill_4 FILLER_179_529 ();
 sg13g2_fill_1 FILLER_179_533 ();
 sg13g2_fill_8 FILLER_179_567 ();
 sg13g2_fill_8 FILLER_179_575 ();
 sg13g2_fill_4 FILLER_179_583 ();
 sg13g2_fill_2 FILLER_179_587 ();
 sg13g2_fill_1 FILLER_179_589 ();
 sg13g2_fill_8 FILLER_179_624 ();
 sg13g2_fill_4 FILLER_179_632 ();
 sg13g2_fill_2 FILLER_179_636 ();
 sg13g2_fill_1 FILLER_179_638 ();
 sg13g2_fill_4 FILLER_179_733 ();
 sg13g2_fill_4 FILLER_179_747 ();
 sg13g2_fill_2 FILLER_179_751 ();
 sg13g2_fill_2 FILLER_179_790 ();
 sg13g2_fill_1 FILLER_179_792 ();
 sg13g2_fill_8 FILLER_179_813 ();
 sg13g2_fill_8 FILLER_179_821 ();
 sg13g2_fill_8 FILLER_179_829 ();
 sg13g2_fill_8 FILLER_179_837 ();
 sg13g2_fill_8 FILLER_179_845 ();
 sg13g2_fill_8 FILLER_179_853 ();
 sg13g2_fill_8 FILLER_179_861 ();
 sg13g2_fill_8 FILLER_179_869 ();
 sg13g2_fill_8 FILLER_179_877 ();
 sg13g2_fill_8 FILLER_179_885 ();
 sg13g2_fill_8 FILLER_179_893 ();
 sg13g2_fill_8 FILLER_179_901 ();
 sg13g2_fill_8 FILLER_179_909 ();
 sg13g2_fill_8 FILLER_179_917 ();
 sg13g2_fill_8 FILLER_179_925 ();
 sg13g2_fill_8 FILLER_179_933 ();
 sg13g2_fill_8 FILLER_179_941 ();
 sg13g2_fill_8 FILLER_179_949 ();
 sg13g2_fill_8 FILLER_179_957 ();
 sg13g2_fill_8 FILLER_179_965 ();
 sg13g2_fill_1 FILLER_179_973 ();
 sg13g2_fill_2 FILLER_179_982 ();
 sg13g2_fill_1 FILLER_179_984 ();
 sg13g2_fill_8 FILLER_179_1011 ();
 sg13g2_fill_4 FILLER_179_1019 ();
 sg13g2_fill_2 FILLER_179_1023 ();
 sg13g2_fill_1 FILLER_179_1025 ();
 sg13g2_fill_8 FILLER_179_1047 ();
 sg13g2_fill_8 FILLER_179_1055 ();
 sg13g2_fill_8 FILLER_179_1063 ();
 sg13g2_fill_4 FILLER_179_1071 ();
 sg13g2_fill_2 FILLER_179_1075 ();
 sg13g2_fill_1 FILLER_179_1077 ();
 sg13g2_fill_2 FILLER_179_1086 ();
 sg13g2_fill_1 FILLER_179_1088 ();
 sg13g2_fill_4 FILLER_179_1103 ();
 sg13g2_fill_1 FILLER_179_1107 ();
 sg13g2_fill_4 FILLER_179_1113 ();
 sg13g2_fill_2 FILLER_179_1117 ();
 sg13g2_fill_4 FILLER_179_1149 ();
 sg13g2_fill_4 FILLER_179_1161 ();
 sg13g2_fill_1 FILLER_179_1173 ();
 sg13g2_fill_2 FILLER_179_1182 ();
 sg13g2_fill_1 FILLER_179_1184 ();
 sg13g2_fill_8 FILLER_179_1190 ();
 sg13g2_fill_8 FILLER_179_1198 ();
 sg13g2_fill_2 FILLER_179_1206 ();
 sg13g2_fill_4 FILLER_179_1216 ();
 sg13g2_fill_2 FILLER_179_1241 ();
 sg13g2_fill_2 FILLER_179_1264 ();
 sg13g2_fill_1 FILLER_179_1287 ();
 sg13g2_fill_4 FILLER_179_1294 ();
 sg13g2_fill_2 FILLER_179_1298 ();
 sg13g2_fill_1 FILLER_179_1300 ();
 sg13g2_fill_8 FILLER_179_1309 ();
 sg13g2_fill_4 FILLER_179_1317 ();
 sg13g2_fill_2 FILLER_179_1321 ();
 sg13g2_fill_8 FILLER_179_1339 ();
 sg13g2_fill_4 FILLER_179_1347 ();
 sg13g2_fill_2 FILLER_179_1361 ();
 sg13g2_fill_1 FILLER_179_1367 ();
 sg13g2_fill_4 FILLER_179_1373 ();
 sg13g2_fill_2 FILLER_179_1385 ();
 sg13g2_fill_1 FILLER_179_1387 ();
 sg13g2_fill_1 FILLER_179_1392 ();
 sg13g2_fill_4 FILLER_179_1398 ();
 sg13g2_fill_1 FILLER_179_1430 ();
 sg13g2_fill_8 FILLER_179_1451 ();
 sg13g2_fill_8 FILLER_179_1459 ();
 sg13g2_fill_8 FILLER_179_1467 ();
 sg13g2_fill_8 FILLER_179_1475 ();
 sg13g2_fill_8 FILLER_179_1483 ();
 sg13g2_fill_8 FILLER_179_1491 ();
 sg13g2_fill_8 FILLER_179_1499 ();
 sg13g2_fill_8 FILLER_179_1507 ();
 sg13g2_fill_8 FILLER_179_1515 ();
 sg13g2_fill_8 FILLER_179_1523 ();
 sg13g2_fill_8 FILLER_179_1531 ();
 sg13g2_fill_8 FILLER_179_1539 ();
 sg13g2_fill_8 FILLER_179_1547 ();
 sg13g2_fill_8 FILLER_179_1555 ();
 sg13g2_fill_8 FILLER_179_1563 ();
 sg13g2_fill_8 FILLER_179_1571 ();
 sg13g2_fill_8 FILLER_179_1579 ();
 sg13g2_fill_4 FILLER_179_1587 ();
 sg13g2_fill_1 FILLER_179_1591 ();
 sg13g2_fill_8 FILLER_180_0 ();
 sg13g2_fill_8 FILLER_180_8 ();
 sg13g2_fill_8 FILLER_180_16 ();
 sg13g2_fill_8 FILLER_180_24 ();
 sg13g2_fill_8 FILLER_180_32 ();
 sg13g2_fill_8 FILLER_180_40 ();
 sg13g2_fill_8 FILLER_180_48 ();
 sg13g2_fill_8 FILLER_180_56 ();
 sg13g2_fill_8 FILLER_180_64 ();
 sg13g2_fill_8 FILLER_180_72 ();
 sg13g2_fill_8 FILLER_180_80 ();
 sg13g2_fill_8 FILLER_180_88 ();
 sg13g2_fill_4 FILLER_180_96 ();
 sg13g2_fill_1 FILLER_180_100 ();
 sg13g2_fill_2 FILLER_180_173 ();
 sg13g2_fill_4 FILLER_180_201 ();
 sg13g2_fill_2 FILLER_180_205 ();
 sg13g2_fill_8 FILLER_180_236 ();
 sg13g2_fill_8 FILLER_180_244 ();
 sg13g2_fill_4 FILLER_180_262 ();
 sg13g2_fill_1 FILLER_180_266 ();
 sg13g2_fill_4 FILLER_180_297 ();
 sg13g2_fill_2 FILLER_180_301 ();
 sg13g2_fill_1 FILLER_180_303 ();
 sg13g2_fill_8 FILLER_180_325 ();
 sg13g2_fill_4 FILLER_180_333 ();
 sg13g2_fill_1 FILLER_180_337 ();
 sg13g2_fill_1 FILLER_180_369 ();
 sg13g2_fill_4 FILLER_180_380 ();
 sg13g2_fill_8 FILLER_180_410 ();
 sg13g2_fill_8 FILLER_180_418 ();
 sg13g2_fill_8 FILLER_180_426 ();
 sg13g2_fill_8 FILLER_180_434 ();
 sg13g2_fill_8 FILLER_180_442 ();
 sg13g2_fill_8 FILLER_180_450 ();
 sg13g2_fill_8 FILLER_180_458 ();
 sg13g2_fill_8 FILLER_180_466 ();
 sg13g2_fill_8 FILLER_180_474 ();
 sg13g2_fill_8 FILLER_180_482 ();
 sg13g2_fill_8 FILLER_180_490 ();
 sg13g2_fill_8 FILLER_180_498 ();
 sg13g2_fill_8 FILLER_180_506 ();
 sg13g2_fill_4 FILLER_180_514 ();
 sg13g2_fill_8 FILLER_180_528 ();
 sg13g2_fill_8 FILLER_180_536 ();
 sg13g2_fill_4 FILLER_180_544 ();
 sg13g2_fill_1 FILLER_180_548 ();
 sg13g2_fill_8 FILLER_180_559 ();
 sg13g2_fill_4 FILLER_180_567 ();
 sg13g2_fill_2 FILLER_180_571 ();
 sg13g2_fill_1 FILLER_180_573 ();
 sg13g2_fill_8 FILLER_180_595 ();
 sg13g2_fill_8 FILLER_180_603 ();
 sg13g2_fill_2 FILLER_180_611 ();
 sg13g2_fill_1 FILLER_180_613 ();
 sg13g2_fill_8 FILLER_180_624 ();
 sg13g2_fill_4 FILLER_180_632 ();
 sg13g2_fill_4 FILLER_180_646 ();
 sg13g2_fill_2 FILLER_180_650 ();
 sg13g2_fill_4 FILLER_180_656 ();
 sg13g2_fill_2 FILLER_180_660 ();
 sg13g2_fill_2 FILLER_180_670 ();
 sg13g2_fill_4 FILLER_180_708 ();
 sg13g2_fill_2 FILLER_180_712 ();
 sg13g2_fill_2 FILLER_180_750 ();
 sg13g2_fill_4 FILLER_180_763 ();
 sg13g2_fill_2 FILLER_180_767 ();
 sg13g2_fill_1 FILLER_180_769 ();
 sg13g2_fill_2 FILLER_180_780 ();
 sg13g2_fill_1 FILLER_180_782 ();
 sg13g2_fill_2 FILLER_180_793 ();
 sg13g2_fill_8 FILLER_180_805 ();
 sg13g2_fill_4 FILLER_180_813 ();
 sg13g2_fill_2 FILLER_180_817 ();
 sg13g2_fill_8 FILLER_180_848 ();
 sg13g2_fill_8 FILLER_180_856 ();
 sg13g2_fill_8 FILLER_180_864 ();
 sg13g2_fill_8 FILLER_180_872 ();
 sg13g2_fill_8 FILLER_180_880 ();
 sg13g2_fill_8 FILLER_180_888 ();
 sg13g2_fill_8 FILLER_180_896 ();
 sg13g2_fill_8 FILLER_180_904 ();
 sg13g2_fill_8 FILLER_180_912 ();
 sg13g2_fill_8 FILLER_180_920 ();
 sg13g2_fill_8 FILLER_180_928 ();
 sg13g2_fill_8 FILLER_180_936 ();
 sg13g2_fill_8 FILLER_180_944 ();
 sg13g2_fill_8 FILLER_180_952 ();
 sg13g2_fill_8 FILLER_180_960 ();
 sg13g2_fill_8 FILLER_180_968 ();
 sg13g2_fill_2 FILLER_180_976 ();
 sg13g2_fill_4 FILLER_180_1001 ();
 sg13g2_fill_1 FILLER_180_1005 ();
 sg13g2_fill_8 FILLER_180_1014 ();
 sg13g2_fill_8 FILLER_180_1022 ();
 sg13g2_fill_1 FILLER_180_1030 ();
 sg13g2_fill_2 FILLER_180_1035 ();
 sg13g2_fill_8 FILLER_180_1040 ();
 sg13g2_fill_4 FILLER_180_1048 ();
 sg13g2_fill_1 FILLER_180_1068 ();
 sg13g2_fill_8 FILLER_180_1088 ();
 sg13g2_fill_4 FILLER_180_1096 ();
 sg13g2_fill_1 FILLER_180_1109 ();
 sg13g2_fill_4 FILLER_180_1121 ();
 sg13g2_fill_2 FILLER_180_1125 ();
 sg13g2_fill_1 FILLER_180_1127 ();
 sg13g2_fill_4 FILLER_180_1138 ();
 sg13g2_fill_1 FILLER_180_1142 ();
 sg13g2_fill_2 FILLER_180_1151 ();
 sg13g2_fill_8 FILLER_180_1161 ();
 sg13g2_fill_8 FILLER_180_1169 ();
 sg13g2_fill_4 FILLER_180_1177 ();
 sg13g2_fill_1 FILLER_180_1181 ();
 sg13g2_fill_4 FILLER_180_1197 ();
 sg13g2_fill_1 FILLER_180_1201 ();
 sg13g2_fill_4 FILLER_180_1218 ();
 sg13g2_fill_2 FILLER_180_1222 ();
 sg13g2_fill_1 FILLER_180_1232 ();
 sg13g2_fill_8 FILLER_180_1262 ();
 sg13g2_fill_4 FILLER_180_1270 ();
 sg13g2_fill_2 FILLER_180_1274 ();
 sg13g2_fill_1 FILLER_180_1276 ();
 sg13g2_fill_4 FILLER_180_1291 ();
 sg13g2_fill_2 FILLER_180_1295 ();
 sg13g2_fill_1 FILLER_180_1297 ();
 sg13g2_fill_8 FILLER_180_1304 ();
 sg13g2_fill_2 FILLER_180_1312 ();
 sg13g2_fill_1 FILLER_180_1314 ();
 sg13g2_fill_8 FILLER_180_1331 ();
 sg13g2_fill_8 FILLER_180_1339 ();
 sg13g2_fill_1 FILLER_180_1347 ();
 sg13g2_fill_2 FILLER_180_1364 ();
 sg13g2_fill_4 FILLER_180_1382 ();
 sg13g2_fill_8 FILLER_180_1398 ();
 sg13g2_fill_4 FILLER_180_1406 ();
 sg13g2_fill_2 FILLER_180_1410 ();
 sg13g2_fill_1 FILLER_180_1412 ();
 sg13g2_fill_8 FILLER_180_1416 ();
 sg13g2_fill_4 FILLER_180_1424 ();
 sg13g2_fill_1 FILLER_180_1433 ();
 sg13g2_fill_8 FILLER_180_1446 ();
 sg13g2_fill_8 FILLER_180_1454 ();
 sg13g2_fill_8 FILLER_180_1462 ();
 sg13g2_fill_8 FILLER_180_1470 ();
 sg13g2_fill_8 FILLER_180_1478 ();
 sg13g2_fill_8 FILLER_180_1486 ();
 sg13g2_fill_8 FILLER_180_1494 ();
 sg13g2_fill_8 FILLER_180_1502 ();
 sg13g2_fill_8 FILLER_180_1510 ();
 sg13g2_fill_8 FILLER_180_1518 ();
 sg13g2_fill_8 FILLER_180_1526 ();
 sg13g2_fill_8 FILLER_180_1534 ();
 sg13g2_fill_8 FILLER_180_1542 ();
 sg13g2_fill_8 FILLER_180_1550 ();
 sg13g2_fill_8 FILLER_180_1558 ();
 sg13g2_fill_8 FILLER_180_1566 ();
 sg13g2_fill_8 FILLER_180_1574 ();
 sg13g2_fill_8 FILLER_180_1582 ();
 sg13g2_fill_2 FILLER_180_1590 ();
 sg13g2_fill_8 FILLER_181_0 ();
 sg13g2_fill_8 FILLER_181_8 ();
 sg13g2_fill_8 FILLER_181_16 ();
 sg13g2_fill_8 FILLER_181_24 ();
 sg13g2_fill_8 FILLER_181_32 ();
 sg13g2_fill_8 FILLER_181_40 ();
 sg13g2_fill_8 FILLER_181_48 ();
 sg13g2_fill_8 FILLER_181_56 ();
 sg13g2_fill_8 FILLER_181_64 ();
 sg13g2_fill_8 FILLER_181_72 ();
 sg13g2_fill_8 FILLER_181_80 ();
 sg13g2_fill_8 FILLER_181_88 ();
 sg13g2_fill_8 FILLER_181_96 ();
 sg13g2_fill_8 FILLER_181_104 ();
 sg13g2_fill_4 FILLER_181_112 ();
 sg13g2_fill_8 FILLER_181_141 ();
 sg13g2_fill_8 FILLER_181_149 ();
 sg13g2_fill_1 FILLER_181_167 ();
 sg13g2_fill_8 FILLER_181_204 ();
 sg13g2_fill_8 FILLER_181_212 ();
 sg13g2_fill_2 FILLER_181_220 ();
 sg13g2_fill_4 FILLER_181_274 ();
 sg13g2_fill_2 FILLER_181_278 ();
 sg13g2_fill_1 FILLER_181_280 ();
 sg13g2_fill_8 FILLER_181_317 ();
 sg13g2_fill_1 FILLER_181_325 ();
 sg13g2_fill_8 FILLER_181_334 ();
 sg13g2_fill_8 FILLER_181_342 ();
 sg13g2_fill_8 FILLER_181_350 ();
 sg13g2_fill_4 FILLER_181_358 ();
 sg13g2_fill_2 FILLER_181_362 ();
 sg13g2_fill_1 FILLER_181_364 ();
 sg13g2_fill_8 FILLER_181_391 ();
 sg13g2_fill_8 FILLER_181_399 ();
 sg13g2_fill_8 FILLER_181_407 ();
 sg13g2_fill_8 FILLER_181_415 ();
 sg13g2_fill_8 FILLER_181_423 ();
 sg13g2_fill_8 FILLER_181_431 ();
 sg13g2_fill_8 FILLER_181_439 ();
 sg13g2_fill_8 FILLER_181_447 ();
 sg13g2_fill_8 FILLER_181_455 ();
 sg13g2_fill_8 FILLER_181_463 ();
 sg13g2_fill_8 FILLER_181_471 ();
 sg13g2_fill_8 FILLER_181_479 ();
 sg13g2_fill_8 FILLER_181_487 ();
 sg13g2_fill_8 FILLER_181_495 ();
 sg13g2_fill_1 FILLER_181_503 ();
 sg13g2_fill_8 FILLER_181_514 ();
 sg13g2_fill_2 FILLER_181_548 ();
 sg13g2_fill_1 FILLER_181_550 ();
 sg13g2_fill_8 FILLER_181_577 ();
 sg13g2_fill_4 FILLER_181_605 ();
 sg13g2_fill_2 FILLER_181_609 ();
 sg13g2_fill_4 FILLER_181_621 ();
 sg13g2_fill_2 FILLER_181_625 ();
 sg13g2_fill_1 FILLER_181_627 ();
 sg13g2_fill_8 FILLER_181_674 ();
 sg13g2_fill_2 FILLER_181_682 ();
 sg13g2_fill_1 FILLER_181_684 ();
 sg13g2_fill_8 FILLER_181_695 ();
 sg13g2_fill_2 FILLER_181_703 ();
 sg13g2_fill_1 FILLER_181_705 ();
 sg13g2_fill_8 FILLER_181_716 ();
 sg13g2_fill_8 FILLER_181_724 ();
 sg13g2_fill_8 FILLER_181_742 ();
 sg13g2_fill_2 FILLER_181_750 ();
 sg13g2_fill_8 FILLER_181_762 ();
 sg13g2_fill_8 FILLER_181_770 ();
 sg13g2_fill_8 FILLER_181_778 ();
 sg13g2_fill_8 FILLER_181_786 ();
 sg13g2_fill_2 FILLER_181_804 ();
 sg13g2_fill_8 FILLER_181_832 ();
 sg13g2_fill_8 FILLER_181_840 ();
 sg13g2_fill_8 FILLER_181_848 ();
 sg13g2_fill_8 FILLER_181_856 ();
 sg13g2_fill_8 FILLER_181_864 ();
 sg13g2_fill_8 FILLER_181_872 ();
 sg13g2_fill_8 FILLER_181_880 ();
 sg13g2_fill_8 FILLER_181_888 ();
 sg13g2_fill_8 FILLER_181_896 ();
 sg13g2_fill_8 FILLER_181_904 ();
 sg13g2_fill_8 FILLER_181_912 ();
 sg13g2_fill_8 FILLER_181_920 ();
 sg13g2_fill_8 FILLER_181_928 ();
 sg13g2_fill_8 FILLER_181_936 ();
 sg13g2_fill_8 FILLER_181_944 ();
 sg13g2_fill_8 FILLER_181_952 ();
 sg13g2_fill_8 FILLER_181_960 ();
 sg13g2_fill_8 FILLER_181_968 ();
 sg13g2_fill_8 FILLER_181_976 ();
 sg13g2_fill_1 FILLER_181_984 ();
 sg13g2_fill_8 FILLER_181_994 ();
 sg13g2_fill_2 FILLER_181_1025 ();
 sg13g2_fill_1 FILLER_181_1027 ();
 sg13g2_fill_8 FILLER_181_1031 ();
 sg13g2_fill_8 FILLER_181_1039 ();
 sg13g2_fill_4 FILLER_181_1047 ();
 sg13g2_fill_2 FILLER_181_1051 ();
 sg13g2_fill_8 FILLER_181_1061 ();
 sg13g2_fill_4 FILLER_181_1069 ();
 sg13g2_fill_1 FILLER_181_1073 ();
 sg13g2_fill_2 FILLER_181_1080 ();
 sg13g2_fill_8 FILLER_181_1090 ();
 sg13g2_fill_8 FILLER_181_1118 ();
 sg13g2_fill_1 FILLER_181_1126 ();
 sg13g2_fill_8 FILLER_181_1132 ();
 sg13g2_fill_8 FILLER_181_1140 ();
 sg13g2_fill_8 FILLER_181_1148 ();
 sg13g2_fill_1 FILLER_181_1156 ();
 sg13g2_fill_8 FILLER_181_1162 ();
 sg13g2_fill_2 FILLER_181_1175 ();
 sg13g2_fill_8 FILLER_181_1185 ();
 sg13g2_fill_2 FILLER_181_1193 ();
 sg13g2_fill_1 FILLER_181_1195 ();
 sg13g2_fill_1 FILLER_181_1220 ();
 sg13g2_fill_8 FILLER_181_1237 ();
 sg13g2_fill_8 FILLER_181_1245 ();
 sg13g2_fill_8 FILLER_181_1253 ();
 sg13g2_fill_4 FILLER_181_1261 ();
 sg13g2_fill_2 FILLER_181_1265 ();
 sg13g2_fill_1 FILLER_181_1267 ();
 sg13g2_fill_8 FILLER_181_1273 ();
 sg13g2_fill_4 FILLER_181_1285 ();
 sg13g2_fill_2 FILLER_181_1289 ();
 sg13g2_fill_1 FILLER_181_1291 ();
 sg13g2_fill_4 FILLER_181_1300 ();
 sg13g2_fill_2 FILLER_181_1304 ();
 sg13g2_fill_1 FILLER_181_1306 ();
 sg13g2_fill_8 FILLER_181_1315 ();
 sg13g2_fill_8 FILLER_181_1328 ();
 sg13g2_fill_4 FILLER_181_1365 ();
 sg13g2_fill_2 FILLER_181_1369 ();
 sg13g2_fill_1 FILLER_181_1371 ();
 sg13g2_fill_8 FILLER_181_1380 ();
 sg13g2_fill_8 FILLER_181_1404 ();
 sg13g2_fill_8 FILLER_181_1412 ();
 sg13g2_fill_8 FILLER_181_1420 ();
 sg13g2_fill_8 FILLER_181_1445 ();
 sg13g2_fill_8 FILLER_181_1453 ();
 sg13g2_fill_8 FILLER_181_1461 ();
 sg13g2_fill_8 FILLER_181_1469 ();
 sg13g2_fill_8 FILLER_181_1477 ();
 sg13g2_fill_8 FILLER_181_1485 ();
 sg13g2_fill_8 FILLER_181_1493 ();
 sg13g2_fill_8 FILLER_181_1501 ();
 sg13g2_fill_8 FILLER_181_1509 ();
 sg13g2_fill_8 FILLER_181_1517 ();
 sg13g2_fill_8 FILLER_181_1525 ();
 sg13g2_fill_8 FILLER_181_1533 ();
 sg13g2_fill_8 FILLER_181_1541 ();
 sg13g2_fill_8 FILLER_181_1549 ();
 sg13g2_fill_8 FILLER_181_1557 ();
 sg13g2_fill_8 FILLER_181_1565 ();
 sg13g2_fill_8 FILLER_181_1573 ();
 sg13g2_fill_8 FILLER_181_1581 ();
 sg13g2_fill_2 FILLER_181_1589 ();
 sg13g2_fill_1 FILLER_181_1591 ();
 sg13g2_fill_8 FILLER_182_0 ();
 sg13g2_fill_8 FILLER_182_8 ();
 sg13g2_fill_8 FILLER_182_16 ();
 sg13g2_fill_8 FILLER_182_24 ();
 sg13g2_fill_8 FILLER_182_32 ();
 sg13g2_fill_8 FILLER_182_40 ();
 sg13g2_fill_8 FILLER_182_48 ();
 sg13g2_fill_8 FILLER_182_56 ();
 sg13g2_fill_8 FILLER_182_64 ();
 sg13g2_fill_8 FILLER_182_72 ();
 sg13g2_fill_8 FILLER_182_80 ();
 sg13g2_fill_8 FILLER_182_88 ();
 sg13g2_fill_8 FILLER_182_96 ();
 sg13g2_fill_8 FILLER_182_104 ();
 sg13g2_fill_4 FILLER_182_112 ();
 sg13g2_fill_2 FILLER_182_116 ();
 sg13g2_fill_8 FILLER_182_126 ();
 sg13g2_fill_4 FILLER_182_134 ();
 sg13g2_fill_8 FILLER_182_197 ();
 sg13g2_fill_1 FILLER_182_205 ();
 sg13g2_fill_4 FILLER_182_216 ();
 sg13g2_fill_1 FILLER_182_220 ();
 sg13g2_fill_8 FILLER_182_256 ();
 sg13g2_fill_4 FILLER_182_264 ();
 sg13g2_fill_1 FILLER_182_268 ();
 sg13g2_fill_8 FILLER_182_304 ();
 sg13g2_fill_8 FILLER_182_312 ();
 sg13g2_fill_4 FILLER_182_320 ();
 sg13g2_fill_2 FILLER_182_360 ();
 sg13g2_fill_8 FILLER_182_388 ();
 sg13g2_fill_8 FILLER_182_396 ();
 sg13g2_fill_8 FILLER_182_404 ();
 sg13g2_fill_8 FILLER_182_412 ();
 sg13g2_fill_8 FILLER_182_420 ();
 sg13g2_fill_8 FILLER_182_428 ();
 sg13g2_fill_8 FILLER_182_436 ();
 sg13g2_fill_8 FILLER_182_444 ();
 sg13g2_fill_8 FILLER_182_452 ();
 sg13g2_fill_8 FILLER_182_460 ();
 sg13g2_fill_8 FILLER_182_468 ();
 sg13g2_fill_8 FILLER_182_476 ();
 sg13g2_fill_8 FILLER_182_484 ();
 sg13g2_fill_2 FILLER_182_492 ();
 sg13g2_fill_1 FILLER_182_494 ();
 sg13g2_fill_2 FILLER_182_521 ();
 sg13g2_fill_8 FILLER_182_553 ();
 sg13g2_fill_1 FILLER_182_561 ();
 sg13g2_fill_2 FILLER_182_570 ();
 sg13g2_fill_1 FILLER_182_572 ();
 sg13g2_fill_4 FILLER_182_625 ();
 sg13g2_fill_4 FILLER_182_639 ();
 sg13g2_fill_2 FILLER_182_643 ();
 sg13g2_fill_1 FILLER_182_645 ();
 sg13g2_fill_8 FILLER_182_656 ();
 sg13g2_fill_8 FILLER_182_664 ();
 sg13g2_fill_8 FILLER_182_672 ();
 sg13g2_fill_2 FILLER_182_680 ();
 sg13g2_fill_1 FILLER_182_682 ();
 sg13g2_fill_2 FILLER_182_709 ();
 sg13g2_fill_4 FILLER_182_737 ();
 sg13g2_fill_2 FILLER_182_741 ();
 sg13g2_fill_1 FILLER_182_743 ();
 sg13g2_fill_8 FILLER_182_770 ();
 sg13g2_fill_8 FILLER_182_778 ();
 sg13g2_fill_2 FILLER_182_786 ();
 sg13g2_fill_8 FILLER_182_808 ();
 sg13g2_fill_8 FILLER_182_816 ();
 sg13g2_fill_8 FILLER_182_824 ();
 sg13g2_fill_8 FILLER_182_832 ();
 sg13g2_fill_8 FILLER_182_840 ();
 sg13g2_fill_8 FILLER_182_848 ();
 sg13g2_fill_8 FILLER_182_856 ();
 sg13g2_fill_8 FILLER_182_864 ();
 sg13g2_fill_8 FILLER_182_872 ();
 sg13g2_fill_8 FILLER_182_880 ();
 sg13g2_fill_8 FILLER_182_888 ();
 sg13g2_fill_8 FILLER_182_896 ();
 sg13g2_fill_8 FILLER_182_904 ();
 sg13g2_fill_8 FILLER_182_912 ();
 sg13g2_fill_8 FILLER_182_920 ();
 sg13g2_fill_8 FILLER_182_928 ();
 sg13g2_fill_8 FILLER_182_936 ();
 sg13g2_fill_8 FILLER_182_944 ();
 sg13g2_fill_8 FILLER_182_952 ();
 sg13g2_fill_8 FILLER_182_960 ();
 sg13g2_fill_8 FILLER_182_968 ();
 sg13g2_fill_2 FILLER_182_976 ();
 sg13g2_fill_8 FILLER_182_984 ();
 sg13g2_fill_4 FILLER_182_992 ();
 sg13g2_fill_2 FILLER_182_996 ();
 sg13g2_fill_1 FILLER_182_998 ();
 sg13g2_fill_1 FILLER_182_1021 ();
 sg13g2_fill_4 FILLER_182_1048 ();
 sg13g2_fill_2 FILLER_182_1052 ();
 sg13g2_fill_4 FILLER_182_1070 ();
 sg13g2_fill_2 FILLER_182_1074 ();
 sg13g2_fill_8 FILLER_182_1093 ();
 sg13g2_fill_8 FILLER_182_1109 ();
 sg13g2_fill_2 FILLER_182_1117 ();
 sg13g2_fill_1 FILLER_182_1119 ();
 sg13g2_fill_8 FILLER_182_1136 ();
 sg13g2_fill_4 FILLER_182_1144 ();
 sg13g2_fill_1 FILLER_182_1148 ();
 sg13g2_fill_1 FILLER_182_1165 ();
 sg13g2_fill_8 FILLER_182_1189 ();
 sg13g2_fill_4 FILLER_182_1202 ();
 sg13g2_fill_8 FILLER_182_1214 ();
 sg13g2_fill_8 FILLER_182_1222 ();
 sg13g2_fill_8 FILLER_182_1230 ();
 sg13g2_fill_8 FILLER_182_1238 ();
 sg13g2_fill_4 FILLER_182_1246 ();
 sg13g2_fill_2 FILLER_182_1250 ();
 sg13g2_fill_2 FILLER_182_1264 ();
 sg13g2_fill_4 FILLER_182_1280 ();
 sg13g2_fill_2 FILLER_182_1284 ();
 sg13g2_fill_1 FILLER_182_1286 ();
 sg13g2_fill_4 FILLER_182_1321 ();
 sg13g2_fill_4 FILLER_182_1341 ();
 sg13g2_fill_2 FILLER_182_1345 ();
 sg13g2_fill_8 FILLER_182_1353 ();
 sg13g2_fill_8 FILLER_182_1376 ();
 sg13g2_fill_8 FILLER_182_1384 ();
 sg13g2_fill_4 FILLER_182_1392 ();
 sg13g2_fill_2 FILLER_182_1404 ();
 sg13g2_fill_8 FILLER_182_1414 ();
 sg13g2_fill_2 FILLER_182_1422 ();
 sg13g2_fill_1 FILLER_182_1424 ();
 sg13g2_fill_8 FILLER_182_1448 ();
 sg13g2_fill_8 FILLER_182_1456 ();
 sg13g2_fill_8 FILLER_182_1464 ();
 sg13g2_fill_8 FILLER_182_1472 ();
 sg13g2_fill_8 FILLER_182_1480 ();
 sg13g2_fill_8 FILLER_182_1488 ();
 sg13g2_fill_8 FILLER_182_1496 ();
 sg13g2_fill_8 FILLER_182_1504 ();
 sg13g2_fill_8 FILLER_182_1512 ();
 sg13g2_fill_8 FILLER_182_1520 ();
 sg13g2_fill_8 FILLER_182_1528 ();
 sg13g2_fill_8 FILLER_182_1536 ();
 sg13g2_fill_8 FILLER_182_1544 ();
 sg13g2_fill_8 FILLER_182_1552 ();
 sg13g2_fill_8 FILLER_182_1560 ();
 sg13g2_fill_8 FILLER_182_1568 ();
 sg13g2_fill_8 FILLER_182_1576 ();
 sg13g2_fill_8 FILLER_182_1584 ();
 sg13g2_fill_8 FILLER_183_0 ();
 sg13g2_fill_8 FILLER_183_8 ();
 sg13g2_fill_8 FILLER_183_16 ();
 sg13g2_fill_8 FILLER_183_24 ();
 sg13g2_fill_8 FILLER_183_32 ();
 sg13g2_fill_8 FILLER_183_40 ();
 sg13g2_fill_8 FILLER_183_48 ();
 sg13g2_fill_8 FILLER_183_56 ();
 sg13g2_fill_8 FILLER_183_64 ();
 sg13g2_fill_8 FILLER_183_72 ();
 sg13g2_fill_8 FILLER_183_80 ();
 sg13g2_fill_8 FILLER_183_88 ();
 sg13g2_fill_8 FILLER_183_96 ();
 sg13g2_fill_8 FILLER_183_104 ();
 sg13g2_fill_8 FILLER_183_112 ();
 sg13g2_fill_8 FILLER_183_120 ();
 sg13g2_fill_8 FILLER_183_128 ();
 sg13g2_fill_8 FILLER_183_136 ();
 sg13g2_fill_8 FILLER_183_144 ();
 sg13g2_fill_8 FILLER_183_152 ();
 sg13g2_fill_8 FILLER_183_160 ();
 sg13g2_fill_4 FILLER_183_168 ();
 sg13g2_fill_1 FILLER_183_172 ();
 sg13g2_fill_4 FILLER_183_203 ();
 sg13g2_fill_1 FILLER_183_207 ();
 sg13g2_fill_4 FILLER_183_234 ();
 sg13g2_fill_1 FILLER_183_279 ();
 sg13g2_fill_4 FILLER_183_316 ();
 sg13g2_fill_2 FILLER_183_320 ();
 sg13g2_fill_1 FILLER_183_322 ();
 sg13g2_fill_8 FILLER_183_333 ();
 sg13g2_fill_4 FILLER_183_341 ();
 sg13g2_fill_2 FILLER_183_345 ();
 sg13g2_fill_1 FILLER_183_347 ();
 sg13g2_fill_8 FILLER_183_394 ();
 sg13g2_fill_8 FILLER_183_402 ();
 sg13g2_fill_8 FILLER_183_410 ();
 sg13g2_fill_8 FILLER_183_418 ();
 sg13g2_fill_8 FILLER_183_426 ();
 sg13g2_fill_8 FILLER_183_434 ();
 sg13g2_fill_8 FILLER_183_442 ();
 sg13g2_fill_8 FILLER_183_450 ();
 sg13g2_fill_8 FILLER_183_458 ();
 sg13g2_fill_8 FILLER_183_466 ();
 sg13g2_fill_8 FILLER_183_474 ();
 sg13g2_fill_8 FILLER_183_482 ();
 sg13g2_fill_8 FILLER_183_490 ();
 sg13g2_fill_8 FILLER_183_498 ();
 sg13g2_fill_2 FILLER_183_506 ();
 sg13g2_fill_2 FILLER_183_524 ();
 sg13g2_fill_8 FILLER_183_561 ();
 sg13g2_fill_4 FILLER_183_569 ();
 sg13g2_fill_8 FILLER_183_583 ();
 sg13g2_fill_1 FILLER_183_591 ();
 sg13g2_fill_8 FILLER_183_605 ();
 sg13g2_fill_8 FILLER_183_613 ();
 sg13g2_fill_4 FILLER_183_621 ();
 sg13g2_fill_8 FILLER_183_635 ();
 sg13g2_fill_4 FILLER_183_643 ();
 sg13g2_fill_1 FILLER_183_647 ();
 sg13g2_fill_8 FILLER_183_674 ();
 sg13g2_fill_8 FILLER_183_682 ();
 sg13g2_fill_8 FILLER_183_715 ();
 sg13g2_fill_8 FILLER_183_723 ();
 sg13g2_fill_8 FILLER_183_731 ();
 sg13g2_fill_8 FILLER_183_739 ();
 sg13g2_fill_8 FILLER_183_747 ();
 sg13g2_fill_2 FILLER_183_755 ();
 sg13g2_fill_2 FILLER_183_767 ();
 sg13g2_fill_1 FILLER_183_769 ();
 sg13g2_fill_4 FILLER_183_796 ();
 sg13g2_fill_2 FILLER_183_800 ();
 sg13g2_fill_1 FILLER_183_802 ();
 sg13g2_fill_8 FILLER_183_829 ();
 sg13g2_fill_8 FILLER_183_837 ();
 sg13g2_fill_8 FILLER_183_845 ();
 sg13g2_fill_8 FILLER_183_853 ();
 sg13g2_fill_8 FILLER_183_861 ();
 sg13g2_fill_8 FILLER_183_869 ();
 sg13g2_fill_8 FILLER_183_877 ();
 sg13g2_fill_8 FILLER_183_885 ();
 sg13g2_fill_8 FILLER_183_893 ();
 sg13g2_fill_8 FILLER_183_901 ();
 sg13g2_fill_8 FILLER_183_909 ();
 sg13g2_fill_8 FILLER_183_917 ();
 sg13g2_fill_8 FILLER_183_925 ();
 sg13g2_fill_8 FILLER_183_933 ();
 sg13g2_fill_8 FILLER_183_941 ();
 sg13g2_fill_8 FILLER_183_949 ();
 sg13g2_fill_8 FILLER_183_957 ();
 sg13g2_fill_8 FILLER_183_965 ();
 sg13g2_fill_4 FILLER_183_973 ();
 sg13g2_fill_1 FILLER_183_977 ();
 sg13g2_fill_4 FILLER_183_995 ();
 sg13g2_fill_2 FILLER_183_999 ();
 sg13g2_fill_2 FILLER_183_1009 ();
 sg13g2_fill_2 FILLER_183_1024 ();
 sg13g2_fill_1 FILLER_183_1026 ();
 sg13g2_fill_2 FILLER_183_1050 ();
 sg13g2_fill_1 FILLER_183_1052 ();
 sg13g2_fill_8 FILLER_183_1069 ();
 sg13g2_fill_1 FILLER_183_1077 ();
 sg13g2_fill_8 FILLER_183_1084 ();
 sg13g2_fill_4 FILLER_183_1092 ();
 sg13g2_fill_2 FILLER_183_1096 ();
 sg13g2_fill_1 FILLER_183_1098 ();
 sg13g2_fill_4 FILLER_183_1113 ();
 sg13g2_fill_2 FILLER_183_1146 ();
 sg13g2_fill_4 FILLER_183_1152 ();
 sg13g2_fill_1 FILLER_183_1156 ();
 sg13g2_fill_8 FILLER_183_1162 ();
 sg13g2_fill_2 FILLER_183_1170 ();
 sg13g2_fill_4 FILLER_183_1183 ();
 sg13g2_fill_2 FILLER_183_1192 ();
 sg13g2_fill_1 FILLER_183_1199 ();
 sg13g2_fill_8 FILLER_183_1206 ();
 sg13g2_fill_8 FILLER_183_1214 ();
 sg13g2_fill_8 FILLER_183_1230 ();
 sg13g2_fill_1 FILLER_183_1238 ();
 sg13g2_fill_2 FILLER_183_1247 ();
 sg13g2_fill_1 FILLER_183_1249 ();
 sg13g2_fill_4 FILLER_183_1261 ();
 sg13g2_fill_8 FILLER_183_1270 ();
 sg13g2_fill_8 FILLER_183_1278 ();
 sg13g2_fill_4 FILLER_183_1286 ();
 sg13g2_fill_1 FILLER_183_1290 ();
 sg13g2_fill_8 FILLER_183_1297 ();
 sg13g2_fill_1 FILLER_183_1309 ();
 sg13g2_fill_1 FILLER_183_1322 ();
 sg13g2_fill_4 FILLER_183_1327 ();
 sg13g2_fill_8 FILLER_183_1336 ();
 sg13g2_fill_4 FILLER_183_1344 ();
 sg13g2_fill_2 FILLER_183_1348 ();
 sg13g2_fill_4 FILLER_183_1382 ();
 sg13g2_fill_2 FILLER_183_1386 ();
 sg13g2_fill_1 FILLER_183_1388 ();
 sg13g2_fill_8 FILLER_183_1410 ();
 sg13g2_fill_8 FILLER_183_1418 ();
 sg13g2_fill_2 FILLER_183_1426 ();
 sg13g2_fill_2 FILLER_183_1433 ();
 sg13g2_fill_8 FILLER_183_1447 ();
 sg13g2_fill_8 FILLER_183_1455 ();
 sg13g2_fill_8 FILLER_183_1463 ();
 sg13g2_fill_8 FILLER_183_1471 ();
 sg13g2_fill_8 FILLER_183_1479 ();
 sg13g2_fill_8 FILLER_183_1487 ();
 sg13g2_fill_8 FILLER_183_1495 ();
 sg13g2_fill_8 FILLER_183_1503 ();
 sg13g2_fill_8 FILLER_183_1511 ();
 sg13g2_fill_8 FILLER_183_1519 ();
 sg13g2_fill_8 FILLER_183_1527 ();
 sg13g2_fill_8 FILLER_183_1535 ();
 sg13g2_fill_8 FILLER_183_1543 ();
 sg13g2_fill_8 FILLER_183_1551 ();
 sg13g2_fill_8 FILLER_183_1559 ();
 sg13g2_fill_8 FILLER_183_1567 ();
 sg13g2_fill_8 FILLER_183_1575 ();
 sg13g2_fill_8 FILLER_183_1583 ();
 sg13g2_fill_1 FILLER_183_1591 ();
 sg13g2_fill_8 FILLER_184_0 ();
 sg13g2_fill_8 FILLER_184_8 ();
 sg13g2_fill_8 FILLER_184_16 ();
 sg13g2_fill_8 FILLER_184_24 ();
 sg13g2_fill_8 FILLER_184_32 ();
 sg13g2_fill_8 FILLER_184_40 ();
 sg13g2_fill_8 FILLER_184_48 ();
 sg13g2_fill_8 FILLER_184_56 ();
 sg13g2_fill_8 FILLER_184_64 ();
 sg13g2_fill_8 FILLER_184_72 ();
 sg13g2_fill_8 FILLER_184_80 ();
 sg13g2_fill_8 FILLER_184_88 ();
 sg13g2_fill_8 FILLER_184_96 ();
 sg13g2_fill_8 FILLER_184_104 ();
 sg13g2_fill_8 FILLER_184_112 ();
 sg13g2_fill_8 FILLER_184_120 ();
 sg13g2_fill_8 FILLER_184_128 ();
 sg13g2_fill_8 FILLER_184_136 ();
 sg13g2_fill_8 FILLER_184_144 ();
 sg13g2_fill_4 FILLER_184_152 ();
 sg13g2_fill_2 FILLER_184_156 ();
 sg13g2_fill_8 FILLER_184_168 ();
 sg13g2_fill_4 FILLER_184_202 ();
 sg13g2_fill_1 FILLER_184_206 ();
 sg13g2_fill_4 FILLER_184_243 ();
 sg13g2_fill_2 FILLER_184_247 ();
 sg13g2_fill_1 FILLER_184_249 ();
 sg13g2_fill_4 FILLER_184_276 ();
 sg13g2_fill_1 FILLER_184_280 ();
 sg13g2_fill_4 FILLER_184_307 ();
 sg13g2_fill_4 FILLER_184_321 ();
 sg13g2_fill_2 FILLER_184_351 ();
 sg13g2_fill_8 FILLER_184_381 ();
 sg13g2_fill_8 FILLER_184_389 ();
 sg13g2_fill_8 FILLER_184_397 ();
 sg13g2_fill_8 FILLER_184_405 ();
 sg13g2_fill_8 FILLER_184_413 ();
 sg13g2_fill_8 FILLER_184_421 ();
 sg13g2_fill_8 FILLER_184_429 ();
 sg13g2_fill_8 FILLER_184_437 ();
 sg13g2_fill_8 FILLER_184_445 ();
 sg13g2_fill_8 FILLER_184_453 ();
 sg13g2_fill_8 FILLER_184_461 ();
 sg13g2_fill_8 FILLER_184_469 ();
 sg13g2_fill_8 FILLER_184_477 ();
 sg13g2_fill_8 FILLER_184_485 ();
 sg13g2_fill_8 FILLER_184_493 ();
 sg13g2_fill_8 FILLER_184_501 ();
 sg13g2_fill_8 FILLER_184_509 ();
 sg13g2_fill_4 FILLER_184_517 ();
 sg13g2_fill_2 FILLER_184_573 ();
 sg13g2_fill_4 FILLER_184_636 ();
 sg13g2_fill_4 FILLER_184_650 ();
 sg13g2_fill_1 FILLER_184_654 ();
 sg13g2_fill_8 FILLER_184_691 ();
 sg13g2_fill_8 FILLER_184_709 ();
 sg13g2_fill_2 FILLER_184_717 ();
 sg13g2_fill_4 FILLER_184_765 ();
 sg13g2_fill_4 FILLER_184_779 ();
 sg13g2_fill_2 FILLER_184_783 ();
 sg13g2_fill_1 FILLER_184_795 ();
 sg13g2_fill_8 FILLER_184_806 ();
 sg13g2_fill_8 FILLER_184_814 ();
 sg13g2_fill_8 FILLER_184_822 ();
 sg13g2_fill_8 FILLER_184_830 ();
 sg13g2_fill_8 FILLER_184_838 ();
 sg13g2_fill_8 FILLER_184_846 ();
 sg13g2_fill_8 FILLER_184_854 ();
 sg13g2_fill_8 FILLER_184_862 ();
 sg13g2_fill_8 FILLER_184_870 ();
 sg13g2_fill_8 FILLER_184_878 ();
 sg13g2_fill_8 FILLER_184_886 ();
 sg13g2_fill_8 FILLER_184_894 ();
 sg13g2_fill_8 FILLER_184_902 ();
 sg13g2_fill_8 FILLER_184_910 ();
 sg13g2_fill_8 FILLER_184_918 ();
 sg13g2_fill_8 FILLER_184_926 ();
 sg13g2_fill_8 FILLER_184_934 ();
 sg13g2_fill_8 FILLER_184_942 ();
 sg13g2_fill_8 FILLER_184_950 ();
 sg13g2_fill_8 FILLER_184_958 ();
 sg13g2_fill_4 FILLER_184_966 ();
 sg13g2_fill_8 FILLER_184_989 ();
 sg13g2_fill_8 FILLER_184_997 ();
 sg13g2_fill_8 FILLER_184_1005 ();
 sg13g2_fill_8 FILLER_184_1013 ();
 sg13g2_fill_2 FILLER_184_1021 ();
 sg13g2_fill_4 FILLER_184_1031 ();
 sg13g2_fill_1 FILLER_184_1040 ();
 sg13g2_fill_2 FILLER_184_1049 ();
 sg13g2_fill_1 FILLER_184_1051 ();
 sg13g2_fill_4 FILLER_184_1068 ();
 sg13g2_fill_2 FILLER_184_1084 ();
 sg13g2_fill_1 FILLER_184_1086 ();
 sg13g2_fill_8 FILLER_184_1095 ();
 sg13g2_fill_1 FILLER_184_1103 ();
 sg13g2_fill_8 FILLER_184_1110 ();
 sg13g2_fill_4 FILLER_184_1118 ();
 sg13g2_fill_1 FILLER_184_1122 ();
 sg13g2_fill_1 FILLER_184_1129 ();
 sg13g2_fill_8 FILLER_184_1135 ();
 sg13g2_fill_4 FILLER_184_1143 ();
 sg13g2_fill_8 FILLER_184_1152 ();
 sg13g2_fill_4 FILLER_184_1160 ();
 sg13g2_fill_2 FILLER_184_1164 ();
 sg13g2_fill_8 FILLER_184_1194 ();
 sg13g2_fill_2 FILLER_184_1202 ();
 sg13g2_fill_4 FILLER_184_1216 ();
 sg13g2_fill_2 FILLER_184_1220 ();
 sg13g2_fill_1 FILLER_184_1222 ();
 sg13g2_fill_2 FILLER_184_1237 ();
 sg13g2_fill_1 FILLER_184_1239 ();
 sg13g2_fill_8 FILLER_184_1256 ();
 sg13g2_fill_4 FILLER_184_1272 ();
 sg13g2_fill_8 FILLER_184_1300 ();
 sg13g2_fill_8 FILLER_184_1308 ();
 sg13g2_fill_2 FILLER_184_1316 ();
 sg13g2_fill_8 FILLER_184_1350 ();
 sg13g2_fill_8 FILLER_184_1358 ();
 sg13g2_fill_8 FILLER_184_1374 ();
 sg13g2_fill_2 FILLER_184_1382 ();
 sg13g2_fill_2 FILLER_184_1418 ();
 sg13g2_fill_8 FILLER_184_1447 ();
 sg13g2_fill_8 FILLER_184_1455 ();
 sg13g2_fill_8 FILLER_184_1463 ();
 sg13g2_fill_8 FILLER_184_1471 ();
 sg13g2_fill_8 FILLER_184_1479 ();
 sg13g2_fill_8 FILLER_184_1487 ();
 sg13g2_fill_8 FILLER_184_1495 ();
 sg13g2_fill_8 FILLER_184_1503 ();
 sg13g2_fill_8 FILLER_184_1511 ();
 sg13g2_fill_8 FILLER_184_1519 ();
 sg13g2_fill_8 FILLER_184_1527 ();
 sg13g2_fill_8 FILLER_184_1535 ();
 sg13g2_fill_8 FILLER_184_1543 ();
 sg13g2_fill_8 FILLER_184_1551 ();
 sg13g2_fill_8 FILLER_184_1559 ();
 sg13g2_fill_8 FILLER_184_1567 ();
 sg13g2_fill_8 FILLER_184_1575 ();
 sg13g2_fill_8 FILLER_184_1583 ();
 sg13g2_fill_1 FILLER_184_1591 ();
 sg13g2_fill_8 FILLER_185_0 ();
 sg13g2_fill_8 FILLER_185_8 ();
 sg13g2_fill_8 FILLER_185_16 ();
 sg13g2_fill_8 FILLER_185_24 ();
 sg13g2_fill_8 FILLER_185_32 ();
 sg13g2_fill_8 FILLER_185_40 ();
 sg13g2_fill_8 FILLER_185_48 ();
 sg13g2_fill_8 FILLER_185_56 ();
 sg13g2_fill_8 FILLER_185_64 ();
 sg13g2_fill_8 FILLER_185_72 ();
 sg13g2_fill_8 FILLER_185_80 ();
 sg13g2_fill_8 FILLER_185_88 ();
 sg13g2_fill_8 FILLER_185_96 ();
 sg13g2_fill_8 FILLER_185_104 ();
 sg13g2_fill_8 FILLER_185_112 ();
 sg13g2_fill_8 FILLER_185_120 ();
 sg13g2_fill_8 FILLER_185_128 ();
 sg13g2_fill_8 FILLER_185_136 ();
 sg13g2_fill_8 FILLER_185_144 ();
 sg13g2_fill_2 FILLER_185_152 ();
 sg13g2_fill_1 FILLER_185_154 ();
 sg13g2_fill_8 FILLER_185_207 ();
 sg13g2_fill_8 FILLER_185_215 ();
 sg13g2_fill_8 FILLER_185_223 ();
 sg13g2_fill_8 FILLER_185_231 ();
 sg13g2_fill_2 FILLER_185_239 ();
 sg13g2_fill_1 FILLER_185_241 ();
 sg13g2_fill_8 FILLER_185_252 ();
 sg13g2_fill_8 FILLER_185_260 ();
 sg13g2_fill_8 FILLER_185_268 ();
 sg13g2_fill_8 FILLER_185_276 ();
 sg13g2_fill_8 FILLER_185_284 ();
 sg13g2_fill_8 FILLER_185_292 ();
 sg13g2_fill_4 FILLER_185_300 ();
 sg13g2_fill_4 FILLER_185_314 ();
 sg13g2_fill_8 FILLER_185_344 ();
 sg13g2_fill_8 FILLER_185_352 ();
 sg13g2_fill_8 FILLER_185_360 ();
 sg13g2_fill_8 FILLER_185_368 ();
 sg13g2_fill_8 FILLER_185_376 ();
 sg13g2_fill_8 FILLER_185_384 ();
 sg13g2_fill_8 FILLER_185_392 ();
 sg13g2_fill_8 FILLER_185_400 ();
 sg13g2_fill_8 FILLER_185_408 ();
 sg13g2_fill_8 FILLER_185_416 ();
 sg13g2_fill_8 FILLER_185_424 ();
 sg13g2_fill_8 FILLER_185_432 ();
 sg13g2_fill_8 FILLER_185_440 ();
 sg13g2_fill_8 FILLER_185_448 ();
 sg13g2_fill_8 FILLER_185_456 ();
 sg13g2_fill_8 FILLER_185_464 ();
 sg13g2_fill_8 FILLER_185_472 ();
 sg13g2_fill_8 FILLER_185_480 ();
 sg13g2_fill_8 FILLER_185_488 ();
 sg13g2_fill_8 FILLER_185_496 ();
 sg13g2_fill_8 FILLER_185_504 ();
 sg13g2_fill_8 FILLER_185_512 ();
 sg13g2_fill_8 FILLER_185_530 ();
 sg13g2_fill_8 FILLER_185_538 ();
 sg13g2_fill_8 FILLER_185_546 ();
 sg13g2_fill_8 FILLER_185_554 ();
 sg13g2_fill_4 FILLER_185_562 ();
 sg13g2_fill_2 FILLER_185_566 ();
 sg13g2_fill_1 FILLER_185_568 ();
 sg13g2_fill_8 FILLER_185_579 ();
 sg13g2_fill_1 FILLER_185_587 ();
 sg13g2_fill_2 FILLER_185_624 ();
 sg13g2_fill_8 FILLER_185_652 ();
 sg13g2_fill_2 FILLER_185_660 ();
 sg13g2_fill_8 FILLER_185_672 ();
 sg13g2_fill_8 FILLER_185_680 ();
 sg13g2_fill_8 FILLER_185_732 ();
 sg13g2_fill_4 FILLER_185_768 ();
 sg13g2_fill_2 FILLER_185_772 ();
 sg13g2_fill_1 FILLER_185_774 ();
 sg13g2_fill_2 FILLER_185_783 ();
 sg13g2_fill_1 FILLER_185_785 ();
 sg13g2_fill_4 FILLER_185_796 ();
 sg13g2_fill_8 FILLER_185_826 ();
 sg13g2_fill_8 FILLER_185_834 ();
 sg13g2_fill_8 FILLER_185_842 ();
 sg13g2_fill_8 FILLER_185_850 ();
 sg13g2_fill_8 FILLER_185_858 ();
 sg13g2_fill_8 FILLER_185_866 ();
 sg13g2_fill_8 FILLER_185_874 ();
 sg13g2_fill_8 FILLER_185_882 ();
 sg13g2_fill_8 FILLER_185_890 ();
 sg13g2_fill_8 FILLER_185_898 ();
 sg13g2_fill_8 FILLER_185_906 ();
 sg13g2_fill_8 FILLER_185_914 ();
 sg13g2_fill_8 FILLER_185_922 ();
 sg13g2_fill_8 FILLER_185_930 ();
 sg13g2_fill_8 FILLER_185_938 ();
 sg13g2_fill_8 FILLER_185_946 ();
 sg13g2_fill_8 FILLER_185_954 ();
 sg13g2_fill_8 FILLER_185_962 ();
 sg13g2_fill_4 FILLER_185_970 ();
 sg13g2_fill_2 FILLER_185_1001 ();
 sg13g2_fill_8 FILLER_185_1011 ();
 sg13g2_fill_8 FILLER_185_1019 ();
 sg13g2_fill_2 FILLER_185_1027 ();
 sg13g2_fill_1 FILLER_185_1029 ();
 sg13g2_fill_8 FILLER_185_1034 ();
 sg13g2_fill_8 FILLER_185_1042 ();
 sg13g2_fill_4 FILLER_185_1050 ();
 sg13g2_fill_2 FILLER_185_1054 ();
 sg13g2_fill_2 FILLER_185_1072 ();
 sg13g2_fill_4 FILLER_185_1088 ();
 sg13g2_fill_8 FILLER_185_1097 ();
 sg13g2_fill_4 FILLER_185_1105 ();
 sg13g2_fill_2 FILLER_185_1109 ();
 sg13g2_fill_1 FILLER_185_1111 ();
 sg13g2_fill_8 FILLER_185_1117 ();
 sg13g2_fill_8 FILLER_185_1125 ();
 sg13g2_fill_4 FILLER_185_1133 ();
 sg13g2_fill_8 FILLER_185_1171 ();
 sg13g2_fill_4 FILLER_185_1179 ();
 sg13g2_fill_2 FILLER_185_1194 ();
 sg13g2_fill_1 FILLER_185_1196 ();
 sg13g2_fill_2 FILLER_185_1203 ();
 sg13g2_fill_1 FILLER_185_1205 ();
 sg13g2_fill_8 FILLER_185_1222 ();
 sg13g2_fill_1 FILLER_185_1230 ();
 sg13g2_fill_8 FILLER_185_1247 ();
 sg13g2_fill_2 FILLER_185_1255 ();
 sg13g2_fill_1 FILLER_185_1302 ();
 sg13g2_fill_8 FILLER_185_1315 ();
 sg13g2_fill_4 FILLER_185_1323 ();
 sg13g2_fill_2 FILLER_185_1327 ();
 sg13g2_fill_1 FILLER_185_1329 ();
 sg13g2_fill_1 FILLER_185_1334 ();
 sg13g2_fill_2 FILLER_185_1343 ();
 sg13g2_fill_1 FILLER_185_1345 ();
 sg13g2_fill_8 FILLER_185_1365 ();
 sg13g2_fill_8 FILLER_185_1373 ();
 sg13g2_fill_8 FILLER_185_1381 ();
 sg13g2_fill_4 FILLER_185_1409 ();
 sg13g2_fill_2 FILLER_185_1413 ();
 sg13g2_fill_8 FILLER_185_1438 ();
 sg13g2_fill_8 FILLER_185_1446 ();
 sg13g2_fill_8 FILLER_185_1454 ();
 sg13g2_fill_8 FILLER_185_1462 ();
 sg13g2_fill_8 FILLER_185_1470 ();
 sg13g2_fill_8 FILLER_185_1478 ();
 sg13g2_fill_8 FILLER_185_1486 ();
 sg13g2_fill_8 FILLER_185_1494 ();
 sg13g2_fill_8 FILLER_185_1502 ();
 sg13g2_fill_8 FILLER_185_1510 ();
 sg13g2_fill_8 FILLER_185_1518 ();
 sg13g2_fill_8 FILLER_185_1526 ();
 sg13g2_fill_8 FILLER_185_1534 ();
 sg13g2_fill_8 FILLER_185_1542 ();
 sg13g2_fill_8 FILLER_185_1550 ();
 sg13g2_fill_8 FILLER_185_1558 ();
 sg13g2_fill_8 FILLER_185_1566 ();
 sg13g2_fill_8 FILLER_185_1574 ();
 sg13g2_fill_8 FILLER_185_1582 ();
 sg13g2_fill_2 FILLER_185_1590 ();
 sg13g2_fill_8 FILLER_186_0 ();
 sg13g2_fill_8 FILLER_186_8 ();
 sg13g2_fill_8 FILLER_186_16 ();
 sg13g2_fill_8 FILLER_186_24 ();
 sg13g2_fill_8 FILLER_186_32 ();
 sg13g2_fill_8 FILLER_186_40 ();
 sg13g2_fill_8 FILLER_186_48 ();
 sg13g2_fill_8 FILLER_186_56 ();
 sg13g2_fill_8 FILLER_186_64 ();
 sg13g2_fill_8 FILLER_186_72 ();
 sg13g2_fill_8 FILLER_186_80 ();
 sg13g2_fill_8 FILLER_186_88 ();
 sg13g2_fill_8 FILLER_186_96 ();
 sg13g2_fill_8 FILLER_186_104 ();
 sg13g2_fill_8 FILLER_186_112 ();
 sg13g2_fill_8 FILLER_186_120 ();
 sg13g2_fill_8 FILLER_186_128 ();
 sg13g2_fill_8 FILLER_186_136 ();
 sg13g2_fill_8 FILLER_186_144 ();
 sg13g2_fill_8 FILLER_186_152 ();
 sg13g2_fill_8 FILLER_186_160 ();
 sg13g2_fill_8 FILLER_186_168 ();
 sg13g2_fill_8 FILLER_186_176 ();
 sg13g2_fill_8 FILLER_186_184 ();
 sg13g2_fill_8 FILLER_186_192 ();
 sg13g2_fill_8 FILLER_186_200 ();
 sg13g2_fill_8 FILLER_186_208 ();
 sg13g2_fill_8 FILLER_186_216 ();
 sg13g2_fill_8 FILLER_186_224 ();
 sg13g2_fill_8 FILLER_186_232 ();
 sg13g2_fill_8 FILLER_186_240 ();
 sg13g2_fill_8 FILLER_186_248 ();
 sg13g2_fill_8 FILLER_186_256 ();
 sg13g2_fill_8 FILLER_186_264 ();
 sg13g2_fill_8 FILLER_186_272 ();
 sg13g2_fill_8 FILLER_186_280 ();
 sg13g2_fill_8 FILLER_186_288 ();
 sg13g2_fill_8 FILLER_186_296 ();
 sg13g2_fill_8 FILLER_186_304 ();
 sg13g2_fill_8 FILLER_186_312 ();
 sg13g2_fill_8 FILLER_186_320 ();
 sg13g2_fill_8 FILLER_186_328 ();
 sg13g2_fill_8 FILLER_186_336 ();
 sg13g2_fill_8 FILLER_186_344 ();
 sg13g2_fill_8 FILLER_186_352 ();
 sg13g2_fill_8 FILLER_186_360 ();
 sg13g2_fill_8 FILLER_186_368 ();
 sg13g2_fill_8 FILLER_186_376 ();
 sg13g2_fill_8 FILLER_186_384 ();
 sg13g2_fill_8 FILLER_186_392 ();
 sg13g2_fill_8 FILLER_186_400 ();
 sg13g2_fill_8 FILLER_186_408 ();
 sg13g2_fill_8 FILLER_186_416 ();
 sg13g2_fill_8 FILLER_186_424 ();
 sg13g2_fill_8 FILLER_186_432 ();
 sg13g2_fill_8 FILLER_186_440 ();
 sg13g2_fill_8 FILLER_186_448 ();
 sg13g2_fill_8 FILLER_186_456 ();
 sg13g2_fill_8 FILLER_186_464 ();
 sg13g2_fill_8 FILLER_186_472 ();
 sg13g2_fill_8 FILLER_186_480 ();
 sg13g2_fill_8 FILLER_186_488 ();
 sg13g2_fill_8 FILLER_186_496 ();
 sg13g2_fill_8 FILLER_186_504 ();
 sg13g2_fill_8 FILLER_186_512 ();
 sg13g2_fill_8 FILLER_186_520 ();
 sg13g2_fill_8 FILLER_186_528 ();
 sg13g2_fill_8 FILLER_186_536 ();
 sg13g2_fill_8 FILLER_186_544 ();
 sg13g2_fill_4 FILLER_186_552 ();
 sg13g2_fill_4 FILLER_186_566 ();
 sg13g2_fill_1 FILLER_186_570 ();
 sg13g2_fill_4 FILLER_186_597 ();
 sg13g2_fill_2 FILLER_186_601 ();
 sg13g2_fill_1 FILLER_186_625 ();
 sg13g2_fill_8 FILLER_186_652 ();
 sg13g2_fill_2 FILLER_186_660 ();
 sg13g2_fill_8 FILLER_186_682 ();
 sg13g2_fill_8 FILLER_186_690 ();
 sg13g2_fill_1 FILLER_186_698 ();
 sg13g2_fill_8 FILLER_186_709 ();
 sg13g2_fill_4 FILLER_186_717 ();
 sg13g2_fill_1 FILLER_186_721 ();
 sg13g2_fill_4 FILLER_186_742 ();
 sg13g2_fill_2 FILLER_186_746 ();
 sg13g2_fill_1 FILLER_186_748 ();
 sg13g2_fill_2 FILLER_186_759 ();
 sg13g2_fill_8 FILLER_186_807 ();
 sg13g2_fill_8 FILLER_186_815 ();
 sg13g2_fill_8 FILLER_186_823 ();
 sg13g2_fill_8 FILLER_186_831 ();
 sg13g2_fill_8 FILLER_186_839 ();
 sg13g2_fill_8 FILLER_186_847 ();
 sg13g2_fill_8 FILLER_186_855 ();
 sg13g2_fill_8 FILLER_186_863 ();
 sg13g2_fill_8 FILLER_186_871 ();
 sg13g2_fill_8 FILLER_186_879 ();
 sg13g2_fill_8 FILLER_186_887 ();
 sg13g2_fill_8 FILLER_186_895 ();
 sg13g2_fill_8 FILLER_186_903 ();
 sg13g2_fill_8 FILLER_186_911 ();
 sg13g2_fill_8 FILLER_186_919 ();
 sg13g2_fill_8 FILLER_186_927 ();
 sg13g2_fill_8 FILLER_186_935 ();
 sg13g2_fill_8 FILLER_186_943 ();
 sg13g2_fill_8 FILLER_186_951 ();
 sg13g2_fill_8 FILLER_186_959 ();
 sg13g2_fill_8 FILLER_186_967 ();
 sg13g2_fill_8 FILLER_186_975 ();
 sg13g2_fill_8 FILLER_186_983 ();
 sg13g2_fill_4 FILLER_186_996 ();
 sg13g2_fill_2 FILLER_186_1000 ();
 sg13g2_fill_1 FILLER_186_1002 ();
 sg13g2_fill_1 FILLER_186_1027 ();
 sg13g2_fill_4 FILLER_186_1040 ();
 sg13g2_fill_1 FILLER_186_1044 ();
 sg13g2_fill_1 FILLER_186_1050 ();
 sg13g2_fill_1 FILLER_186_1055 ();
 sg13g2_fill_8 FILLER_186_1064 ();
 sg13g2_fill_4 FILLER_186_1072 ();
 sg13g2_fill_2 FILLER_186_1076 ();
 sg13g2_fill_1 FILLER_186_1078 ();
 sg13g2_fill_8 FILLER_186_1085 ();
 sg13g2_fill_4 FILLER_186_1093 ();
 sg13g2_fill_2 FILLER_186_1097 ();
 sg13g2_fill_1 FILLER_186_1099 ();
 sg13g2_fill_4 FILLER_186_1131 ();
 sg13g2_fill_2 FILLER_186_1135 ();
 sg13g2_fill_1 FILLER_186_1137 ();
 sg13g2_fill_4 FILLER_186_1146 ();
 sg13g2_fill_2 FILLER_186_1150 ();
 sg13g2_fill_4 FILLER_186_1162 ();
 sg13g2_fill_4 FILLER_186_1172 ();
 sg13g2_fill_8 FILLER_186_1188 ();
 sg13g2_fill_4 FILLER_186_1196 ();
 sg13g2_fill_2 FILLER_186_1200 ();
 sg13g2_fill_1 FILLER_186_1202 ();
 sg13g2_fill_8 FILLER_186_1219 ();
 sg13g2_fill_8 FILLER_186_1227 ();
 sg13g2_fill_4 FILLER_186_1235 ();
 sg13g2_fill_4 FILLER_186_1255 ();
 sg13g2_fill_8 FILLER_186_1280 ();
 sg13g2_fill_1 FILLER_186_1288 ();
 sg13g2_fill_2 FILLER_186_1297 ();
 sg13g2_fill_2 FILLER_186_1304 ();
 sg13g2_fill_4 FILLER_186_1322 ();
 sg13g2_fill_1 FILLER_186_1326 ();
 sg13g2_fill_4 FILLER_186_1331 ();
 sg13g2_fill_1 FILLER_186_1335 ();
 sg13g2_fill_1 FILLER_186_1344 ();
 sg13g2_fill_8 FILLER_186_1349 ();
 sg13g2_fill_8 FILLER_186_1357 ();
 sg13g2_fill_1 FILLER_186_1365 ();
 sg13g2_fill_4 FILLER_186_1380 ();
 sg13g2_fill_4 FILLER_186_1393 ();
 sg13g2_fill_8 FILLER_186_1402 ();
 sg13g2_fill_1 FILLER_186_1410 ();
 sg13g2_fill_2 FILLER_186_1421 ();
 sg13g2_fill_1 FILLER_186_1423 ();
 sg13g2_fill_8 FILLER_186_1429 ();
 sg13g2_fill_8 FILLER_186_1437 ();
 sg13g2_fill_8 FILLER_186_1445 ();
 sg13g2_fill_8 FILLER_186_1453 ();
 sg13g2_fill_8 FILLER_186_1461 ();
 sg13g2_fill_8 FILLER_186_1469 ();
 sg13g2_fill_8 FILLER_186_1477 ();
 sg13g2_fill_8 FILLER_186_1485 ();
 sg13g2_fill_8 FILLER_186_1493 ();
 sg13g2_fill_8 FILLER_186_1501 ();
 sg13g2_fill_8 FILLER_186_1509 ();
 sg13g2_fill_8 FILLER_186_1517 ();
 sg13g2_fill_8 FILLER_186_1525 ();
 sg13g2_fill_8 FILLER_186_1533 ();
 sg13g2_fill_8 FILLER_186_1541 ();
 sg13g2_fill_8 FILLER_186_1549 ();
 sg13g2_fill_8 FILLER_186_1557 ();
 sg13g2_fill_8 FILLER_186_1565 ();
 sg13g2_fill_8 FILLER_186_1573 ();
 sg13g2_fill_8 FILLER_186_1581 ();
 sg13g2_fill_2 FILLER_186_1589 ();
 sg13g2_fill_1 FILLER_186_1591 ();
 sg13g2_fill_8 FILLER_187_0 ();
 sg13g2_fill_8 FILLER_187_8 ();
 sg13g2_fill_8 FILLER_187_16 ();
 sg13g2_fill_8 FILLER_187_24 ();
 sg13g2_fill_8 FILLER_187_32 ();
 sg13g2_fill_8 FILLER_187_40 ();
 sg13g2_fill_8 FILLER_187_48 ();
 sg13g2_fill_8 FILLER_187_56 ();
 sg13g2_fill_8 FILLER_187_64 ();
 sg13g2_fill_8 FILLER_187_72 ();
 sg13g2_fill_8 FILLER_187_80 ();
 sg13g2_fill_8 FILLER_187_88 ();
 sg13g2_fill_8 FILLER_187_96 ();
 sg13g2_fill_8 FILLER_187_104 ();
 sg13g2_fill_8 FILLER_187_112 ();
 sg13g2_fill_8 FILLER_187_120 ();
 sg13g2_fill_8 FILLER_187_128 ();
 sg13g2_fill_8 FILLER_187_136 ();
 sg13g2_fill_8 FILLER_187_144 ();
 sg13g2_fill_8 FILLER_187_152 ();
 sg13g2_fill_8 FILLER_187_160 ();
 sg13g2_fill_8 FILLER_187_168 ();
 sg13g2_fill_8 FILLER_187_176 ();
 sg13g2_fill_8 FILLER_187_184 ();
 sg13g2_fill_8 FILLER_187_192 ();
 sg13g2_fill_8 FILLER_187_200 ();
 sg13g2_fill_8 FILLER_187_208 ();
 sg13g2_fill_8 FILLER_187_216 ();
 sg13g2_fill_8 FILLER_187_224 ();
 sg13g2_fill_8 FILLER_187_232 ();
 sg13g2_fill_8 FILLER_187_240 ();
 sg13g2_fill_8 FILLER_187_248 ();
 sg13g2_fill_8 FILLER_187_256 ();
 sg13g2_fill_8 FILLER_187_264 ();
 sg13g2_fill_8 FILLER_187_272 ();
 sg13g2_fill_8 FILLER_187_280 ();
 sg13g2_fill_8 FILLER_187_288 ();
 sg13g2_fill_8 FILLER_187_296 ();
 sg13g2_fill_8 FILLER_187_304 ();
 sg13g2_fill_8 FILLER_187_312 ();
 sg13g2_fill_8 FILLER_187_320 ();
 sg13g2_fill_8 FILLER_187_328 ();
 sg13g2_fill_8 FILLER_187_336 ();
 sg13g2_fill_8 FILLER_187_344 ();
 sg13g2_fill_8 FILLER_187_352 ();
 sg13g2_fill_8 FILLER_187_360 ();
 sg13g2_fill_8 FILLER_187_368 ();
 sg13g2_fill_8 FILLER_187_376 ();
 sg13g2_fill_8 FILLER_187_384 ();
 sg13g2_fill_8 FILLER_187_392 ();
 sg13g2_fill_8 FILLER_187_400 ();
 sg13g2_fill_8 FILLER_187_408 ();
 sg13g2_fill_8 FILLER_187_416 ();
 sg13g2_fill_8 FILLER_187_424 ();
 sg13g2_fill_8 FILLER_187_432 ();
 sg13g2_fill_8 FILLER_187_440 ();
 sg13g2_fill_8 FILLER_187_448 ();
 sg13g2_fill_8 FILLER_187_456 ();
 sg13g2_fill_8 FILLER_187_464 ();
 sg13g2_fill_8 FILLER_187_472 ();
 sg13g2_fill_8 FILLER_187_480 ();
 sg13g2_fill_8 FILLER_187_488 ();
 sg13g2_fill_8 FILLER_187_496 ();
 sg13g2_fill_8 FILLER_187_504 ();
 sg13g2_fill_8 FILLER_187_512 ();
 sg13g2_fill_8 FILLER_187_520 ();
 sg13g2_fill_8 FILLER_187_528 ();
 sg13g2_fill_8 FILLER_187_536 ();
 sg13g2_fill_8 FILLER_187_544 ();
 sg13g2_fill_2 FILLER_187_552 ();
 sg13g2_fill_1 FILLER_187_554 ();
 sg13g2_fill_8 FILLER_187_575 ();
 sg13g2_fill_8 FILLER_187_583 ();
 sg13g2_fill_2 FILLER_187_591 ();
 sg13g2_fill_4 FILLER_187_603 ();
 sg13g2_fill_1 FILLER_187_607 ();
 sg13g2_fill_2 FILLER_187_669 ();
 sg13g2_fill_1 FILLER_187_671 ();
 sg13g2_fill_4 FILLER_187_698 ();
 sg13g2_fill_8 FILLER_187_728 ();
 sg13g2_fill_1 FILLER_187_736 ();
 sg13g2_fill_8 FILLER_187_763 ();
 sg13g2_fill_8 FILLER_187_771 ();
 sg13g2_fill_8 FILLER_187_779 ();
 sg13g2_fill_8 FILLER_187_787 ();
 sg13g2_fill_8 FILLER_187_795 ();
 sg13g2_fill_8 FILLER_187_803 ();
 sg13g2_fill_8 FILLER_187_811 ();
 sg13g2_fill_8 FILLER_187_819 ();
 sg13g2_fill_8 FILLER_187_827 ();
 sg13g2_fill_8 FILLER_187_835 ();
 sg13g2_fill_8 FILLER_187_843 ();
 sg13g2_fill_8 FILLER_187_851 ();
 sg13g2_fill_8 FILLER_187_859 ();
 sg13g2_fill_8 FILLER_187_867 ();
 sg13g2_fill_8 FILLER_187_875 ();
 sg13g2_fill_8 FILLER_187_883 ();
 sg13g2_fill_8 FILLER_187_891 ();
 sg13g2_fill_8 FILLER_187_899 ();
 sg13g2_fill_8 FILLER_187_907 ();
 sg13g2_fill_8 FILLER_187_915 ();
 sg13g2_fill_8 FILLER_187_923 ();
 sg13g2_fill_8 FILLER_187_931 ();
 sg13g2_fill_8 FILLER_187_939 ();
 sg13g2_fill_8 FILLER_187_947 ();
 sg13g2_fill_8 FILLER_187_955 ();
 sg13g2_fill_8 FILLER_187_963 ();
 sg13g2_fill_8 FILLER_187_971 ();
 sg13g2_fill_8 FILLER_187_979 ();
 sg13g2_fill_8 FILLER_187_987 ();
 sg13g2_fill_8 FILLER_187_995 ();
 sg13g2_fill_4 FILLER_187_1003 ();
 sg13g2_fill_1 FILLER_187_1007 ();
 sg13g2_fill_1 FILLER_187_1017 ();
 sg13g2_fill_1 FILLER_187_1044 ();
 sg13g2_fill_2 FILLER_187_1050 ();
 sg13g2_fill_1 FILLER_187_1052 ();
 sg13g2_fill_1 FILLER_187_1077 ();
 sg13g2_fill_8 FILLER_187_1090 ();
 sg13g2_fill_1 FILLER_187_1098 ();
 sg13g2_fill_1 FILLER_187_1123 ();
 sg13g2_fill_4 FILLER_187_1143 ();
 sg13g2_fill_8 FILLER_187_1152 ();
 sg13g2_fill_4 FILLER_187_1160 ();
 sg13g2_fill_1 FILLER_187_1164 ();
 sg13g2_fill_8 FILLER_187_1170 ();
 sg13g2_fill_2 FILLER_187_1178 ();
 sg13g2_fill_8 FILLER_187_1199 ();
 sg13g2_fill_8 FILLER_187_1215 ();
 sg13g2_fill_2 FILLER_187_1223 ();
 sg13g2_fill_1 FILLER_187_1225 ();
 sg13g2_fill_8 FILLER_187_1243 ();
 sg13g2_fill_8 FILLER_187_1251 ();
 sg13g2_fill_8 FILLER_187_1259 ();
 sg13g2_fill_4 FILLER_187_1273 ();
 sg13g2_fill_1 FILLER_187_1277 ();
 sg13g2_fill_8 FILLER_187_1283 ();
 sg13g2_fill_4 FILLER_187_1297 ();
 sg13g2_fill_2 FILLER_187_1308 ();
 sg13g2_fill_2 FILLER_187_1331 ();
 sg13g2_fill_1 FILLER_187_1333 ();
 sg13g2_fill_8 FILLER_187_1342 ();
 sg13g2_fill_4 FILLER_187_1350 ();
 sg13g2_fill_2 FILLER_187_1354 ();
 sg13g2_fill_1 FILLER_187_1356 ();
 sg13g2_fill_1 FILLER_187_1373 ();
 sg13g2_fill_4 FILLER_187_1405 ();
 sg13g2_fill_1 FILLER_187_1409 ();
 sg13g2_fill_8 FILLER_187_1415 ();
 sg13g2_fill_2 FILLER_187_1423 ();
 sg13g2_fill_8 FILLER_187_1430 ();
 sg13g2_fill_8 FILLER_187_1438 ();
 sg13g2_fill_8 FILLER_187_1446 ();
 sg13g2_fill_8 FILLER_187_1454 ();
 sg13g2_fill_8 FILLER_187_1462 ();
 sg13g2_fill_8 FILLER_187_1470 ();
 sg13g2_fill_8 FILLER_187_1478 ();
 sg13g2_fill_8 FILLER_187_1486 ();
 sg13g2_fill_8 FILLER_187_1494 ();
 sg13g2_fill_8 FILLER_187_1502 ();
 sg13g2_fill_8 FILLER_187_1510 ();
 sg13g2_fill_8 FILLER_187_1518 ();
 sg13g2_fill_8 FILLER_187_1526 ();
 sg13g2_fill_8 FILLER_187_1534 ();
 sg13g2_fill_8 FILLER_187_1542 ();
 sg13g2_fill_8 FILLER_187_1550 ();
 sg13g2_fill_8 FILLER_187_1558 ();
 sg13g2_fill_8 FILLER_187_1566 ();
 sg13g2_fill_8 FILLER_187_1574 ();
 sg13g2_fill_8 FILLER_187_1582 ();
 sg13g2_fill_2 FILLER_187_1590 ();
 sg13g2_fill_8 FILLER_188_0 ();
 sg13g2_fill_8 FILLER_188_8 ();
 sg13g2_fill_8 FILLER_188_16 ();
 sg13g2_fill_8 FILLER_188_24 ();
 sg13g2_fill_8 FILLER_188_32 ();
 sg13g2_fill_8 FILLER_188_40 ();
 sg13g2_fill_8 FILLER_188_48 ();
 sg13g2_fill_8 FILLER_188_56 ();
 sg13g2_fill_8 FILLER_188_64 ();
 sg13g2_fill_8 FILLER_188_72 ();
 sg13g2_fill_8 FILLER_188_80 ();
 sg13g2_fill_8 FILLER_188_88 ();
 sg13g2_fill_8 FILLER_188_96 ();
 sg13g2_fill_8 FILLER_188_104 ();
 sg13g2_fill_8 FILLER_188_112 ();
 sg13g2_fill_8 FILLER_188_120 ();
 sg13g2_fill_8 FILLER_188_128 ();
 sg13g2_fill_8 FILLER_188_136 ();
 sg13g2_fill_8 FILLER_188_144 ();
 sg13g2_fill_8 FILLER_188_152 ();
 sg13g2_fill_8 FILLER_188_160 ();
 sg13g2_fill_8 FILLER_188_168 ();
 sg13g2_fill_8 FILLER_188_176 ();
 sg13g2_fill_8 FILLER_188_184 ();
 sg13g2_fill_8 FILLER_188_192 ();
 sg13g2_fill_8 FILLER_188_200 ();
 sg13g2_fill_8 FILLER_188_208 ();
 sg13g2_fill_8 FILLER_188_216 ();
 sg13g2_fill_8 FILLER_188_224 ();
 sg13g2_fill_8 FILLER_188_232 ();
 sg13g2_fill_8 FILLER_188_240 ();
 sg13g2_fill_8 FILLER_188_248 ();
 sg13g2_fill_8 FILLER_188_256 ();
 sg13g2_fill_8 FILLER_188_264 ();
 sg13g2_fill_8 FILLER_188_272 ();
 sg13g2_fill_8 FILLER_188_280 ();
 sg13g2_fill_8 FILLER_188_288 ();
 sg13g2_fill_8 FILLER_188_296 ();
 sg13g2_fill_8 FILLER_188_304 ();
 sg13g2_fill_8 FILLER_188_312 ();
 sg13g2_fill_8 FILLER_188_320 ();
 sg13g2_fill_8 FILLER_188_328 ();
 sg13g2_fill_8 FILLER_188_336 ();
 sg13g2_fill_8 FILLER_188_344 ();
 sg13g2_fill_8 FILLER_188_352 ();
 sg13g2_fill_8 FILLER_188_360 ();
 sg13g2_fill_8 FILLER_188_368 ();
 sg13g2_fill_8 FILLER_188_376 ();
 sg13g2_fill_8 FILLER_188_384 ();
 sg13g2_fill_8 FILLER_188_392 ();
 sg13g2_fill_8 FILLER_188_400 ();
 sg13g2_fill_8 FILLER_188_408 ();
 sg13g2_fill_8 FILLER_188_416 ();
 sg13g2_fill_8 FILLER_188_424 ();
 sg13g2_fill_8 FILLER_188_432 ();
 sg13g2_fill_8 FILLER_188_440 ();
 sg13g2_fill_8 FILLER_188_448 ();
 sg13g2_fill_8 FILLER_188_456 ();
 sg13g2_fill_8 FILLER_188_464 ();
 sg13g2_fill_8 FILLER_188_472 ();
 sg13g2_fill_8 FILLER_188_480 ();
 sg13g2_fill_8 FILLER_188_488 ();
 sg13g2_fill_8 FILLER_188_496 ();
 sg13g2_fill_8 FILLER_188_504 ();
 sg13g2_fill_8 FILLER_188_512 ();
 sg13g2_fill_8 FILLER_188_520 ();
 sg13g2_fill_8 FILLER_188_528 ();
 sg13g2_fill_8 FILLER_188_536 ();
 sg13g2_fill_8 FILLER_188_544 ();
 sg13g2_fill_8 FILLER_188_552 ();
 sg13g2_fill_2 FILLER_188_560 ();
 sg13g2_fill_8 FILLER_188_588 ();
 sg13g2_fill_1 FILLER_188_596 ();
 sg13g2_fill_2 FILLER_188_633 ();
 sg13g2_fill_8 FILLER_188_643 ();
 sg13g2_fill_8 FILLER_188_651 ();
 sg13g2_fill_4 FILLER_188_659 ();
 sg13g2_fill_8 FILLER_188_673 ();
 sg13g2_fill_8 FILLER_188_681 ();
 sg13g2_fill_8 FILLER_188_689 ();
 sg13g2_fill_8 FILLER_188_697 ();
 sg13g2_fill_8 FILLER_188_705 ();
 sg13g2_fill_8 FILLER_188_713 ();
 sg13g2_fill_8 FILLER_188_721 ();
 sg13g2_fill_8 FILLER_188_729 ();
 sg13g2_fill_8 FILLER_188_737 ();
 sg13g2_fill_8 FILLER_188_745 ();
 sg13g2_fill_8 FILLER_188_753 ();
 sg13g2_fill_8 FILLER_188_761 ();
 sg13g2_fill_8 FILLER_188_769 ();
 sg13g2_fill_8 FILLER_188_777 ();
 sg13g2_fill_8 FILLER_188_785 ();
 sg13g2_fill_8 FILLER_188_793 ();
 sg13g2_fill_8 FILLER_188_801 ();
 sg13g2_fill_8 FILLER_188_809 ();
 sg13g2_fill_8 FILLER_188_817 ();
 sg13g2_fill_8 FILLER_188_825 ();
 sg13g2_fill_8 FILLER_188_833 ();
 sg13g2_fill_8 FILLER_188_841 ();
 sg13g2_fill_8 FILLER_188_849 ();
 sg13g2_fill_8 FILLER_188_857 ();
 sg13g2_fill_8 FILLER_188_865 ();
 sg13g2_fill_8 FILLER_188_873 ();
 sg13g2_fill_8 FILLER_188_881 ();
 sg13g2_fill_8 FILLER_188_889 ();
 sg13g2_fill_8 FILLER_188_897 ();
 sg13g2_fill_8 FILLER_188_905 ();
 sg13g2_fill_8 FILLER_188_913 ();
 sg13g2_fill_8 FILLER_188_921 ();
 sg13g2_fill_8 FILLER_188_929 ();
 sg13g2_fill_8 FILLER_188_937 ();
 sg13g2_fill_8 FILLER_188_945 ();
 sg13g2_fill_8 FILLER_188_953 ();
 sg13g2_fill_8 FILLER_188_961 ();
 sg13g2_fill_8 FILLER_188_969 ();
 sg13g2_fill_8 FILLER_188_977 ();
 sg13g2_fill_8 FILLER_188_985 ();
 sg13g2_fill_8 FILLER_188_993 ();
 sg13g2_fill_2 FILLER_188_1001 ();
 sg13g2_fill_8 FILLER_188_1020 ();
 sg13g2_fill_8 FILLER_188_1028 ();
 sg13g2_fill_8 FILLER_188_1036 ();
 sg13g2_fill_2 FILLER_188_1044 ();
 sg13g2_fill_1 FILLER_188_1046 ();
 sg13g2_fill_1 FILLER_188_1059 ();
 sg13g2_fill_8 FILLER_188_1068 ();
 sg13g2_fill_2 FILLER_188_1076 ();
 sg13g2_fill_2 FILLER_188_1101 ();
 sg13g2_fill_2 FILLER_188_1108 ();
 sg13g2_fill_1 FILLER_188_1110 ();
 sg13g2_fill_2 FILLER_188_1125 ();
 sg13g2_fill_4 FILLER_188_1132 ();
 sg13g2_fill_1 FILLER_188_1136 ();
 sg13g2_fill_8 FILLER_188_1147 ();
 sg13g2_fill_4 FILLER_188_1155 ();
 sg13g2_fill_2 FILLER_188_1159 ();
 sg13g2_fill_1 FILLER_188_1161 ();
 sg13g2_fill_8 FILLER_188_1176 ();
 sg13g2_fill_4 FILLER_188_1184 ();
 sg13g2_fill_1 FILLER_188_1188 ();
 sg13g2_fill_4 FILLER_188_1202 ();
 sg13g2_fill_2 FILLER_188_1206 ();
 sg13g2_fill_4 FILLER_188_1224 ();
 sg13g2_fill_2 FILLER_188_1228 ();
 sg13g2_fill_4 FILLER_188_1262 ();
 sg13g2_fill_1 FILLER_188_1266 ();
 sg13g2_fill_4 FILLER_188_1273 ();
 sg13g2_fill_4 FILLER_188_1295 ();
 sg13g2_fill_8 FILLER_188_1311 ();
 sg13g2_fill_2 FILLER_188_1319 ();
 sg13g2_fill_4 FILLER_188_1330 ();
 sg13g2_fill_2 FILLER_188_1334 ();
 sg13g2_fill_1 FILLER_188_1341 ();
 sg13g2_fill_2 FILLER_188_1350 ();
 sg13g2_fill_8 FILLER_188_1356 ();
 sg13g2_fill_1 FILLER_188_1364 ();
 sg13g2_fill_4 FILLER_188_1370 ();
 sg13g2_fill_2 FILLER_188_1374 ();
 sg13g2_fill_2 FILLER_188_1380 ();
 sg13g2_fill_1 FILLER_188_1382 ();
 sg13g2_fill_8 FILLER_188_1393 ();
 sg13g2_fill_1 FILLER_188_1401 ();
 sg13g2_fill_8 FILLER_188_1422 ();
 sg13g2_fill_8 FILLER_188_1430 ();
 sg13g2_fill_8 FILLER_188_1438 ();
 sg13g2_fill_8 FILLER_188_1446 ();
 sg13g2_fill_8 FILLER_188_1454 ();
 sg13g2_fill_8 FILLER_188_1462 ();
 sg13g2_fill_8 FILLER_188_1470 ();
 sg13g2_fill_8 FILLER_188_1478 ();
 sg13g2_fill_8 FILLER_188_1486 ();
 sg13g2_fill_8 FILLER_188_1494 ();
 sg13g2_fill_8 FILLER_188_1502 ();
 sg13g2_fill_8 FILLER_188_1510 ();
 sg13g2_fill_8 FILLER_188_1518 ();
 sg13g2_fill_8 FILLER_188_1526 ();
 sg13g2_fill_8 FILLER_188_1534 ();
 sg13g2_fill_8 FILLER_188_1542 ();
 sg13g2_fill_8 FILLER_188_1550 ();
 sg13g2_fill_8 FILLER_188_1558 ();
 sg13g2_fill_8 FILLER_188_1566 ();
 sg13g2_fill_8 FILLER_188_1574 ();
 sg13g2_fill_8 FILLER_188_1582 ();
 sg13g2_fill_2 FILLER_188_1590 ();
 sg13g2_fill_8 FILLER_189_0 ();
 sg13g2_fill_8 FILLER_189_8 ();
 sg13g2_fill_8 FILLER_189_16 ();
 sg13g2_fill_8 FILLER_189_24 ();
 sg13g2_fill_8 FILLER_189_32 ();
 sg13g2_fill_8 FILLER_189_40 ();
 sg13g2_fill_8 FILLER_189_48 ();
 sg13g2_fill_8 FILLER_189_56 ();
 sg13g2_fill_8 FILLER_189_64 ();
 sg13g2_fill_8 FILLER_189_72 ();
 sg13g2_fill_8 FILLER_189_80 ();
 sg13g2_fill_8 FILLER_189_88 ();
 sg13g2_fill_8 FILLER_189_96 ();
 sg13g2_fill_8 FILLER_189_104 ();
 sg13g2_fill_8 FILLER_189_112 ();
 sg13g2_fill_8 FILLER_189_120 ();
 sg13g2_fill_8 FILLER_189_128 ();
 sg13g2_fill_8 FILLER_189_136 ();
 sg13g2_fill_8 FILLER_189_144 ();
 sg13g2_fill_8 FILLER_189_152 ();
 sg13g2_fill_8 FILLER_189_160 ();
 sg13g2_fill_8 FILLER_189_168 ();
 sg13g2_fill_8 FILLER_189_176 ();
 sg13g2_fill_8 FILLER_189_184 ();
 sg13g2_fill_8 FILLER_189_192 ();
 sg13g2_fill_8 FILLER_189_200 ();
 sg13g2_fill_8 FILLER_189_208 ();
 sg13g2_fill_8 FILLER_189_216 ();
 sg13g2_fill_8 FILLER_189_224 ();
 sg13g2_fill_8 FILLER_189_232 ();
 sg13g2_fill_8 FILLER_189_240 ();
 sg13g2_fill_8 FILLER_189_248 ();
 sg13g2_fill_8 FILLER_189_256 ();
 sg13g2_fill_8 FILLER_189_264 ();
 sg13g2_fill_8 FILLER_189_272 ();
 sg13g2_fill_8 FILLER_189_280 ();
 sg13g2_fill_8 FILLER_189_288 ();
 sg13g2_fill_8 FILLER_189_296 ();
 sg13g2_fill_8 FILLER_189_304 ();
 sg13g2_fill_8 FILLER_189_312 ();
 sg13g2_fill_8 FILLER_189_320 ();
 sg13g2_fill_8 FILLER_189_328 ();
 sg13g2_fill_8 FILLER_189_336 ();
 sg13g2_fill_8 FILLER_189_344 ();
 sg13g2_fill_8 FILLER_189_352 ();
 sg13g2_fill_8 FILLER_189_360 ();
 sg13g2_fill_8 FILLER_189_368 ();
 sg13g2_fill_8 FILLER_189_376 ();
 sg13g2_fill_8 FILLER_189_384 ();
 sg13g2_fill_8 FILLER_189_392 ();
 sg13g2_fill_8 FILLER_189_400 ();
 sg13g2_fill_8 FILLER_189_408 ();
 sg13g2_fill_8 FILLER_189_416 ();
 sg13g2_fill_8 FILLER_189_424 ();
 sg13g2_fill_8 FILLER_189_432 ();
 sg13g2_fill_8 FILLER_189_440 ();
 sg13g2_fill_8 FILLER_189_448 ();
 sg13g2_fill_8 FILLER_189_456 ();
 sg13g2_fill_8 FILLER_189_464 ();
 sg13g2_fill_8 FILLER_189_472 ();
 sg13g2_fill_8 FILLER_189_480 ();
 sg13g2_fill_8 FILLER_189_488 ();
 sg13g2_fill_8 FILLER_189_496 ();
 sg13g2_fill_8 FILLER_189_504 ();
 sg13g2_fill_8 FILLER_189_512 ();
 sg13g2_fill_8 FILLER_189_520 ();
 sg13g2_fill_8 FILLER_189_528 ();
 sg13g2_fill_8 FILLER_189_536 ();
 sg13g2_fill_8 FILLER_189_544 ();
 sg13g2_fill_8 FILLER_189_552 ();
 sg13g2_fill_8 FILLER_189_560 ();
 sg13g2_fill_8 FILLER_189_568 ();
 sg13g2_fill_8 FILLER_189_576 ();
 sg13g2_fill_8 FILLER_189_584 ();
 sg13g2_fill_8 FILLER_189_592 ();
 sg13g2_fill_8 FILLER_189_600 ();
 sg13g2_fill_8 FILLER_189_608 ();
 sg13g2_fill_8 FILLER_189_616 ();
 sg13g2_fill_8 FILLER_189_624 ();
 sg13g2_fill_8 FILLER_189_632 ();
 sg13g2_fill_8 FILLER_189_640 ();
 sg13g2_fill_8 FILLER_189_648 ();
 sg13g2_fill_8 FILLER_189_656 ();
 sg13g2_fill_8 FILLER_189_664 ();
 sg13g2_fill_8 FILLER_189_672 ();
 sg13g2_fill_8 FILLER_189_680 ();
 sg13g2_fill_8 FILLER_189_688 ();
 sg13g2_fill_8 FILLER_189_696 ();
 sg13g2_fill_8 FILLER_189_704 ();
 sg13g2_fill_8 FILLER_189_712 ();
 sg13g2_fill_8 FILLER_189_720 ();
 sg13g2_fill_8 FILLER_189_728 ();
 sg13g2_fill_8 FILLER_189_736 ();
 sg13g2_fill_8 FILLER_189_744 ();
 sg13g2_fill_8 FILLER_189_752 ();
 sg13g2_fill_8 FILLER_189_760 ();
 sg13g2_fill_8 FILLER_189_768 ();
 sg13g2_fill_8 FILLER_189_776 ();
 sg13g2_fill_8 FILLER_189_784 ();
 sg13g2_fill_8 FILLER_189_792 ();
 sg13g2_fill_8 FILLER_189_800 ();
 sg13g2_fill_8 FILLER_189_808 ();
 sg13g2_fill_8 FILLER_189_816 ();
 sg13g2_fill_8 FILLER_189_824 ();
 sg13g2_fill_8 FILLER_189_832 ();
 sg13g2_fill_8 FILLER_189_840 ();
 sg13g2_fill_8 FILLER_189_848 ();
 sg13g2_fill_8 FILLER_189_856 ();
 sg13g2_fill_8 FILLER_189_864 ();
 sg13g2_fill_8 FILLER_189_872 ();
 sg13g2_fill_8 FILLER_189_880 ();
 sg13g2_fill_8 FILLER_189_888 ();
 sg13g2_fill_8 FILLER_189_896 ();
 sg13g2_fill_8 FILLER_189_904 ();
 sg13g2_fill_8 FILLER_189_912 ();
 sg13g2_fill_8 FILLER_189_920 ();
 sg13g2_fill_8 FILLER_189_928 ();
 sg13g2_fill_8 FILLER_189_936 ();
 sg13g2_fill_8 FILLER_189_944 ();
 sg13g2_fill_8 FILLER_189_952 ();
 sg13g2_fill_8 FILLER_189_960 ();
 sg13g2_fill_8 FILLER_189_968 ();
 sg13g2_fill_8 FILLER_189_976 ();
 sg13g2_fill_8 FILLER_189_984 ();
 sg13g2_fill_8 FILLER_189_992 ();
 sg13g2_fill_4 FILLER_189_1000 ();
 sg13g2_fill_2 FILLER_189_1004 ();
 sg13g2_fill_1 FILLER_189_1006 ();
 sg13g2_fill_8 FILLER_189_1027 ();
 sg13g2_fill_8 FILLER_189_1035 ();
 sg13g2_fill_8 FILLER_189_1051 ();
 sg13g2_fill_8 FILLER_189_1059 ();
 sg13g2_fill_2 FILLER_189_1067 ();
 sg13g2_fill_1 FILLER_189_1069 ();
 sg13g2_fill_4 FILLER_189_1078 ();
 sg13g2_fill_2 FILLER_189_1082 ();
 sg13g2_fill_1 FILLER_189_1084 ();
 sg13g2_fill_8 FILLER_189_1092 ();
 sg13g2_fill_8 FILLER_189_1104 ();
 sg13g2_fill_8 FILLER_189_1112 ();
 sg13g2_fill_4 FILLER_189_1120 ();
 sg13g2_fill_1 FILLER_189_1124 ();
 sg13g2_fill_2 FILLER_189_1131 ();
 sg13g2_fill_1 FILLER_189_1133 ();
 sg13g2_fill_4 FILLER_189_1154 ();
 sg13g2_fill_8 FILLER_189_1179 ();
 sg13g2_fill_4 FILLER_189_1195 ();
 sg13g2_fill_1 FILLER_189_1199 ();
 sg13g2_fill_8 FILLER_189_1223 ();
 sg13g2_fill_8 FILLER_189_1231 ();
 sg13g2_fill_8 FILLER_189_1239 ();
 sg13g2_fill_1 FILLER_189_1247 ();
 sg13g2_fill_8 FILLER_189_1273 ();
 sg13g2_fill_1 FILLER_189_1281 ();
 sg13g2_fill_8 FILLER_189_1288 ();
 sg13g2_fill_8 FILLER_189_1301 ();
 sg13g2_fill_8 FILLER_189_1309 ();
 sg13g2_fill_8 FILLER_189_1317 ();
 sg13g2_fill_8 FILLER_189_1325 ();
 sg13g2_fill_8 FILLER_189_1333 ();
 sg13g2_fill_8 FILLER_189_1341 ();
 sg13g2_fill_8 FILLER_189_1349 ();
 sg13g2_fill_8 FILLER_189_1357 ();
 sg13g2_fill_8 FILLER_189_1365 ();
 sg13g2_fill_8 FILLER_189_1373 ();
 sg13g2_fill_8 FILLER_189_1381 ();
 sg13g2_fill_8 FILLER_189_1389 ();
 sg13g2_fill_1 FILLER_189_1397 ();
 sg13g2_fill_1 FILLER_189_1408 ();
 sg13g2_fill_8 FILLER_189_1422 ();
 sg13g2_fill_8 FILLER_189_1430 ();
 sg13g2_fill_8 FILLER_189_1438 ();
 sg13g2_fill_8 FILLER_189_1446 ();
 sg13g2_fill_8 FILLER_189_1454 ();
 sg13g2_fill_8 FILLER_189_1462 ();
 sg13g2_fill_8 FILLER_189_1470 ();
 sg13g2_fill_8 FILLER_189_1478 ();
 sg13g2_fill_8 FILLER_189_1486 ();
 sg13g2_fill_8 FILLER_189_1494 ();
 sg13g2_fill_8 FILLER_189_1502 ();
 sg13g2_fill_8 FILLER_189_1510 ();
 sg13g2_fill_8 FILLER_189_1518 ();
 sg13g2_fill_8 FILLER_189_1526 ();
 sg13g2_fill_8 FILLER_189_1534 ();
 sg13g2_fill_8 FILLER_189_1542 ();
 sg13g2_fill_8 FILLER_189_1550 ();
 sg13g2_fill_8 FILLER_189_1558 ();
 sg13g2_fill_8 FILLER_189_1566 ();
 sg13g2_fill_8 FILLER_189_1574 ();
 sg13g2_fill_8 FILLER_189_1582 ();
 sg13g2_fill_2 FILLER_189_1590 ();
 sg13g2_fill_8 FILLER_190_0 ();
 sg13g2_fill_8 FILLER_190_8 ();
 sg13g2_fill_8 FILLER_190_16 ();
 sg13g2_fill_8 FILLER_190_24 ();
 sg13g2_fill_8 FILLER_190_32 ();
 sg13g2_fill_8 FILLER_190_40 ();
 sg13g2_fill_8 FILLER_190_48 ();
 sg13g2_fill_8 FILLER_190_56 ();
 sg13g2_fill_8 FILLER_190_64 ();
 sg13g2_fill_8 FILLER_190_72 ();
 sg13g2_fill_8 FILLER_190_80 ();
 sg13g2_fill_8 FILLER_190_88 ();
 sg13g2_fill_8 FILLER_190_96 ();
 sg13g2_fill_8 FILLER_190_104 ();
 sg13g2_fill_8 FILLER_190_112 ();
 sg13g2_fill_8 FILLER_190_120 ();
 sg13g2_fill_8 FILLER_190_128 ();
 sg13g2_fill_8 FILLER_190_136 ();
 sg13g2_fill_8 FILLER_190_144 ();
 sg13g2_fill_8 FILLER_190_152 ();
 sg13g2_fill_8 FILLER_190_160 ();
 sg13g2_fill_8 FILLER_190_168 ();
 sg13g2_fill_8 FILLER_190_176 ();
 sg13g2_fill_8 FILLER_190_184 ();
 sg13g2_fill_8 FILLER_190_192 ();
 sg13g2_fill_8 FILLER_190_200 ();
 sg13g2_fill_8 FILLER_190_208 ();
 sg13g2_fill_8 FILLER_190_216 ();
 sg13g2_fill_8 FILLER_190_224 ();
 sg13g2_fill_8 FILLER_190_232 ();
 sg13g2_fill_8 FILLER_190_240 ();
 sg13g2_fill_8 FILLER_190_248 ();
 sg13g2_fill_8 FILLER_190_256 ();
 sg13g2_fill_8 FILLER_190_264 ();
 sg13g2_fill_8 FILLER_190_272 ();
 sg13g2_fill_8 FILLER_190_280 ();
 sg13g2_fill_8 FILLER_190_288 ();
 sg13g2_fill_8 FILLER_190_296 ();
 sg13g2_fill_8 FILLER_190_304 ();
 sg13g2_fill_8 FILLER_190_312 ();
 sg13g2_fill_8 FILLER_190_320 ();
 sg13g2_fill_8 FILLER_190_328 ();
 sg13g2_fill_8 FILLER_190_336 ();
 sg13g2_fill_8 FILLER_190_344 ();
 sg13g2_fill_8 FILLER_190_352 ();
 sg13g2_fill_8 FILLER_190_360 ();
 sg13g2_fill_8 FILLER_190_368 ();
 sg13g2_fill_8 FILLER_190_376 ();
 sg13g2_fill_8 FILLER_190_384 ();
 sg13g2_fill_8 FILLER_190_392 ();
 sg13g2_fill_8 FILLER_190_400 ();
 sg13g2_fill_8 FILLER_190_408 ();
 sg13g2_fill_8 FILLER_190_416 ();
 sg13g2_fill_8 FILLER_190_424 ();
 sg13g2_fill_8 FILLER_190_432 ();
 sg13g2_fill_8 FILLER_190_440 ();
 sg13g2_fill_8 FILLER_190_448 ();
 sg13g2_fill_8 FILLER_190_456 ();
 sg13g2_fill_8 FILLER_190_464 ();
 sg13g2_fill_8 FILLER_190_472 ();
 sg13g2_fill_8 FILLER_190_480 ();
 sg13g2_fill_8 FILLER_190_488 ();
 sg13g2_fill_8 FILLER_190_496 ();
 sg13g2_fill_8 FILLER_190_504 ();
 sg13g2_fill_8 FILLER_190_512 ();
 sg13g2_fill_8 FILLER_190_520 ();
 sg13g2_fill_8 FILLER_190_528 ();
 sg13g2_fill_8 FILLER_190_536 ();
 sg13g2_fill_8 FILLER_190_544 ();
 sg13g2_fill_8 FILLER_190_552 ();
 sg13g2_fill_8 FILLER_190_560 ();
 sg13g2_fill_8 FILLER_190_568 ();
 sg13g2_fill_8 FILLER_190_576 ();
 sg13g2_fill_8 FILLER_190_584 ();
 sg13g2_fill_8 FILLER_190_592 ();
 sg13g2_fill_8 FILLER_190_600 ();
 sg13g2_fill_8 FILLER_190_608 ();
 sg13g2_fill_8 FILLER_190_616 ();
 sg13g2_fill_8 FILLER_190_624 ();
 sg13g2_fill_8 FILLER_190_632 ();
 sg13g2_fill_8 FILLER_190_640 ();
 sg13g2_fill_8 FILLER_190_648 ();
 sg13g2_fill_8 FILLER_190_656 ();
 sg13g2_fill_8 FILLER_190_664 ();
 sg13g2_fill_8 FILLER_190_672 ();
 sg13g2_fill_8 FILLER_190_680 ();
 sg13g2_fill_8 FILLER_190_688 ();
 sg13g2_fill_8 FILLER_190_696 ();
 sg13g2_fill_8 FILLER_190_704 ();
 sg13g2_fill_8 FILLER_190_712 ();
 sg13g2_fill_8 FILLER_190_720 ();
 sg13g2_fill_8 FILLER_190_728 ();
 sg13g2_fill_8 FILLER_190_736 ();
 sg13g2_fill_8 FILLER_190_744 ();
 sg13g2_fill_8 FILLER_190_752 ();
 sg13g2_fill_8 FILLER_190_760 ();
 sg13g2_fill_8 FILLER_190_768 ();
 sg13g2_fill_8 FILLER_190_776 ();
 sg13g2_fill_8 FILLER_190_784 ();
 sg13g2_fill_8 FILLER_190_792 ();
 sg13g2_fill_8 FILLER_190_800 ();
 sg13g2_fill_8 FILLER_190_808 ();
 sg13g2_fill_8 FILLER_190_816 ();
 sg13g2_fill_8 FILLER_190_824 ();
 sg13g2_fill_8 FILLER_190_832 ();
 sg13g2_fill_8 FILLER_190_840 ();
 sg13g2_fill_8 FILLER_190_848 ();
 sg13g2_fill_8 FILLER_190_856 ();
 sg13g2_fill_8 FILLER_190_864 ();
 sg13g2_fill_8 FILLER_190_872 ();
 sg13g2_fill_8 FILLER_190_880 ();
 sg13g2_fill_8 FILLER_190_888 ();
 sg13g2_fill_8 FILLER_190_896 ();
 sg13g2_fill_8 FILLER_190_904 ();
 sg13g2_fill_8 FILLER_190_912 ();
 sg13g2_fill_8 FILLER_190_920 ();
 sg13g2_fill_8 FILLER_190_928 ();
 sg13g2_fill_8 FILLER_190_936 ();
 sg13g2_fill_8 FILLER_190_944 ();
 sg13g2_fill_8 FILLER_190_952 ();
 sg13g2_fill_8 FILLER_190_960 ();
 sg13g2_fill_8 FILLER_190_968 ();
 sg13g2_fill_8 FILLER_190_976 ();
 sg13g2_fill_8 FILLER_190_984 ();
 sg13g2_fill_8 FILLER_190_992 ();
 sg13g2_fill_4 FILLER_190_1000 ();
 sg13g2_fill_2 FILLER_190_1004 ();
 sg13g2_fill_1 FILLER_190_1006 ();
 sg13g2_fill_8 FILLER_190_1012 ();
 sg13g2_fill_1 FILLER_190_1020 ();
 sg13g2_fill_2 FILLER_190_1035 ();
 sg13g2_fill_1 FILLER_190_1037 ();
 sg13g2_fill_4 FILLER_190_1058 ();
 sg13g2_fill_1 FILLER_190_1062 ();
 sg13g2_fill_8 FILLER_190_1083 ();
 sg13g2_fill_2 FILLER_190_1091 ();
 sg13g2_fill_1 FILLER_190_1093 ();
 sg13g2_fill_4 FILLER_190_1113 ();
 sg13g2_fill_1 FILLER_190_1134 ();
 sg13g2_fill_4 FILLER_190_1147 ();
 sg13g2_fill_2 FILLER_190_1151 ();
 sg13g2_fill_2 FILLER_190_1183 ();
 sg13g2_fill_1 FILLER_190_1185 ();
 sg13g2_fill_8 FILLER_190_1199 ();
 sg13g2_fill_8 FILLER_190_1207 ();
 sg13g2_fill_2 FILLER_190_1215 ();
 sg13g2_fill_1 FILLER_190_1217 ();
 sg13g2_fill_2 FILLER_190_1246 ();
 sg13g2_fill_8 FILLER_190_1256 ();
 sg13g2_fill_1 FILLER_190_1279 ();
 sg13g2_fill_8 FILLER_190_1292 ();
 sg13g2_fill_1 FILLER_190_1300 ();
 sg13g2_fill_2 FILLER_190_1308 ();
 sg13g2_fill_1 FILLER_190_1310 ();
 sg13g2_fill_1 FILLER_190_1352 ();
 sg13g2_fill_8 FILLER_190_1371 ();
 sg13g2_fill_2 FILLER_190_1379 ();
 sg13g2_fill_1 FILLER_190_1381 ();
 sg13g2_fill_2 FILLER_190_1398 ();
 sg13g2_fill_4 FILLER_190_1405 ();
 sg13g2_fill_8 FILLER_190_1418 ();
 sg13g2_fill_8 FILLER_190_1426 ();
 sg13g2_fill_8 FILLER_190_1434 ();
 sg13g2_fill_8 FILLER_190_1442 ();
 sg13g2_fill_8 FILLER_190_1450 ();
 sg13g2_fill_8 FILLER_190_1458 ();
 sg13g2_fill_8 FILLER_190_1466 ();
 sg13g2_fill_8 FILLER_190_1474 ();
 sg13g2_fill_8 FILLER_190_1482 ();
 sg13g2_fill_8 FILLER_190_1490 ();
 sg13g2_fill_8 FILLER_190_1498 ();
 sg13g2_fill_8 FILLER_190_1506 ();
 sg13g2_fill_8 FILLER_190_1514 ();
 sg13g2_fill_8 FILLER_190_1522 ();
 sg13g2_fill_8 FILLER_190_1530 ();
 sg13g2_fill_8 FILLER_190_1538 ();
 sg13g2_fill_8 FILLER_190_1546 ();
 sg13g2_fill_8 FILLER_190_1554 ();
 sg13g2_fill_8 FILLER_190_1562 ();
 sg13g2_fill_8 FILLER_190_1570 ();
 sg13g2_fill_8 FILLER_190_1578 ();
 sg13g2_fill_4 FILLER_190_1586 ();
 sg13g2_fill_2 FILLER_190_1590 ();
 sg13g2_fill_8 FILLER_191_0 ();
 sg13g2_fill_8 FILLER_191_8 ();
 sg13g2_fill_8 FILLER_191_16 ();
 sg13g2_fill_8 FILLER_191_24 ();
 sg13g2_fill_8 FILLER_191_32 ();
 sg13g2_fill_8 FILLER_191_40 ();
 sg13g2_fill_8 FILLER_191_48 ();
 sg13g2_fill_8 FILLER_191_56 ();
 sg13g2_fill_8 FILLER_191_64 ();
 sg13g2_fill_8 FILLER_191_72 ();
 sg13g2_fill_8 FILLER_191_80 ();
 sg13g2_fill_8 FILLER_191_88 ();
 sg13g2_fill_8 FILLER_191_96 ();
 sg13g2_fill_8 FILLER_191_104 ();
 sg13g2_fill_8 FILLER_191_112 ();
 sg13g2_fill_8 FILLER_191_120 ();
 sg13g2_fill_8 FILLER_191_128 ();
 sg13g2_fill_8 FILLER_191_136 ();
 sg13g2_fill_8 FILLER_191_144 ();
 sg13g2_fill_8 FILLER_191_152 ();
 sg13g2_fill_8 FILLER_191_160 ();
 sg13g2_fill_8 FILLER_191_168 ();
 sg13g2_fill_8 FILLER_191_176 ();
 sg13g2_fill_8 FILLER_191_184 ();
 sg13g2_fill_8 FILLER_191_192 ();
 sg13g2_fill_8 FILLER_191_200 ();
 sg13g2_fill_8 FILLER_191_208 ();
 sg13g2_fill_8 FILLER_191_216 ();
 sg13g2_fill_8 FILLER_191_224 ();
 sg13g2_fill_8 FILLER_191_232 ();
 sg13g2_fill_8 FILLER_191_240 ();
 sg13g2_fill_8 FILLER_191_248 ();
 sg13g2_fill_8 FILLER_191_256 ();
 sg13g2_fill_8 FILLER_191_264 ();
 sg13g2_fill_8 FILLER_191_272 ();
 sg13g2_fill_8 FILLER_191_280 ();
 sg13g2_fill_8 FILLER_191_288 ();
 sg13g2_fill_8 FILLER_191_296 ();
 sg13g2_fill_8 FILLER_191_304 ();
 sg13g2_fill_8 FILLER_191_312 ();
 sg13g2_fill_8 FILLER_191_320 ();
 sg13g2_fill_8 FILLER_191_328 ();
 sg13g2_fill_8 FILLER_191_336 ();
 sg13g2_fill_8 FILLER_191_344 ();
 sg13g2_fill_8 FILLER_191_352 ();
 sg13g2_fill_8 FILLER_191_360 ();
 sg13g2_fill_8 FILLER_191_368 ();
 sg13g2_fill_8 FILLER_191_376 ();
 sg13g2_fill_8 FILLER_191_384 ();
 sg13g2_fill_8 FILLER_191_392 ();
 sg13g2_fill_8 FILLER_191_400 ();
 sg13g2_fill_8 FILLER_191_408 ();
 sg13g2_fill_8 FILLER_191_416 ();
 sg13g2_fill_8 FILLER_191_424 ();
 sg13g2_fill_8 FILLER_191_432 ();
 sg13g2_fill_8 FILLER_191_440 ();
 sg13g2_fill_8 FILLER_191_448 ();
 sg13g2_fill_8 FILLER_191_456 ();
 sg13g2_fill_8 FILLER_191_464 ();
 sg13g2_fill_8 FILLER_191_472 ();
 sg13g2_fill_8 FILLER_191_480 ();
 sg13g2_fill_8 FILLER_191_488 ();
 sg13g2_fill_8 FILLER_191_496 ();
 sg13g2_fill_8 FILLER_191_504 ();
 sg13g2_fill_8 FILLER_191_512 ();
 sg13g2_fill_8 FILLER_191_520 ();
 sg13g2_fill_8 FILLER_191_528 ();
 sg13g2_fill_8 FILLER_191_536 ();
 sg13g2_fill_8 FILLER_191_544 ();
 sg13g2_fill_8 FILLER_191_552 ();
 sg13g2_fill_8 FILLER_191_560 ();
 sg13g2_fill_8 FILLER_191_568 ();
 sg13g2_fill_8 FILLER_191_576 ();
 sg13g2_fill_8 FILLER_191_584 ();
 sg13g2_fill_8 FILLER_191_592 ();
 sg13g2_fill_8 FILLER_191_600 ();
 sg13g2_fill_8 FILLER_191_608 ();
 sg13g2_fill_8 FILLER_191_616 ();
 sg13g2_fill_8 FILLER_191_624 ();
 sg13g2_fill_8 FILLER_191_632 ();
 sg13g2_fill_8 FILLER_191_640 ();
 sg13g2_fill_8 FILLER_191_648 ();
 sg13g2_fill_8 FILLER_191_656 ();
 sg13g2_fill_8 FILLER_191_664 ();
 sg13g2_fill_8 FILLER_191_672 ();
 sg13g2_fill_8 FILLER_191_680 ();
 sg13g2_fill_8 FILLER_191_688 ();
 sg13g2_fill_8 FILLER_191_696 ();
 sg13g2_fill_8 FILLER_191_704 ();
 sg13g2_fill_8 FILLER_191_712 ();
 sg13g2_fill_8 FILLER_191_720 ();
 sg13g2_fill_8 FILLER_191_728 ();
 sg13g2_fill_8 FILLER_191_736 ();
 sg13g2_fill_8 FILLER_191_744 ();
 sg13g2_fill_8 FILLER_191_752 ();
 sg13g2_fill_8 FILLER_191_760 ();
 sg13g2_fill_8 FILLER_191_768 ();
 sg13g2_fill_8 FILLER_191_776 ();
 sg13g2_fill_8 FILLER_191_784 ();
 sg13g2_fill_8 FILLER_191_792 ();
 sg13g2_fill_8 FILLER_191_800 ();
 sg13g2_fill_8 FILLER_191_808 ();
 sg13g2_fill_8 FILLER_191_816 ();
 sg13g2_fill_8 FILLER_191_824 ();
 sg13g2_fill_8 FILLER_191_832 ();
 sg13g2_fill_8 FILLER_191_840 ();
 sg13g2_fill_8 FILLER_191_848 ();
 sg13g2_fill_8 FILLER_191_856 ();
 sg13g2_fill_8 FILLER_191_864 ();
 sg13g2_fill_8 FILLER_191_872 ();
 sg13g2_fill_8 FILLER_191_880 ();
 sg13g2_fill_8 FILLER_191_888 ();
 sg13g2_fill_8 FILLER_191_896 ();
 sg13g2_fill_8 FILLER_191_904 ();
 sg13g2_fill_8 FILLER_191_912 ();
 sg13g2_fill_8 FILLER_191_920 ();
 sg13g2_fill_8 FILLER_191_928 ();
 sg13g2_fill_8 FILLER_191_936 ();
 sg13g2_fill_8 FILLER_191_944 ();
 sg13g2_fill_8 FILLER_191_952 ();
 sg13g2_fill_8 FILLER_191_960 ();
 sg13g2_fill_8 FILLER_191_968 ();
 sg13g2_fill_8 FILLER_191_976 ();
 sg13g2_fill_8 FILLER_191_984 ();
 sg13g2_fill_8 FILLER_191_992 ();
 sg13g2_fill_4 FILLER_191_1000 ();
 sg13g2_fill_2 FILLER_191_1004 ();
 sg13g2_fill_4 FILLER_191_1030 ();
 sg13g2_fill_2 FILLER_191_1034 ();
 sg13g2_fill_1 FILLER_191_1058 ();
 sg13g2_fill_8 FILLER_191_1084 ();
 sg13g2_fill_2 FILLER_191_1092 ();
 sg13g2_fill_1 FILLER_191_1114 ();
 sg13g2_fill_8 FILLER_191_1135 ();
 sg13g2_fill_1 FILLER_191_1143 ();
 sg13g2_fill_4 FILLER_191_1150 ();
 sg13g2_fill_2 FILLER_191_1154 ();
 sg13g2_fill_1 FILLER_191_1156 ();
 sg13g2_fill_8 FILLER_191_1167 ();
 sg13g2_fill_4 FILLER_191_1175 ();
 sg13g2_fill_2 FILLER_191_1179 ();
 sg13g2_fill_4 FILLER_191_1189 ();
 sg13g2_fill_1 FILLER_191_1199 ();
 sg13g2_fill_8 FILLER_191_1206 ();
 sg13g2_fill_8 FILLER_191_1214 ();
 sg13g2_fill_4 FILLER_191_1222 ();
 sg13g2_fill_2 FILLER_191_1226 ();
 sg13g2_fill_8 FILLER_191_1246 ();
 sg13g2_fill_8 FILLER_191_1254 ();
 sg13g2_fill_8 FILLER_191_1262 ();
 sg13g2_fill_2 FILLER_191_1279 ();
 sg13g2_fill_1 FILLER_191_1281 ();
 sg13g2_fill_1 FILLER_191_1288 ();
 sg13g2_fill_4 FILLER_191_1308 ();
 sg13g2_fill_1 FILLER_191_1312 ();
 sg13g2_fill_2 FILLER_191_1356 ();
 sg13g2_fill_4 FILLER_191_1374 ();
 sg13g2_fill_8 FILLER_191_1386 ();
 sg13g2_fill_4 FILLER_191_1394 ();
 sg13g2_fill_2 FILLER_191_1398 ();
 sg13g2_fill_8 FILLER_191_1412 ();
 sg13g2_fill_8 FILLER_191_1420 ();
 sg13g2_fill_8 FILLER_191_1428 ();
 sg13g2_fill_8 FILLER_191_1436 ();
 sg13g2_fill_8 FILLER_191_1444 ();
 sg13g2_fill_8 FILLER_191_1452 ();
 sg13g2_fill_8 FILLER_191_1460 ();
 sg13g2_fill_8 FILLER_191_1468 ();
 sg13g2_fill_8 FILLER_191_1476 ();
 sg13g2_fill_8 FILLER_191_1484 ();
 sg13g2_fill_8 FILLER_191_1492 ();
 sg13g2_fill_8 FILLER_191_1500 ();
 sg13g2_fill_8 FILLER_191_1508 ();
 sg13g2_fill_8 FILLER_191_1516 ();
 sg13g2_fill_8 FILLER_191_1524 ();
 sg13g2_fill_8 FILLER_191_1532 ();
 sg13g2_fill_8 FILLER_191_1540 ();
 sg13g2_fill_8 FILLER_191_1548 ();
 sg13g2_fill_8 FILLER_191_1556 ();
 sg13g2_fill_8 FILLER_191_1564 ();
 sg13g2_fill_8 FILLER_191_1572 ();
 sg13g2_fill_8 FILLER_191_1580 ();
 sg13g2_fill_4 FILLER_191_1588 ();
 sg13g2_fill_8 FILLER_192_0 ();
 sg13g2_fill_8 FILLER_192_8 ();
 sg13g2_fill_8 FILLER_192_16 ();
 sg13g2_fill_8 FILLER_192_24 ();
 sg13g2_fill_8 FILLER_192_32 ();
 sg13g2_fill_8 FILLER_192_40 ();
 sg13g2_fill_8 FILLER_192_48 ();
 sg13g2_fill_8 FILLER_192_56 ();
 sg13g2_fill_8 FILLER_192_64 ();
 sg13g2_fill_8 FILLER_192_72 ();
 sg13g2_fill_8 FILLER_192_80 ();
 sg13g2_fill_8 FILLER_192_88 ();
 sg13g2_fill_8 FILLER_192_96 ();
 sg13g2_fill_8 FILLER_192_104 ();
 sg13g2_fill_8 FILLER_192_112 ();
 sg13g2_fill_8 FILLER_192_120 ();
 sg13g2_fill_8 FILLER_192_128 ();
 sg13g2_fill_8 FILLER_192_136 ();
 sg13g2_fill_8 FILLER_192_144 ();
 sg13g2_fill_8 FILLER_192_152 ();
 sg13g2_fill_8 FILLER_192_160 ();
 sg13g2_fill_8 FILLER_192_168 ();
 sg13g2_fill_8 FILLER_192_176 ();
 sg13g2_fill_8 FILLER_192_184 ();
 sg13g2_fill_8 FILLER_192_192 ();
 sg13g2_fill_8 FILLER_192_200 ();
 sg13g2_fill_8 FILLER_192_208 ();
 sg13g2_fill_8 FILLER_192_216 ();
 sg13g2_fill_8 FILLER_192_224 ();
 sg13g2_fill_8 FILLER_192_232 ();
 sg13g2_fill_8 FILLER_192_240 ();
 sg13g2_fill_8 FILLER_192_248 ();
 sg13g2_fill_8 FILLER_192_256 ();
 sg13g2_fill_8 FILLER_192_264 ();
 sg13g2_fill_8 FILLER_192_272 ();
 sg13g2_fill_8 FILLER_192_280 ();
 sg13g2_fill_8 FILLER_192_288 ();
 sg13g2_fill_8 FILLER_192_296 ();
 sg13g2_fill_8 FILLER_192_304 ();
 sg13g2_fill_8 FILLER_192_312 ();
 sg13g2_fill_8 FILLER_192_320 ();
 sg13g2_fill_8 FILLER_192_328 ();
 sg13g2_fill_8 FILLER_192_336 ();
 sg13g2_fill_8 FILLER_192_344 ();
 sg13g2_fill_8 FILLER_192_352 ();
 sg13g2_fill_8 FILLER_192_360 ();
 sg13g2_fill_8 FILLER_192_368 ();
 sg13g2_fill_8 FILLER_192_376 ();
 sg13g2_fill_8 FILLER_192_384 ();
 sg13g2_fill_8 FILLER_192_392 ();
 sg13g2_fill_8 FILLER_192_400 ();
 sg13g2_fill_8 FILLER_192_408 ();
 sg13g2_fill_8 FILLER_192_416 ();
 sg13g2_fill_8 FILLER_192_424 ();
 sg13g2_fill_8 FILLER_192_432 ();
 sg13g2_fill_8 FILLER_192_440 ();
 sg13g2_fill_8 FILLER_192_448 ();
 sg13g2_fill_8 FILLER_192_456 ();
 sg13g2_fill_8 FILLER_192_464 ();
 sg13g2_fill_8 FILLER_192_472 ();
 sg13g2_fill_8 FILLER_192_480 ();
 sg13g2_fill_8 FILLER_192_488 ();
 sg13g2_fill_8 FILLER_192_496 ();
 sg13g2_fill_8 FILLER_192_504 ();
 sg13g2_fill_8 FILLER_192_512 ();
 sg13g2_fill_8 FILLER_192_520 ();
 sg13g2_fill_8 FILLER_192_528 ();
 sg13g2_fill_8 FILLER_192_536 ();
 sg13g2_fill_8 FILLER_192_544 ();
 sg13g2_fill_8 FILLER_192_552 ();
 sg13g2_fill_8 FILLER_192_560 ();
 sg13g2_fill_8 FILLER_192_568 ();
 sg13g2_fill_8 FILLER_192_576 ();
 sg13g2_fill_8 FILLER_192_584 ();
 sg13g2_fill_8 FILLER_192_592 ();
 sg13g2_fill_8 FILLER_192_600 ();
 sg13g2_fill_8 FILLER_192_608 ();
 sg13g2_fill_8 FILLER_192_616 ();
 sg13g2_fill_8 FILLER_192_624 ();
 sg13g2_fill_8 FILLER_192_632 ();
 sg13g2_fill_8 FILLER_192_640 ();
 sg13g2_fill_8 FILLER_192_648 ();
 sg13g2_fill_8 FILLER_192_656 ();
 sg13g2_fill_8 FILLER_192_664 ();
 sg13g2_fill_8 FILLER_192_672 ();
 sg13g2_fill_8 FILLER_192_680 ();
 sg13g2_fill_8 FILLER_192_688 ();
 sg13g2_fill_8 FILLER_192_696 ();
 sg13g2_fill_8 FILLER_192_704 ();
 sg13g2_fill_8 FILLER_192_712 ();
 sg13g2_fill_8 FILLER_192_720 ();
 sg13g2_fill_8 FILLER_192_728 ();
 sg13g2_fill_8 FILLER_192_736 ();
 sg13g2_fill_8 FILLER_192_744 ();
 sg13g2_fill_8 FILLER_192_752 ();
 sg13g2_fill_8 FILLER_192_760 ();
 sg13g2_fill_8 FILLER_192_768 ();
 sg13g2_fill_8 FILLER_192_776 ();
 sg13g2_fill_8 FILLER_192_784 ();
 sg13g2_fill_8 FILLER_192_792 ();
 sg13g2_fill_8 FILLER_192_800 ();
 sg13g2_fill_8 FILLER_192_808 ();
 sg13g2_fill_8 FILLER_192_816 ();
 sg13g2_fill_8 FILLER_192_824 ();
 sg13g2_fill_8 FILLER_192_832 ();
 sg13g2_fill_8 FILLER_192_840 ();
 sg13g2_fill_8 FILLER_192_848 ();
 sg13g2_fill_8 FILLER_192_856 ();
 sg13g2_fill_8 FILLER_192_864 ();
 sg13g2_fill_8 FILLER_192_872 ();
 sg13g2_fill_8 FILLER_192_880 ();
 sg13g2_fill_8 FILLER_192_888 ();
 sg13g2_fill_8 FILLER_192_896 ();
 sg13g2_fill_8 FILLER_192_904 ();
 sg13g2_fill_8 FILLER_192_912 ();
 sg13g2_fill_8 FILLER_192_920 ();
 sg13g2_fill_8 FILLER_192_928 ();
 sg13g2_fill_8 FILLER_192_936 ();
 sg13g2_fill_8 FILLER_192_944 ();
 sg13g2_fill_8 FILLER_192_952 ();
 sg13g2_fill_8 FILLER_192_960 ();
 sg13g2_fill_8 FILLER_192_968 ();
 sg13g2_fill_8 FILLER_192_976 ();
 sg13g2_fill_8 FILLER_192_984 ();
 sg13g2_fill_8 FILLER_192_992 ();
 sg13g2_fill_8 FILLER_192_1000 ();
 sg13g2_fill_8 FILLER_192_1008 ();
 sg13g2_fill_2 FILLER_192_1016 ();
 sg13g2_fill_8 FILLER_192_1023 ();
 sg13g2_fill_8 FILLER_192_1031 ();
 sg13g2_fill_8 FILLER_192_1039 ();
 sg13g2_fill_8 FILLER_192_1047 ();
 sg13g2_fill_2 FILLER_192_1055 ();
 sg13g2_fill_4 FILLER_192_1062 ();
 sg13g2_fill_2 FILLER_192_1066 ();
 sg13g2_fill_1 FILLER_192_1068 ();
 sg13g2_fill_8 FILLER_192_1077 ();
 sg13g2_fill_8 FILLER_192_1085 ();
 sg13g2_fill_8 FILLER_192_1093 ();
 sg13g2_fill_8 FILLER_192_1101 ();
 sg13g2_fill_8 FILLER_192_1122 ();
 sg13g2_fill_8 FILLER_192_1130 ();
 sg13g2_fill_2 FILLER_192_1150 ();
 sg13g2_fill_2 FILLER_192_1157 ();
 sg13g2_fill_1 FILLER_192_1159 ();
 sg13g2_fill_2 FILLER_192_1168 ();
 sg13g2_fill_8 FILLER_192_1175 ();
 sg13g2_fill_8 FILLER_192_1183 ();
 sg13g2_fill_2 FILLER_192_1191 ();
 sg13g2_fill_2 FILLER_192_1227 ();
 sg13g2_fill_1 FILLER_192_1229 ();
 sg13g2_fill_2 FILLER_192_1238 ();
 sg13g2_fill_8 FILLER_192_1248 ();
 sg13g2_fill_2 FILLER_192_1256 ();
 sg13g2_fill_1 FILLER_192_1258 ();
 sg13g2_fill_2 FILLER_192_1276 ();
 sg13g2_fill_1 FILLER_192_1278 ();
 sg13g2_fill_8 FILLER_192_1287 ();
 sg13g2_fill_4 FILLER_192_1295 ();
 sg13g2_fill_2 FILLER_192_1299 ();
 sg13g2_fill_8 FILLER_192_1308 ();
 sg13g2_fill_8 FILLER_192_1321 ();
 sg13g2_fill_4 FILLER_192_1329 ();
 sg13g2_fill_2 FILLER_192_1333 ();
 sg13g2_fill_1 FILLER_192_1335 ();
 sg13g2_fill_2 FILLER_192_1342 ();
 sg13g2_fill_1 FILLER_192_1344 ();
 sg13g2_fill_2 FILLER_192_1354 ();
 sg13g2_fill_1 FILLER_192_1356 ();
 sg13g2_fill_2 FILLER_192_1362 ();
 sg13g2_fill_1 FILLER_192_1364 ();
 sg13g2_fill_8 FILLER_192_1374 ();
 sg13g2_fill_8 FILLER_192_1382 ();
 sg13g2_fill_4 FILLER_192_1390 ();
 sg13g2_fill_1 FILLER_192_1394 ();
 sg13g2_fill_8 FILLER_192_1408 ();
 sg13g2_fill_8 FILLER_192_1416 ();
 sg13g2_fill_8 FILLER_192_1424 ();
 sg13g2_fill_8 FILLER_192_1432 ();
 sg13g2_fill_8 FILLER_192_1440 ();
 sg13g2_fill_8 FILLER_192_1448 ();
 sg13g2_fill_8 FILLER_192_1456 ();
 sg13g2_fill_8 FILLER_192_1464 ();
 sg13g2_fill_8 FILLER_192_1472 ();
 sg13g2_fill_8 FILLER_192_1480 ();
 sg13g2_fill_8 FILLER_192_1488 ();
 sg13g2_fill_8 FILLER_192_1496 ();
 sg13g2_fill_8 FILLER_192_1504 ();
 sg13g2_fill_8 FILLER_192_1512 ();
 sg13g2_fill_8 FILLER_192_1520 ();
 sg13g2_fill_8 FILLER_192_1528 ();
 sg13g2_fill_8 FILLER_192_1536 ();
 sg13g2_fill_8 FILLER_192_1544 ();
 sg13g2_fill_8 FILLER_192_1552 ();
 sg13g2_fill_8 FILLER_192_1560 ();
 sg13g2_fill_8 FILLER_192_1568 ();
 sg13g2_fill_8 FILLER_192_1576 ();
 sg13g2_fill_8 FILLER_192_1584 ();
 sg13g2_fill_8 FILLER_193_0 ();
 sg13g2_fill_8 FILLER_193_8 ();
 sg13g2_fill_8 FILLER_193_16 ();
 sg13g2_fill_8 FILLER_193_24 ();
 sg13g2_fill_8 FILLER_193_32 ();
 sg13g2_fill_8 FILLER_193_40 ();
 sg13g2_fill_8 FILLER_193_48 ();
 sg13g2_fill_8 FILLER_193_56 ();
 sg13g2_fill_8 FILLER_193_64 ();
 sg13g2_fill_8 FILLER_193_72 ();
 sg13g2_fill_8 FILLER_193_80 ();
 sg13g2_fill_8 FILLER_193_88 ();
 sg13g2_fill_8 FILLER_193_96 ();
 sg13g2_fill_8 FILLER_193_104 ();
 sg13g2_fill_8 FILLER_193_112 ();
 sg13g2_fill_8 FILLER_193_120 ();
 sg13g2_fill_8 FILLER_193_128 ();
 sg13g2_fill_8 FILLER_193_136 ();
 sg13g2_fill_8 FILLER_193_144 ();
 sg13g2_fill_8 FILLER_193_152 ();
 sg13g2_fill_8 FILLER_193_160 ();
 sg13g2_fill_8 FILLER_193_168 ();
 sg13g2_fill_8 FILLER_193_176 ();
 sg13g2_fill_8 FILLER_193_184 ();
 sg13g2_fill_8 FILLER_193_192 ();
 sg13g2_fill_8 FILLER_193_200 ();
 sg13g2_fill_8 FILLER_193_208 ();
 sg13g2_fill_8 FILLER_193_216 ();
 sg13g2_fill_8 FILLER_193_224 ();
 sg13g2_fill_8 FILLER_193_232 ();
 sg13g2_fill_8 FILLER_193_240 ();
 sg13g2_fill_8 FILLER_193_248 ();
 sg13g2_fill_8 FILLER_193_256 ();
 sg13g2_fill_8 FILLER_193_264 ();
 sg13g2_fill_8 FILLER_193_272 ();
 sg13g2_fill_8 FILLER_193_280 ();
 sg13g2_fill_8 FILLER_193_288 ();
 sg13g2_fill_8 FILLER_193_296 ();
 sg13g2_fill_8 FILLER_193_304 ();
 sg13g2_fill_8 FILLER_193_312 ();
 sg13g2_fill_8 FILLER_193_320 ();
 sg13g2_fill_8 FILLER_193_328 ();
 sg13g2_fill_8 FILLER_193_336 ();
 sg13g2_fill_8 FILLER_193_344 ();
 sg13g2_fill_8 FILLER_193_352 ();
 sg13g2_fill_8 FILLER_193_360 ();
 sg13g2_fill_8 FILLER_193_368 ();
 sg13g2_fill_8 FILLER_193_376 ();
 sg13g2_fill_8 FILLER_193_384 ();
 sg13g2_fill_8 FILLER_193_392 ();
 sg13g2_fill_8 FILLER_193_400 ();
 sg13g2_fill_8 FILLER_193_408 ();
 sg13g2_fill_8 FILLER_193_416 ();
 sg13g2_fill_8 FILLER_193_424 ();
 sg13g2_fill_8 FILLER_193_432 ();
 sg13g2_fill_8 FILLER_193_440 ();
 sg13g2_fill_8 FILLER_193_448 ();
 sg13g2_fill_8 FILLER_193_456 ();
 sg13g2_fill_8 FILLER_193_464 ();
 sg13g2_fill_8 FILLER_193_472 ();
 sg13g2_fill_8 FILLER_193_480 ();
 sg13g2_fill_8 FILLER_193_488 ();
 sg13g2_fill_8 FILLER_193_496 ();
 sg13g2_fill_8 FILLER_193_504 ();
 sg13g2_fill_8 FILLER_193_512 ();
 sg13g2_fill_8 FILLER_193_520 ();
 sg13g2_fill_8 FILLER_193_528 ();
 sg13g2_fill_8 FILLER_193_536 ();
 sg13g2_fill_8 FILLER_193_544 ();
 sg13g2_fill_8 FILLER_193_552 ();
 sg13g2_fill_8 FILLER_193_560 ();
 sg13g2_fill_8 FILLER_193_568 ();
 sg13g2_fill_8 FILLER_193_576 ();
 sg13g2_fill_8 FILLER_193_584 ();
 sg13g2_fill_8 FILLER_193_592 ();
 sg13g2_fill_8 FILLER_193_600 ();
 sg13g2_fill_8 FILLER_193_608 ();
 sg13g2_fill_8 FILLER_193_616 ();
 sg13g2_fill_8 FILLER_193_624 ();
 sg13g2_fill_8 FILLER_193_632 ();
 sg13g2_fill_8 FILLER_193_640 ();
 sg13g2_fill_8 FILLER_193_648 ();
 sg13g2_fill_8 FILLER_193_656 ();
 sg13g2_fill_8 FILLER_193_664 ();
 sg13g2_fill_8 FILLER_193_672 ();
 sg13g2_fill_8 FILLER_193_680 ();
 sg13g2_fill_8 FILLER_193_688 ();
 sg13g2_fill_8 FILLER_193_696 ();
 sg13g2_fill_8 FILLER_193_704 ();
 sg13g2_fill_8 FILLER_193_712 ();
 sg13g2_fill_8 FILLER_193_720 ();
 sg13g2_fill_8 FILLER_193_728 ();
 sg13g2_fill_8 FILLER_193_736 ();
 sg13g2_fill_8 FILLER_193_744 ();
 sg13g2_fill_8 FILLER_193_752 ();
 sg13g2_fill_8 FILLER_193_760 ();
 sg13g2_fill_8 FILLER_193_768 ();
 sg13g2_fill_8 FILLER_193_776 ();
 sg13g2_fill_8 FILLER_193_784 ();
 sg13g2_fill_8 FILLER_193_792 ();
 sg13g2_fill_8 FILLER_193_800 ();
 sg13g2_fill_8 FILLER_193_808 ();
 sg13g2_fill_8 FILLER_193_816 ();
 sg13g2_fill_8 FILLER_193_824 ();
 sg13g2_fill_8 FILLER_193_832 ();
 sg13g2_fill_8 FILLER_193_840 ();
 sg13g2_fill_8 FILLER_193_848 ();
 sg13g2_fill_8 FILLER_193_856 ();
 sg13g2_fill_8 FILLER_193_864 ();
 sg13g2_fill_8 FILLER_193_872 ();
 sg13g2_fill_8 FILLER_193_880 ();
 sg13g2_fill_8 FILLER_193_888 ();
 sg13g2_fill_8 FILLER_193_896 ();
 sg13g2_fill_8 FILLER_193_904 ();
 sg13g2_fill_8 FILLER_193_912 ();
 sg13g2_fill_8 FILLER_193_920 ();
 sg13g2_fill_8 FILLER_193_928 ();
 sg13g2_fill_8 FILLER_193_936 ();
 sg13g2_fill_8 FILLER_193_944 ();
 sg13g2_fill_8 FILLER_193_952 ();
 sg13g2_fill_8 FILLER_193_960 ();
 sg13g2_fill_8 FILLER_193_968 ();
 sg13g2_fill_8 FILLER_193_976 ();
 sg13g2_fill_8 FILLER_193_984 ();
 sg13g2_fill_8 FILLER_193_992 ();
 sg13g2_fill_8 FILLER_193_1000 ();
 sg13g2_fill_4 FILLER_193_1008 ();
 sg13g2_fill_2 FILLER_193_1012 ();
 sg13g2_fill_1 FILLER_193_1018 ();
 sg13g2_fill_8 FILLER_193_1040 ();
 sg13g2_fill_2 FILLER_193_1048 ();
 sg13g2_fill_1 FILLER_193_1050 ();
 sg13g2_fill_2 FILLER_193_1059 ();
 sg13g2_fill_8 FILLER_193_1071 ();
 sg13g2_fill_4 FILLER_193_1079 ();
 sg13g2_fill_2 FILLER_193_1083 ();
 sg13g2_fill_8 FILLER_193_1097 ();
 sg13g2_fill_1 FILLER_193_1105 ();
 sg13g2_fill_1 FILLER_193_1119 ();
 sg13g2_fill_4 FILLER_193_1138 ();
 sg13g2_fill_2 FILLER_193_1142 ();
 sg13g2_fill_1 FILLER_193_1144 ();
 sg13g2_fill_8 FILLER_193_1153 ();
 sg13g2_fill_2 FILLER_193_1171 ();
 sg13g2_fill_8 FILLER_193_1193 ();
 sg13g2_fill_8 FILLER_193_1201 ();
 sg13g2_fill_4 FILLER_193_1223 ();
 sg13g2_fill_2 FILLER_193_1227 ();
 sg13g2_fill_2 FILLER_193_1258 ();
 sg13g2_fill_1 FILLER_193_1260 ();
 sg13g2_fill_8 FILLER_193_1273 ();
 sg13g2_fill_1 FILLER_193_1281 ();
 sg13g2_fill_1 FILLER_193_1292 ();
 sg13g2_fill_4 FILLER_193_1315 ();
 sg13g2_fill_8 FILLER_193_1326 ();
 sg13g2_fill_8 FILLER_193_1334 ();
 sg13g2_fill_2 FILLER_193_1342 ();
 sg13g2_fill_2 FILLER_193_1387 ();
 sg13g2_fill_8 FILLER_193_1415 ();
 sg13g2_fill_8 FILLER_193_1423 ();
 sg13g2_fill_8 FILLER_193_1431 ();
 sg13g2_fill_8 FILLER_193_1439 ();
 sg13g2_fill_8 FILLER_193_1447 ();
 sg13g2_fill_8 FILLER_193_1455 ();
 sg13g2_fill_8 FILLER_193_1463 ();
 sg13g2_fill_8 FILLER_193_1471 ();
 sg13g2_fill_8 FILLER_193_1479 ();
 sg13g2_fill_8 FILLER_193_1487 ();
 sg13g2_fill_8 FILLER_193_1495 ();
 sg13g2_fill_8 FILLER_193_1503 ();
 sg13g2_fill_8 FILLER_193_1511 ();
 sg13g2_fill_8 FILLER_193_1519 ();
 sg13g2_fill_8 FILLER_193_1527 ();
 sg13g2_fill_8 FILLER_193_1535 ();
 sg13g2_fill_8 FILLER_193_1543 ();
 sg13g2_fill_8 FILLER_193_1551 ();
 sg13g2_fill_8 FILLER_193_1559 ();
 sg13g2_fill_8 FILLER_193_1567 ();
 sg13g2_fill_8 FILLER_193_1575 ();
 sg13g2_fill_8 FILLER_193_1583 ();
 sg13g2_fill_1 FILLER_193_1591 ();
 sg13g2_fill_8 FILLER_194_0 ();
 sg13g2_fill_8 FILLER_194_8 ();
 sg13g2_fill_8 FILLER_194_16 ();
 sg13g2_fill_8 FILLER_194_24 ();
 sg13g2_fill_8 FILLER_194_32 ();
 sg13g2_fill_8 FILLER_194_40 ();
 sg13g2_fill_8 FILLER_194_48 ();
 sg13g2_fill_8 FILLER_194_56 ();
 sg13g2_fill_8 FILLER_194_64 ();
 sg13g2_fill_8 FILLER_194_72 ();
 sg13g2_fill_8 FILLER_194_80 ();
 sg13g2_fill_8 FILLER_194_88 ();
 sg13g2_fill_8 FILLER_194_96 ();
 sg13g2_fill_8 FILLER_194_104 ();
 sg13g2_fill_8 FILLER_194_112 ();
 sg13g2_fill_8 FILLER_194_120 ();
 sg13g2_fill_8 FILLER_194_128 ();
 sg13g2_fill_8 FILLER_194_136 ();
 sg13g2_fill_8 FILLER_194_144 ();
 sg13g2_fill_8 FILLER_194_152 ();
 sg13g2_fill_8 FILLER_194_160 ();
 sg13g2_fill_8 FILLER_194_168 ();
 sg13g2_fill_8 FILLER_194_176 ();
 sg13g2_fill_8 FILLER_194_184 ();
 sg13g2_fill_8 FILLER_194_192 ();
 sg13g2_fill_8 FILLER_194_200 ();
 sg13g2_fill_8 FILLER_194_208 ();
 sg13g2_fill_8 FILLER_194_216 ();
 sg13g2_fill_8 FILLER_194_224 ();
 sg13g2_fill_8 FILLER_194_232 ();
 sg13g2_fill_8 FILLER_194_240 ();
 sg13g2_fill_8 FILLER_194_248 ();
 sg13g2_fill_8 FILLER_194_256 ();
 sg13g2_fill_8 FILLER_194_264 ();
 sg13g2_fill_8 FILLER_194_272 ();
 sg13g2_fill_8 FILLER_194_280 ();
 sg13g2_fill_8 FILLER_194_288 ();
 sg13g2_fill_8 FILLER_194_296 ();
 sg13g2_fill_8 FILLER_194_304 ();
 sg13g2_fill_8 FILLER_194_312 ();
 sg13g2_fill_8 FILLER_194_320 ();
 sg13g2_fill_8 FILLER_194_328 ();
 sg13g2_fill_8 FILLER_194_336 ();
 sg13g2_fill_8 FILLER_194_344 ();
 sg13g2_fill_8 FILLER_194_352 ();
 sg13g2_fill_8 FILLER_194_360 ();
 sg13g2_fill_8 FILLER_194_368 ();
 sg13g2_fill_8 FILLER_194_376 ();
 sg13g2_fill_8 FILLER_194_384 ();
 sg13g2_fill_8 FILLER_194_392 ();
 sg13g2_fill_8 FILLER_194_400 ();
 sg13g2_fill_8 FILLER_194_408 ();
 sg13g2_fill_8 FILLER_194_416 ();
 sg13g2_fill_8 FILLER_194_424 ();
 sg13g2_fill_8 FILLER_194_432 ();
 sg13g2_fill_8 FILLER_194_440 ();
 sg13g2_fill_8 FILLER_194_448 ();
 sg13g2_fill_8 FILLER_194_456 ();
 sg13g2_fill_8 FILLER_194_464 ();
 sg13g2_fill_8 FILLER_194_472 ();
 sg13g2_fill_8 FILLER_194_480 ();
 sg13g2_fill_8 FILLER_194_488 ();
 sg13g2_fill_8 FILLER_194_496 ();
 sg13g2_fill_8 FILLER_194_504 ();
 sg13g2_fill_8 FILLER_194_512 ();
 sg13g2_fill_8 FILLER_194_520 ();
 sg13g2_fill_8 FILLER_194_528 ();
 sg13g2_fill_8 FILLER_194_536 ();
 sg13g2_fill_8 FILLER_194_544 ();
 sg13g2_fill_8 FILLER_194_552 ();
 sg13g2_fill_8 FILLER_194_560 ();
 sg13g2_fill_8 FILLER_194_568 ();
 sg13g2_fill_8 FILLER_194_576 ();
 sg13g2_fill_8 FILLER_194_584 ();
 sg13g2_fill_8 FILLER_194_592 ();
 sg13g2_fill_8 FILLER_194_600 ();
 sg13g2_fill_8 FILLER_194_608 ();
 sg13g2_fill_8 FILLER_194_616 ();
 sg13g2_fill_8 FILLER_194_624 ();
 sg13g2_fill_8 FILLER_194_632 ();
 sg13g2_fill_8 FILLER_194_640 ();
 sg13g2_fill_8 FILLER_194_648 ();
 sg13g2_fill_8 FILLER_194_656 ();
 sg13g2_fill_8 FILLER_194_664 ();
 sg13g2_fill_8 FILLER_194_672 ();
 sg13g2_fill_8 FILLER_194_680 ();
 sg13g2_fill_8 FILLER_194_688 ();
 sg13g2_fill_8 FILLER_194_696 ();
 sg13g2_fill_8 FILLER_194_704 ();
 sg13g2_fill_8 FILLER_194_712 ();
 sg13g2_fill_8 FILLER_194_720 ();
 sg13g2_fill_8 FILLER_194_728 ();
 sg13g2_fill_8 FILLER_194_736 ();
 sg13g2_fill_8 FILLER_194_744 ();
 sg13g2_fill_8 FILLER_194_752 ();
 sg13g2_fill_8 FILLER_194_760 ();
 sg13g2_fill_8 FILLER_194_768 ();
 sg13g2_fill_8 FILLER_194_776 ();
 sg13g2_fill_8 FILLER_194_784 ();
 sg13g2_fill_8 FILLER_194_792 ();
 sg13g2_fill_8 FILLER_194_800 ();
 sg13g2_fill_8 FILLER_194_808 ();
 sg13g2_fill_8 FILLER_194_816 ();
 sg13g2_fill_8 FILLER_194_824 ();
 sg13g2_fill_8 FILLER_194_832 ();
 sg13g2_fill_8 FILLER_194_840 ();
 sg13g2_fill_8 FILLER_194_848 ();
 sg13g2_fill_8 FILLER_194_856 ();
 sg13g2_fill_8 FILLER_194_864 ();
 sg13g2_fill_8 FILLER_194_872 ();
 sg13g2_fill_8 FILLER_194_880 ();
 sg13g2_fill_8 FILLER_194_888 ();
 sg13g2_fill_8 FILLER_194_896 ();
 sg13g2_fill_8 FILLER_194_904 ();
 sg13g2_fill_8 FILLER_194_912 ();
 sg13g2_fill_8 FILLER_194_920 ();
 sg13g2_fill_8 FILLER_194_928 ();
 sg13g2_fill_8 FILLER_194_936 ();
 sg13g2_fill_8 FILLER_194_944 ();
 sg13g2_fill_8 FILLER_194_952 ();
 sg13g2_fill_8 FILLER_194_960 ();
 sg13g2_fill_8 FILLER_194_968 ();
 sg13g2_fill_8 FILLER_194_976 ();
 sg13g2_fill_8 FILLER_194_984 ();
 sg13g2_fill_8 FILLER_194_992 ();
 sg13g2_fill_8 FILLER_194_1000 ();
 sg13g2_fill_4 FILLER_194_1008 ();
 sg13g2_fill_1 FILLER_194_1012 ();
 sg13g2_fill_1 FILLER_194_1064 ();
 sg13g2_fill_1 FILLER_194_1078 ();
 sg13g2_fill_4 FILLER_194_1138 ();
 sg13g2_fill_2 FILLER_194_1142 ();
 sg13g2_fill_1 FILLER_194_1144 ();
 sg13g2_fill_8 FILLER_194_1161 ();
 sg13g2_fill_1 FILLER_194_1169 ();
 sg13g2_fill_8 FILLER_194_1178 ();
 sg13g2_fill_8 FILLER_194_1186 ();
 sg13g2_fill_4 FILLER_194_1194 ();
 sg13g2_fill_8 FILLER_194_1228 ();
 sg13g2_fill_4 FILLER_194_1236 ();
 sg13g2_fill_2 FILLER_194_1256 ();
 sg13g2_fill_1 FILLER_194_1258 ();
 sg13g2_fill_8 FILLER_194_1267 ();
 sg13g2_fill_8 FILLER_194_1275 ();
 sg13g2_fill_1 FILLER_194_1283 ();
 sg13g2_fill_8 FILLER_194_1291 ();
 sg13g2_fill_4 FILLER_194_1299 ();
 sg13g2_fill_1 FILLER_194_1303 ();
 sg13g2_fill_4 FILLER_194_1311 ();
 sg13g2_fill_2 FILLER_194_1315 ();
 sg13g2_fill_1 FILLER_194_1317 ();
 sg13g2_fill_2 FILLER_194_1358 ();
 sg13g2_fill_4 FILLER_194_1372 ();
 sg13g2_fill_1 FILLER_194_1376 ();
 sg13g2_fill_8 FILLER_194_1411 ();
 sg13g2_fill_8 FILLER_194_1419 ();
 sg13g2_fill_8 FILLER_194_1427 ();
 sg13g2_fill_8 FILLER_194_1435 ();
 sg13g2_fill_8 FILLER_194_1443 ();
 sg13g2_fill_8 FILLER_194_1451 ();
 sg13g2_fill_8 FILLER_194_1459 ();
 sg13g2_fill_8 FILLER_194_1467 ();
 sg13g2_fill_8 FILLER_194_1475 ();
 sg13g2_fill_8 FILLER_194_1483 ();
 sg13g2_fill_8 FILLER_194_1491 ();
 sg13g2_fill_8 FILLER_194_1499 ();
 sg13g2_fill_8 FILLER_194_1507 ();
 sg13g2_fill_8 FILLER_194_1515 ();
 sg13g2_fill_8 FILLER_194_1523 ();
 sg13g2_fill_8 FILLER_194_1531 ();
 sg13g2_fill_8 FILLER_194_1539 ();
 sg13g2_fill_8 FILLER_194_1547 ();
 sg13g2_fill_8 FILLER_194_1555 ();
 sg13g2_fill_8 FILLER_194_1563 ();
 sg13g2_fill_8 FILLER_194_1571 ();
 sg13g2_fill_8 FILLER_194_1579 ();
 sg13g2_fill_4 FILLER_194_1587 ();
 sg13g2_fill_1 FILLER_194_1591 ();
 sg13g2_fill_2 FILLER_195_0 ();
 sg13g2_fill_8 FILLER_195_15 ();
 sg13g2_fill_8 FILLER_195_23 ();
 sg13g2_fill_8 FILLER_195_31 ();
 sg13g2_fill_8 FILLER_195_39 ();
 sg13g2_fill_8 FILLER_195_47 ();
 sg13g2_fill_8 FILLER_195_55 ();
 sg13g2_fill_8 FILLER_195_63 ();
 sg13g2_fill_8 FILLER_195_71 ();
 sg13g2_fill_8 FILLER_195_79 ();
 sg13g2_fill_8 FILLER_195_87 ();
 sg13g2_fill_8 FILLER_195_95 ();
 sg13g2_fill_8 FILLER_195_103 ();
 sg13g2_fill_8 FILLER_195_111 ();
 sg13g2_fill_8 FILLER_195_119 ();
 sg13g2_fill_8 FILLER_195_127 ();
 sg13g2_fill_8 FILLER_195_135 ();
 sg13g2_fill_8 FILLER_195_143 ();
 sg13g2_fill_8 FILLER_195_151 ();
 sg13g2_fill_8 FILLER_195_159 ();
 sg13g2_fill_8 FILLER_195_167 ();
 sg13g2_fill_8 FILLER_195_175 ();
 sg13g2_fill_8 FILLER_195_183 ();
 sg13g2_fill_8 FILLER_195_191 ();
 sg13g2_fill_8 FILLER_195_199 ();
 sg13g2_fill_8 FILLER_195_207 ();
 sg13g2_fill_8 FILLER_195_215 ();
 sg13g2_fill_8 FILLER_195_223 ();
 sg13g2_fill_8 FILLER_195_231 ();
 sg13g2_fill_8 FILLER_195_239 ();
 sg13g2_fill_8 FILLER_195_247 ();
 sg13g2_fill_8 FILLER_195_255 ();
 sg13g2_fill_8 FILLER_195_263 ();
 sg13g2_fill_8 FILLER_195_271 ();
 sg13g2_fill_8 FILLER_195_279 ();
 sg13g2_fill_8 FILLER_195_287 ();
 sg13g2_fill_8 FILLER_195_295 ();
 sg13g2_fill_8 FILLER_195_303 ();
 sg13g2_fill_8 FILLER_195_311 ();
 sg13g2_fill_8 FILLER_195_319 ();
 sg13g2_fill_8 FILLER_195_327 ();
 sg13g2_fill_8 FILLER_195_335 ();
 sg13g2_fill_8 FILLER_195_343 ();
 sg13g2_fill_8 FILLER_195_351 ();
 sg13g2_fill_8 FILLER_195_359 ();
 sg13g2_fill_8 FILLER_195_367 ();
 sg13g2_fill_8 FILLER_195_375 ();
 sg13g2_fill_8 FILLER_195_383 ();
 sg13g2_fill_8 FILLER_195_391 ();
 sg13g2_fill_8 FILLER_195_399 ();
 sg13g2_fill_8 FILLER_195_407 ();
 sg13g2_fill_8 FILLER_195_415 ();
 sg13g2_fill_8 FILLER_195_423 ();
 sg13g2_fill_8 FILLER_195_431 ();
 sg13g2_fill_8 FILLER_195_439 ();
 sg13g2_fill_8 FILLER_195_447 ();
 sg13g2_fill_8 FILLER_195_455 ();
 sg13g2_fill_8 FILLER_195_463 ();
 sg13g2_fill_8 FILLER_195_471 ();
 sg13g2_fill_8 FILLER_195_479 ();
 sg13g2_fill_8 FILLER_195_487 ();
 sg13g2_fill_8 FILLER_195_495 ();
 sg13g2_fill_8 FILLER_195_503 ();
 sg13g2_fill_8 FILLER_195_511 ();
 sg13g2_fill_8 FILLER_195_519 ();
 sg13g2_fill_8 FILLER_195_527 ();
 sg13g2_fill_8 FILLER_195_535 ();
 sg13g2_fill_8 FILLER_195_543 ();
 sg13g2_fill_8 FILLER_195_551 ();
 sg13g2_fill_8 FILLER_195_559 ();
 sg13g2_fill_8 FILLER_195_567 ();
 sg13g2_fill_8 FILLER_195_575 ();
 sg13g2_fill_8 FILLER_195_583 ();
 sg13g2_fill_8 FILLER_195_591 ();
 sg13g2_fill_8 FILLER_195_599 ();
 sg13g2_fill_8 FILLER_195_607 ();
 sg13g2_fill_8 FILLER_195_615 ();
 sg13g2_fill_8 FILLER_195_623 ();
 sg13g2_fill_8 FILLER_195_631 ();
 sg13g2_fill_8 FILLER_195_639 ();
 sg13g2_fill_8 FILLER_195_647 ();
 sg13g2_fill_8 FILLER_195_655 ();
 sg13g2_fill_8 FILLER_195_663 ();
 sg13g2_fill_8 FILLER_195_671 ();
 sg13g2_fill_8 FILLER_195_679 ();
 sg13g2_fill_8 FILLER_195_687 ();
 sg13g2_fill_8 FILLER_195_695 ();
 sg13g2_fill_8 FILLER_195_703 ();
 sg13g2_fill_8 FILLER_195_711 ();
 sg13g2_fill_8 FILLER_195_719 ();
 sg13g2_fill_8 FILLER_195_727 ();
 sg13g2_fill_8 FILLER_195_735 ();
 sg13g2_fill_8 FILLER_195_743 ();
 sg13g2_fill_8 FILLER_195_751 ();
 sg13g2_fill_8 FILLER_195_759 ();
 sg13g2_fill_8 FILLER_195_767 ();
 sg13g2_fill_8 FILLER_195_775 ();
 sg13g2_fill_8 FILLER_195_783 ();
 sg13g2_fill_8 FILLER_195_791 ();
 sg13g2_fill_8 FILLER_195_799 ();
 sg13g2_fill_8 FILLER_195_807 ();
 sg13g2_fill_8 FILLER_195_815 ();
 sg13g2_fill_8 FILLER_195_823 ();
 sg13g2_fill_8 FILLER_195_831 ();
 sg13g2_fill_8 FILLER_195_839 ();
 sg13g2_fill_8 FILLER_195_847 ();
 sg13g2_fill_8 FILLER_195_855 ();
 sg13g2_fill_8 FILLER_195_863 ();
 sg13g2_fill_8 FILLER_195_871 ();
 sg13g2_fill_8 FILLER_195_879 ();
 sg13g2_fill_8 FILLER_195_887 ();
 sg13g2_fill_8 FILLER_195_895 ();
 sg13g2_fill_8 FILLER_195_903 ();
 sg13g2_fill_8 FILLER_195_911 ();
 sg13g2_fill_8 FILLER_195_919 ();
 sg13g2_fill_8 FILLER_195_927 ();
 sg13g2_fill_8 FILLER_195_935 ();
 sg13g2_fill_8 FILLER_195_943 ();
 sg13g2_fill_8 FILLER_195_951 ();
 sg13g2_fill_8 FILLER_195_959 ();
 sg13g2_fill_8 FILLER_195_967 ();
 sg13g2_fill_8 FILLER_195_975 ();
 sg13g2_fill_8 FILLER_195_983 ();
 sg13g2_fill_8 FILLER_195_991 ();
 sg13g2_fill_8 FILLER_195_999 ();
 sg13g2_fill_8 FILLER_195_1007 ();
 sg13g2_fill_4 FILLER_195_1015 ();
 sg13g2_fill_2 FILLER_195_1019 ();
 sg13g2_fill_1 FILLER_195_1021 ();
 sg13g2_fill_2 FILLER_195_1041 ();
 sg13g2_fill_1 FILLER_195_1043 ();
 sg13g2_fill_8 FILLER_195_1052 ();
 sg13g2_fill_4 FILLER_195_1060 ();
 sg13g2_fill_8 FILLER_195_1075 ();
 sg13g2_fill_1 FILLER_195_1083 ();
 sg13g2_fill_8 FILLER_195_1089 ();
 sg13g2_fill_8 FILLER_195_1097 ();
 sg13g2_fill_4 FILLER_195_1105 ();
 sg13g2_fill_2 FILLER_195_1109 ();
 sg13g2_fill_4 FILLER_195_1115 ();
 sg13g2_fill_1 FILLER_195_1119 ();
 sg13g2_fill_8 FILLER_195_1124 ();
 sg13g2_fill_4 FILLER_195_1132 ();
 sg13g2_fill_1 FILLER_195_1136 ();
 sg13g2_fill_4 FILLER_195_1162 ();
 sg13g2_fill_2 FILLER_195_1166 ();
 sg13g2_fill_1 FILLER_195_1168 ();
 sg13g2_fill_4 FILLER_195_1193 ();
 sg13g2_fill_1 FILLER_195_1197 ();
 sg13g2_fill_4 FILLER_195_1214 ();
 sg13g2_fill_2 FILLER_195_1218 ();
 sg13g2_fill_1 FILLER_195_1220 ();
 sg13g2_fill_8 FILLER_195_1229 ();
 sg13g2_fill_8 FILLER_195_1237 ();
 sg13g2_fill_8 FILLER_195_1245 ();
 sg13g2_fill_4 FILLER_195_1253 ();
 sg13g2_fill_2 FILLER_195_1281 ();
 sg13g2_fill_1 FILLER_195_1283 ();
 sg13g2_fill_4 FILLER_195_1300 ();
 sg13g2_fill_2 FILLER_195_1304 ();
 sg13g2_fill_1 FILLER_195_1306 ();
 sg13g2_fill_8 FILLER_195_1315 ();
 sg13g2_fill_8 FILLER_195_1323 ();
 sg13g2_fill_8 FILLER_195_1331 ();
 sg13g2_fill_8 FILLER_195_1339 ();
 sg13g2_fill_2 FILLER_195_1347 ();
 sg13g2_fill_8 FILLER_195_1356 ();
 sg13g2_fill_8 FILLER_195_1364 ();
 sg13g2_fill_8 FILLER_195_1372 ();
 sg13g2_fill_8 FILLER_195_1380 ();
 sg13g2_fill_4 FILLER_195_1388 ();
 sg13g2_fill_1 FILLER_195_1395 ();
 sg13g2_fill_8 FILLER_195_1404 ();
 sg13g2_fill_8 FILLER_195_1412 ();
 sg13g2_fill_8 FILLER_195_1420 ();
 sg13g2_fill_8 FILLER_195_1428 ();
 sg13g2_fill_8 FILLER_195_1436 ();
 sg13g2_fill_8 FILLER_195_1444 ();
 sg13g2_fill_8 FILLER_195_1452 ();
 sg13g2_fill_8 FILLER_195_1460 ();
 sg13g2_fill_8 FILLER_195_1468 ();
 sg13g2_fill_8 FILLER_195_1476 ();
 sg13g2_fill_8 FILLER_195_1484 ();
 sg13g2_fill_8 FILLER_195_1492 ();
 sg13g2_fill_8 FILLER_195_1500 ();
 sg13g2_fill_8 FILLER_195_1508 ();
 sg13g2_fill_8 FILLER_195_1516 ();
 sg13g2_fill_8 FILLER_195_1524 ();
 sg13g2_fill_8 FILLER_195_1532 ();
 sg13g2_fill_8 FILLER_195_1540 ();
 sg13g2_fill_8 FILLER_195_1548 ();
 sg13g2_fill_8 FILLER_195_1556 ();
 sg13g2_fill_8 FILLER_195_1564 ();
 sg13g2_fill_8 FILLER_195_1572 ();
 sg13g2_fill_8 FILLER_195_1580 ();
 sg13g2_fill_4 FILLER_195_1588 ();
 sg13g2_fill_8 FILLER_196_0 ();
 sg13g2_fill_8 FILLER_196_8 ();
 sg13g2_fill_8 FILLER_196_16 ();
 sg13g2_fill_8 FILLER_196_24 ();
 sg13g2_fill_8 FILLER_196_32 ();
 sg13g2_fill_8 FILLER_196_40 ();
 sg13g2_fill_8 FILLER_196_48 ();
 sg13g2_fill_8 FILLER_196_56 ();
 sg13g2_fill_8 FILLER_196_64 ();
 sg13g2_fill_8 FILLER_196_72 ();
 sg13g2_fill_8 FILLER_196_80 ();
 sg13g2_fill_8 FILLER_196_88 ();
 sg13g2_fill_8 FILLER_196_96 ();
 sg13g2_fill_8 FILLER_196_104 ();
 sg13g2_fill_8 FILLER_196_112 ();
 sg13g2_fill_8 FILLER_196_120 ();
 sg13g2_fill_8 FILLER_196_128 ();
 sg13g2_fill_8 FILLER_196_136 ();
 sg13g2_fill_8 FILLER_196_144 ();
 sg13g2_fill_8 FILLER_196_152 ();
 sg13g2_fill_8 FILLER_196_160 ();
 sg13g2_fill_8 FILLER_196_168 ();
 sg13g2_fill_8 FILLER_196_176 ();
 sg13g2_fill_8 FILLER_196_184 ();
 sg13g2_fill_8 FILLER_196_192 ();
 sg13g2_fill_8 FILLER_196_200 ();
 sg13g2_fill_8 FILLER_196_208 ();
 sg13g2_fill_8 FILLER_196_216 ();
 sg13g2_fill_8 FILLER_196_224 ();
 sg13g2_fill_8 FILLER_196_232 ();
 sg13g2_fill_8 FILLER_196_240 ();
 sg13g2_fill_8 FILLER_196_248 ();
 sg13g2_fill_8 FILLER_196_256 ();
 sg13g2_fill_8 FILLER_196_264 ();
 sg13g2_fill_8 FILLER_196_272 ();
 sg13g2_fill_8 FILLER_196_280 ();
 sg13g2_fill_8 FILLER_196_288 ();
 sg13g2_fill_8 FILLER_196_296 ();
 sg13g2_fill_8 FILLER_196_304 ();
 sg13g2_fill_8 FILLER_196_312 ();
 sg13g2_fill_8 FILLER_196_320 ();
 sg13g2_fill_8 FILLER_196_328 ();
 sg13g2_fill_8 FILLER_196_336 ();
 sg13g2_fill_8 FILLER_196_344 ();
 sg13g2_fill_8 FILLER_196_352 ();
 sg13g2_fill_8 FILLER_196_360 ();
 sg13g2_fill_8 FILLER_196_368 ();
 sg13g2_fill_8 FILLER_196_376 ();
 sg13g2_fill_8 FILLER_196_384 ();
 sg13g2_fill_8 FILLER_196_392 ();
 sg13g2_fill_8 FILLER_196_400 ();
 sg13g2_fill_8 FILLER_196_408 ();
 sg13g2_fill_8 FILLER_196_416 ();
 sg13g2_fill_8 FILLER_196_424 ();
 sg13g2_fill_8 FILLER_196_432 ();
 sg13g2_fill_8 FILLER_196_440 ();
 sg13g2_fill_8 FILLER_196_448 ();
 sg13g2_fill_8 FILLER_196_456 ();
 sg13g2_fill_8 FILLER_196_464 ();
 sg13g2_fill_8 FILLER_196_472 ();
 sg13g2_fill_8 FILLER_196_480 ();
 sg13g2_fill_8 FILLER_196_488 ();
 sg13g2_fill_8 FILLER_196_496 ();
 sg13g2_fill_8 FILLER_196_504 ();
 sg13g2_fill_8 FILLER_196_512 ();
 sg13g2_fill_8 FILLER_196_520 ();
 sg13g2_fill_8 FILLER_196_528 ();
 sg13g2_fill_8 FILLER_196_536 ();
 sg13g2_fill_8 FILLER_196_544 ();
 sg13g2_fill_8 FILLER_196_552 ();
 sg13g2_fill_8 FILLER_196_560 ();
 sg13g2_fill_8 FILLER_196_568 ();
 sg13g2_fill_8 FILLER_196_576 ();
 sg13g2_fill_8 FILLER_196_584 ();
 sg13g2_fill_8 FILLER_196_592 ();
 sg13g2_fill_8 FILLER_196_600 ();
 sg13g2_fill_8 FILLER_196_608 ();
 sg13g2_fill_8 FILLER_196_616 ();
 sg13g2_fill_8 FILLER_196_624 ();
 sg13g2_fill_8 FILLER_196_632 ();
 sg13g2_fill_8 FILLER_196_640 ();
 sg13g2_fill_8 FILLER_196_648 ();
 sg13g2_fill_8 FILLER_196_656 ();
 sg13g2_fill_8 FILLER_196_664 ();
 sg13g2_fill_8 FILLER_196_672 ();
 sg13g2_fill_8 FILLER_196_680 ();
 sg13g2_fill_8 FILLER_196_688 ();
 sg13g2_fill_8 FILLER_196_696 ();
 sg13g2_fill_8 FILLER_196_704 ();
 sg13g2_fill_8 FILLER_196_712 ();
 sg13g2_fill_8 FILLER_196_720 ();
 sg13g2_fill_8 FILLER_196_728 ();
 sg13g2_fill_8 FILLER_196_736 ();
 sg13g2_fill_8 FILLER_196_744 ();
 sg13g2_fill_8 FILLER_196_752 ();
 sg13g2_fill_8 FILLER_196_760 ();
 sg13g2_fill_8 FILLER_196_768 ();
 sg13g2_fill_8 FILLER_196_776 ();
 sg13g2_fill_8 FILLER_196_784 ();
 sg13g2_fill_8 FILLER_196_792 ();
 sg13g2_fill_8 FILLER_196_800 ();
 sg13g2_fill_8 FILLER_196_808 ();
 sg13g2_fill_8 FILLER_196_816 ();
 sg13g2_fill_8 FILLER_196_824 ();
 sg13g2_fill_8 FILLER_196_832 ();
 sg13g2_fill_8 FILLER_196_840 ();
 sg13g2_fill_8 FILLER_196_848 ();
 sg13g2_fill_8 FILLER_196_856 ();
 sg13g2_fill_8 FILLER_196_864 ();
 sg13g2_fill_8 FILLER_196_872 ();
 sg13g2_fill_8 FILLER_196_880 ();
 sg13g2_fill_8 FILLER_196_888 ();
 sg13g2_fill_8 FILLER_196_896 ();
 sg13g2_fill_8 FILLER_196_904 ();
 sg13g2_fill_8 FILLER_196_912 ();
 sg13g2_fill_8 FILLER_196_920 ();
 sg13g2_fill_8 FILLER_196_928 ();
 sg13g2_fill_8 FILLER_196_936 ();
 sg13g2_fill_8 FILLER_196_944 ();
 sg13g2_fill_8 FILLER_196_952 ();
 sg13g2_fill_8 FILLER_196_960 ();
 sg13g2_fill_8 FILLER_196_968 ();
 sg13g2_fill_8 FILLER_196_976 ();
 sg13g2_fill_8 FILLER_196_984 ();
 sg13g2_fill_8 FILLER_196_992 ();
 sg13g2_fill_8 FILLER_196_1000 ();
 sg13g2_fill_8 FILLER_196_1008 ();
 sg13g2_fill_8 FILLER_196_1016 ();
 sg13g2_fill_8 FILLER_196_1024 ();
 sg13g2_fill_8 FILLER_196_1032 ();
 sg13g2_fill_8 FILLER_196_1040 ();
 sg13g2_fill_8 FILLER_196_1064 ();
 sg13g2_fill_2 FILLER_196_1072 ();
 sg13g2_fill_1 FILLER_196_1074 ();
 sg13g2_fill_2 FILLER_196_1079 ();
 sg13g2_fill_2 FILLER_196_1085 ();
 sg13g2_fill_1 FILLER_196_1087 ();
 sg13g2_fill_4 FILLER_196_1092 ();
 sg13g2_fill_2 FILLER_196_1096 ();
 sg13g2_fill_1 FILLER_196_1098 ();
 sg13g2_fill_8 FILLER_196_1107 ();
 sg13g2_fill_1 FILLER_196_1115 ();
 sg13g2_fill_8 FILLER_196_1130 ();
 sg13g2_fill_8 FILLER_196_1138 ();
 sg13g2_fill_2 FILLER_196_1146 ();
 sg13g2_fill_8 FILLER_196_1152 ();
 sg13g2_fill_8 FILLER_196_1160 ();
 sg13g2_fill_4 FILLER_196_1168 ();
 sg13g2_fill_1 FILLER_196_1172 ();
 sg13g2_fill_8 FILLER_196_1181 ();
 sg13g2_fill_8 FILLER_196_1189 ();
 sg13g2_fill_4 FILLER_196_1197 ();
 sg13g2_fill_2 FILLER_196_1201 ();
 sg13g2_fill_1 FILLER_196_1203 ();
 sg13g2_fill_2 FILLER_196_1212 ();
 sg13g2_fill_1 FILLER_196_1214 ();
 sg13g2_fill_8 FILLER_196_1219 ();
 sg13g2_fill_2 FILLER_196_1227 ();
 sg13g2_fill_1 FILLER_196_1229 ();
 sg13g2_fill_8 FILLER_196_1233 ();
 sg13g2_fill_8 FILLER_196_1241 ();
 sg13g2_fill_8 FILLER_196_1249 ();
 sg13g2_fill_4 FILLER_196_1257 ();
 sg13g2_fill_4 FILLER_196_1277 ();
 sg13g2_fill_1 FILLER_196_1281 ();
 sg13g2_fill_8 FILLER_196_1293 ();
 sg13g2_fill_4 FILLER_196_1301 ();
 sg13g2_fill_4 FILLER_196_1321 ();
 sg13g2_fill_1 FILLER_196_1325 ();
 sg13g2_fill_8 FILLER_196_1334 ();
 sg13g2_fill_1 FILLER_196_1342 ();
 sg13g2_fill_8 FILLER_196_1351 ();
 sg13g2_fill_2 FILLER_196_1359 ();
 sg13g2_fill_1 FILLER_196_1361 ();
 sg13g2_fill_8 FILLER_196_1386 ();
 sg13g2_fill_8 FILLER_196_1394 ();
 sg13g2_fill_2 FILLER_196_1402 ();
 sg13g2_fill_2 FILLER_196_1408 ();
 sg13g2_fill_8 FILLER_196_1423 ();
 sg13g2_fill_8 FILLER_196_1431 ();
 sg13g2_fill_8 FILLER_196_1439 ();
 sg13g2_fill_8 FILLER_196_1447 ();
 sg13g2_fill_8 FILLER_196_1455 ();
 sg13g2_fill_8 FILLER_196_1463 ();
 sg13g2_fill_8 FILLER_196_1471 ();
 sg13g2_fill_8 FILLER_196_1479 ();
 sg13g2_fill_8 FILLER_196_1487 ();
 sg13g2_fill_8 FILLER_196_1495 ();
 sg13g2_fill_8 FILLER_196_1503 ();
 sg13g2_fill_8 FILLER_196_1511 ();
 sg13g2_fill_8 FILLER_196_1519 ();
 sg13g2_fill_8 FILLER_196_1527 ();
 sg13g2_fill_8 FILLER_196_1535 ();
 sg13g2_fill_8 FILLER_196_1543 ();
 sg13g2_fill_8 FILLER_196_1551 ();
 sg13g2_fill_8 FILLER_196_1559 ();
 sg13g2_fill_8 FILLER_196_1567 ();
 sg13g2_fill_8 FILLER_196_1575 ();
 sg13g2_fill_8 FILLER_196_1583 ();
 sg13g2_fill_1 FILLER_196_1591 ();
 sg13g2_fill_8 FILLER_197_0 ();
 sg13g2_fill_8 FILLER_197_8 ();
 sg13g2_fill_8 FILLER_197_16 ();
 sg13g2_fill_8 FILLER_197_24 ();
 sg13g2_fill_8 FILLER_197_32 ();
 sg13g2_fill_8 FILLER_197_40 ();
 sg13g2_fill_8 FILLER_197_48 ();
 sg13g2_fill_8 FILLER_197_56 ();
 sg13g2_fill_8 FILLER_197_64 ();
 sg13g2_fill_8 FILLER_197_72 ();
 sg13g2_fill_8 FILLER_197_80 ();
 sg13g2_fill_8 FILLER_197_88 ();
 sg13g2_fill_8 FILLER_197_96 ();
 sg13g2_fill_8 FILLER_197_104 ();
 sg13g2_fill_8 FILLER_197_112 ();
 sg13g2_fill_8 FILLER_197_120 ();
 sg13g2_fill_8 FILLER_197_128 ();
 sg13g2_fill_8 FILLER_197_136 ();
 sg13g2_fill_8 FILLER_197_144 ();
 sg13g2_fill_8 FILLER_197_152 ();
 sg13g2_fill_8 FILLER_197_160 ();
 sg13g2_fill_8 FILLER_197_168 ();
 sg13g2_fill_8 FILLER_197_176 ();
 sg13g2_fill_8 FILLER_197_184 ();
 sg13g2_fill_8 FILLER_197_192 ();
 sg13g2_fill_8 FILLER_197_200 ();
 sg13g2_fill_8 FILLER_197_208 ();
 sg13g2_fill_8 FILLER_197_216 ();
 sg13g2_fill_8 FILLER_197_224 ();
 sg13g2_fill_8 FILLER_197_232 ();
 sg13g2_fill_8 FILLER_197_240 ();
 sg13g2_fill_8 FILLER_197_248 ();
 sg13g2_fill_8 FILLER_197_256 ();
 sg13g2_fill_8 FILLER_197_264 ();
 sg13g2_fill_8 FILLER_197_272 ();
 sg13g2_fill_8 FILLER_197_280 ();
 sg13g2_fill_8 FILLER_197_288 ();
 sg13g2_fill_8 FILLER_197_296 ();
 sg13g2_fill_8 FILLER_197_304 ();
 sg13g2_fill_8 FILLER_197_312 ();
 sg13g2_fill_8 FILLER_197_320 ();
 sg13g2_fill_8 FILLER_197_328 ();
 sg13g2_fill_8 FILLER_197_336 ();
 sg13g2_fill_8 FILLER_197_344 ();
 sg13g2_fill_8 FILLER_197_352 ();
 sg13g2_fill_8 FILLER_197_360 ();
 sg13g2_fill_8 FILLER_197_368 ();
 sg13g2_fill_8 FILLER_197_376 ();
 sg13g2_fill_8 FILLER_197_384 ();
 sg13g2_fill_8 FILLER_197_392 ();
 sg13g2_fill_8 FILLER_197_400 ();
 sg13g2_fill_8 FILLER_197_408 ();
 sg13g2_fill_8 FILLER_197_416 ();
 sg13g2_fill_8 FILLER_197_424 ();
 sg13g2_fill_8 FILLER_197_432 ();
 sg13g2_fill_8 FILLER_197_440 ();
 sg13g2_fill_8 FILLER_197_448 ();
 sg13g2_fill_8 FILLER_197_456 ();
 sg13g2_fill_8 FILLER_197_464 ();
 sg13g2_fill_8 FILLER_197_472 ();
 sg13g2_fill_8 FILLER_197_480 ();
 sg13g2_fill_8 FILLER_197_488 ();
 sg13g2_fill_8 FILLER_197_496 ();
 sg13g2_fill_8 FILLER_197_504 ();
 sg13g2_fill_8 FILLER_197_512 ();
 sg13g2_fill_8 FILLER_197_520 ();
 sg13g2_fill_8 FILLER_197_528 ();
 sg13g2_fill_8 FILLER_197_536 ();
 sg13g2_fill_8 FILLER_197_544 ();
 sg13g2_fill_8 FILLER_197_552 ();
 sg13g2_fill_8 FILLER_197_560 ();
 sg13g2_fill_8 FILLER_197_568 ();
 sg13g2_fill_8 FILLER_197_576 ();
 sg13g2_fill_8 FILLER_197_584 ();
 sg13g2_fill_8 FILLER_197_592 ();
 sg13g2_fill_8 FILLER_197_600 ();
 sg13g2_fill_8 FILLER_197_608 ();
 sg13g2_fill_8 FILLER_197_616 ();
 sg13g2_fill_8 FILLER_197_624 ();
 sg13g2_fill_8 FILLER_197_632 ();
 sg13g2_fill_8 FILLER_197_640 ();
 sg13g2_fill_8 FILLER_197_648 ();
 sg13g2_fill_8 FILLER_197_656 ();
 sg13g2_fill_8 FILLER_197_664 ();
 sg13g2_fill_8 FILLER_197_672 ();
 sg13g2_fill_8 FILLER_197_680 ();
 sg13g2_fill_8 FILLER_197_688 ();
 sg13g2_fill_8 FILLER_197_696 ();
 sg13g2_fill_8 FILLER_197_704 ();
 sg13g2_fill_8 FILLER_197_712 ();
 sg13g2_fill_8 FILLER_197_720 ();
 sg13g2_fill_8 FILLER_197_728 ();
 sg13g2_fill_8 FILLER_197_736 ();
 sg13g2_fill_8 FILLER_197_744 ();
 sg13g2_fill_8 FILLER_197_752 ();
 sg13g2_fill_8 FILLER_197_760 ();
 sg13g2_fill_8 FILLER_197_768 ();
 sg13g2_fill_8 FILLER_197_776 ();
 sg13g2_fill_8 FILLER_197_784 ();
 sg13g2_fill_8 FILLER_197_792 ();
 sg13g2_fill_8 FILLER_197_800 ();
 sg13g2_fill_8 FILLER_197_808 ();
 sg13g2_fill_8 FILLER_197_816 ();
 sg13g2_fill_8 FILLER_197_824 ();
 sg13g2_fill_8 FILLER_197_832 ();
 sg13g2_fill_8 FILLER_197_840 ();
 sg13g2_fill_8 FILLER_197_848 ();
 sg13g2_fill_8 FILLER_197_856 ();
 sg13g2_fill_8 FILLER_197_864 ();
 sg13g2_fill_8 FILLER_197_872 ();
 sg13g2_fill_8 FILLER_197_880 ();
 sg13g2_fill_8 FILLER_197_888 ();
 sg13g2_fill_8 FILLER_197_896 ();
 sg13g2_fill_8 FILLER_197_904 ();
 sg13g2_fill_8 FILLER_197_912 ();
 sg13g2_fill_8 FILLER_197_920 ();
 sg13g2_fill_8 FILLER_197_928 ();
 sg13g2_fill_8 FILLER_197_936 ();
 sg13g2_fill_8 FILLER_197_944 ();
 sg13g2_fill_8 FILLER_197_952 ();
 sg13g2_fill_8 FILLER_197_960 ();
 sg13g2_fill_8 FILLER_197_968 ();
 sg13g2_fill_8 FILLER_197_976 ();
 sg13g2_fill_8 FILLER_197_984 ();
 sg13g2_fill_8 FILLER_197_992 ();
 sg13g2_fill_8 FILLER_197_1000 ();
 sg13g2_fill_8 FILLER_197_1008 ();
 sg13g2_fill_8 FILLER_197_1016 ();
 sg13g2_fill_8 FILLER_197_1024 ();
 sg13g2_fill_8 FILLER_197_1032 ();
 sg13g2_fill_8 FILLER_197_1040 ();
 sg13g2_fill_2 FILLER_197_1048 ();
 sg13g2_fill_1 FILLER_197_1050 ();
 sg13g2_fill_1 FILLER_197_1063 ();
 sg13g2_fill_2 FILLER_197_1086 ();
 sg13g2_fill_4 FILLER_197_1109 ();
 sg13g2_fill_4 FILLER_197_1123 ();
 sg13g2_fill_2 FILLER_197_1139 ();
 sg13g2_fill_8 FILLER_197_1165 ();
 sg13g2_fill_2 FILLER_197_1173 ();
 sg13g2_fill_8 FILLER_197_1196 ();
 sg13g2_fill_4 FILLER_197_1204 ();
 sg13g2_fill_1 FILLER_197_1208 ();
 sg13g2_fill_1 FILLER_197_1230 ();
 sg13g2_fill_1 FILLER_197_1247 ();
 sg13g2_fill_8 FILLER_197_1256 ();
 sg13g2_fill_2 FILLER_197_1264 ();
 sg13g2_fill_2 FILLER_197_1271 ();
 sg13g2_fill_8 FILLER_197_1278 ();
 sg13g2_fill_1 FILLER_197_1286 ();
 sg13g2_fill_8 FILLER_197_1295 ();
 sg13g2_fill_1 FILLER_197_1303 ();
 sg13g2_fill_2 FILLER_197_1320 ();
 sg13g2_fill_2 FILLER_197_1349 ();
 sg13g2_fill_1 FILLER_197_1351 ();
 sg13g2_fill_4 FILLER_197_1357 ();
 sg13g2_fill_2 FILLER_197_1361 ();
 sg13g2_fill_8 FILLER_197_1376 ();
 sg13g2_fill_4 FILLER_197_1384 ();
 sg13g2_fill_2 FILLER_197_1388 ();
 sg13g2_fill_8 FILLER_197_1427 ();
 sg13g2_fill_8 FILLER_197_1435 ();
 sg13g2_fill_8 FILLER_197_1443 ();
 sg13g2_fill_8 FILLER_197_1451 ();
 sg13g2_fill_8 FILLER_197_1459 ();
 sg13g2_fill_8 FILLER_197_1467 ();
 sg13g2_fill_8 FILLER_197_1475 ();
 sg13g2_fill_8 FILLER_197_1483 ();
 sg13g2_fill_8 FILLER_197_1491 ();
 sg13g2_fill_8 FILLER_197_1499 ();
 sg13g2_fill_8 FILLER_197_1507 ();
 sg13g2_fill_8 FILLER_197_1515 ();
 sg13g2_fill_8 FILLER_197_1523 ();
 sg13g2_fill_8 FILLER_197_1531 ();
 sg13g2_fill_8 FILLER_197_1539 ();
 sg13g2_fill_8 FILLER_197_1547 ();
 sg13g2_fill_8 FILLER_197_1555 ();
 sg13g2_fill_8 FILLER_197_1563 ();
 sg13g2_fill_8 FILLER_197_1571 ();
 sg13g2_fill_8 FILLER_197_1579 ();
 sg13g2_fill_4 FILLER_197_1587 ();
 sg13g2_fill_1 FILLER_197_1591 ();
 sg13g2_fill_8 FILLER_198_0 ();
 sg13g2_fill_8 FILLER_198_8 ();
 sg13g2_fill_8 FILLER_198_16 ();
 sg13g2_fill_8 FILLER_198_24 ();
 sg13g2_fill_8 FILLER_198_32 ();
 sg13g2_fill_8 FILLER_198_40 ();
 sg13g2_fill_8 FILLER_198_48 ();
 sg13g2_fill_8 FILLER_198_56 ();
 sg13g2_fill_8 FILLER_198_64 ();
 sg13g2_fill_8 FILLER_198_72 ();
 sg13g2_fill_8 FILLER_198_80 ();
 sg13g2_fill_8 FILLER_198_88 ();
 sg13g2_fill_8 FILLER_198_96 ();
 sg13g2_fill_8 FILLER_198_104 ();
 sg13g2_fill_8 FILLER_198_112 ();
 sg13g2_fill_8 FILLER_198_120 ();
 sg13g2_fill_8 FILLER_198_128 ();
 sg13g2_fill_8 FILLER_198_136 ();
 sg13g2_fill_8 FILLER_198_144 ();
 sg13g2_fill_8 FILLER_198_152 ();
 sg13g2_fill_8 FILLER_198_160 ();
 sg13g2_fill_8 FILLER_198_168 ();
 sg13g2_fill_8 FILLER_198_176 ();
 sg13g2_fill_8 FILLER_198_184 ();
 sg13g2_fill_8 FILLER_198_192 ();
 sg13g2_fill_8 FILLER_198_200 ();
 sg13g2_fill_8 FILLER_198_208 ();
 sg13g2_fill_8 FILLER_198_216 ();
 sg13g2_fill_8 FILLER_198_224 ();
 sg13g2_fill_8 FILLER_198_232 ();
 sg13g2_fill_8 FILLER_198_240 ();
 sg13g2_fill_8 FILLER_198_248 ();
 sg13g2_fill_8 FILLER_198_256 ();
 sg13g2_fill_8 FILLER_198_264 ();
 sg13g2_fill_8 FILLER_198_272 ();
 sg13g2_fill_8 FILLER_198_280 ();
 sg13g2_fill_8 FILLER_198_288 ();
 sg13g2_fill_8 FILLER_198_296 ();
 sg13g2_fill_8 FILLER_198_304 ();
 sg13g2_fill_8 FILLER_198_312 ();
 sg13g2_fill_8 FILLER_198_320 ();
 sg13g2_fill_8 FILLER_198_328 ();
 sg13g2_fill_8 FILLER_198_336 ();
 sg13g2_fill_8 FILLER_198_344 ();
 sg13g2_fill_8 FILLER_198_352 ();
 sg13g2_fill_8 FILLER_198_360 ();
 sg13g2_fill_8 FILLER_198_368 ();
 sg13g2_fill_8 FILLER_198_376 ();
 sg13g2_fill_8 FILLER_198_384 ();
 sg13g2_fill_8 FILLER_198_392 ();
 sg13g2_fill_8 FILLER_198_400 ();
 sg13g2_fill_8 FILLER_198_408 ();
 sg13g2_fill_8 FILLER_198_416 ();
 sg13g2_fill_8 FILLER_198_424 ();
 sg13g2_fill_8 FILLER_198_432 ();
 sg13g2_fill_8 FILLER_198_440 ();
 sg13g2_fill_8 FILLER_198_448 ();
 sg13g2_fill_8 FILLER_198_456 ();
 sg13g2_fill_8 FILLER_198_464 ();
 sg13g2_fill_8 FILLER_198_472 ();
 sg13g2_fill_8 FILLER_198_480 ();
 sg13g2_fill_8 FILLER_198_488 ();
 sg13g2_fill_8 FILLER_198_496 ();
 sg13g2_fill_8 FILLER_198_504 ();
 sg13g2_fill_8 FILLER_198_512 ();
 sg13g2_fill_8 FILLER_198_520 ();
 sg13g2_fill_8 FILLER_198_528 ();
 sg13g2_fill_8 FILLER_198_536 ();
 sg13g2_fill_8 FILLER_198_544 ();
 sg13g2_fill_8 FILLER_198_552 ();
 sg13g2_fill_8 FILLER_198_560 ();
 sg13g2_fill_8 FILLER_198_568 ();
 sg13g2_fill_8 FILLER_198_576 ();
 sg13g2_fill_8 FILLER_198_584 ();
 sg13g2_fill_8 FILLER_198_592 ();
 sg13g2_fill_8 FILLER_198_600 ();
 sg13g2_fill_8 FILLER_198_608 ();
 sg13g2_fill_8 FILLER_198_616 ();
 sg13g2_fill_8 FILLER_198_624 ();
 sg13g2_fill_8 FILLER_198_632 ();
 sg13g2_fill_8 FILLER_198_640 ();
 sg13g2_fill_8 FILLER_198_648 ();
 sg13g2_fill_8 FILLER_198_656 ();
 sg13g2_fill_8 FILLER_198_664 ();
 sg13g2_fill_8 FILLER_198_672 ();
 sg13g2_fill_8 FILLER_198_680 ();
 sg13g2_fill_8 FILLER_198_688 ();
 sg13g2_fill_8 FILLER_198_696 ();
 sg13g2_fill_8 FILLER_198_704 ();
 sg13g2_fill_8 FILLER_198_712 ();
 sg13g2_fill_8 FILLER_198_720 ();
 sg13g2_fill_8 FILLER_198_728 ();
 sg13g2_fill_8 FILLER_198_736 ();
 sg13g2_fill_8 FILLER_198_744 ();
 sg13g2_fill_8 FILLER_198_752 ();
 sg13g2_fill_8 FILLER_198_760 ();
 sg13g2_fill_8 FILLER_198_768 ();
 sg13g2_fill_8 FILLER_198_776 ();
 sg13g2_fill_8 FILLER_198_784 ();
 sg13g2_fill_8 FILLER_198_792 ();
 sg13g2_fill_8 FILLER_198_800 ();
 sg13g2_fill_8 FILLER_198_808 ();
 sg13g2_fill_8 FILLER_198_816 ();
 sg13g2_fill_8 FILLER_198_824 ();
 sg13g2_fill_8 FILLER_198_832 ();
 sg13g2_fill_8 FILLER_198_840 ();
 sg13g2_fill_8 FILLER_198_848 ();
 sg13g2_fill_8 FILLER_198_856 ();
 sg13g2_fill_8 FILLER_198_864 ();
 sg13g2_fill_8 FILLER_198_872 ();
 sg13g2_fill_8 FILLER_198_880 ();
 sg13g2_fill_8 FILLER_198_888 ();
 sg13g2_fill_8 FILLER_198_896 ();
 sg13g2_fill_8 FILLER_198_904 ();
 sg13g2_fill_8 FILLER_198_912 ();
 sg13g2_fill_8 FILLER_198_920 ();
 sg13g2_fill_8 FILLER_198_928 ();
 sg13g2_fill_8 FILLER_198_936 ();
 sg13g2_fill_8 FILLER_198_944 ();
 sg13g2_fill_8 FILLER_198_952 ();
 sg13g2_fill_8 FILLER_198_960 ();
 sg13g2_fill_8 FILLER_198_968 ();
 sg13g2_fill_8 FILLER_198_976 ();
 sg13g2_fill_8 FILLER_198_984 ();
 sg13g2_fill_8 FILLER_198_992 ();
 sg13g2_fill_8 FILLER_198_1000 ();
 sg13g2_fill_8 FILLER_198_1008 ();
 sg13g2_fill_8 FILLER_198_1016 ();
 sg13g2_fill_8 FILLER_198_1024 ();
 sg13g2_fill_8 FILLER_198_1032 ();
 sg13g2_fill_8 FILLER_198_1040 ();
 sg13g2_fill_4 FILLER_198_1048 ();
 sg13g2_fill_2 FILLER_198_1052 ();
 sg13g2_fill_1 FILLER_198_1054 ();
 sg13g2_fill_8 FILLER_198_1059 ();
 sg13g2_fill_1 FILLER_198_1071 ();
 sg13g2_fill_8 FILLER_198_1086 ();
 sg13g2_fill_4 FILLER_198_1094 ();
 sg13g2_fill_8 FILLER_198_1106 ();
 sg13g2_fill_4 FILLER_198_1114 ();
 sg13g2_fill_1 FILLER_198_1118 ();
 sg13g2_fill_8 FILLER_198_1135 ();
 sg13g2_fill_8 FILLER_198_1143 ();
 sg13g2_fill_8 FILLER_198_1151 ();
 sg13g2_fill_8 FILLER_198_1159 ();
 sg13g2_fill_4 FILLER_198_1167 ();
 sg13g2_fill_2 FILLER_198_1187 ();
 sg13g2_fill_8 FILLER_198_1218 ();
 sg13g2_fill_8 FILLER_198_1226 ();
 sg13g2_fill_1 FILLER_198_1234 ();
 sg13g2_fill_8 FILLER_198_1259 ();
 sg13g2_fill_2 FILLER_198_1281 ();
 sg13g2_fill_4 FILLER_198_1299 ();
 sg13g2_fill_2 FILLER_198_1303 ();
 sg13g2_fill_1 FILLER_198_1305 ();
 sg13g2_fill_8 FILLER_198_1314 ();
 sg13g2_fill_2 FILLER_198_1322 ();
 sg13g2_fill_1 FILLER_198_1324 ();
 sg13g2_fill_2 FILLER_198_1353 ();
 sg13g2_fill_2 FILLER_198_1362 ();
 sg13g2_fill_4 FILLER_198_1386 ();
 sg13g2_fill_4 FILLER_198_1405 ();
 sg13g2_fill_1 FILLER_198_1409 ();
 sg13g2_fill_8 FILLER_198_1420 ();
 sg13g2_fill_8 FILLER_198_1428 ();
 sg13g2_fill_8 FILLER_198_1436 ();
 sg13g2_fill_8 FILLER_198_1444 ();
 sg13g2_fill_8 FILLER_198_1452 ();
 sg13g2_fill_8 FILLER_198_1460 ();
 sg13g2_fill_8 FILLER_198_1468 ();
 sg13g2_fill_8 FILLER_198_1476 ();
 sg13g2_fill_8 FILLER_198_1484 ();
 sg13g2_fill_8 FILLER_198_1492 ();
 sg13g2_fill_8 FILLER_198_1500 ();
 sg13g2_fill_8 FILLER_198_1508 ();
 sg13g2_fill_8 FILLER_198_1516 ();
 sg13g2_fill_8 FILLER_198_1524 ();
 sg13g2_fill_8 FILLER_198_1532 ();
 sg13g2_fill_8 FILLER_198_1540 ();
 sg13g2_fill_8 FILLER_198_1548 ();
 sg13g2_fill_8 FILLER_198_1556 ();
 sg13g2_fill_8 FILLER_198_1564 ();
 sg13g2_fill_8 FILLER_198_1572 ();
 sg13g2_fill_8 FILLER_198_1580 ();
 sg13g2_fill_4 FILLER_198_1588 ();
 sg13g2_fill_8 FILLER_199_0 ();
 sg13g2_fill_8 FILLER_199_8 ();
 sg13g2_fill_8 FILLER_199_16 ();
 sg13g2_fill_8 FILLER_199_24 ();
 sg13g2_fill_8 FILLER_199_32 ();
 sg13g2_fill_8 FILLER_199_40 ();
 sg13g2_fill_8 FILLER_199_48 ();
 sg13g2_fill_8 FILLER_199_56 ();
 sg13g2_fill_8 FILLER_199_64 ();
 sg13g2_fill_8 FILLER_199_72 ();
 sg13g2_fill_8 FILLER_199_80 ();
 sg13g2_fill_8 FILLER_199_88 ();
 sg13g2_fill_8 FILLER_199_96 ();
 sg13g2_fill_8 FILLER_199_104 ();
 sg13g2_fill_8 FILLER_199_112 ();
 sg13g2_fill_8 FILLER_199_120 ();
 sg13g2_fill_8 FILLER_199_128 ();
 sg13g2_fill_8 FILLER_199_136 ();
 sg13g2_fill_8 FILLER_199_144 ();
 sg13g2_fill_8 FILLER_199_152 ();
 sg13g2_fill_8 FILLER_199_160 ();
 sg13g2_fill_8 FILLER_199_168 ();
 sg13g2_fill_8 FILLER_199_176 ();
 sg13g2_fill_8 FILLER_199_184 ();
 sg13g2_fill_8 FILLER_199_192 ();
 sg13g2_fill_8 FILLER_199_200 ();
 sg13g2_fill_8 FILLER_199_208 ();
 sg13g2_fill_8 FILLER_199_216 ();
 sg13g2_fill_8 FILLER_199_224 ();
 sg13g2_fill_8 FILLER_199_232 ();
 sg13g2_fill_8 FILLER_199_240 ();
 sg13g2_fill_8 FILLER_199_248 ();
 sg13g2_fill_8 FILLER_199_256 ();
 sg13g2_fill_8 FILLER_199_264 ();
 sg13g2_fill_8 FILLER_199_272 ();
 sg13g2_fill_8 FILLER_199_280 ();
 sg13g2_fill_8 FILLER_199_288 ();
 sg13g2_fill_8 FILLER_199_296 ();
 sg13g2_fill_8 FILLER_199_304 ();
 sg13g2_fill_8 FILLER_199_312 ();
 sg13g2_fill_8 FILLER_199_320 ();
 sg13g2_fill_8 FILLER_199_328 ();
 sg13g2_fill_8 FILLER_199_336 ();
 sg13g2_fill_8 FILLER_199_344 ();
 sg13g2_fill_8 FILLER_199_352 ();
 sg13g2_fill_8 FILLER_199_360 ();
 sg13g2_fill_8 FILLER_199_368 ();
 sg13g2_fill_8 FILLER_199_376 ();
 sg13g2_fill_8 FILLER_199_384 ();
 sg13g2_fill_8 FILLER_199_392 ();
 sg13g2_fill_8 FILLER_199_400 ();
 sg13g2_fill_8 FILLER_199_408 ();
 sg13g2_fill_8 FILLER_199_416 ();
 sg13g2_fill_8 FILLER_199_424 ();
 sg13g2_fill_8 FILLER_199_432 ();
 sg13g2_fill_8 FILLER_199_440 ();
 sg13g2_fill_8 FILLER_199_448 ();
 sg13g2_fill_8 FILLER_199_456 ();
 sg13g2_fill_8 FILLER_199_464 ();
 sg13g2_fill_8 FILLER_199_472 ();
 sg13g2_fill_8 FILLER_199_480 ();
 sg13g2_fill_8 FILLER_199_488 ();
 sg13g2_fill_8 FILLER_199_496 ();
 sg13g2_fill_8 FILLER_199_504 ();
 sg13g2_fill_8 FILLER_199_512 ();
 sg13g2_fill_8 FILLER_199_520 ();
 sg13g2_fill_8 FILLER_199_528 ();
 sg13g2_fill_8 FILLER_199_536 ();
 sg13g2_fill_8 FILLER_199_544 ();
 sg13g2_fill_8 FILLER_199_552 ();
 sg13g2_fill_8 FILLER_199_560 ();
 sg13g2_fill_8 FILLER_199_568 ();
 sg13g2_fill_8 FILLER_199_576 ();
 sg13g2_fill_8 FILLER_199_584 ();
 sg13g2_fill_8 FILLER_199_592 ();
 sg13g2_fill_8 FILLER_199_600 ();
 sg13g2_fill_8 FILLER_199_608 ();
 sg13g2_fill_8 FILLER_199_616 ();
 sg13g2_fill_8 FILLER_199_624 ();
 sg13g2_fill_8 FILLER_199_632 ();
 sg13g2_fill_8 FILLER_199_640 ();
 sg13g2_fill_8 FILLER_199_648 ();
 sg13g2_fill_8 FILLER_199_656 ();
 sg13g2_fill_8 FILLER_199_664 ();
 sg13g2_fill_8 FILLER_199_672 ();
 sg13g2_fill_8 FILLER_199_680 ();
 sg13g2_fill_8 FILLER_199_688 ();
 sg13g2_fill_8 FILLER_199_696 ();
 sg13g2_fill_8 FILLER_199_704 ();
 sg13g2_fill_8 FILLER_199_712 ();
 sg13g2_fill_8 FILLER_199_720 ();
 sg13g2_fill_8 FILLER_199_728 ();
 sg13g2_fill_8 FILLER_199_736 ();
 sg13g2_fill_8 FILLER_199_744 ();
 sg13g2_fill_8 FILLER_199_752 ();
 sg13g2_fill_8 FILLER_199_760 ();
 sg13g2_fill_8 FILLER_199_768 ();
 sg13g2_fill_8 FILLER_199_776 ();
 sg13g2_fill_8 FILLER_199_784 ();
 sg13g2_fill_8 FILLER_199_792 ();
 sg13g2_fill_8 FILLER_199_800 ();
 sg13g2_fill_8 FILLER_199_808 ();
 sg13g2_fill_8 FILLER_199_816 ();
 sg13g2_fill_8 FILLER_199_824 ();
 sg13g2_fill_8 FILLER_199_832 ();
 sg13g2_fill_8 FILLER_199_840 ();
 sg13g2_fill_8 FILLER_199_848 ();
 sg13g2_fill_8 FILLER_199_856 ();
 sg13g2_fill_8 FILLER_199_864 ();
 sg13g2_fill_8 FILLER_199_872 ();
 sg13g2_fill_8 FILLER_199_880 ();
 sg13g2_fill_8 FILLER_199_888 ();
 sg13g2_fill_8 FILLER_199_896 ();
 sg13g2_fill_8 FILLER_199_904 ();
 sg13g2_fill_8 FILLER_199_912 ();
 sg13g2_fill_8 FILLER_199_920 ();
 sg13g2_fill_8 FILLER_199_928 ();
 sg13g2_fill_8 FILLER_199_936 ();
 sg13g2_fill_8 FILLER_199_944 ();
 sg13g2_fill_8 FILLER_199_952 ();
 sg13g2_fill_8 FILLER_199_960 ();
 sg13g2_fill_8 FILLER_199_968 ();
 sg13g2_fill_8 FILLER_199_976 ();
 sg13g2_fill_8 FILLER_199_984 ();
 sg13g2_fill_8 FILLER_199_992 ();
 sg13g2_fill_8 FILLER_199_1000 ();
 sg13g2_fill_8 FILLER_199_1008 ();
 sg13g2_fill_8 FILLER_199_1016 ();
 sg13g2_fill_8 FILLER_199_1024 ();
 sg13g2_fill_8 FILLER_199_1032 ();
 sg13g2_fill_8 FILLER_199_1040 ();
 sg13g2_fill_8 FILLER_199_1048 ();
 sg13g2_fill_8 FILLER_199_1056 ();
 sg13g2_fill_4 FILLER_199_1064 ();
 sg13g2_fill_1 FILLER_199_1068 ();
 sg13g2_fill_8 FILLER_199_1077 ();
 sg13g2_fill_8 FILLER_199_1085 ();
 sg13g2_fill_8 FILLER_199_1093 ();
 sg13g2_fill_8 FILLER_199_1101 ();
 sg13g2_fill_8 FILLER_199_1109 ();
 sg13g2_fill_4 FILLER_199_1117 ();
 sg13g2_fill_2 FILLER_199_1121 ();
 sg13g2_fill_1 FILLER_199_1123 ();
 sg13g2_fill_2 FILLER_199_1137 ();
 sg13g2_fill_1 FILLER_199_1139 ();
 sg13g2_fill_8 FILLER_199_1148 ();
 sg13g2_fill_1 FILLER_199_1156 ();
 sg13g2_fill_8 FILLER_199_1182 ();
 sg13g2_fill_8 FILLER_199_1190 ();
 sg13g2_fill_8 FILLER_199_1198 ();
 sg13g2_fill_2 FILLER_199_1206 ();
 sg13g2_fill_1 FILLER_199_1208 ();
 sg13g2_fill_8 FILLER_199_1218 ();
 sg13g2_fill_4 FILLER_199_1226 ();
 sg13g2_fill_2 FILLER_199_1230 ();
 sg13g2_fill_2 FILLER_199_1236 ();
 sg13g2_fill_8 FILLER_199_1250 ();
 sg13g2_fill_2 FILLER_199_1274 ();
 sg13g2_fill_4 FILLER_199_1284 ();
 sg13g2_fill_2 FILLER_199_1288 ();
 sg13g2_fill_8 FILLER_199_1298 ();
 sg13g2_fill_4 FILLER_199_1306 ();
 sg13g2_fill_8 FILLER_199_1327 ();
 sg13g2_fill_4 FILLER_199_1335 ();
 sg13g2_fill_4 FILLER_199_1344 ();
 sg13g2_fill_1 FILLER_199_1348 ();
 sg13g2_fill_8 FILLER_199_1377 ();
 sg13g2_fill_8 FILLER_199_1385 ();
 sg13g2_fill_8 FILLER_199_1393 ();
 sg13g2_fill_8 FILLER_199_1401 ();
 sg13g2_fill_8 FILLER_199_1409 ();
 sg13g2_fill_8 FILLER_199_1417 ();
 sg13g2_fill_8 FILLER_199_1425 ();
 sg13g2_fill_8 FILLER_199_1433 ();
 sg13g2_fill_8 FILLER_199_1441 ();
 sg13g2_fill_8 FILLER_199_1449 ();
 sg13g2_fill_8 FILLER_199_1457 ();
 sg13g2_fill_8 FILLER_199_1465 ();
 sg13g2_fill_8 FILLER_199_1473 ();
 sg13g2_fill_8 FILLER_199_1481 ();
 sg13g2_fill_8 FILLER_199_1489 ();
 sg13g2_fill_8 FILLER_199_1497 ();
 sg13g2_fill_8 FILLER_199_1505 ();
 sg13g2_fill_8 FILLER_199_1513 ();
 sg13g2_fill_8 FILLER_199_1521 ();
 sg13g2_fill_8 FILLER_199_1529 ();
 sg13g2_fill_8 FILLER_199_1537 ();
 sg13g2_fill_8 FILLER_199_1545 ();
 sg13g2_fill_8 FILLER_199_1553 ();
 sg13g2_fill_8 FILLER_199_1561 ();
 sg13g2_fill_8 FILLER_199_1569 ();
 sg13g2_fill_8 FILLER_199_1577 ();
 sg13g2_fill_4 FILLER_199_1585 ();
 sg13g2_fill_2 FILLER_199_1589 ();
 sg13g2_fill_1 FILLER_199_1591 ();
 sg13g2_fill_8 FILLER_200_0 ();
 sg13g2_fill_8 FILLER_200_8 ();
 sg13g2_fill_8 FILLER_200_16 ();
 sg13g2_fill_8 FILLER_200_24 ();
 sg13g2_fill_8 FILLER_200_32 ();
 sg13g2_fill_8 FILLER_200_40 ();
 sg13g2_fill_8 FILLER_200_48 ();
 sg13g2_fill_8 FILLER_200_56 ();
 sg13g2_fill_8 FILLER_200_64 ();
 sg13g2_fill_8 FILLER_200_72 ();
 sg13g2_fill_8 FILLER_200_80 ();
 sg13g2_fill_8 FILLER_200_88 ();
 sg13g2_fill_8 FILLER_200_96 ();
 sg13g2_fill_8 FILLER_200_104 ();
 sg13g2_fill_8 FILLER_200_112 ();
 sg13g2_fill_8 FILLER_200_120 ();
 sg13g2_fill_8 FILLER_200_128 ();
 sg13g2_fill_8 FILLER_200_136 ();
 sg13g2_fill_8 FILLER_200_144 ();
 sg13g2_fill_8 FILLER_200_152 ();
 sg13g2_fill_8 FILLER_200_160 ();
 sg13g2_fill_8 FILLER_200_168 ();
 sg13g2_fill_8 FILLER_200_176 ();
 sg13g2_fill_8 FILLER_200_184 ();
 sg13g2_fill_8 FILLER_200_192 ();
 sg13g2_fill_8 FILLER_200_200 ();
 sg13g2_fill_8 FILLER_200_208 ();
 sg13g2_fill_8 FILLER_200_216 ();
 sg13g2_fill_8 FILLER_200_224 ();
 sg13g2_fill_8 FILLER_200_232 ();
 sg13g2_fill_8 FILLER_200_240 ();
 sg13g2_fill_8 FILLER_200_248 ();
 sg13g2_fill_8 FILLER_200_256 ();
 sg13g2_fill_8 FILLER_200_264 ();
 sg13g2_fill_8 FILLER_200_272 ();
 sg13g2_fill_8 FILLER_200_280 ();
 sg13g2_fill_8 FILLER_200_288 ();
 sg13g2_fill_8 FILLER_200_296 ();
 sg13g2_fill_8 FILLER_200_304 ();
 sg13g2_fill_8 FILLER_200_312 ();
 sg13g2_fill_8 FILLER_200_320 ();
 sg13g2_fill_8 FILLER_200_328 ();
 sg13g2_fill_8 FILLER_200_336 ();
 sg13g2_fill_8 FILLER_200_344 ();
 sg13g2_fill_8 FILLER_200_352 ();
 sg13g2_fill_8 FILLER_200_360 ();
 sg13g2_fill_8 FILLER_200_368 ();
 sg13g2_fill_8 FILLER_200_376 ();
 sg13g2_fill_8 FILLER_200_384 ();
 sg13g2_fill_8 FILLER_200_392 ();
 sg13g2_fill_8 FILLER_200_400 ();
 sg13g2_fill_8 FILLER_200_408 ();
 sg13g2_fill_8 FILLER_200_416 ();
 sg13g2_fill_8 FILLER_200_424 ();
 sg13g2_fill_8 FILLER_200_432 ();
 sg13g2_fill_8 FILLER_200_440 ();
 sg13g2_fill_8 FILLER_200_448 ();
 sg13g2_fill_8 FILLER_200_456 ();
 sg13g2_fill_8 FILLER_200_464 ();
 sg13g2_fill_8 FILLER_200_472 ();
 sg13g2_fill_8 FILLER_200_480 ();
 sg13g2_fill_8 FILLER_200_488 ();
 sg13g2_fill_8 FILLER_200_496 ();
 sg13g2_fill_8 FILLER_200_504 ();
 sg13g2_fill_8 FILLER_200_512 ();
 sg13g2_fill_8 FILLER_200_520 ();
 sg13g2_fill_8 FILLER_200_528 ();
 sg13g2_fill_8 FILLER_200_536 ();
 sg13g2_fill_8 FILLER_200_544 ();
 sg13g2_fill_8 FILLER_200_552 ();
 sg13g2_fill_8 FILLER_200_560 ();
 sg13g2_fill_8 FILLER_200_568 ();
 sg13g2_fill_8 FILLER_200_576 ();
 sg13g2_fill_8 FILLER_200_584 ();
 sg13g2_fill_8 FILLER_200_592 ();
 sg13g2_fill_8 FILLER_200_600 ();
 sg13g2_fill_8 FILLER_200_608 ();
 sg13g2_fill_8 FILLER_200_616 ();
 sg13g2_fill_8 FILLER_200_624 ();
 sg13g2_fill_8 FILLER_200_632 ();
 sg13g2_fill_8 FILLER_200_640 ();
 sg13g2_fill_8 FILLER_200_648 ();
 sg13g2_fill_8 FILLER_200_656 ();
 sg13g2_fill_8 FILLER_200_664 ();
 sg13g2_fill_8 FILLER_200_672 ();
 sg13g2_fill_8 FILLER_200_680 ();
 sg13g2_fill_8 FILLER_200_688 ();
 sg13g2_fill_8 FILLER_200_696 ();
 sg13g2_fill_8 FILLER_200_704 ();
 sg13g2_fill_8 FILLER_200_712 ();
 sg13g2_fill_8 FILLER_200_720 ();
 sg13g2_fill_8 FILLER_200_728 ();
 sg13g2_fill_8 FILLER_200_736 ();
 sg13g2_fill_8 FILLER_200_744 ();
 sg13g2_fill_8 FILLER_200_752 ();
 sg13g2_fill_8 FILLER_200_760 ();
 sg13g2_fill_8 FILLER_200_768 ();
 sg13g2_fill_8 FILLER_200_776 ();
 sg13g2_fill_8 FILLER_200_784 ();
 sg13g2_fill_8 FILLER_200_792 ();
 sg13g2_fill_8 FILLER_200_800 ();
 sg13g2_fill_8 FILLER_200_808 ();
 sg13g2_fill_8 FILLER_200_816 ();
 sg13g2_fill_8 FILLER_200_824 ();
 sg13g2_fill_8 FILLER_200_832 ();
 sg13g2_fill_8 FILLER_200_840 ();
 sg13g2_fill_8 FILLER_200_848 ();
 sg13g2_fill_8 FILLER_200_856 ();
 sg13g2_fill_8 FILLER_200_864 ();
 sg13g2_fill_8 FILLER_200_872 ();
 sg13g2_fill_8 FILLER_200_880 ();
 sg13g2_fill_8 FILLER_200_888 ();
 sg13g2_fill_8 FILLER_200_896 ();
 sg13g2_fill_8 FILLER_200_904 ();
 sg13g2_fill_8 FILLER_200_912 ();
 sg13g2_fill_8 FILLER_200_920 ();
 sg13g2_fill_8 FILLER_200_928 ();
 sg13g2_fill_8 FILLER_200_936 ();
 sg13g2_fill_8 FILLER_200_944 ();
 sg13g2_fill_8 FILLER_200_952 ();
 sg13g2_fill_8 FILLER_200_960 ();
 sg13g2_fill_8 FILLER_200_968 ();
 sg13g2_fill_8 FILLER_200_976 ();
 sg13g2_fill_8 FILLER_200_984 ();
 sg13g2_fill_8 FILLER_200_992 ();
 sg13g2_fill_8 FILLER_200_1000 ();
 sg13g2_fill_8 FILLER_200_1008 ();
 sg13g2_fill_8 FILLER_200_1016 ();
 sg13g2_fill_8 FILLER_200_1024 ();
 sg13g2_fill_8 FILLER_200_1032 ();
 sg13g2_fill_8 FILLER_200_1040 ();
 sg13g2_fill_8 FILLER_200_1048 ();
 sg13g2_fill_8 FILLER_200_1056 ();
 sg13g2_fill_8 FILLER_200_1064 ();
 sg13g2_fill_8 FILLER_200_1072 ();
 sg13g2_fill_4 FILLER_200_1080 ();
 sg13g2_fill_1 FILLER_200_1084 ();
 sg13g2_fill_1 FILLER_200_1088 ();
 sg13g2_fill_1 FILLER_200_1101 ();
 sg13g2_fill_2 FILLER_200_1116 ();
 sg13g2_fill_4 FILLER_200_1123 ();
 sg13g2_fill_2 FILLER_200_1127 ();
 sg13g2_fill_1 FILLER_200_1139 ();
 sg13g2_fill_8 FILLER_200_1172 ();
 sg13g2_fill_2 FILLER_200_1180 ();
 sg13g2_fill_1 FILLER_200_1182 ();
 sg13g2_fill_8 FILLER_200_1191 ();
 sg13g2_fill_2 FILLER_200_1199 ();
 sg13g2_fill_4 FILLER_200_1226 ();
 sg13g2_fill_2 FILLER_200_1235 ();
 sg13g2_fill_1 FILLER_200_1237 ();
 sg13g2_fill_2 FILLER_200_1243 ();
 sg13g2_fill_2 FILLER_200_1249 ();
 sg13g2_fill_4 FILLER_200_1255 ();
 sg13g2_fill_2 FILLER_200_1275 ();
 sg13g2_fill_8 FILLER_200_1285 ();
 sg13g2_fill_8 FILLER_200_1293 ();
 sg13g2_fill_1 FILLER_200_1301 ();
 sg13g2_fill_2 FILLER_200_1322 ();
 sg13g2_fill_1 FILLER_200_1324 ();
 sg13g2_fill_8 FILLER_200_1333 ();
 sg13g2_fill_8 FILLER_200_1341 ();
 sg13g2_fill_8 FILLER_200_1354 ();
 sg13g2_fill_2 FILLER_200_1362 ();
 sg13g2_fill_8 FILLER_200_1370 ();
 sg13g2_fill_8 FILLER_200_1378 ();
 sg13g2_fill_8 FILLER_200_1386 ();
 sg13g2_fill_8 FILLER_200_1394 ();
 sg13g2_fill_8 FILLER_200_1402 ();
 sg13g2_fill_8 FILLER_200_1410 ();
 sg13g2_fill_8 FILLER_200_1418 ();
 sg13g2_fill_8 FILLER_200_1426 ();
 sg13g2_fill_8 FILLER_200_1434 ();
 sg13g2_fill_8 FILLER_200_1442 ();
 sg13g2_fill_8 FILLER_200_1450 ();
 sg13g2_fill_8 FILLER_200_1458 ();
 sg13g2_fill_8 FILLER_200_1466 ();
 sg13g2_fill_8 FILLER_200_1474 ();
 sg13g2_fill_8 FILLER_200_1482 ();
 sg13g2_fill_8 FILLER_200_1490 ();
 sg13g2_fill_8 FILLER_200_1498 ();
 sg13g2_fill_8 FILLER_200_1506 ();
 sg13g2_fill_8 FILLER_200_1514 ();
 sg13g2_fill_8 FILLER_200_1522 ();
 sg13g2_fill_8 FILLER_200_1530 ();
 sg13g2_fill_8 FILLER_200_1538 ();
 sg13g2_fill_8 FILLER_200_1546 ();
 sg13g2_fill_8 FILLER_200_1554 ();
 sg13g2_fill_8 FILLER_200_1562 ();
 sg13g2_fill_8 FILLER_200_1570 ();
 sg13g2_fill_8 FILLER_200_1578 ();
 sg13g2_fill_4 FILLER_200_1586 ();
 sg13g2_fill_2 FILLER_200_1590 ();
 sg13g2_fill_8 FILLER_201_0 ();
 sg13g2_fill_8 FILLER_201_8 ();
 sg13g2_fill_8 FILLER_201_16 ();
 sg13g2_fill_8 FILLER_201_24 ();
 sg13g2_fill_8 FILLER_201_32 ();
 sg13g2_fill_8 FILLER_201_40 ();
 sg13g2_fill_8 FILLER_201_48 ();
 sg13g2_fill_8 FILLER_201_56 ();
 sg13g2_fill_8 FILLER_201_64 ();
 sg13g2_fill_8 FILLER_201_72 ();
 sg13g2_fill_8 FILLER_201_80 ();
 sg13g2_fill_8 FILLER_201_88 ();
 sg13g2_fill_8 FILLER_201_96 ();
 sg13g2_fill_8 FILLER_201_104 ();
 sg13g2_fill_8 FILLER_201_112 ();
 sg13g2_fill_8 FILLER_201_120 ();
 sg13g2_fill_8 FILLER_201_128 ();
 sg13g2_fill_8 FILLER_201_136 ();
 sg13g2_fill_8 FILLER_201_144 ();
 sg13g2_fill_8 FILLER_201_152 ();
 sg13g2_fill_8 FILLER_201_160 ();
 sg13g2_fill_8 FILLER_201_168 ();
 sg13g2_fill_8 FILLER_201_176 ();
 sg13g2_fill_8 FILLER_201_184 ();
 sg13g2_fill_8 FILLER_201_192 ();
 sg13g2_fill_8 FILLER_201_200 ();
 sg13g2_fill_8 FILLER_201_208 ();
 sg13g2_fill_8 FILLER_201_216 ();
 sg13g2_fill_8 FILLER_201_224 ();
 sg13g2_fill_8 FILLER_201_232 ();
 sg13g2_fill_8 FILLER_201_240 ();
 sg13g2_fill_8 FILLER_201_248 ();
 sg13g2_fill_8 FILLER_201_256 ();
 sg13g2_fill_8 FILLER_201_264 ();
 sg13g2_fill_8 FILLER_201_272 ();
 sg13g2_fill_8 FILLER_201_280 ();
 sg13g2_fill_8 FILLER_201_288 ();
 sg13g2_fill_8 FILLER_201_296 ();
 sg13g2_fill_8 FILLER_201_304 ();
 sg13g2_fill_8 FILLER_201_312 ();
 sg13g2_fill_8 FILLER_201_320 ();
 sg13g2_fill_8 FILLER_201_328 ();
 sg13g2_fill_8 FILLER_201_336 ();
 sg13g2_fill_8 FILLER_201_344 ();
 sg13g2_fill_8 FILLER_201_352 ();
 sg13g2_fill_8 FILLER_201_360 ();
 sg13g2_fill_8 FILLER_201_368 ();
 sg13g2_fill_8 FILLER_201_376 ();
 sg13g2_fill_8 FILLER_201_384 ();
 sg13g2_fill_8 FILLER_201_392 ();
 sg13g2_fill_8 FILLER_201_400 ();
 sg13g2_fill_8 FILLER_201_408 ();
 sg13g2_fill_8 FILLER_201_416 ();
 sg13g2_fill_8 FILLER_201_424 ();
 sg13g2_fill_8 FILLER_201_432 ();
 sg13g2_fill_8 FILLER_201_440 ();
 sg13g2_fill_8 FILLER_201_448 ();
 sg13g2_fill_8 FILLER_201_456 ();
 sg13g2_fill_8 FILLER_201_464 ();
 sg13g2_fill_8 FILLER_201_472 ();
 sg13g2_fill_8 FILLER_201_480 ();
 sg13g2_fill_8 FILLER_201_488 ();
 sg13g2_fill_8 FILLER_201_496 ();
 sg13g2_fill_8 FILLER_201_504 ();
 sg13g2_fill_8 FILLER_201_512 ();
 sg13g2_fill_8 FILLER_201_520 ();
 sg13g2_fill_8 FILLER_201_528 ();
 sg13g2_fill_8 FILLER_201_536 ();
 sg13g2_fill_8 FILLER_201_544 ();
 sg13g2_fill_8 FILLER_201_552 ();
 sg13g2_fill_8 FILLER_201_560 ();
 sg13g2_fill_8 FILLER_201_568 ();
 sg13g2_fill_8 FILLER_201_576 ();
 sg13g2_fill_8 FILLER_201_584 ();
 sg13g2_fill_8 FILLER_201_592 ();
 sg13g2_fill_8 FILLER_201_600 ();
 sg13g2_fill_8 FILLER_201_608 ();
 sg13g2_fill_8 FILLER_201_616 ();
 sg13g2_fill_8 FILLER_201_624 ();
 sg13g2_fill_8 FILLER_201_632 ();
 sg13g2_fill_8 FILLER_201_640 ();
 sg13g2_fill_8 FILLER_201_648 ();
 sg13g2_fill_8 FILLER_201_656 ();
 sg13g2_fill_8 FILLER_201_664 ();
 sg13g2_fill_8 FILLER_201_672 ();
 sg13g2_fill_8 FILLER_201_680 ();
 sg13g2_fill_8 FILLER_201_688 ();
 sg13g2_fill_8 FILLER_201_696 ();
 sg13g2_fill_8 FILLER_201_704 ();
 sg13g2_fill_8 FILLER_201_712 ();
 sg13g2_fill_8 FILLER_201_720 ();
 sg13g2_fill_8 FILLER_201_728 ();
 sg13g2_fill_8 FILLER_201_736 ();
 sg13g2_fill_8 FILLER_201_744 ();
 sg13g2_fill_8 FILLER_201_752 ();
 sg13g2_fill_8 FILLER_201_760 ();
 sg13g2_fill_8 FILLER_201_768 ();
 sg13g2_fill_8 FILLER_201_776 ();
 sg13g2_fill_8 FILLER_201_784 ();
 sg13g2_fill_8 FILLER_201_792 ();
 sg13g2_fill_8 FILLER_201_800 ();
 sg13g2_fill_8 FILLER_201_808 ();
 sg13g2_fill_8 FILLER_201_816 ();
 sg13g2_fill_8 FILLER_201_824 ();
 sg13g2_fill_8 FILLER_201_832 ();
 sg13g2_fill_8 FILLER_201_840 ();
 sg13g2_fill_8 FILLER_201_848 ();
 sg13g2_fill_8 FILLER_201_856 ();
 sg13g2_fill_8 FILLER_201_864 ();
 sg13g2_fill_8 FILLER_201_872 ();
 sg13g2_fill_8 FILLER_201_880 ();
 sg13g2_fill_8 FILLER_201_888 ();
 sg13g2_fill_8 FILLER_201_896 ();
 sg13g2_fill_8 FILLER_201_904 ();
 sg13g2_fill_8 FILLER_201_912 ();
 sg13g2_fill_8 FILLER_201_920 ();
 sg13g2_fill_8 FILLER_201_928 ();
 sg13g2_fill_8 FILLER_201_936 ();
 sg13g2_fill_8 FILLER_201_944 ();
 sg13g2_fill_8 FILLER_201_952 ();
 sg13g2_fill_8 FILLER_201_960 ();
 sg13g2_fill_8 FILLER_201_968 ();
 sg13g2_fill_8 FILLER_201_976 ();
 sg13g2_fill_8 FILLER_201_984 ();
 sg13g2_fill_8 FILLER_201_992 ();
 sg13g2_fill_8 FILLER_201_1000 ();
 sg13g2_fill_8 FILLER_201_1008 ();
 sg13g2_fill_8 FILLER_201_1016 ();
 sg13g2_fill_8 FILLER_201_1024 ();
 sg13g2_fill_8 FILLER_201_1032 ();
 sg13g2_fill_8 FILLER_201_1040 ();
 sg13g2_fill_8 FILLER_201_1048 ();
 sg13g2_fill_8 FILLER_201_1056 ();
 sg13g2_fill_4 FILLER_201_1064 ();
 sg13g2_fill_2 FILLER_201_1068 ();
 sg13g2_fill_1 FILLER_201_1070 ();
 sg13g2_fill_2 FILLER_201_1079 ();
 sg13g2_fill_8 FILLER_201_1134 ();
 sg13g2_fill_8 FILLER_201_1142 ();
 sg13g2_fill_8 FILLER_201_1150 ();
 sg13g2_fill_8 FILLER_201_1158 ();
 sg13g2_fill_2 FILLER_201_1166 ();
 sg13g2_fill_1 FILLER_201_1168 ();
 sg13g2_fill_1 FILLER_201_1181 ();
 sg13g2_fill_4 FILLER_201_1196 ();
 sg13g2_fill_2 FILLER_201_1200 ();
 sg13g2_fill_1 FILLER_201_1202 ();
 sg13g2_fill_8 FILLER_201_1214 ();
 sg13g2_fill_2 FILLER_201_1259 ();
 sg13g2_fill_8 FILLER_201_1267 ();
 sg13g2_fill_8 FILLER_201_1275 ();
 sg13g2_fill_2 FILLER_201_1287 ();
 sg13g2_fill_1 FILLER_201_1289 ();
 sg13g2_fill_2 FILLER_201_1299 ();
 sg13g2_fill_1 FILLER_201_1301 ();
 sg13g2_fill_1 FILLER_201_1314 ();
 sg13g2_fill_8 FILLER_201_1320 ();
 sg13g2_fill_8 FILLER_201_1328 ();
 sg13g2_fill_8 FILLER_201_1336 ();
 sg13g2_fill_8 FILLER_201_1344 ();
 sg13g2_fill_8 FILLER_201_1352 ();
 sg13g2_fill_8 FILLER_201_1360 ();
 sg13g2_fill_8 FILLER_201_1368 ();
 sg13g2_fill_8 FILLER_201_1376 ();
 sg13g2_fill_8 FILLER_201_1384 ();
 sg13g2_fill_8 FILLER_201_1392 ();
 sg13g2_fill_8 FILLER_201_1400 ();
 sg13g2_fill_8 FILLER_201_1408 ();
 sg13g2_fill_8 FILLER_201_1416 ();
 sg13g2_fill_8 FILLER_201_1424 ();
 sg13g2_fill_8 FILLER_201_1432 ();
 sg13g2_fill_8 FILLER_201_1440 ();
 sg13g2_fill_8 FILLER_201_1448 ();
 sg13g2_fill_8 FILLER_201_1456 ();
 sg13g2_fill_8 FILLER_201_1464 ();
 sg13g2_fill_8 FILLER_201_1472 ();
 sg13g2_fill_8 FILLER_201_1480 ();
 sg13g2_fill_8 FILLER_201_1488 ();
 sg13g2_fill_8 FILLER_201_1496 ();
 sg13g2_fill_8 FILLER_201_1504 ();
 sg13g2_fill_8 FILLER_201_1512 ();
 sg13g2_fill_8 FILLER_201_1520 ();
 sg13g2_fill_8 FILLER_201_1528 ();
 sg13g2_fill_8 FILLER_201_1536 ();
 sg13g2_fill_8 FILLER_201_1544 ();
 sg13g2_fill_8 FILLER_201_1552 ();
 sg13g2_fill_8 FILLER_201_1560 ();
 sg13g2_fill_8 FILLER_201_1568 ();
 sg13g2_fill_8 FILLER_201_1576 ();
 sg13g2_fill_8 FILLER_201_1584 ();
 sg13g2_fill_8 FILLER_202_0 ();
 sg13g2_fill_8 FILLER_202_8 ();
 sg13g2_fill_8 FILLER_202_16 ();
 sg13g2_fill_8 FILLER_202_24 ();
 sg13g2_fill_8 FILLER_202_32 ();
 sg13g2_fill_8 FILLER_202_40 ();
 sg13g2_fill_8 FILLER_202_48 ();
 sg13g2_fill_8 FILLER_202_56 ();
 sg13g2_fill_8 FILLER_202_64 ();
 sg13g2_fill_8 FILLER_202_72 ();
 sg13g2_fill_8 FILLER_202_80 ();
 sg13g2_fill_8 FILLER_202_88 ();
 sg13g2_fill_8 FILLER_202_96 ();
 sg13g2_fill_8 FILLER_202_104 ();
 sg13g2_fill_8 FILLER_202_112 ();
 sg13g2_fill_8 FILLER_202_120 ();
 sg13g2_fill_8 FILLER_202_128 ();
 sg13g2_fill_8 FILLER_202_136 ();
 sg13g2_fill_8 FILLER_202_144 ();
 sg13g2_fill_8 FILLER_202_152 ();
 sg13g2_fill_8 FILLER_202_160 ();
 sg13g2_fill_8 FILLER_202_168 ();
 sg13g2_fill_8 FILLER_202_176 ();
 sg13g2_fill_8 FILLER_202_184 ();
 sg13g2_fill_8 FILLER_202_192 ();
 sg13g2_fill_8 FILLER_202_200 ();
 sg13g2_fill_8 FILLER_202_208 ();
 sg13g2_fill_8 FILLER_202_216 ();
 sg13g2_fill_8 FILLER_202_224 ();
 sg13g2_fill_8 FILLER_202_232 ();
 sg13g2_fill_8 FILLER_202_240 ();
 sg13g2_fill_8 FILLER_202_248 ();
 sg13g2_fill_8 FILLER_202_256 ();
 sg13g2_fill_8 FILLER_202_264 ();
 sg13g2_fill_8 FILLER_202_272 ();
 sg13g2_fill_8 FILLER_202_280 ();
 sg13g2_fill_8 FILLER_202_288 ();
 sg13g2_fill_8 FILLER_202_296 ();
 sg13g2_fill_8 FILLER_202_304 ();
 sg13g2_fill_8 FILLER_202_312 ();
 sg13g2_fill_8 FILLER_202_320 ();
 sg13g2_fill_8 FILLER_202_328 ();
 sg13g2_fill_8 FILLER_202_336 ();
 sg13g2_fill_8 FILLER_202_344 ();
 sg13g2_fill_8 FILLER_202_352 ();
 sg13g2_fill_8 FILLER_202_360 ();
 sg13g2_fill_8 FILLER_202_368 ();
 sg13g2_fill_8 FILLER_202_376 ();
 sg13g2_fill_8 FILLER_202_384 ();
 sg13g2_fill_8 FILLER_202_392 ();
 sg13g2_fill_8 FILLER_202_400 ();
 sg13g2_fill_8 FILLER_202_408 ();
 sg13g2_fill_8 FILLER_202_416 ();
 sg13g2_fill_8 FILLER_202_424 ();
 sg13g2_fill_8 FILLER_202_432 ();
 sg13g2_fill_8 FILLER_202_440 ();
 sg13g2_fill_8 FILLER_202_448 ();
 sg13g2_fill_8 FILLER_202_456 ();
 sg13g2_fill_8 FILLER_202_464 ();
 sg13g2_fill_8 FILLER_202_472 ();
 sg13g2_fill_8 FILLER_202_480 ();
 sg13g2_fill_8 FILLER_202_488 ();
 sg13g2_fill_8 FILLER_202_496 ();
 sg13g2_fill_8 FILLER_202_504 ();
 sg13g2_fill_8 FILLER_202_512 ();
 sg13g2_fill_8 FILLER_202_520 ();
 sg13g2_fill_8 FILLER_202_528 ();
 sg13g2_fill_8 FILLER_202_536 ();
 sg13g2_fill_8 FILLER_202_544 ();
 sg13g2_fill_8 FILLER_202_552 ();
 sg13g2_fill_8 FILLER_202_560 ();
 sg13g2_fill_8 FILLER_202_568 ();
 sg13g2_fill_8 FILLER_202_576 ();
 sg13g2_fill_8 FILLER_202_584 ();
 sg13g2_fill_8 FILLER_202_592 ();
 sg13g2_fill_8 FILLER_202_600 ();
 sg13g2_fill_8 FILLER_202_608 ();
 sg13g2_fill_8 FILLER_202_616 ();
 sg13g2_fill_8 FILLER_202_624 ();
 sg13g2_fill_8 FILLER_202_632 ();
 sg13g2_fill_8 FILLER_202_640 ();
 sg13g2_fill_8 FILLER_202_648 ();
 sg13g2_fill_8 FILLER_202_656 ();
 sg13g2_fill_8 FILLER_202_664 ();
 sg13g2_fill_8 FILLER_202_672 ();
 sg13g2_fill_8 FILLER_202_680 ();
 sg13g2_fill_8 FILLER_202_688 ();
 sg13g2_fill_8 FILLER_202_696 ();
 sg13g2_fill_8 FILLER_202_704 ();
 sg13g2_fill_8 FILLER_202_712 ();
 sg13g2_fill_8 FILLER_202_720 ();
 sg13g2_fill_8 FILLER_202_728 ();
 sg13g2_fill_8 FILLER_202_736 ();
 sg13g2_fill_8 FILLER_202_744 ();
 sg13g2_fill_8 FILLER_202_752 ();
 sg13g2_fill_8 FILLER_202_760 ();
 sg13g2_fill_8 FILLER_202_768 ();
 sg13g2_fill_8 FILLER_202_776 ();
 sg13g2_fill_8 FILLER_202_784 ();
 sg13g2_fill_8 FILLER_202_792 ();
 sg13g2_fill_8 FILLER_202_800 ();
 sg13g2_fill_8 FILLER_202_808 ();
 sg13g2_fill_8 FILLER_202_816 ();
 sg13g2_fill_8 FILLER_202_824 ();
 sg13g2_fill_8 FILLER_202_832 ();
 sg13g2_fill_8 FILLER_202_840 ();
 sg13g2_fill_8 FILLER_202_848 ();
 sg13g2_fill_8 FILLER_202_856 ();
 sg13g2_fill_8 FILLER_202_864 ();
 sg13g2_fill_8 FILLER_202_872 ();
 sg13g2_fill_8 FILLER_202_880 ();
 sg13g2_fill_8 FILLER_202_888 ();
 sg13g2_fill_8 FILLER_202_896 ();
 sg13g2_fill_8 FILLER_202_904 ();
 sg13g2_fill_8 FILLER_202_912 ();
 sg13g2_fill_8 FILLER_202_920 ();
 sg13g2_fill_8 FILLER_202_928 ();
 sg13g2_fill_8 FILLER_202_936 ();
 sg13g2_fill_8 FILLER_202_944 ();
 sg13g2_fill_8 FILLER_202_952 ();
 sg13g2_fill_8 FILLER_202_960 ();
 sg13g2_fill_8 FILLER_202_968 ();
 sg13g2_fill_8 FILLER_202_976 ();
 sg13g2_fill_8 FILLER_202_984 ();
 sg13g2_fill_8 FILLER_202_992 ();
 sg13g2_fill_8 FILLER_202_1000 ();
 sg13g2_fill_8 FILLER_202_1008 ();
 sg13g2_fill_8 FILLER_202_1016 ();
 sg13g2_fill_8 FILLER_202_1024 ();
 sg13g2_fill_8 FILLER_202_1032 ();
 sg13g2_fill_8 FILLER_202_1040 ();
 sg13g2_fill_8 FILLER_202_1048 ();
 sg13g2_fill_8 FILLER_202_1056 ();
 sg13g2_fill_8 FILLER_202_1064 ();
 sg13g2_fill_8 FILLER_202_1072 ();
 sg13g2_fill_4 FILLER_202_1080 ();
 sg13g2_fill_2 FILLER_202_1110 ();
 sg13g2_fill_4 FILLER_202_1136 ();
 sg13g2_fill_2 FILLER_202_1140 ();
 sg13g2_fill_8 FILLER_202_1155 ();
 sg13g2_fill_2 FILLER_202_1205 ();
 sg13g2_fill_1 FILLER_202_1207 ();
 sg13g2_fill_8 FILLER_202_1216 ();
 sg13g2_fill_2 FILLER_202_1224 ();
 sg13g2_fill_4 FILLER_202_1231 ();
 sg13g2_fill_2 FILLER_202_1235 ();
 sg13g2_fill_1 FILLER_202_1237 ();
 sg13g2_fill_8 FILLER_202_1241 ();
 sg13g2_fill_8 FILLER_202_1249 ();
 sg13g2_fill_8 FILLER_202_1257 ();
 sg13g2_fill_8 FILLER_202_1265 ();
 sg13g2_fill_4 FILLER_202_1273 ();
 sg13g2_fill_2 FILLER_202_1277 ();
 sg13g2_fill_8 FILLER_202_1290 ();
 sg13g2_fill_1 FILLER_202_1298 ();
 sg13g2_fill_8 FILLER_202_1324 ();
 sg13g2_fill_8 FILLER_202_1332 ();
 sg13g2_fill_8 FILLER_202_1340 ();
 sg13g2_fill_8 FILLER_202_1348 ();
 sg13g2_fill_8 FILLER_202_1356 ();
 sg13g2_fill_8 FILLER_202_1364 ();
 sg13g2_fill_8 FILLER_202_1372 ();
 sg13g2_fill_8 FILLER_202_1380 ();
 sg13g2_fill_8 FILLER_202_1388 ();
 sg13g2_fill_8 FILLER_202_1396 ();
 sg13g2_fill_8 FILLER_202_1404 ();
 sg13g2_fill_8 FILLER_202_1412 ();
 sg13g2_fill_8 FILLER_202_1420 ();
 sg13g2_fill_8 FILLER_202_1428 ();
 sg13g2_fill_8 FILLER_202_1436 ();
 sg13g2_fill_8 FILLER_202_1444 ();
 sg13g2_fill_8 FILLER_202_1452 ();
 sg13g2_fill_8 FILLER_202_1460 ();
 sg13g2_fill_8 FILLER_202_1468 ();
 sg13g2_fill_8 FILLER_202_1476 ();
 sg13g2_fill_8 FILLER_202_1484 ();
 sg13g2_fill_8 FILLER_202_1492 ();
 sg13g2_fill_8 FILLER_202_1500 ();
 sg13g2_fill_8 FILLER_202_1508 ();
 sg13g2_fill_8 FILLER_202_1516 ();
 sg13g2_fill_8 FILLER_202_1524 ();
 sg13g2_fill_8 FILLER_202_1532 ();
 sg13g2_fill_8 FILLER_202_1540 ();
 sg13g2_fill_8 FILLER_202_1548 ();
 sg13g2_fill_8 FILLER_202_1556 ();
 sg13g2_fill_8 FILLER_202_1564 ();
 sg13g2_fill_8 FILLER_202_1572 ();
 sg13g2_fill_8 FILLER_202_1580 ();
 sg13g2_fill_4 FILLER_202_1588 ();
 sg13g2_fill_8 FILLER_203_0 ();
 sg13g2_fill_8 FILLER_203_8 ();
 sg13g2_fill_8 FILLER_203_16 ();
 sg13g2_fill_8 FILLER_203_24 ();
 sg13g2_fill_8 FILLER_203_32 ();
 sg13g2_fill_8 FILLER_203_40 ();
 sg13g2_fill_8 FILLER_203_48 ();
 sg13g2_fill_8 FILLER_203_56 ();
 sg13g2_fill_8 FILLER_203_64 ();
 sg13g2_fill_8 FILLER_203_72 ();
 sg13g2_fill_8 FILLER_203_80 ();
 sg13g2_fill_8 FILLER_203_88 ();
 sg13g2_fill_8 FILLER_203_96 ();
 sg13g2_fill_8 FILLER_203_104 ();
 sg13g2_fill_8 FILLER_203_112 ();
 sg13g2_fill_8 FILLER_203_120 ();
 sg13g2_fill_8 FILLER_203_128 ();
 sg13g2_fill_8 FILLER_203_136 ();
 sg13g2_fill_8 FILLER_203_144 ();
 sg13g2_fill_8 FILLER_203_152 ();
 sg13g2_fill_8 FILLER_203_160 ();
 sg13g2_fill_8 FILLER_203_168 ();
 sg13g2_fill_8 FILLER_203_176 ();
 sg13g2_fill_8 FILLER_203_184 ();
 sg13g2_fill_8 FILLER_203_192 ();
 sg13g2_fill_8 FILLER_203_200 ();
 sg13g2_fill_8 FILLER_203_208 ();
 sg13g2_fill_8 FILLER_203_216 ();
 sg13g2_fill_8 FILLER_203_224 ();
 sg13g2_fill_8 FILLER_203_232 ();
 sg13g2_fill_8 FILLER_203_240 ();
 sg13g2_fill_8 FILLER_203_248 ();
 sg13g2_fill_8 FILLER_203_256 ();
 sg13g2_fill_8 FILLER_203_264 ();
 sg13g2_fill_8 FILLER_203_272 ();
 sg13g2_fill_8 FILLER_203_280 ();
 sg13g2_fill_8 FILLER_203_288 ();
 sg13g2_fill_8 FILLER_203_296 ();
 sg13g2_fill_8 FILLER_203_304 ();
 sg13g2_fill_8 FILLER_203_312 ();
 sg13g2_fill_8 FILLER_203_320 ();
 sg13g2_fill_8 FILLER_203_328 ();
 sg13g2_fill_8 FILLER_203_336 ();
 sg13g2_fill_8 FILLER_203_344 ();
 sg13g2_fill_8 FILLER_203_352 ();
 sg13g2_fill_8 FILLER_203_360 ();
 sg13g2_fill_8 FILLER_203_368 ();
 sg13g2_fill_8 FILLER_203_376 ();
 sg13g2_fill_8 FILLER_203_384 ();
 sg13g2_fill_8 FILLER_203_392 ();
 sg13g2_fill_8 FILLER_203_400 ();
 sg13g2_fill_8 FILLER_203_408 ();
 sg13g2_fill_8 FILLER_203_416 ();
 sg13g2_fill_8 FILLER_203_424 ();
 sg13g2_fill_8 FILLER_203_432 ();
 sg13g2_fill_8 FILLER_203_440 ();
 sg13g2_fill_8 FILLER_203_448 ();
 sg13g2_fill_8 FILLER_203_456 ();
 sg13g2_fill_8 FILLER_203_464 ();
 sg13g2_fill_8 FILLER_203_472 ();
 sg13g2_fill_8 FILLER_203_480 ();
 sg13g2_fill_8 FILLER_203_488 ();
 sg13g2_fill_8 FILLER_203_496 ();
 sg13g2_fill_8 FILLER_203_504 ();
 sg13g2_fill_8 FILLER_203_512 ();
 sg13g2_fill_8 FILLER_203_520 ();
 sg13g2_fill_8 FILLER_203_528 ();
 sg13g2_fill_8 FILLER_203_536 ();
 sg13g2_fill_8 FILLER_203_544 ();
 sg13g2_fill_8 FILLER_203_552 ();
 sg13g2_fill_8 FILLER_203_560 ();
 sg13g2_fill_8 FILLER_203_568 ();
 sg13g2_fill_8 FILLER_203_576 ();
 sg13g2_fill_8 FILLER_203_584 ();
 sg13g2_fill_8 FILLER_203_592 ();
 sg13g2_fill_8 FILLER_203_600 ();
 sg13g2_fill_8 FILLER_203_608 ();
 sg13g2_fill_8 FILLER_203_616 ();
 sg13g2_fill_8 FILLER_203_624 ();
 sg13g2_fill_8 FILLER_203_632 ();
 sg13g2_fill_8 FILLER_203_640 ();
 sg13g2_fill_8 FILLER_203_648 ();
 sg13g2_fill_8 FILLER_203_656 ();
 sg13g2_fill_8 FILLER_203_664 ();
 sg13g2_fill_8 FILLER_203_672 ();
 sg13g2_fill_8 FILLER_203_680 ();
 sg13g2_fill_8 FILLER_203_688 ();
 sg13g2_fill_8 FILLER_203_696 ();
 sg13g2_fill_8 FILLER_203_704 ();
 sg13g2_fill_8 FILLER_203_712 ();
 sg13g2_fill_8 FILLER_203_720 ();
 sg13g2_fill_8 FILLER_203_728 ();
 sg13g2_fill_8 FILLER_203_736 ();
 sg13g2_fill_8 FILLER_203_744 ();
 sg13g2_fill_8 FILLER_203_752 ();
 sg13g2_fill_8 FILLER_203_760 ();
 sg13g2_fill_8 FILLER_203_768 ();
 sg13g2_fill_8 FILLER_203_776 ();
 sg13g2_fill_8 FILLER_203_784 ();
 sg13g2_fill_8 FILLER_203_792 ();
 sg13g2_fill_8 FILLER_203_800 ();
 sg13g2_fill_8 FILLER_203_808 ();
 sg13g2_fill_8 FILLER_203_816 ();
 sg13g2_fill_8 FILLER_203_824 ();
 sg13g2_fill_8 FILLER_203_832 ();
 sg13g2_fill_8 FILLER_203_840 ();
 sg13g2_fill_8 FILLER_203_848 ();
 sg13g2_fill_8 FILLER_203_856 ();
 sg13g2_fill_8 FILLER_203_864 ();
 sg13g2_fill_8 FILLER_203_872 ();
 sg13g2_fill_8 FILLER_203_880 ();
 sg13g2_fill_8 FILLER_203_888 ();
 sg13g2_fill_8 FILLER_203_896 ();
 sg13g2_fill_8 FILLER_203_904 ();
 sg13g2_fill_8 FILLER_203_912 ();
 sg13g2_fill_8 FILLER_203_920 ();
 sg13g2_fill_8 FILLER_203_928 ();
 sg13g2_fill_8 FILLER_203_936 ();
 sg13g2_fill_8 FILLER_203_944 ();
 sg13g2_fill_8 FILLER_203_952 ();
 sg13g2_fill_8 FILLER_203_960 ();
 sg13g2_fill_8 FILLER_203_968 ();
 sg13g2_fill_8 FILLER_203_976 ();
 sg13g2_fill_8 FILLER_203_984 ();
 sg13g2_fill_8 FILLER_203_992 ();
 sg13g2_fill_8 FILLER_203_1000 ();
 sg13g2_fill_8 FILLER_203_1008 ();
 sg13g2_fill_8 FILLER_203_1016 ();
 sg13g2_fill_8 FILLER_203_1024 ();
 sg13g2_fill_8 FILLER_203_1032 ();
 sg13g2_fill_8 FILLER_203_1040 ();
 sg13g2_fill_8 FILLER_203_1048 ();
 sg13g2_fill_8 FILLER_203_1056 ();
 sg13g2_fill_8 FILLER_203_1064 ();
 sg13g2_fill_8 FILLER_203_1072 ();
 sg13g2_fill_8 FILLER_203_1080 ();
 sg13g2_fill_4 FILLER_203_1088 ();
 sg13g2_fill_8 FILLER_203_1100 ();
 sg13g2_fill_8 FILLER_203_1108 ();
 sg13g2_fill_8 FILLER_203_1116 ();
 sg13g2_fill_8 FILLER_203_1124 ();
 sg13g2_fill_2 FILLER_203_1132 ();
 sg13g2_fill_1 FILLER_203_1142 ();
 sg13g2_fill_8 FILLER_203_1164 ();
 sg13g2_fill_1 FILLER_203_1172 ();
 sg13g2_fill_1 FILLER_203_1197 ();
 sg13g2_fill_8 FILLER_203_1213 ();
 sg13g2_fill_8 FILLER_203_1221 ();
 sg13g2_fill_4 FILLER_203_1229 ();
 sg13g2_fill_2 FILLER_203_1233 ();
 sg13g2_fill_1 FILLER_203_1235 ();
 sg13g2_fill_1 FILLER_203_1241 ();
 sg13g2_fill_1 FILLER_203_1251 ();
 sg13g2_fill_2 FILLER_203_1257 ();
 sg13g2_fill_2 FILLER_203_1268 ();
 sg13g2_fill_1 FILLER_203_1270 ();
 sg13g2_fill_1 FILLER_203_1275 ();
 sg13g2_fill_1 FILLER_203_1279 ();
 sg13g2_fill_8 FILLER_203_1285 ();
 sg13g2_fill_8 FILLER_203_1293 ();
 sg13g2_fill_2 FILLER_203_1301 ();
 sg13g2_fill_1 FILLER_203_1303 ();
 sg13g2_fill_8 FILLER_203_1308 ();
 sg13g2_fill_8 FILLER_203_1316 ();
 sg13g2_fill_8 FILLER_203_1324 ();
 sg13g2_fill_8 FILLER_203_1332 ();
 sg13g2_fill_8 FILLER_203_1340 ();
 sg13g2_fill_8 FILLER_203_1348 ();
 sg13g2_fill_8 FILLER_203_1356 ();
 sg13g2_fill_8 FILLER_203_1364 ();
 sg13g2_fill_8 FILLER_203_1372 ();
 sg13g2_fill_8 FILLER_203_1380 ();
 sg13g2_fill_8 FILLER_203_1388 ();
 sg13g2_fill_8 FILLER_203_1396 ();
 sg13g2_fill_8 FILLER_203_1404 ();
 sg13g2_fill_8 FILLER_203_1412 ();
 sg13g2_fill_8 FILLER_203_1420 ();
 sg13g2_fill_8 FILLER_203_1428 ();
 sg13g2_fill_8 FILLER_203_1436 ();
 sg13g2_fill_8 FILLER_203_1444 ();
 sg13g2_fill_8 FILLER_203_1452 ();
 sg13g2_fill_8 FILLER_203_1460 ();
 sg13g2_fill_8 FILLER_203_1468 ();
 sg13g2_fill_8 FILLER_203_1476 ();
 sg13g2_fill_8 FILLER_203_1484 ();
 sg13g2_fill_8 FILLER_203_1492 ();
 sg13g2_fill_8 FILLER_203_1500 ();
 sg13g2_fill_8 FILLER_203_1508 ();
 sg13g2_fill_8 FILLER_203_1516 ();
 sg13g2_fill_8 FILLER_203_1524 ();
 sg13g2_fill_8 FILLER_203_1532 ();
 sg13g2_fill_8 FILLER_203_1540 ();
 sg13g2_fill_8 FILLER_203_1548 ();
 sg13g2_fill_8 FILLER_203_1556 ();
 sg13g2_fill_8 FILLER_203_1564 ();
 sg13g2_fill_8 FILLER_203_1572 ();
 sg13g2_fill_8 FILLER_203_1580 ();
 sg13g2_fill_4 FILLER_203_1588 ();
 sg13g2_fill_8 FILLER_204_0 ();
 sg13g2_fill_8 FILLER_204_8 ();
 sg13g2_fill_8 FILLER_204_16 ();
 sg13g2_fill_8 FILLER_204_24 ();
 sg13g2_fill_8 FILLER_204_32 ();
 sg13g2_fill_8 FILLER_204_40 ();
 sg13g2_fill_8 FILLER_204_48 ();
 sg13g2_fill_8 FILLER_204_56 ();
 sg13g2_fill_8 FILLER_204_64 ();
 sg13g2_fill_8 FILLER_204_72 ();
 sg13g2_fill_8 FILLER_204_80 ();
 sg13g2_fill_8 FILLER_204_88 ();
 sg13g2_fill_8 FILLER_204_96 ();
 sg13g2_fill_8 FILLER_204_104 ();
 sg13g2_fill_8 FILLER_204_112 ();
 sg13g2_fill_8 FILLER_204_120 ();
 sg13g2_fill_8 FILLER_204_128 ();
 sg13g2_fill_8 FILLER_204_136 ();
 sg13g2_fill_8 FILLER_204_144 ();
 sg13g2_fill_8 FILLER_204_152 ();
 sg13g2_fill_8 FILLER_204_160 ();
 sg13g2_fill_8 FILLER_204_168 ();
 sg13g2_fill_8 FILLER_204_176 ();
 sg13g2_fill_8 FILLER_204_184 ();
 sg13g2_fill_8 FILLER_204_192 ();
 sg13g2_fill_8 FILLER_204_200 ();
 sg13g2_fill_8 FILLER_204_208 ();
 sg13g2_fill_8 FILLER_204_216 ();
 sg13g2_fill_8 FILLER_204_224 ();
 sg13g2_fill_8 FILLER_204_232 ();
 sg13g2_fill_8 FILLER_204_240 ();
 sg13g2_fill_8 FILLER_204_248 ();
 sg13g2_fill_8 FILLER_204_256 ();
 sg13g2_fill_8 FILLER_204_264 ();
 sg13g2_fill_8 FILLER_204_272 ();
 sg13g2_fill_8 FILLER_204_280 ();
 sg13g2_fill_8 FILLER_204_288 ();
 sg13g2_fill_8 FILLER_204_296 ();
 sg13g2_fill_8 FILLER_204_304 ();
 sg13g2_fill_8 FILLER_204_312 ();
 sg13g2_fill_8 FILLER_204_320 ();
 sg13g2_fill_8 FILLER_204_328 ();
 sg13g2_fill_8 FILLER_204_336 ();
 sg13g2_fill_8 FILLER_204_344 ();
 sg13g2_fill_8 FILLER_204_352 ();
 sg13g2_fill_8 FILLER_204_360 ();
 sg13g2_fill_8 FILLER_204_368 ();
 sg13g2_fill_8 FILLER_204_376 ();
 sg13g2_fill_8 FILLER_204_384 ();
 sg13g2_fill_8 FILLER_204_392 ();
 sg13g2_fill_8 FILLER_204_400 ();
 sg13g2_fill_8 FILLER_204_408 ();
 sg13g2_fill_8 FILLER_204_416 ();
 sg13g2_fill_8 FILLER_204_424 ();
 sg13g2_fill_8 FILLER_204_432 ();
 sg13g2_fill_8 FILLER_204_440 ();
 sg13g2_fill_8 FILLER_204_448 ();
 sg13g2_fill_8 FILLER_204_456 ();
 sg13g2_fill_8 FILLER_204_464 ();
 sg13g2_fill_8 FILLER_204_472 ();
 sg13g2_fill_8 FILLER_204_480 ();
 sg13g2_fill_8 FILLER_204_488 ();
 sg13g2_fill_8 FILLER_204_496 ();
 sg13g2_fill_8 FILLER_204_504 ();
 sg13g2_fill_8 FILLER_204_512 ();
 sg13g2_fill_8 FILLER_204_520 ();
 sg13g2_fill_8 FILLER_204_528 ();
 sg13g2_fill_8 FILLER_204_536 ();
 sg13g2_fill_8 FILLER_204_544 ();
 sg13g2_fill_8 FILLER_204_552 ();
 sg13g2_fill_8 FILLER_204_560 ();
 sg13g2_fill_8 FILLER_204_568 ();
 sg13g2_fill_8 FILLER_204_576 ();
 sg13g2_fill_8 FILLER_204_584 ();
 sg13g2_fill_8 FILLER_204_592 ();
 sg13g2_fill_8 FILLER_204_600 ();
 sg13g2_fill_8 FILLER_204_608 ();
 sg13g2_fill_8 FILLER_204_616 ();
 sg13g2_fill_8 FILLER_204_624 ();
 sg13g2_fill_8 FILLER_204_632 ();
 sg13g2_fill_8 FILLER_204_640 ();
 sg13g2_fill_8 FILLER_204_648 ();
 sg13g2_fill_8 FILLER_204_656 ();
 sg13g2_fill_8 FILLER_204_664 ();
 sg13g2_fill_8 FILLER_204_672 ();
 sg13g2_fill_8 FILLER_204_680 ();
 sg13g2_fill_8 FILLER_204_688 ();
 sg13g2_fill_8 FILLER_204_696 ();
 sg13g2_fill_8 FILLER_204_704 ();
 sg13g2_fill_8 FILLER_204_712 ();
 sg13g2_fill_8 FILLER_204_720 ();
 sg13g2_fill_8 FILLER_204_728 ();
 sg13g2_fill_8 FILLER_204_736 ();
 sg13g2_fill_8 FILLER_204_744 ();
 sg13g2_fill_8 FILLER_204_752 ();
 sg13g2_fill_8 FILLER_204_760 ();
 sg13g2_fill_8 FILLER_204_768 ();
 sg13g2_fill_8 FILLER_204_776 ();
 sg13g2_fill_8 FILLER_204_784 ();
 sg13g2_fill_8 FILLER_204_792 ();
 sg13g2_fill_8 FILLER_204_800 ();
 sg13g2_fill_8 FILLER_204_808 ();
 sg13g2_fill_8 FILLER_204_816 ();
 sg13g2_fill_8 FILLER_204_824 ();
 sg13g2_fill_8 FILLER_204_832 ();
 sg13g2_fill_8 FILLER_204_840 ();
 sg13g2_fill_8 FILLER_204_848 ();
 sg13g2_fill_8 FILLER_204_856 ();
 sg13g2_fill_8 FILLER_204_864 ();
 sg13g2_fill_8 FILLER_204_872 ();
 sg13g2_fill_8 FILLER_204_880 ();
 sg13g2_fill_8 FILLER_204_888 ();
 sg13g2_fill_8 FILLER_204_896 ();
 sg13g2_fill_8 FILLER_204_904 ();
 sg13g2_fill_8 FILLER_204_912 ();
 sg13g2_fill_8 FILLER_204_920 ();
 sg13g2_fill_8 FILLER_204_928 ();
 sg13g2_fill_8 FILLER_204_936 ();
 sg13g2_fill_8 FILLER_204_944 ();
 sg13g2_fill_8 FILLER_204_952 ();
 sg13g2_fill_8 FILLER_204_960 ();
 sg13g2_fill_8 FILLER_204_968 ();
 sg13g2_fill_8 FILLER_204_976 ();
 sg13g2_fill_8 FILLER_204_984 ();
 sg13g2_fill_8 FILLER_204_992 ();
 sg13g2_fill_8 FILLER_204_1000 ();
 sg13g2_fill_8 FILLER_204_1008 ();
 sg13g2_fill_8 FILLER_204_1016 ();
 sg13g2_fill_8 FILLER_204_1024 ();
 sg13g2_fill_8 FILLER_204_1032 ();
 sg13g2_fill_8 FILLER_204_1040 ();
 sg13g2_fill_8 FILLER_204_1048 ();
 sg13g2_fill_8 FILLER_204_1056 ();
 sg13g2_fill_8 FILLER_204_1064 ();
 sg13g2_fill_8 FILLER_204_1072 ();
 sg13g2_fill_8 FILLER_204_1080 ();
 sg13g2_fill_8 FILLER_204_1088 ();
 sg13g2_fill_8 FILLER_204_1096 ();
 sg13g2_fill_8 FILLER_204_1104 ();
 sg13g2_fill_8 FILLER_204_1112 ();
 sg13g2_fill_8 FILLER_204_1120 ();
 sg13g2_fill_8 FILLER_204_1128 ();
 sg13g2_fill_4 FILLER_204_1136 ();
 sg13g2_fill_2 FILLER_204_1140 ();
 sg13g2_fill_8 FILLER_204_1159 ();
 sg13g2_fill_4 FILLER_204_1167 ();
 sg13g2_fill_4 FILLER_204_1204 ();
 sg13g2_fill_4 FILLER_204_1226 ();
 sg13g2_fill_1 FILLER_204_1248 ();
 sg13g2_fill_8 FILLER_204_1293 ();
 sg13g2_fill_8 FILLER_204_1301 ();
 sg13g2_fill_8 FILLER_204_1317 ();
 sg13g2_fill_8 FILLER_204_1325 ();
 sg13g2_fill_8 FILLER_204_1333 ();
 sg13g2_fill_8 FILLER_204_1341 ();
 sg13g2_fill_8 FILLER_204_1349 ();
 sg13g2_fill_8 FILLER_204_1357 ();
 sg13g2_fill_8 FILLER_204_1365 ();
 sg13g2_fill_8 FILLER_204_1373 ();
 sg13g2_fill_8 FILLER_204_1381 ();
 sg13g2_fill_8 FILLER_204_1389 ();
 sg13g2_fill_8 FILLER_204_1397 ();
 sg13g2_fill_8 FILLER_204_1405 ();
 sg13g2_fill_8 FILLER_204_1413 ();
 sg13g2_fill_8 FILLER_204_1421 ();
 sg13g2_fill_8 FILLER_204_1429 ();
 sg13g2_fill_8 FILLER_204_1437 ();
 sg13g2_fill_8 FILLER_204_1445 ();
 sg13g2_fill_8 FILLER_204_1453 ();
 sg13g2_fill_8 FILLER_204_1461 ();
 sg13g2_fill_8 FILLER_204_1469 ();
 sg13g2_fill_8 FILLER_204_1477 ();
 sg13g2_fill_8 FILLER_204_1485 ();
 sg13g2_fill_8 FILLER_204_1493 ();
 sg13g2_fill_8 FILLER_204_1501 ();
 sg13g2_fill_8 FILLER_204_1509 ();
 sg13g2_fill_8 FILLER_204_1517 ();
 sg13g2_fill_8 FILLER_204_1525 ();
 sg13g2_fill_8 FILLER_204_1533 ();
 sg13g2_fill_8 FILLER_204_1541 ();
 sg13g2_fill_8 FILLER_204_1549 ();
 sg13g2_fill_8 FILLER_204_1557 ();
 sg13g2_fill_8 FILLER_204_1565 ();
 sg13g2_fill_8 FILLER_204_1573 ();
 sg13g2_fill_8 FILLER_204_1581 ();
 sg13g2_fill_2 FILLER_204_1589 ();
 sg13g2_fill_1 FILLER_204_1591 ();
 sg13g2_fill_8 FILLER_205_0 ();
 sg13g2_fill_8 FILLER_205_8 ();
 sg13g2_fill_8 FILLER_205_16 ();
 sg13g2_fill_8 FILLER_205_24 ();
 sg13g2_fill_8 FILLER_205_32 ();
 sg13g2_fill_8 FILLER_205_40 ();
 sg13g2_fill_8 FILLER_205_48 ();
 sg13g2_fill_8 FILLER_205_56 ();
 sg13g2_fill_8 FILLER_205_64 ();
 sg13g2_fill_8 FILLER_205_72 ();
 sg13g2_fill_8 FILLER_205_80 ();
 sg13g2_fill_8 FILLER_205_88 ();
 sg13g2_fill_8 FILLER_205_96 ();
 sg13g2_fill_8 FILLER_205_104 ();
 sg13g2_fill_8 FILLER_205_112 ();
 sg13g2_fill_8 FILLER_205_120 ();
 sg13g2_fill_8 FILLER_205_128 ();
 sg13g2_fill_8 FILLER_205_136 ();
 sg13g2_fill_8 FILLER_205_144 ();
 sg13g2_fill_8 FILLER_205_152 ();
 sg13g2_fill_8 FILLER_205_160 ();
 sg13g2_fill_8 FILLER_205_168 ();
 sg13g2_fill_8 FILLER_205_176 ();
 sg13g2_fill_8 FILLER_205_184 ();
 sg13g2_fill_8 FILLER_205_192 ();
 sg13g2_fill_8 FILLER_205_200 ();
 sg13g2_fill_8 FILLER_205_208 ();
 sg13g2_fill_8 FILLER_205_216 ();
 sg13g2_fill_8 FILLER_205_224 ();
 sg13g2_fill_8 FILLER_205_232 ();
 sg13g2_fill_8 FILLER_205_240 ();
 sg13g2_fill_8 FILLER_205_248 ();
 sg13g2_fill_8 FILLER_205_256 ();
 sg13g2_fill_8 FILLER_205_264 ();
 sg13g2_fill_8 FILLER_205_272 ();
 sg13g2_fill_8 FILLER_205_280 ();
 sg13g2_fill_8 FILLER_205_288 ();
 sg13g2_fill_8 FILLER_205_296 ();
 sg13g2_fill_8 FILLER_205_304 ();
 sg13g2_fill_8 FILLER_205_312 ();
 sg13g2_fill_8 FILLER_205_320 ();
 sg13g2_fill_8 FILLER_205_328 ();
 sg13g2_fill_8 FILLER_205_336 ();
 sg13g2_fill_8 FILLER_205_344 ();
 sg13g2_fill_8 FILLER_205_352 ();
 sg13g2_fill_8 FILLER_205_360 ();
 sg13g2_fill_8 FILLER_205_368 ();
 sg13g2_fill_8 FILLER_205_376 ();
 sg13g2_fill_8 FILLER_205_384 ();
 sg13g2_fill_8 FILLER_205_392 ();
 sg13g2_fill_8 FILLER_205_400 ();
 sg13g2_fill_8 FILLER_205_408 ();
 sg13g2_fill_8 FILLER_205_416 ();
 sg13g2_fill_8 FILLER_205_424 ();
 sg13g2_fill_8 FILLER_205_432 ();
 sg13g2_fill_8 FILLER_205_440 ();
 sg13g2_fill_8 FILLER_205_448 ();
 sg13g2_fill_8 FILLER_205_456 ();
 sg13g2_fill_8 FILLER_205_464 ();
 sg13g2_fill_8 FILLER_205_472 ();
 sg13g2_fill_8 FILLER_205_480 ();
 sg13g2_fill_8 FILLER_205_488 ();
 sg13g2_fill_8 FILLER_205_496 ();
 sg13g2_fill_8 FILLER_205_504 ();
 sg13g2_fill_8 FILLER_205_512 ();
 sg13g2_fill_8 FILLER_205_520 ();
 sg13g2_fill_8 FILLER_205_528 ();
 sg13g2_fill_8 FILLER_205_536 ();
 sg13g2_fill_8 FILLER_205_544 ();
 sg13g2_fill_8 FILLER_205_552 ();
 sg13g2_fill_8 FILLER_205_560 ();
 sg13g2_fill_8 FILLER_205_568 ();
 sg13g2_fill_8 FILLER_205_576 ();
 sg13g2_fill_8 FILLER_205_584 ();
 sg13g2_fill_8 FILLER_205_592 ();
 sg13g2_fill_8 FILLER_205_600 ();
 sg13g2_fill_8 FILLER_205_608 ();
 sg13g2_fill_8 FILLER_205_616 ();
 sg13g2_fill_8 FILLER_205_624 ();
 sg13g2_fill_8 FILLER_205_632 ();
 sg13g2_fill_8 FILLER_205_640 ();
 sg13g2_fill_8 FILLER_205_648 ();
 sg13g2_fill_8 FILLER_205_656 ();
 sg13g2_fill_8 FILLER_205_664 ();
 sg13g2_fill_8 FILLER_205_672 ();
 sg13g2_fill_8 FILLER_205_680 ();
 sg13g2_fill_8 FILLER_205_688 ();
 sg13g2_fill_8 FILLER_205_696 ();
 sg13g2_fill_8 FILLER_205_704 ();
 sg13g2_fill_8 FILLER_205_712 ();
 sg13g2_fill_8 FILLER_205_720 ();
 sg13g2_fill_8 FILLER_205_728 ();
 sg13g2_fill_8 FILLER_205_736 ();
 sg13g2_fill_8 FILLER_205_744 ();
 sg13g2_fill_8 FILLER_205_752 ();
 sg13g2_fill_8 FILLER_205_760 ();
 sg13g2_fill_8 FILLER_205_768 ();
 sg13g2_fill_8 FILLER_205_776 ();
 sg13g2_fill_8 FILLER_205_784 ();
 sg13g2_fill_8 FILLER_205_792 ();
 sg13g2_fill_8 FILLER_205_800 ();
 sg13g2_fill_8 FILLER_205_808 ();
 sg13g2_fill_8 FILLER_205_816 ();
 sg13g2_fill_8 FILLER_205_824 ();
 sg13g2_fill_8 FILLER_205_832 ();
 sg13g2_fill_8 FILLER_205_840 ();
 sg13g2_fill_8 FILLER_205_848 ();
 sg13g2_fill_8 FILLER_205_856 ();
 sg13g2_fill_8 FILLER_205_864 ();
 sg13g2_fill_8 FILLER_205_872 ();
 sg13g2_fill_8 FILLER_205_880 ();
 sg13g2_fill_8 FILLER_205_888 ();
 sg13g2_fill_8 FILLER_205_896 ();
 sg13g2_fill_8 FILLER_205_904 ();
 sg13g2_fill_8 FILLER_205_912 ();
 sg13g2_fill_8 FILLER_205_920 ();
 sg13g2_fill_8 FILLER_205_928 ();
 sg13g2_fill_8 FILLER_205_936 ();
 sg13g2_fill_8 FILLER_205_944 ();
 sg13g2_fill_8 FILLER_205_952 ();
 sg13g2_fill_8 FILLER_205_960 ();
 sg13g2_fill_8 FILLER_205_968 ();
 sg13g2_fill_8 FILLER_205_976 ();
 sg13g2_fill_8 FILLER_205_984 ();
 sg13g2_fill_8 FILLER_205_992 ();
 sg13g2_fill_8 FILLER_205_1000 ();
 sg13g2_fill_8 FILLER_205_1008 ();
 sg13g2_fill_8 FILLER_205_1016 ();
 sg13g2_fill_8 FILLER_205_1024 ();
 sg13g2_fill_8 FILLER_205_1032 ();
 sg13g2_fill_8 FILLER_205_1040 ();
 sg13g2_fill_8 FILLER_205_1048 ();
 sg13g2_fill_8 FILLER_205_1056 ();
 sg13g2_fill_8 FILLER_205_1064 ();
 sg13g2_fill_8 FILLER_205_1072 ();
 sg13g2_fill_8 FILLER_205_1080 ();
 sg13g2_fill_8 FILLER_205_1088 ();
 sg13g2_fill_8 FILLER_205_1096 ();
 sg13g2_fill_8 FILLER_205_1104 ();
 sg13g2_fill_8 FILLER_205_1112 ();
 sg13g2_fill_8 FILLER_205_1120 ();
 sg13g2_fill_8 FILLER_205_1128 ();
 sg13g2_fill_8 FILLER_205_1168 ();
 sg13g2_fill_8 FILLER_205_1176 ();
 sg13g2_fill_8 FILLER_205_1184 ();
 sg13g2_fill_8 FILLER_205_1200 ();
 sg13g2_fill_4 FILLER_205_1208 ();
 sg13g2_fill_2 FILLER_205_1212 ();
 sg13g2_fill_1 FILLER_205_1214 ();
 sg13g2_fill_2 FILLER_205_1231 ();
 sg13g2_fill_2 FILLER_205_1238 ();
 sg13g2_fill_2 FILLER_205_1244 ();
 sg13g2_fill_1 FILLER_205_1246 ();
 sg13g2_fill_8 FILLER_205_1269 ();
 sg13g2_fill_4 FILLER_205_1277 ();
 sg13g2_fill_2 FILLER_205_1281 ();
 sg13g2_fill_2 FILLER_205_1287 ();
 sg13g2_fill_8 FILLER_205_1329 ();
 sg13g2_fill_8 FILLER_205_1337 ();
 sg13g2_fill_8 FILLER_205_1345 ();
 sg13g2_fill_8 FILLER_205_1353 ();
 sg13g2_fill_8 FILLER_205_1361 ();
 sg13g2_fill_8 FILLER_205_1369 ();
 sg13g2_fill_8 FILLER_205_1377 ();
 sg13g2_fill_8 FILLER_205_1385 ();
 sg13g2_fill_8 FILLER_205_1393 ();
 sg13g2_fill_8 FILLER_205_1401 ();
 sg13g2_fill_8 FILLER_205_1409 ();
 sg13g2_fill_8 FILLER_205_1417 ();
 sg13g2_fill_8 FILLER_205_1425 ();
 sg13g2_fill_8 FILLER_205_1433 ();
 sg13g2_fill_8 FILLER_205_1441 ();
 sg13g2_fill_8 FILLER_205_1449 ();
 sg13g2_fill_8 FILLER_205_1457 ();
 sg13g2_fill_8 FILLER_205_1465 ();
 sg13g2_fill_8 FILLER_205_1473 ();
 sg13g2_fill_8 FILLER_205_1481 ();
 sg13g2_fill_8 FILLER_205_1489 ();
 sg13g2_fill_8 FILLER_205_1497 ();
 sg13g2_fill_8 FILLER_205_1505 ();
 sg13g2_fill_8 FILLER_205_1513 ();
 sg13g2_fill_8 FILLER_205_1521 ();
 sg13g2_fill_8 FILLER_205_1529 ();
 sg13g2_fill_8 FILLER_205_1537 ();
 sg13g2_fill_8 FILLER_205_1545 ();
 sg13g2_fill_8 FILLER_205_1553 ();
 sg13g2_fill_8 FILLER_205_1561 ();
 sg13g2_fill_8 FILLER_205_1569 ();
 sg13g2_fill_8 FILLER_205_1577 ();
 sg13g2_fill_4 FILLER_205_1585 ();
 sg13g2_fill_2 FILLER_205_1589 ();
 sg13g2_fill_1 FILLER_205_1591 ();
 sg13g2_fill_8 FILLER_206_0 ();
 sg13g2_fill_8 FILLER_206_8 ();
 sg13g2_fill_8 FILLER_206_16 ();
 sg13g2_fill_8 FILLER_206_24 ();
 sg13g2_fill_8 FILLER_206_32 ();
 sg13g2_fill_8 FILLER_206_40 ();
 sg13g2_fill_8 FILLER_206_48 ();
 sg13g2_fill_8 FILLER_206_56 ();
 sg13g2_fill_8 FILLER_206_64 ();
 sg13g2_fill_8 FILLER_206_72 ();
 sg13g2_fill_8 FILLER_206_80 ();
 sg13g2_fill_8 FILLER_206_88 ();
 sg13g2_fill_8 FILLER_206_96 ();
 sg13g2_fill_8 FILLER_206_104 ();
 sg13g2_fill_8 FILLER_206_112 ();
 sg13g2_fill_8 FILLER_206_120 ();
 sg13g2_fill_8 FILLER_206_128 ();
 sg13g2_fill_8 FILLER_206_136 ();
 sg13g2_fill_8 FILLER_206_144 ();
 sg13g2_fill_8 FILLER_206_152 ();
 sg13g2_fill_8 FILLER_206_160 ();
 sg13g2_fill_8 FILLER_206_168 ();
 sg13g2_fill_8 FILLER_206_176 ();
 sg13g2_fill_8 FILLER_206_184 ();
 sg13g2_fill_8 FILLER_206_192 ();
 sg13g2_fill_8 FILLER_206_200 ();
 sg13g2_fill_8 FILLER_206_208 ();
 sg13g2_fill_8 FILLER_206_216 ();
 sg13g2_fill_8 FILLER_206_224 ();
 sg13g2_fill_8 FILLER_206_232 ();
 sg13g2_fill_8 FILLER_206_240 ();
 sg13g2_fill_8 FILLER_206_248 ();
 sg13g2_fill_8 FILLER_206_256 ();
 sg13g2_fill_8 FILLER_206_264 ();
 sg13g2_fill_8 FILLER_206_272 ();
 sg13g2_fill_8 FILLER_206_280 ();
 sg13g2_fill_8 FILLER_206_288 ();
 sg13g2_fill_8 FILLER_206_296 ();
 sg13g2_fill_8 FILLER_206_304 ();
 sg13g2_fill_8 FILLER_206_312 ();
 sg13g2_fill_8 FILLER_206_320 ();
 sg13g2_fill_8 FILLER_206_328 ();
 sg13g2_fill_8 FILLER_206_336 ();
 sg13g2_fill_8 FILLER_206_344 ();
 sg13g2_fill_8 FILLER_206_352 ();
 sg13g2_fill_8 FILLER_206_360 ();
 sg13g2_fill_8 FILLER_206_368 ();
 sg13g2_fill_8 FILLER_206_376 ();
 sg13g2_fill_8 FILLER_206_384 ();
 sg13g2_fill_8 FILLER_206_392 ();
 sg13g2_fill_8 FILLER_206_400 ();
 sg13g2_fill_8 FILLER_206_408 ();
 sg13g2_fill_8 FILLER_206_416 ();
 sg13g2_fill_8 FILLER_206_424 ();
 sg13g2_fill_8 FILLER_206_432 ();
 sg13g2_fill_8 FILLER_206_440 ();
 sg13g2_fill_8 FILLER_206_448 ();
 sg13g2_fill_8 FILLER_206_456 ();
 sg13g2_fill_8 FILLER_206_464 ();
 sg13g2_fill_8 FILLER_206_472 ();
 sg13g2_fill_8 FILLER_206_480 ();
 sg13g2_fill_8 FILLER_206_488 ();
 sg13g2_fill_8 FILLER_206_496 ();
 sg13g2_fill_8 FILLER_206_504 ();
 sg13g2_fill_8 FILLER_206_512 ();
 sg13g2_fill_8 FILLER_206_520 ();
 sg13g2_fill_8 FILLER_206_528 ();
 sg13g2_fill_8 FILLER_206_536 ();
 sg13g2_fill_8 FILLER_206_544 ();
 sg13g2_fill_8 FILLER_206_552 ();
 sg13g2_fill_8 FILLER_206_560 ();
 sg13g2_fill_8 FILLER_206_568 ();
 sg13g2_fill_8 FILLER_206_576 ();
 sg13g2_fill_8 FILLER_206_584 ();
 sg13g2_fill_8 FILLER_206_592 ();
 sg13g2_fill_8 FILLER_206_600 ();
 sg13g2_fill_8 FILLER_206_608 ();
 sg13g2_fill_8 FILLER_206_616 ();
 sg13g2_fill_8 FILLER_206_624 ();
 sg13g2_fill_8 FILLER_206_632 ();
 sg13g2_fill_8 FILLER_206_640 ();
 sg13g2_fill_8 FILLER_206_648 ();
 sg13g2_fill_8 FILLER_206_656 ();
 sg13g2_fill_8 FILLER_206_664 ();
 sg13g2_fill_8 FILLER_206_672 ();
 sg13g2_fill_8 FILLER_206_680 ();
 sg13g2_fill_8 FILLER_206_688 ();
 sg13g2_fill_8 FILLER_206_696 ();
 sg13g2_fill_8 FILLER_206_704 ();
 sg13g2_fill_8 FILLER_206_712 ();
 sg13g2_fill_8 FILLER_206_720 ();
 sg13g2_fill_8 FILLER_206_728 ();
 sg13g2_fill_8 FILLER_206_736 ();
 sg13g2_fill_8 FILLER_206_744 ();
 sg13g2_fill_8 FILLER_206_752 ();
 sg13g2_fill_8 FILLER_206_760 ();
 sg13g2_fill_8 FILLER_206_768 ();
 sg13g2_fill_8 FILLER_206_776 ();
 sg13g2_fill_8 FILLER_206_784 ();
 sg13g2_fill_8 FILLER_206_792 ();
 sg13g2_fill_8 FILLER_206_800 ();
 sg13g2_fill_8 FILLER_206_808 ();
 sg13g2_fill_8 FILLER_206_816 ();
 sg13g2_fill_8 FILLER_206_824 ();
 sg13g2_fill_8 FILLER_206_832 ();
 sg13g2_fill_8 FILLER_206_840 ();
 sg13g2_fill_8 FILLER_206_848 ();
 sg13g2_fill_8 FILLER_206_856 ();
 sg13g2_fill_8 FILLER_206_864 ();
 sg13g2_fill_8 FILLER_206_872 ();
 sg13g2_fill_8 FILLER_206_880 ();
 sg13g2_fill_8 FILLER_206_888 ();
 sg13g2_fill_8 FILLER_206_896 ();
 sg13g2_fill_8 FILLER_206_904 ();
 sg13g2_fill_8 FILLER_206_912 ();
 sg13g2_fill_8 FILLER_206_920 ();
 sg13g2_fill_8 FILLER_206_928 ();
 sg13g2_fill_8 FILLER_206_936 ();
 sg13g2_fill_8 FILLER_206_944 ();
 sg13g2_fill_8 FILLER_206_952 ();
 sg13g2_fill_8 FILLER_206_960 ();
 sg13g2_fill_8 FILLER_206_968 ();
 sg13g2_fill_8 FILLER_206_976 ();
 sg13g2_fill_8 FILLER_206_984 ();
 sg13g2_fill_8 FILLER_206_992 ();
 sg13g2_fill_8 FILLER_206_1000 ();
 sg13g2_fill_8 FILLER_206_1008 ();
 sg13g2_fill_8 FILLER_206_1016 ();
 sg13g2_fill_8 FILLER_206_1024 ();
 sg13g2_fill_8 FILLER_206_1032 ();
 sg13g2_fill_8 FILLER_206_1040 ();
 sg13g2_fill_8 FILLER_206_1048 ();
 sg13g2_fill_8 FILLER_206_1056 ();
 sg13g2_fill_8 FILLER_206_1064 ();
 sg13g2_fill_8 FILLER_206_1072 ();
 sg13g2_fill_8 FILLER_206_1080 ();
 sg13g2_fill_8 FILLER_206_1088 ();
 sg13g2_fill_8 FILLER_206_1096 ();
 sg13g2_fill_8 FILLER_206_1104 ();
 sg13g2_fill_8 FILLER_206_1112 ();
 sg13g2_fill_8 FILLER_206_1120 ();
 sg13g2_fill_8 FILLER_206_1128 ();
 sg13g2_fill_4 FILLER_206_1136 ();
 sg13g2_fill_2 FILLER_206_1140 ();
 sg13g2_fill_1 FILLER_206_1150 ();
 sg13g2_fill_8 FILLER_206_1175 ();
 sg13g2_fill_4 FILLER_206_1183 ();
 sg13g2_fill_2 FILLER_206_1187 ();
 sg13g2_fill_8 FILLER_206_1194 ();
 sg13g2_fill_4 FILLER_206_1202 ();
 sg13g2_fill_8 FILLER_206_1232 ();
 sg13g2_fill_8 FILLER_206_1240 ();
 sg13g2_fill_4 FILLER_206_1248 ();
 sg13g2_fill_8 FILLER_206_1273 ();
 sg13g2_fill_8 FILLER_206_1281 ();
 sg13g2_fill_4 FILLER_206_1289 ();
 sg13g2_fill_2 FILLER_206_1293 ();
 sg13g2_fill_8 FILLER_206_1298 ();
 sg13g2_fill_8 FILLER_206_1306 ();
 sg13g2_fill_8 FILLER_206_1314 ();
 sg13g2_fill_8 FILLER_206_1322 ();
 sg13g2_fill_8 FILLER_206_1330 ();
 sg13g2_fill_8 FILLER_206_1338 ();
 sg13g2_fill_8 FILLER_206_1346 ();
 sg13g2_fill_8 FILLER_206_1354 ();
 sg13g2_fill_8 FILLER_206_1362 ();
 sg13g2_fill_8 FILLER_206_1370 ();
 sg13g2_fill_8 FILLER_206_1378 ();
 sg13g2_fill_8 FILLER_206_1386 ();
 sg13g2_fill_8 FILLER_206_1394 ();
 sg13g2_fill_8 FILLER_206_1402 ();
 sg13g2_fill_8 FILLER_206_1410 ();
 sg13g2_fill_8 FILLER_206_1418 ();
 sg13g2_fill_8 FILLER_206_1426 ();
 sg13g2_fill_8 FILLER_206_1434 ();
 sg13g2_fill_8 FILLER_206_1442 ();
 sg13g2_fill_8 FILLER_206_1450 ();
 sg13g2_fill_8 FILLER_206_1458 ();
 sg13g2_fill_8 FILLER_206_1466 ();
 sg13g2_fill_8 FILLER_206_1474 ();
 sg13g2_fill_8 FILLER_206_1482 ();
 sg13g2_fill_8 FILLER_206_1490 ();
 sg13g2_fill_8 FILLER_206_1498 ();
 sg13g2_fill_8 FILLER_206_1506 ();
 sg13g2_fill_8 FILLER_206_1514 ();
 sg13g2_fill_8 FILLER_206_1522 ();
 sg13g2_fill_8 FILLER_206_1530 ();
 sg13g2_fill_8 FILLER_206_1538 ();
 sg13g2_fill_8 FILLER_206_1546 ();
 sg13g2_fill_8 FILLER_206_1554 ();
 sg13g2_fill_8 FILLER_206_1562 ();
 sg13g2_fill_8 FILLER_206_1570 ();
 sg13g2_fill_8 FILLER_206_1578 ();
 sg13g2_fill_4 FILLER_206_1586 ();
 sg13g2_fill_2 FILLER_206_1590 ();
 sg13g2_fill_8 FILLER_207_0 ();
 sg13g2_fill_8 FILLER_207_8 ();
 sg13g2_fill_8 FILLER_207_16 ();
 sg13g2_fill_8 FILLER_207_24 ();
 sg13g2_fill_8 FILLER_207_32 ();
 sg13g2_fill_8 FILLER_207_40 ();
 sg13g2_fill_8 FILLER_207_48 ();
 sg13g2_fill_8 FILLER_207_56 ();
 sg13g2_fill_8 FILLER_207_64 ();
 sg13g2_fill_8 FILLER_207_72 ();
 sg13g2_fill_8 FILLER_207_80 ();
 sg13g2_fill_8 FILLER_207_88 ();
 sg13g2_fill_8 FILLER_207_96 ();
 sg13g2_fill_8 FILLER_207_104 ();
 sg13g2_fill_8 FILLER_207_112 ();
 sg13g2_fill_8 FILLER_207_120 ();
 sg13g2_fill_8 FILLER_207_128 ();
 sg13g2_fill_8 FILLER_207_136 ();
 sg13g2_fill_8 FILLER_207_144 ();
 sg13g2_fill_8 FILLER_207_152 ();
 sg13g2_fill_8 FILLER_207_160 ();
 sg13g2_fill_8 FILLER_207_168 ();
 sg13g2_fill_8 FILLER_207_176 ();
 sg13g2_fill_8 FILLER_207_184 ();
 sg13g2_fill_8 FILLER_207_192 ();
 sg13g2_fill_8 FILLER_207_200 ();
 sg13g2_fill_8 FILLER_207_208 ();
 sg13g2_fill_8 FILLER_207_216 ();
 sg13g2_fill_8 FILLER_207_224 ();
 sg13g2_fill_8 FILLER_207_232 ();
 sg13g2_fill_8 FILLER_207_240 ();
 sg13g2_fill_8 FILLER_207_248 ();
 sg13g2_fill_8 FILLER_207_256 ();
 sg13g2_fill_8 FILLER_207_264 ();
 sg13g2_fill_8 FILLER_207_272 ();
 sg13g2_fill_8 FILLER_207_280 ();
 sg13g2_fill_8 FILLER_207_288 ();
 sg13g2_fill_8 FILLER_207_296 ();
 sg13g2_fill_8 FILLER_207_304 ();
 sg13g2_fill_8 FILLER_207_312 ();
 sg13g2_fill_8 FILLER_207_320 ();
 sg13g2_fill_8 FILLER_207_328 ();
 sg13g2_fill_8 FILLER_207_336 ();
 sg13g2_fill_8 FILLER_207_344 ();
 sg13g2_fill_8 FILLER_207_352 ();
 sg13g2_fill_8 FILLER_207_360 ();
 sg13g2_fill_8 FILLER_207_368 ();
 sg13g2_fill_8 FILLER_207_376 ();
 sg13g2_fill_8 FILLER_207_384 ();
 sg13g2_fill_8 FILLER_207_392 ();
 sg13g2_fill_8 FILLER_207_400 ();
 sg13g2_fill_8 FILLER_207_408 ();
 sg13g2_fill_8 FILLER_207_416 ();
 sg13g2_fill_8 FILLER_207_424 ();
 sg13g2_fill_8 FILLER_207_432 ();
 sg13g2_fill_8 FILLER_207_440 ();
 sg13g2_fill_8 FILLER_207_448 ();
 sg13g2_fill_8 FILLER_207_456 ();
 sg13g2_fill_8 FILLER_207_464 ();
 sg13g2_fill_8 FILLER_207_472 ();
 sg13g2_fill_8 FILLER_207_480 ();
 sg13g2_fill_8 FILLER_207_488 ();
 sg13g2_fill_8 FILLER_207_496 ();
 sg13g2_fill_8 FILLER_207_504 ();
 sg13g2_fill_8 FILLER_207_512 ();
 sg13g2_fill_8 FILLER_207_520 ();
 sg13g2_fill_8 FILLER_207_528 ();
 sg13g2_fill_8 FILLER_207_536 ();
 sg13g2_fill_8 FILLER_207_544 ();
 sg13g2_fill_8 FILLER_207_552 ();
 sg13g2_fill_8 FILLER_207_560 ();
 sg13g2_fill_8 FILLER_207_568 ();
 sg13g2_fill_8 FILLER_207_576 ();
 sg13g2_fill_8 FILLER_207_584 ();
 sg13g2_fill_8 FILLER_207_592 ();
 sg13g2_fill_8 FILLER_207_600 ();
 sg13g2_fill_8 FILLER_207_608 ();
 sg13g2_fill_8 FILLER_207_616 ();
 sg13g2_fill_8 FILLER_207_624 ();
 sg13g2_fill_8 FILLER_207_632 ();
 sg13g2_fill_8 FILLER_207_640 ();
 sg13g2_fill_8 FILLER_207_648 ();
 sg13g2_fill_8 FILLER_207_656 ();
 sg13g2_fill_8 FILLER_207_664 ();
 sg13g2_fill_8 FILLER_207_672 ();
 sg13g2_fill_8 FILLER_207_680 ();
 sg13g2_fill_8 FILLER_207_688 ();
 sg13g2_fill_8 FILLER_207_696 ();
 sg13g2_fill_8 FILLER_207_704 ();
 sg13g2_fill_8 FILLER_207_712 ();
 sg13g2_fill_8 FILLER_207_720 ();
 sg13g2_fill_8 FILLER_207_728 ();
 sg13g2_fill_8 FILLER_207_736 ();
 sg13g2_fill_8 FILLER_207_744 ();
 sg13g2_fill_8 FILLER_207_752 ();
 sg13g2_fill_8 FILLER_207_760 ();
 sg13g2_fill_8 FILLER_207_768 ();
 sg13g2_fill_8 FILLER_207_776 ();
 sg13g2_fill_8 FILLER_207_784 ();
 sg13g2_fill_8 FILLER_207_792 ();
 sg13g2_fill_8 FILLER_207_800 ();
 sg13g2_fill_8 FILLER_207_808 ();
 sg13g2_fill_8 FILLER_207_816 ();
 sg13g2_fill_8 FILLER_207_824 ();
 sg13g2_fill_8 FILLER_207_832 ();
 sg13g2_fill_8 FILLER_207_840 ();
 sg13g2_fill_8 FILLER_207_848 ();
 sg13g2_fill_8 FILLER_207_856 ();
 sg13g2_fill_8 FILLER_207_864 ();
 sg13g2_fill_8 FILLER_207_872 ();
 sg13g2_fill_8 FILLER_207_880 ();
 sg13g2_fill_8 FILLER_207_888 ();
 sg13g2_fill_8 FILLER_207_896 ();
 sg13g2_fill_8 FILLER_207_904 ();
 sg13g2_fill_8 FILLER_207_912 ();
 sg13g2_fill_8 FILLER_207_920 ();
 sg13g2_fill_8 FILLER_207_928 ();
 sg13g2_fill_8 FILLER_207_936 ();
 sg13g2_fill_8 FILLER_207_944 ();
 sg13g2_fill_8 FILLER_207_952 ();
 sg13g2_fill_8 FILLER_207_960 ();
 sg13g2_fill_8 FILLER_207_968 ();
 sg13g2_fill_8 FILLER_207_976 ();
 sg13g2_fill_8 FILLER_207_984 ();
 sg13g2_fill_8 FILLER_207_992 ();
 sg13g2_fill_8 FILLER_207_1000 ();
 sg13g2_fill_8 FILLER_207_1008 ();
 sg13g2_fill_8 FILLER_207_1016 ();
 sg13g2_fill_8 FILLER_207_1024 ();
 sg13g2_fill_8 FILLER_207_1032 ();
 sg13g2_fill_8 FILLER_207_1040 ();
 sg13g2_fill_8 FILLER_207_1048 ();
 sg13g2_fill_8 FILLER_207_1056 ();
 sg13g2_fill_8 FILLER_207_1064 ();
 sg13g2_fill_8 FILLER_207_1072 ();
 sg13g2_fill_8 FILLER_207_1080 ();
 sg13g2_fill_8 FILLER_207_1088 ();
 sg13g2_fill_8 FILLER_207_1096 ();
 sg13g2_fill_8 FILLER_207_1104 ();
 sg13g2_fill_8 FILLER_207_1112 ();
 sg13g2_fill_8 FILLER_207_1120 ();
 sg13g2_fill_8 FILLER_207_1128 ();
 sg13g2_fill_8 FILLER_207_1136 ();
 sg13g2_fill_8 FILLER_207_1144 ();
 sg13g2_fill_8 FILLER_207_1152 ();
 sg13g2_fill_8 FILLER_207_1160 ();
 sg13g2_fill_4 FILLER_207_1168 ();
 sg13g2_fill_2 FILLER_207_1172 ();
 sg13g2_fill_1 FILLER_207_1174 ();
 sg13g2_fill_1 FILLER_207_1178 ();
 sg13g2_fill_1 FILLER_207_1184 ();
 sg13g2_fill_4 FILLER_207_1203 ();
 sg13g2_fill_2 FILLER_207_1207 ();
 sg13g2_fill_4 FILLER_207_1213 ();
 sg13g2_fill_2 FILLER_207_1217 ();
 sg13g2_fill_8 FILLER_207_1231 ();
 sg13g2_fill_8 FILLER_207_1239 ();
 sg13g2_fill_8 FILLER_207_1247 ();
 sg13g2_fill_8 FILLER_207_1255 ();
 sg13g2_fill_4 FILLER_207_1263 ();
 sg13g2_fill_2 FILLER_207_1267 ();
 sg13g2_fill_1 FILLER_207_1273 ();
 sg13g2_fill_8 FILLER_207_1285 ();
 sg13g2_fill_2 FILLER_207_1301 ();
 sg13g2_fill_8 FILLER_207_1313 ();
 sg13g2_fill_8 FILLER_207_1321 ();
 sg13g2_fill_8 FILLER_207_1329 ();
 sg13g2_fill_8 FILLER_207_1337 ();
 sg13g2_fill_8 FILLER_207_1345 ();
 sg13g2_fill_8 FILLER_207_1353 ();
 sg13g2_fill_8 FILLER_207_1361 ();
 sg13g2_fill_8 FILLER_207_1369 ();
 sg13g2_fill_8 FILLER_207_1377 ();
 sg13g2_fill_8 FILLER_207_1385 ();
 sg13g2_fill_8 FILLER_207_1393 ();
 sg13g2_fill_8 FILLER_207_1401 ();
 sg13g2_fill_8 FILLER_207_1409 ();
 sg13g2_fill_8 FILLER_207_1417 ();
 sg13g2_fill_8 FILLER_207_1425 ();
 sg13g2_fill_8 FILLER_207_1433 ();
 sg13g2_fill_8 FILLER_207_1441 ();
 sg13g2_fill_8 FILLER_207_1449 ();
 sg13g2_fill_8 FILLER_207_1457 ();
 sg13g2_fill_8 FILLER_207_1465 ();
 sg13g2_fill_8 FILLER_207_1473 ();
 sg13g2_fill_8 FILLER_207_1481 ();
 sg13g2_fill_8 FILLER_207_1489 ();
 sg13g2_fill_8 FILLER_207_1497 ();
 sg13g2_fill_8 FILLER_207_1505 ();
 sg13g2_fill_8 FILLER_207_1513 ();
 sg13g2_fill_8 FILLER_207_1521 ();
 sg13g2_fill_8 FILLER_207_1529 ();
 sg13g2_fill_8 FILLER_207_1537 ();
 sg13g2_fill_8 FILLER_207_1545 ();
 sg13g2_fill_8 FILLER_207_1553 ();
 sg13g2_fill_8 FILLER_207_1561 ();
 sg13g2_fill_8 FILLER_207_1569 ();
 sg13g2_fill_8 FILLER_207_1577 ();
 sg13g2_fill_4 FILLER_207_1585 ();
 sg13g2_fill_2 FILLER_207_1589 ();
 sg13g2_fill_1 FILLER_207_1591 ();
 sg13g2_fill_8 FILLER_208_0 ();
 sg13g2_fill_8 FILLER_208_8 ();
 sg13g2_fill_8 FILLER_208_16 ();
 sg13g2_fill_8 FILLER_208_24 ();
 sg13g2_fill_8 FILLER_208_32 ();
 sg13g2_fill_8 FILLER_208_40 ();
 sg13g2_fill_8 FILLER_208_48 ();
 sg13g2_fill_8 FILLER_208_56 ();
 sg13g2_fill_8 FILLER_208_64 ();
 sg13g2_fill_8 FILLER_208_72 ();
 sg13g2_fill_8 FILLER_208_80 ();
 sg13g2_fill_8 FILLER_208_88 ();
 sg13g2_fill_8 FILLER_208_96 ();
 sg13g2_fill_8 FILLER_208_104 ();
 sg13g2_fill_8 FILLER_208_112 ();
 sg13g2_fill_8 FILLER_208_120 ();
 sg13g2_fill_8 FILLER_208_128 ();
 sg13g2_fill_8 FILLER_208_136 ();
 sg13g2_fill_8 FILLER_208_144 ();
 sg13g2_fill_8 FILLER_208_152 ();
 sg13g2_fill_8 FILLER_208_160 ();
 sg13g2_fill_8 FILLER_208_168 ();
 sg13g2_fill_8 FILLER_208_176 ();
 sg13g2_fill_8 FILLER_208_184 ();
 sg13g2_fill_8 FILLER_208_192 ();
 sg13g2_fill_8 FILLER_208_200 ();
 sg13g2_fill_8 FILLER_208_208 ();
 sg13g2_fill_8 FILLER_208_216 ();
 sg13g2_fill_8 FILLER_208_224 ();
 sg13g2_fill_8 FILLER_208_232 ();
 sg13g2_fill_8 FILLER_208_240 ();
 sg13g2_fill_8 FILLER_208_248 ();
 sg13g2_fill_8 FILLER_208_256 ();
 sg13g2_fill_8 FILLER_208_264 ();
 sg13g2_fill_8 FILLER_208_272 ();
 sg13g2_fill_8 FILLER_208_280 ();
 sg13g2_fill_8 FILLER_208_288 ();
 sg13g2_fill_8 FILLER_208_296 ();
 sg13g2_fill_8 FILLER_208_304 ();
 sg13g2_fill_8 FILLER_208_312 ();
 sg13g2_fill_8 FILLER_208_320 ();
 sg13g2_fill_8 FILLER_208_328 ();
 sg13g2_fill_8 FILLER_208_336 ();
 sg13g2_fill_8 FILLER_208_344 ();
 sg13g2_fill_8 FILLER_208_352 ();
 sg13g2_fill_8 FILLER_208_360 ();
 sg13g2_fill_8 FILLER_208_368 ();
 sg13g2_fill_8 FILLER_208_376 ();
 sg13g2_fill_8 FILLER_208_384 ();
 sg13g2_fill_8 FILLER_208_392 ();
 sg13g2_fill_8 FILLER_208_400 ();
 sg13g2_fill_8 FILLER_208_408 ();
 sg13g2_fill_8 FILLER_208_416 ();
 sg13g2_fill_8 FILLER_208_424 ();
 sg13g2_fill_8 FILLER_208_432 ();
 sg13g2_fill_8 FILLER_208_440 ();
 sg13g2_fill_8 FILLER_208_448 ();
 sg13g2_fill_8 FILLER_208_456 ();
 sg13g2_fill_8 FILLER_208_464 ();
 sg13g2_fill_8 FILLER_208_472 ();
 sg13g2_fill_8 FILLER_208_480 ();
 sg13g2_fill_8 FILLER_208_488 ();
 sg13g2_fill_8 FILLER_208_496 ();
 sg13g2_fill_8 FILLER_208_504 ();
 sg13g2_fill_8 FILLER_208_512 ();
 sg13g2_fill_8 FILLER_208_520 ();
 sg13g2_fill_8 FILLER_208_528 ();
 sg13g2_fill_8 FILLER_208_536 ();
 sg13g2_fill_8 FILLER_208_544 ();
 sg13g2_fill_8 FILLER_208_552 ();
 sg13g2_fill_8 FILLER_208_560 ();
 sg13g2_fill_8 FILLER_208_568 ();
 sg13g2_fill_8 FILLER_208_576 ();
 sg13g2_fill_8 FILLER_208_584 ();
 sg13g2_fill_8 FILLER_208_592 ();
 sg13g2_fill_8 FILLER_208_600 ();
 sg13g2_fill_8 FILLER_208_608 ();
 sg13g2_fill_8 FILLER_208_616 ();
 sg13g2_fill_8 FILLER_208_624 ();
 sg13g2_fill_8 FILLER_208_632 ();
 sg13g2_fill_8 FILLER_208_640 ();
 sg13g2_fill_8 FILLER_208_648 ();
 sg13g2_fill_8 FILLER_208_656 ();
 sg13g2_fill_8 FILLER_208_664 ();
 sg13g2_fill_8 FILLER_208_672 ();
 sg13g2_fill_8 FILLER_208_680 ();
 sg13g2_fill_8 FILLER_208_688 ();
 sg13g2_fill_8 FILLER_208_696 ();
 sg13g2_fill_8 FILLER_208_704 ();
 sg13g2_fill_8 FILLER_208_712 ();
 sg13g2_fill_8 FILLER_208_720 ();
 sg13g2_fill_8 FILLER_208_728 ();
 sg13g2_fill_8 FILLER_208_736 ();
 sg13g2_fill_8 FILLER_208_744 ();
 sg13g2_fill_8 FILLER_208_752 ();
 sg13g2_fill_8 FILLER_208_760 ();
 sg13g2_fill_8 FILLER_208_768 ();
 sg13g2_fill_8 FILLER_208_776 ();
 sg13g2_fill_8 FILLER_208_784 ();
 sg13g2_fill_8 FILLER_208_792 ();
 sg13g2_fill_8 FILLER_208_800 ();
 sg13g2_fill_8 FILLER_208_808 ();
 sg13g2_fill_8 FILLER_208_816 ();
 sg13g2_fill_8 FILLER_208_824 ();
 sg13g2_fill_8 FILLER_208_832 ();
 sg13g2_fill_8 FILLER_208_840 ();
 sg13g2_fill_8 FILLER_208_848 ();
 sg13g2_fill_8 FILLER_208_856 ();
 sg13g2_fill_8 FILLER_208_864 ();
 sg13g2_fill_8 FILLER_208_872 ();
 sg13g2_fill_8 FILLER_208_880 ();
 sg13g2_fill_8 FILLER_208_888 ();
 sg13g2_fill_8 FILLER_208_896 ();
 sg13g2_fill_8 FILLER_208_904 ();
 sg13g2_fill_8 FILLER_208_912 ();
 sg13g2_fill_8 FILLER_208_920 ();
 sg13g2_fill_8 FILLER_208_928 ();
 sg13g2_fill_8 FILLER_208_936 ();
 sg13g2_fill_8 FILLER_208_944 ();
 sg13g2_fill_8 FILLER_208_952 ();
 sg13g2_fill_8 FILLER_208_960 ();
 sg13g2_fill_8 FILLER_208_968 ();
 sg13g2_fill_8 FILLER_208_976 ();
 sg13g2_fill_8 FILLER_208_984 ();
 sg13g2_fill_8 FILLER_208_992 ();
 sg13g2_fill_8 FILLER_208_1000 ();
 sg13g2_fill_8 FILLER_208_1008 ();
 sg13g2_fill_8 FILLER_208_1016 ();
 sg13g2_fill_8 FILLER_208_1024 ();
 sg13g2_fill_8 FILLER_208_1032 ();
 sg13g2_fill_8 FILLER_208_1040 ();
 sg13g2_fill_8 FILLER_208_1048 ();
 sg13g2_fill_8 FILLER_208_1056 ();
 sg13g2_fill_8 FILLER_208_1064 ();
 sg13g2_fill_8 FILLER_208_1072 ();
 sg13g2_fill_8 FILLER_208_1080 ();
 sg13g2_fill_8 FILLER_208_1088 ();
 sg13g2_fill_8 FILLER_208_1096 ();
 sg13g2_fill_8 FILLER_208_1104 ();
 sg13g2_fill_8 FILLER_208_1112 ();
 sg13g2_fill_8 FILLER_208_1120 ();
 sg13g2_fill_8 FILLER_208_1128 ();
 sg13g2_fill_8 FILLER_208_1136 ();
 sg13g2_fill_8 FILLER_208_1144 ();
 sg13g2_fill_8 FILLER_208_1152 ();
 sg13g2_fill_4 FILLER_208_1160 ();
 sg13g2_fill_2 FILLER_208_1164 ();
 sg13g2_fill_2 FILLER_208_1174 ();
 sg13g2_fill_1 FILLER_208_1192 ();
 sg13g2_fill_8 FILLER_208_1201 ();
 sg13g2_fill_8 FILLER_208_1212 ();
 sg13g2_fill_8 FILLER_208_1220 ();
 sg13g2_fill_1 FILLER_208_1228 ();
 sg13g2_fill_4 FILLER_208_1237 ();
 sg13g2_fill_2 FILLER_208_1241 ();
 sg13g2_fill_2 FILLER_208_1251 ();
 sg13g2_fill_2 FILLER_208_1256 ();
 sg13g2_fill_1 FILLER_208_1264 ();
 sg13g2_fill_1 FILLER_208_1274 ();
 sg13g2_fill_4 FILLER_208_1286 ();
 sg13g2_fill_8 FILLER_208_1324 ();
 sg13g2_fill_8 FILLER_208_1332 ();
 sg13g2_fill_8 FILLER_208_1340 ();
 sg13g2_fill_8 FILLER_208_1348 ();
 sg13g2_fill_8 FILLER_208_1356 ();
 sg13g2_fill_8 FILLER_208_1364 ();
 sg13g2_fill_8 FILLER_208_1372 ();
 sg13g2_fill_8 FILLER_208_1380 ();
 sg13g2_fill_8 FILLER_208_1388 ();
 sg13g2_fill_8 FILLER_208_1396 ();
 sg13g2_fill_8 FILLER_208_1404 ();
 sg13g2_fill_8 FILLER_208_1412 ();
 sg13g2_fill_8 FILLER_208_1420 ();
 sg13g2_fill_8 FILLER_208_1428 ();
 sg13g2_fill_8 FILLER_208_1436 ();
 sg13g2_fill_8 FILLER_208_1444 ();
 sg13g2_fill_8 FILLER_208_1452 ();
 sg13g2_fill_8 FILLER_208_1460 ();
 sg13g2_fill_8 FILLER_208_1468 ();
 sg13g2_fill_8 FILLER_208_1476 ();
 sg13g2_fill_8 FILLER_208_1484 ();
 sg13g2_fill_8 FILLER_208_1492 ();
 sg13g2_fill_8 FILLER_208_1500 ();
 sg13g2_fill_8 FILLER_208_1508 ();
 sg13g2_fill_8 FILLER_208_1516 ();
 sg13g2_fill_8 FILLER_208_1524 ();
 sg13g2_fill_8 FILLER_208_1532 ();
 sg13g2_fill_8 FILLER_208_1540 ();
 sg13g2_fill_8 FILLER_208_1548 ();
 sg13g2_fill_8 FILLER_208_1556 ();
 sg13g2_fill_8 FILLER_208_1564 ();
 sg13g2_fill_8 FILLER_208_1572 ();
 sg13g2_fill_8 FILLER_208_1580 ();
 sg13g2_fill_4 FILLER_208_1588 ();
 sg13g2_fill_8 FILLER_209_0 ();
 sg13g2_fill_8 FILLER_209_8 ();
 sg13g2_fill_8 FILLER_209_16 ();
 sg13g2_fill_8 FILLER_209_24 ();
 sg13g2_fill_8 FILLER_209_32 ();
 sg13g2_fill_8 FILLER_209_40 ();
 sg13g2_fill_8 FILLER_209_48 ();
 sg13g2_fill_8 FILLER_209_56 ();
 sg13g2_fill_8 FILLER_209_64 ();
 sg13g2_fill_8 FILLER_209_72 ();
 sg13g2_fill_8 FILLER_209_80 ();
 sg13g2_fill_8 FILLER_209_88 ();
 sg13g2_fill_8 FILLER_209_96 ();
 sg13g2_fill_8 FILLER_209_104 ();
 sg13g2_fill_8 FILLER_209_112 ();
 sg13g2_fill_8 FILLER_209_120 ();
 sg13g2_fill_8 FILLER_209_128 ();
 sg13g2_fill_8 FILLER_209_136 ();
 sg13g2_fill_8 FILLER_209_144 ();
 sg13g2_fill_8 FILLER_209_152 ();
 sg13g2_fill_8 FILLER_209_160 ();
 sg13g2_fill_8 FILLER_209_168 ();
 sg13g2_fill_8 FILLER_209_176 ();
 sg13g2_fill_8 FILLER_209_184 ();
 sg13g2_fill_8 FILLER_209_192 ();
 sg13g2_fill_8 FILLER_209_200 ();
 sg13g2_fill_8 FILLER_209_208 ();
 sg13g2_fill_8 FILLER_209_216 ();
 sg13g2_fill_8 FILLER_209_224 ();
 sg13g2_fill_8 FILLER_209_232 ();
 sg13g2_fill_8 FILLER_209_240 ();
 sg13g2_fill_8 FILLER_209_248 ();
 sg13g2_fill_8 FILLER_209_256 ();
 sg13g2_fill_8 FILLER_209_264 ();
 sg13g2_fill_8 FILLER_209_272 ();
 sg13g2_fill_8 FILLER_209_280 ();
 sg13g2_fill_8 FILLER_209_288 ();
 sg13g2_fill_8 FILLER_209_296 ();
 sg13g2_fill_8 FILLER_209_304 ();
 sg13g2_fill_8 FILLER_209_312 ();
 sg13g2_fill_8 FILLER_209_320 ();
 sg13g2_fill_8 FILLER_209_328 ();
 sg13g2_fill_8 FILLER_209_336 ();
 sg13g2_fill_8 FILLER_209_344 ();
 sg13g2_fill_8 FILLER_209_352 ();
 sg13g2_fill_8 FILLER_209_360 ();
 sg13g2_fill_8 FILLER_209_368 ();
 sg13g2_fill_8 FILLER_209_376 ();
 sg13g2_fill_8 FILLER_209_384 ();
 sg13g2_fill_8 FILLER_209_392 ();
 sg13g2_fill_8 FILLER_209_400 ();
 sg13g2_fill_8 FILLER_209_408 ();
 sg13g2_fill_8 FILLER_209_416 ();
 sg13g2_fill_8 FILLER_209_424 ();
 sg13g2_fill_8 FILLER_209_432 ();
 sg13g2_fill_8 FILLER_209_440 ();
 sg13g2_fill_8 FILLER_209_448 ();
 sg13g2_fill_8 FILLER_209_456 ();
 sg13g2_fill_8 FILLER_209_464 ();
 sg13g2_fill_8 FILLER_209_472 ();
 sg13g2_fill_8 FILLER_209_480 ();
 sg13g2_fill_8 FILLER_209_488 ();
 sg13g2_fill_8 FILLER_209_496 ();
 sg13g2_fill_8 FILLER_209_504 ();
 sg13g2_fill_8 FILLER_209_512 ();
 sg13g2_fill_8 FILLER_209_520 ();
 sg13g2_fill_8 FILLER_209_528 ();
 sg13g2_fill_8 FILLER_209_536 ();
 sg13g2_fill_8 FILLER_209_544 ();
 sg13g2_fill_8 FILLER_209_552 ();
 sg13g2_fill_8 FILLER_209_560 ();
 sg13g2_fill_8 FILLER_209_568 ();
 sg13g2_fill_8 FILLER_209_576 ();
 sg13g2_fill_8 FILLER_209_584 ();
 sg13g2_fill_8 FILLER_209_592 ();
 sg13g2_fill_8 FILLER_209_600 ();
 sg13g2_fill_8 FILLER_209_608 ();
 sg13g2_fill_8 FILLER_209_616 ();
 sg13g2_fill_8 FILLER_209_624 ();
 sg13g2_fill_8 FILLER_209_632 ();
 sg13g2_fill_8 FILLER_209_640 ();
 sg13g2_fill_8 FILLER_209_648 ();
 sg13g2_fill_8 FILLER_209_656 ();
 sg13g2_fill_8 FILLER_209_664 ();
 sg13g2_fill_8 FILLER_209_672 ();
 sg13g2_fill_8 FILLER_209_680 ();
 sg13g2_fill_8 FILLER_209_688 ();
 sg13g2_fill_8 FILLER_209_696 ();
 sg13g2_fill_8 FILLER_209_704 ();
 sg13g2_fill_8 FILLER_209_712 ();
 sg13g2_fill_8 FILLER_209_720 ();
 sg13g2_fill_8 FILLER_209_728 ();
 sg13g2_fill_8 FILLER_209_736 ();
 sg13g2_fill_8 FILLER_209_744 ();
 sg13g2_fill_8 FILLER_209_752 ();
 sg13g2_fill_8 FILLER_209_760 ();
 sg13g2_fill_8 FILLER_209_768 ();
 sg13g2_fill_8 FILLER_209_776 ();
 sg13g2_fill_8 FILLER_209_784 ();
 sg13g2_fill_8 FILLER_209_792 ();
 sg13g2_fill_8 FILLER_209_800 ();
 sg13g2_fill_8 FILLER_209_808 ();
 sg13g2_fill_8 FILLER_209_816 ();
 sg13g2_fill_8 FILLER_209_824 ();
 sg13g2_fill_8 FILLER_209_832 ();
 sg13g2_fill_8 FILLER_209_840 ();
 sg13g2_fill_8 FILLER_209_848 ();
 sg13g2_fill_8 FILLER_209_856 ();
 sg13g2_fill_8 FILLER_209_864 ();
 sg13g2_fill_8 FILLER_209_872 ();
 sg13g2_fill_8 FILLER_209_880 ();
 sg13g2_fill_8 FILLER_209_888 ();
 sg13g2_fill_8 FILLER_209_896 ();
 sg13g2_fill_8 FILLER_209_904 ();
 sg13g2_fill_8 FILLER_209_912 ();
 sg13g2_fill_8 FILLER_209_920 ();
 sg13g2_fill_8 FILLER_209_928 ();
 sg13g2_fill_8 FILLER_209_936 ();
 sg13g2_fill_8 FILLER_209_944 ();
 sg13g2_fill_8 FILLER_209_952 ();
 sg13g2_fill_8 FILLER_209_960 ();
 sg13g2_fill_8 FILLER_209_968 ();
 sg13g2_fill_8 FILLER_209_976 ();
 sg13g2_fill_8 FILLER_209_984 ();
 sg13g2_fill_8 FILLER_209_992 ();
 sg13g2_fill_8 FILLER_209_1000 ();
 sg13g2_fill_8 FILLER_209_1008 ();
 sg13g2_fill_8 FILLER_209_1016 ();
 sg13g2_fill_8 FILLER_209_1024 ();
 sg13g2_fill_8 FILLER_209_1032 ();
 sg13g2_fill_8 FILLER_209_1040 ();
 sg13g2_fill_8 FILLER_209_1048 ();
 sg13g2_fill_8 FILLER_209_1056 ();
 sg13g2_fill_8 FILLER_209_1064 ();
 sg13g2_fill_8 FILLER_209_1072 ();
 sg13g2_fill_8 FILLER_209_1080 ();
 sg13g2_fill_8 FILLER_209_1088 ();
 sg13g2_fill_8 FILLER_209_1096 ();
 sg13g2_fill_8 FILLER_209_1104 ();
 sg13g2_fill_8 FILLER_209_1112 ();
 sg13g2_fill_8 FILLER_209_1120 ();
 sg13g2_fill_8 FILLER_209_1128 ();
 sg13g2_fill_8 FILLER_209_1136 ();
 sg13g2_fill_8 FILLER_209_1144 ();
 sg13g2_fill_4 FILLER_209_1152 ();
 sg13g2_fill_1 FILLER_209_1156 ();
 sg13g2_fill_8 FILLER_209_1173 ();
 sg13g2_fill_4 FILLER_209_1181 ();
 sg13g2_fill_8 FILLER_209_1190 ();
 sg13g2_fill_4 FILLER_209_1198 ();
 sg13g2_fill_1 FILLER_209_1279 ();
 sg13g2_fill_8 FILLER_209_1326 ();
 sg13g2_fill_8 FILLER_209_1334 ();
 sg13g2_fill_8 FILLER_209_1342 ();
 sg13g2_fill_8 FILLER_209_1350 ();
 sg13g2_fill_8 FILLER_209_1358 ();
 sg13g2_fill_8 FILLER_209_1366 ();
 sg13g2_fill_8 FILLER_209_1374 ();
 sg13g2_fill_8 FILLER_209_1382 ();
 sg13g2_fill_8 FILLER_209_1390 ();
 sg13g2_fill_8 FILLER_209_1398 ();
 sg13g2_fill_8 FILLER_209_1406 ();
 sg13g2_fill_8 FILLER_209_1414 ();
 sg13g2_fill_8 FILLER_209_1422 ();
 sg13g2_fill_8 FILLER_209_1430 ();
 sg13g2_fill_8 FILLER_209_1438 ();
 sg13g2_fill_8 FILLER_209_1446 ();
 sg13g2_fill_8 FILLER_209_1454 ();
 sg13g2_fill_8 FILLER_209_1462 ();
 sg13g2_fill_8 FILLER_209_1470 ();
 sg13g2_fill_8 FILLER_209_1478 ();
 sg13g2_fill_8 FILLER_209_1486 ();
 sg13g2_fill_8 FILLER_209_1494 ();
 sg13g2_fill_8 FILLER_209_1502 ();
 sg13g2_fill_8 FILLER_209_1510 ();
 sg13g2_fill_8 FILLER_209_1518 ();
 sg13g2_fill_8 FILLER_209_1526 ();
 sg13g2_fill_8 FILLER_209_1534 ();
 sg13g2_fill_8 FILLER_209_1542 ();
 sg13g2_fill_8 FILLER_209_1550 ();
 sg13g2_fill_8 FILLER_209_1558 ();
 sg13g2_fill_8 FILLER_209_1566 ();
 sg13g2_fill_8 FILLER_209_1574 ();
 sg13g2_fill_8 FILLER_209_1582 ();
 sg13g2_fill_2 FILLER_209_1590 ();
 sg13g2_fill_8 FILLER_210_0 ();
 sg13g2_fill_8 FILLER_210_8 ();
 sg13g2_fill_8 FILLER_210_16 ();
 sg13g2_fill_8 FILLER_210_24 ();
 sg13g2_fill_8 FILLER_210_32 ();
 sg13g2_fill_8 FILLER_210_40 ();
 sg13g2_fill_8 FILLER_210_48 ();
 sg13g2_fill_8 FILLER_210_56 ();
 sg13g2_fill_8 FILLER_210_64 ();
 sg13g2_fill_8 FILLER_210_72 ();
 sg13g2_fill_8 FILLER_210_80 ();
 sg13g2_fill_8 FILLER_210_88 ();
 sg13g2_fill_8 FILLER_210_96 ();
 sg13g2_fill_8 FILLER_210_104 ();
 sg13g2_fill_8 FILLER_210_112 ();
 sg13g2_fill_8 FILLER_210_120 ();
 sg13g2_fill_8 FILLER_210_128 ();
 sg13g2_fill_8 FILLER_210_136 ();
 sg13g2_fill_8 FILLER_210_144 ();
 sg13g2_fill_8 FILLER_210_152 ();
 sg13g2_fill_8 FILLER_210_160 ();
 sg13g2_fill_8 FILLER_210_168 ();
 sg13g2_fill_8 FILLER_210_176 ();
 sg13g2_fill_8 FILLER_210_184 ();
 sg13g2_fill_8 FILLER_210_192 ();
 sg13g2_fill_8 FILLER_210_200 ();
 sg13g2_fill_8 FILLER_210_208 ();
 sg13g2_fill_8 FILLER_210_216 ();
 sg13g2_fill_8 FILLER_210_224 ();
 sg13g2_fill_8 FILLER_210_232 ();
 sg13g2_fill_8 FILLER_210_240 ();
 sg13g2_fill_8 FILLER_210_248 ();
 sg13g2_fill_8 FILLER_210_256 ();
 sg13g2_fill_8 FILLER_210_264 ();
 sg13g2_fill_8 FILLER_210_272 ();
 sg13g2_fill_8 FILLER_210_280 ();
 sg13g2_fill_8 FILLER_210_288 ();
 sg13g2_fill_8 FILLER_210_296 ();
 sg13g2_fill_8 FILLER_210_304 ();
 sg13g2_fill_8 FILLER_210_312 ();
 sg13g2_fill_8 FILLER_210_320 ();
 sg13g2_fill_8 FILLER_210_328 ();
 sg13g2_fill_8 FILLER_210_336 ();
 sg13g2_fill_8 FILLER_210_344 ();
 sg13g2_fill_8 FILLER_210_352 ();
 sg13g2_fill_8 FILLER_210_360 ();
 sg13g2_fill_8 FILLER_210_368 ();
 sg13g2_fill_8 FILLER_210_376 ();
 sg13g2_fill_8 FILLER_210_384 ();
 sg13g2_fill_8 FILLER_210_392 ();
 sg13g2_fill_8 FILLER_210_400 ();
 sg13g2_fill_8 FILLER_210_408 ();
 sg13g2_fill_8 FILLER_210_416 ();
 sg13g2_fill_8 FILLER_210_424 ();
 sg13g2_fill_8 FILLER_210_432 ();
 sg13g2_fill_8 FILLER_210_440 ();
 sg13g2_fill_8 FILLER_210_448 ();
 sg13g2_fill_8 FILLER_210_456 ();
 sg13g2_fill_8 FILLER_210_464 ();
 sg13g2_fill_8 FILLER_210_472 ();
 sg13g2_fill_8 FILLER_210_480 ();
 sg13g2_fill_8 FILLER_210_488 ();
 sg13g2_fill_8 FILLER_210_496 ();
 sg13g2_fill_8 FILLER_210_504 ();
 sg13g2_fill_8 FILLER_210_512 ();
 sg13g2_fill_8 FILLER_210_520 ();
 sg13g2_fill_8 FILLER_210_528 ();
 sg13g2_fill_8 FILLER_210_536 ();
 sg13g2_fill_8 FILLER_210_544 ();
 sg13g2_fill_8 FILLER_210_552 ();
 sg13g2_fill_8 FILLER_210_560 ();
 sg13g2_fill_8 FILLER_210_568 ();
 sg13g2_fill_8 FILLER_210_576 ();
 sg13g2_fill_8 FILLER_210_584 ();
 sg13g2_fill_8 FILLER_210_592 ();
 sg13g2_fill_8 FILLER_210_600 ();
 sg13g2_fill_8 FILLER_210_608 ();
 sg13g2_fill_8 FILLER_210_616 ();
 sg13g2_fill_8 FILLER_210_624 ();
 sg13g2_fill_8 FILLER_210_632 ();
 sg13g2_fill_8 FILLER_210_640 ();
 sg13g2_fill_8 FILLER_210_648 ();
 sg13g2_fill_8 FILLER_210_656 ();
 sg13g2_fill_8 FILLER_210_664 ();
 sg13g2_fill_8 FILLER_210_672 ();
 sg13g2_fill_8 FILLER_210_680 ();
 sg13g2_fill_8 FILLER_210_688 ();
 sg13g2_fill_8 FILLER_210_696 ();
 sg13g2_fill_8 FILLER_210_704 ();
 sg13g2_fill_8 FILLER_210_712 ();
 sg13g2_fill_8 FILLER_210_720 ();
 sg13g2_fill_8 FILLER_210_728 ();
 sg13g2_fill_8 FILLER_210_736 ();
 sg13g2_fill_8 FILLER_210_744 ();
 sg13g2_fill_8 FILLER_210_752 ();
 sg13g2_fill_8 FILLER_210_760 ();
 sg13g2_fill_8 FILLER_210_768 ();
 sg13g2_fill_8 FILLER_210_776 ();
 sg13g2_fill_8 FILLER_210_784 ();
 sg13g2_fill_8 FILLER_210_792 ();
 sg13g2_fill_8 FILLER_210_800 ();
 sg13g2_fill_8 FILLER_210_808 ();
 sg13g2_fill_8 FILLER_210_816 ();
 sg13g2_fill_8 FILLER_210_824 ();
 sg13g2_fill_8 FILLER_210_832 ();
 sg13g2_fill_8 FILLER_210_840 ();
 sg13g2_fill_8 FILLER_210_848 ();
 sg13g2_fill_8 FILLER_210_856 ();
 sg13g2_fill_8 FILLER_210_864 ();
 sg13g2_fill_8 FILLER_210_872 ();
 sg13g2_fill_8 FILLER_210_880 ();
 sg13g2_fill_8 FILLER_210_888 ();
 sg13g2_fill_8 FILLER_210_896 ();
 sg13g2_fill_8 FILLER_210_904 ();
 sg13g2_fill_8 FILLER_210_912 ();
 sg13g2_fill_8 FILLER_210_920 ();
 sg13g2_fill_8 FILLER_210_928 ();
 sg13g2_fill_8 FILLER_210_936 ();
 sg13g2_fill_8 FILLER_210_944 ();
 sg13g2_fill_8 FILLER_210_952 ();
 sg13g2_fill_8 FILLER_210_960 ();
 sg13g2_fill_8 FILLER_210_968 ();
 sg13g2_fill_8 FILLER_210_976 ();
 sg13g2_fill_8 FILLER_210_984 ();
 sg13g2_fill_8 FILLER_210_992 ();
 sg13g2_fill_8 FILLER_210_1000 ();
 sg13g2_fill_8 FILLER_210_1008 ();
 sg13g2_fill_8 FILLER_210_1016 ();
 sg13g2_fill_8 FILLER_210_1024 ();
 sg13g2_fill_8 FILLER_210_1032 ();
 sg13g2_fill_8 FILLER_210_1040 ();
 sg13g2_fill_8 FILLER_210_1048 ();
 sg13g2_fill_8 FILLER_210_1056 ();
 sg13g2_fill_8 FILLER_210_1064 ();
 sg13g2_fill_8 FILLER_210_1072 ();
 sg13g2_fill_8 FILLER_210_1080 ();
 sg13g2_fill_8 FILLER_210_1088 ();
 sg13g2_fill_8 FILLER_210_1096 ();
 sg13g2_fill_8 FILLER_210_1104 ();
 sg13g2_fill_8 FILLER_210_1112 ();
 sg13g2_fill_8 FILLER_210_1120 ();
 sg13g2_fill_8 FILLER_210_1128 ();
 sg13g2_fill_8 FILLER_210_1136 ();
 sg13g2_fill_8 FILLER_210_1144 ();
 sg13g2_fill_4 FILLER_210_1152 ();
 sg13g2_fill_1 FILLER_210_1177 ();
 sg13g2_fill_2 FILLER_210_1186 ();
 sg13g2_fill_1 FILLER_210_1188 ();
 sg13g2_fill_8 FILLER_210_1218 ();
 sg13g2_fill_2 FILLER_210_1226 ();
 sg13g2_fill_1 FILLER_210_1228 ();
 sg13g2_fill_8 FILLER_210_1233 ();
 sg13g2_fill_8 FILLER_210_1241 ();
 sg13g2_fill_4 FILLER_210_1249 ();
 sg13g2_fill_1 FILLER_210_1253 ();
 sg13g2_fill_8 FILLER_210_1262 ();
 sg13g2_fill_8 FILLER_210_1270 ();
 sg13g2_fill_8 FILLER_210_1278 ();
 sg13g2_fill_1 FILLER_210_1286 ();
 sg13g2_fill_2 FILLER_210_1292 ();
 sg13g2_fill_2 FILLER_210_1303 ();
 sg13g2_fill_1 FILLER_210_1305 ();
 sg13g2_fill_1 FILLER_210_1311 ();
 sg13g2_fill_8 FILLER_210_1316 ();
 sg13g2_fill_8 FILLER_210_1324 ();
 sg13g2_fill_8 FILLER_210_1332 ();
 sg13g2_fill_8 FILLER_210_1340 ();
 sg13g2_fill_8 FILLER_210_1348 ();
 sg13g2_fill_8 FILLER_210_1356 ();
 sg13g2_fill_8 FILLER_210_1364 ();
 sg13g2_fill_8 FILLER_210_1372 ();
 sg13g2_fill_8 FILLER_210_1380 ();
 sg13g2_fill_8 FILLER_210_1388 ();
 sg13g2_fill_8 FILLER_210_1396 ();
 sg13g2_fill_8 FILLER_210_1404 ();
 sg13g2_fill_8 FILLER_210_1412 ();
 sg13g2_fill_8 FILLER_210_1420 ();
 sg13g2_fill_8 FILLER_210_1428 ();
 sg13g2_fill_8 FILLER_210_1436 ();
 sg13g2_fill_8 FILLER_210_1444 ();
 sg13g2_fill_8 FILLER_210_1452 ();
 sg13g2_fill_8 FILLER_210_1460 ();
 sg13g2_fill_8 FILLER_210_1468 ();
 sg13g2_fill_8 FILLER_210_1476 ();
 sg13g2_fill_8 FILLER_210_1484 ();
 sg13g2_fill_8 FILLER_210_1492 ();
 sg13g2_fill_8 FILLER_210_1500 ();
 sg13g2_fill_8 FILLER_210_1508 ();
 sg13g2_fill_8 FILLER_210_1516 ();
 sg13g2_fill_8 FILLER_210_1524 ();
 sg13g2_fill_8 FILLER_210_1532 ();
 sg13g2_fill_8 FILLER_210_1540 ();
 sg13g2_fill_8 FILLER_210_1548 ();
 sg13g2_fill_8 FILLER_210_1556 ();
 sg13g2_fill_8 FILLER_210_1564 ();
 sg13g2_fill_8 FILLER_210_1572 ();
 sg13g2_fill_8 FILLER_210_1580 ();
 sg13g2_fill_4 FILLER_210_1588 ();
 sg13g2_fill_8 FILLER_211_0 ();
 sg13g2_fill_8 FILLER_211_8 ();
 sg13g2_fill_8 FILLER_211_16 ();
 sg13g2_fill_8 FILLER_211_24 ();
 sg13g2_fill_8 FILLER_211_32 ();
 sg13g2_fill_8 FILLER_211_40 ();
 sg13g2_fill_8 FILLER_211_48 ();
 sg13g2_fill_8 FILLER_211_56 ();
 sg13g2_fill_8 FILLER_211_64 ();
 sg13g2_fill_8 FILLER_211_72 ();
 sg13g2_fill_8 FILLER_211_80 ();
 sg13g2_fill_8 FILLER_211_88 ();
 sg13g2_fill_8 FILLER_211_96 ();
 sg13g2_fill_8 FILLER_211_104 ();
 sg13g2_fill_8 FILLER_211_112 ();
 sg13g2_fill_8 FILLER_211_120 ();
 sg13g2_fill_8 FILLER_211_128 ();
 sg13g2_fill_8 FILLER_211_136 ();
 sg13g2_fill_8 FILLER_211_144 ();
 sg13g2_fill_8 FILLER_211_152 ();
 sg13g2_fill_8 FILLER_211_160 ();
 sg13g2_fill_8 FILLER_211_168 ();
 sg13g2_fill_8 FILLER_211_176 ();
 sg13g2_fill_8 FILLER_211_184 ();
 sg13g2_fill_8 FILLER_211_192 ();
 sg13g2_fill_8 FILLER_211_200 ();
 sg13g2_fill_8 FILLER_211_208 ();
 sg13g2_fill_8 FILLER_211_216 ();
 sg13g2_fill_8 FILLER_211_224 ();
 sg13g2_fill_8 FILLER_211_232 ();
 sg13g2_fill_8 FILLER_211_240 ();
 sg13g2_fill_8 FILLER_211_248 ();
 sg13g2_fill_8 FILLER_211_256 ();
 sg13g2_fill_8 FILLER_211_264 ();
 sg13g2_fill_8 FILLER_211_272 ();
 sg13g2_fill_8 FILLER_211_280 ();
 sg13g2_fill_8 FILLER_211_288 ();
 sg13g2_fill_8 FILLER_211_296 ();
 sg13g2_fill_8 FILLER_211_304 ();
 sg13g2_fill_8 FILLER_211_312 ();
 sg13g2_fill_8 FILLER_211_320 ();
 sg13g2_fill_8 FILLER_211_328 ();
 sg13g2_fill_8 FILLER_211_336 ();
 sg13g2_fill_8 FILLER_211_344 ();
 sg13g2_fill_8 FILLER_211_352 ();
 sg13g2_fill_8 FILLER_211_360 ();
 sg13g2_fill_8 FILLER_211_368 ();
 sg13g2_fill_8 FILLER_211_376 ();
 sg13g2_fill_8 FILLER_211_384 ();
 sg13g2_fill_8 FILLER_211_392 ();
 sg13g2_fill_8 FILLER_211_400 ();
 sg13g2_fill_8 FILLER_211_408 ();
 sg13g2_fill_8 FILLER_211_416 ();
 sg13g2_fill_8 FILLER_211_424 ();
 sg13g2_fill_8 FILLER_211_432 ();
 sg13g2_fill_8 FILLER_211_440 ();
 sg13g2_fill_8 FILLER_211_448 ();
 sg13g2_fill_8 FILLER_211_456 ();
 sg13g2_fill_8 FILLER_211_464 ();
 sg13g2_fill_8 FILLER_211_472 ();
 sg13g2_fill_8 FILLER_211_480 ();
 sg13g2_fill_8 FILLER_211_488 ();
 sg13g2_fill_8 FILLER_211_496 ();
 sg13g2_fill_8 FILLER_211_504 ();
 sg13g2_fill_8 FILLER_211_512 ();
 sg13g2_fill_8 FILLER_211_520 ();
 sg13g2_fill_8 FILLER_211_528 ();
 sg13g2_fill_8 FILLER_211_536 ();
 sg13g2_fill_8 FILLER_211_544 ();
 sg13g2_fill_8 FILLER_211_552 ();
 sg13g2_fill_8 FILLER_211_560 ();
 sg13g2_fill_8 FILLER_211_568 ();
 sg13g2_fill_8 FILLER_211_576 ();
 sg13g2_fill_8 FILLER_211_584 ();
 sg13g2_fill_8 FILLER_211_592 ();
 sg13g2_fill_8 FILLER_211_600 ();
 sg13g2_fill_8 FILLER_211_608 ();
 sg13g2_fill_8 FILLER_211_616 ();
 sg13g2_fill_8 FILLER_211_624 ();
 sg13g2_fill_8 FILLER_211_632 ();
 sg13g2_fill_8 FILLER_211_640 ();
 sg13g2_fill_8 FILLER_211_648 ();
 sg13g2_fill_8 FILLER_211_656 ();
 sg13g2_fill_8 FILLER_211_664 ();
 sg13g2_fill_8 FILLER_211_672 ();
 sg13g2_fill_8 FILLER_211_680 ();
 sg13g2_fill_8 FILLER_211_688 ();
 sg13g2_fill_8 FILLER_211_696 ();
 sg13g2_fill_8 FILLER_211_704 ();
 sg13g2_fill_8 FILLER_211_712 ();
 sg13g2_fill_8 FILLER_211_720 ();
 sg13g2_fill_8 FILLER_211_728 ();
 sg13g2_fill_8 FILLER_211_736 ();
 sg13g2_fill_8 FILLER_211_744 ();
 sg13g2_fill_8 FILLER_211_752 ();
 sg13g2_fill_8 FILLER_211_760 ();
 sg13g2_fill_8 FILLER_211_768 ();
 sg13g2_fill_8 FILLER_211_776 ();
 sg13g2_fill_8 FILLER_211_784 ();
 sg13g2_fill_8 FILLER_211_792 ();
 sg13g2_fill_8 FILLER_211_800 ();
 sg13g2_fill_8 FILLER_211_808 ();
 sg13g2_fill_8 FILLER_211_816 ();
 sg13g2_fill_8 FILLER_211_824 ();
 sg13g2_fill_8 FILLER_211_832 ();
 sg13g2_fill_8 FILLER_211_840 ();
 sg13g2_fill_8 FILLER_211_848 ();
 sg13g2_fill_8 FILLER_211_856 ();
 sg13g2_fill_8 FILLER_211_864 ();
 sg13g2_fill_8 FILLER_211_872 ();
 sg13g2_fill_8 FILLER_211_880 ();
 sg13g2_fill_8 FILLER_211_888 ();
 sg13g2_fill_8 FILLER_211_896 ();
 sg13g2_fill_8 FILLER_211_904 ();
 sg13g2_fill_8 FILLER_211_912 ();
 sg13g2_fill_8 FILLER_211_920 ();
 sg13g2_fill_8 FILLER_211_928 ();
 sg13g2_fill_8 FILLER_211_936 ();
 sg13g2_fill_8 FILLER_211_944 ();
 sg13g2_fill_8 FILLER_211_952 ();
 sg13g2_fill_8 FILLER_211_960 ();
 sg13g2_fill_8 FILLER_211_968 ();
 sg13g2_fill_8 FILLER_211_976 ();
 sg13g2_fill_8 FILLER_211_984 ();
 sg13g2_fill_8 FILLER_211_992 ();
 sg13g2_fill_8 FILLER_211_1000 ();
 sg13g2_fill_8 FILLER_211_1008 ();
 sg13g2_fill_8 FILLER_211_1016 ();
 sg13g2_fill_8 FILLER_211_1024 ();
 sg13g2_fill_8 FILLER_211_1032 ();
 sg13g2_fill_8 FILLER_211_1040 ();
 sg13g2_fill_8 FILLER_211_1048 ();
 sg13g2_fill_8 FILLER_211_1056 ();
 sg13g2_fill_8 FILLER_211_1064 ();
 sg13g2_fill_8 FILLER_211_1072 ();
 sg13g2_fill_8 FILLER_211_1080 ();
 sg13g2_fill_8 FILLER_211_1088 ();
 sg13g2_fill_8 FILLER_211_1096 ();
 sg13g2_fill_8 FILLER_211_1104 ();
 sg13g2_fill_8 FILLER_211_1112 ();
 sg13g2_fill_8 FILLER_211_1120 ();
 sg13g2_fill_8 FILLER_211_1128 ();
 sg13g2_fill_8 FILLER_211_1136 ();
 sg13g2_fill_8 FILLER_211_1144 ();
 sg13g2_fill_8 FILLER_211_1152 ();
 sg13g2_fill_8 FILLER_211_1160 ();
 sg13g2_fill_8 FILLER_211_1168 ();
 sg13g2_fill_4 FILLER_211_1176 ();
 sg13g2_fill_2 FILLER_211_1180 ();
 sg13g2_fill_1 FILLER_211_1182 ();
 sg13g2_fill_2 FILLER_211_1194 ();
 sg13g2_fill_4 FILLER_211_1209 ();
 sg13g2_fill_2 FILLER_211_1213 ();
 sg13g2_fill_8 FILLER_211_1231 ();
 sg13g2_fill_4 FILLER_211_1239 ();
 sg13g2_fill_1 FILLER_211_1243 ();
 sg13g2_fill_2 FILLER_211_1252 ();
 sg13g2_fill_8 FILLER_211_1267 ();
 sg13g2_fill_8 FILLER_211_1275 ();
 sg13g2_fill_8 FILLER_211_1283 ();
 sg13g2_fill_8 FILLER_211_1291 ();
 sg13g2_fill_8 FILLER_211_1299 ();
 sg13g2_fill_8 FILLER_211_1307 ();
 sg13g2_fill_8 FILLER_211_1315 ();
 sg13g2_fill_8 FILLER_211_1323 ();
 sg13g2_fill_8 FILLER_211_1331 ();
 sg13g2_fill_8 FILLER_211_1339 ();
 sg13g2_fill_8 FILLER_211_1347 ();
 sg13g2_fill_8 FILLER_211_1355 ();
 sg13g2_fill_8 FILLER_211_1363 ();
 sg13g2_fill_8 FILLER_211_1371 ();
 sg13g2_fill_8 FILLER_211_1379 ();
 sg13g2_fill_8 FILLER_211_1387 ();
 sg13g2_fill_8 FILLER_211_1395 ();
 sg13g2_fill_8 FILLER_211_1403 ();
 sg13g2_fill_8 FILLER_211_1411 ();
 sg13g2_fill_8 FILLER_211_1419 ();
 sg13g2_fill_8 FILLER_211_1427 ();
 sg13g2_fill_8 FILLER_211_1435 ();
 sg13g2_fill_8 FILLER_211_1443 ();
 sg13g2_fill_8 FILLER_211_1451 ();
 sg13g2_fill_8 FILLER_211_1459 ();
 sg13g2_fill_8 FILLER_211_1467 ();
 sg13g2_fill_8 FILLER_211_1475 ();
 sg13g2_fill_8 FILLER_211_1483 ();
 sg13g2_fill_8 FILLER_211_1491 ();
 sg13g2_fill_8 FILLER_211_1499 ();
 sg13g2_fill_8 FILLER_211_1507 ();
 sg13g2_fill_8 FILLER_211_1515 ();
 sg13g2_fill_8 FILLER_211_1523 ();
 sg13g2_fill_8 FILLER_211_1531 ();
 sg13g2_fill_8 FILLER_211_1539 ();
 sg13g2_fill_8 FILLER_211_1547 ();
 sg13g2_fill_8 FILLER_211_1555 ();
 sg13g2_fill_8 FILLER_211_1563 ();
 sg13g2_fill_8 FILLER_211_1571 ();
 sg13g2_fill_8 FILLER_211_1579 ();
 sg13g2_fill_4 FILLER_211_1587 ();
 sg13g2_fill_1 FILLER_211_1591 ();
 sg13g2_fill_8 FILLER_212_0 ();
 sg13g2_fill_8 FILLER_212_8 ();
 sg13g2_fill_8 FILLER_212_16 ();
 sg13g2_fill_8 FILLER_212_24 ();
 sg13g2_fill_8 FILLER_212_32 ();
 sg13g2_fill_8 FILLER_212_40 ();
 sg13g2_fill_8 FILLER_212_48 ();
 sg13g2_fill_8 FILLER_212_56 ();
 sg13g2_fill_8 FILLER_212_64 ();
 sg13g2_fill_8 FILLER_212_72 ();
 sg13g2_fill_8 FILLER_212_80 ();
 sg13g2_fill_8 FILLER_212_88 ();
 sg13g2_fill_8 FILLER_212_96 ();
 sg13g2_fill_8 FILLER_212_104 ();
 sg13g2_fill_8 FILLER_212_112 ();
 sg13g2_fill_8 FILLER_212_120 ();
 sg13g2_fill_8 FILLER_212_128 ();
 sg13g2_fill_8 FILLER_212_136 ();
 sg13g2_fill_8 FILLER_212_144 ();
 sg13g2_fill_8 FILLER_212_152 ();
 sg13g2_fill_8 FILLER_212_160 ();
 sg13g2_fill_8 FILLER_212_168 ();
 sg13g2_fill_8 FILLER_212_176 ();
 sg13g2_fill_8 FILLER_212_184 ();
 sg13g2_fill_8 FILLER_212_192 ();
 sg13g2_fill_8 FILLER_212_200 ();
 sg13g2_fill_8 FILLER_212_208 ();
 sg13g2_fill_8 FILLER_212_216 ();
 sg13g2_fill_8 FILLER_212_224 ();
 sg13g2_fill_8 FILLER_212_232 ();
 sg13g2_fill_8 FILLER_212_240 ();
 sg13g2_fill_8 FILLER_212_248 ();
 sg13g2_fill_8 FILLER_212_256 ();
 sg13g2_fill_8 FILLER_212_264 ();
 sg13g2_fill_8 FILLER_212_272 ();
 sg13g2_fill_8 FILLER_212_280 ();
 sg13g2_fill_8 FILLER_212_288 ();
 sg13g2_fill_8 FILLER_212_296 ();
 sg13g2_fill_8 FILLER_212_304 ();
 sg13g2_fill_8 FILLER_212_312 ();
 sg13g2_fill_8 FILLER_212_320 ();
 sg13g2_fill_8 FILLER_212_328 ();
 sg13g2_fill_8 FILLER_212_336 ();
 sg13g2_fill_8 FILLER_212_344 ();
 sg13g2_fill_8 FILLER_212_352 ();
 sg13g2_fill_8 FILLER_212_360 ();
 sg13g2_fill_8 FILLER_212_368 ();
 sg13g2_fill_8 FILLER_212_376 ();
 sg13g2_fill_8 FILLER_212_384 ();
 sg13g2_fill_8 FILLER_212_392 ();
 sg13g2_fill_8 FILLER_212_400 ();
 sg13g2_fill_8 FILLER_212_408 ();
 sg13g2_fill_8 FILLER_212_416 ();
 sg13g2_fill_8 FILLER_212_424 ();
 sg13g2_fill_8 FILLER_212_432 ();
 sg13g2_fill_8 FILLER_212_440 ();
 sg13g2_fill_8 FILLER_212_448 ();
 sg13g2_fill_8 FILLER_212_456 ();
 sg13g2_fill_8 FILLER_212_464 ();
 sg13g2_fill_8 FILLER_212_472 ();
 sg13g2_fill_8 FILLER_212_480 ();
 sg13g2_fill_8 FILLER_212_488 ();
 sg13g2_fill_8 FILLER_212_496 ();
 sg13g2_fill_8 FILLER_212_504 ();
 sg13g2_fill_8 FILLER_212_512 ();
 sg13g2_fill_8 FILLER_212_520 ();
 sg13g2_fill_8 FILLER_212_528 ();
 sg13g2_fill_8 FILLER_212_536 ();
 sg13g2_fill_8 FILLER_212_544 ();
 sg13g2_fill_8 FILLER_212_552 ();
 sg13g2_fill_8 FILLER_212_560 ();
 sg13g2_fill_8 FILLER_212_568 ();
 sg13g2_fill_8 FILLER_212_576 ();
 sg13g2_fill_8 FILLER_212_584 ();
 sg13g2_fill_8 FILLER_212_592 ();
 sg13g2_fill_8 FILLER_212_600 ();
 sg13g2_fill_8 FILLER_212_608 ();
 sg13g2_fill_8 FILLER_212_616 ();
 sg13g2_fill_8 FILLER_212_624 ();
 sg13g2_fill_8 FILLER_212_632 ();
 sg13g2_fill_8 FILLER_212_640 ();
 sg13g2_fill_8 FILLER_212_648 ();
 sg13g2_fill_8 FILLER_212_656 ();
 sg13g2_fill_8 FILLER_212_664 ();
 sg13g2_fill_8 FILLER_212_672 ();
 sg13g2_fill_8 FILLER_212_680 ();
 sg13g2_fill_8 FILLER_212_688 ();
 sg13g2_fill_8 FILLER_212_696 ();
 sg13g2_fill_8 FILLER_212_704 ();
 sg13g2_fill_8 FILLER_212_712 ();
 sg13g2_fill_8 FILLER_212_720 ();
 sg13g2_fill_8 FILLER_212_728 ();
 sg13g2_fill_8 FILLER_212_736 ();
 sg13g2_fill_8 FILLER_212_744 ();
 sg13g2_fill_8 FILLER_212_752 ();
 sg13g2_fill_8 FILLER_212_760 ();
 sg13g2_fill_8 FILLER_212_768 ();
 sg13g2_fill_8 FILLER_212_776 ();
 sg13g2_fill_8 FILLER_212_784 ();
 sg13g2_fill_8 FILLER_212_792 ();
 sg13g2_fill_8 FILLER_212_800 ();
 sg13g2_fill_8 FILLER_212_808 ();
 sg13g2_fill_8 FILLER_212_816 ();
 sg13g2_fill_8 FILLER_212_824 ();
 sg13g2_fill_8 FILLER_212_832 ();
 sg13g2_fill_8 FILLER_212_840 ();
 sg13g2_fill_8 FILLER_212_848 ();
 sg13g2_fill_8 FILLER_212_856 ();
 sg13g2_fill_8 FILLER_212_864 ();
 sg13g2_fill_8 FILLER_212_872 ();
 sg13g2_fill_8 FILLER_212_880 ();
 sg13g2_fill_8 FILLER_212_888 ();
 sg13g2_fill_8 FILLER_212_896 ();
 sg13g2_fill_8 FILLER_212_904 ();
 sg13g2_fill_8 FILLER_212_912 ();
 sg13g2_fill_8 FILLER_212_920 ();
 sg13g2_fill_8 FILLER_212_928 ();
 sg13g2_fill_8 FILLER_212_936 ();
 sg13g2_fill_8 FILLER_212_944 ();
 sg13g2_fill_8 FILLER_212_952 ();
 sg13g2_fill_8 FILLER_212_960 ();
 sg13g2_fill_8 FILLER_212_968 ();
 sg13g2_fill_8 FILLER_212_976 ();
 sg13g2_fill_8 FILLER_212_984 ();
 sg13g2_fill_8 FILLER_212_992 ();
 sg13g2_fill_8 FILLER_212_1000 ();
 sg13g2_fill_8 FILLER_212_1008 ();
 sg13g2_fill_8 FILLER_212_1016 ();
 sg13g2_fill_8 FILLER_212_1024 ();
 sg13g2_fill_8 FILLER_212_1032 ();
 sg13g2_fill_8 FILLER_212_1040 ();
 sg13g2_fill_8 FILLER_212_1048 ();
 sg13g2_fill_8 FILLER_212_1056 ();
 sg13g2_fill_8 FILLER_212_1064 ();
 sg13g2_fill_8 FILLER_212_1072 ();
 sg13g2_fill_8 FILLER_212_1080 ();
 sg13g2_fill_8 FILLER_212_1088 ();
 sg13g2_fill_8 FILLER_212_1096 ();
 sg13g2_fill_8 FILLER_212_1104 ();
 sg13g2_fill_8 FILLER_212_1112 ();
 sg13g2_fill_8 FILLER_212_1120 ();
 sg13g2_fill_8 FILLER_212_1128 ();
 sg13g2_fill_8 FILLER_212_1136 ();
 sg13g2_fill_8 FILLER_212_1144 ();
 sg13g2_fill_8 FILLER_212_1152 ();
 sg13g2_fill_8 FILLER_212_1160 ();
 sg13g2_fill_8 FILLER_212_1168 ();
 sg13g2_fill_8 FILLER_212_1176 ();
 sg13g2_fill_8 FILLER_212_1184 ();
 sg13g2_fill_4 FILLER_212_1197 ();
 sg13g2_fill_8 FILLER_212_1206 ();
 sg13g2_fill_8 FILLER_212_1214 ();
 sg13g2_fill_2 FILLER_212_1222 ();
 sg13g2_fill_8 FILLER_212_1232 ();
 sg13g2_fill_8 FILLER_212_1240 ();
 sg13g2_fill_4 FILLER_212_1248 ();
 sg13g2_fill_1 FILLER_212_1252 ();
 sg13g2_fill_8 FILLER_212_1272 ();
 sg13g2_fill_8 FILLER_212_1280 ();
 sg13g2_fill_8 FILLER_212_1288 ();
 sg13g2_fill_8 FILLER_212_1296 ();
 sg13g2_fill_8 FILLER_212_1304 ();
 sg13g2_fill_8 FILLER_212_1312 ();
 sg13g2_fill_8 FILLER_212_1320 ();
 sg13g2_fill_8 FILLER_212_1328 ();
 sg13g2_fill_8 FILLER_212_1336 ();
 sg13g2_fill_8 FILLER_212_1344 ();
 sg13g2_fill_8 FILLER_212_1352 ();
 sg13g2_fill_8 FILLER_212_1360 ();
 sg13g2_fill_8 FILLER_212_1368 ();
 sg13g2_fill_8 FILLER_212_1376 ();
 sg13g2_fill_8 FILLER_212_1384 ();
 sg13g2_fill_8 FILLER_212_1392 ();
 sg13g2_fill_8 FILLER_212_1400 ();
 sg13g2_fill_8 FILLER_212_1408 ();
 sg13g2_fill_8 FILLER_212_1416 ();
 sg13g2_fill_8 FILLER_212_1424 ();
 sg13g2_fill_8 FILLER_212_1432 ();
 sg13g2_fill_8 FILLER_212_1440 ();
 sg13g2_fill_8 FILLER_212_1448 ();
 sg13g2_fill_8 FILLER_212_1456 ();
 sg13g2_fill_8 FILLER_212_1464 ();
 sg13g2_fill_8 FILLER_212_1472 ();
 sg13g2_fill_8 FILLER_212_1480 ();
 sg13g2_fill_8 FILLER_212_1488 ();
 sg13g2_fill_8 FILLER_212_1496 ();
 sg13g2_fill_8 FILLER_212_1504 ();
 sg13g2_fill_8 FILLER_212_1512 ();
 sg13g2_fill_8 FILLER_212_1520 ();
 sg13g2_fill_8 FILLER_212_1528 ();
 sg13g2_fill_8 FILLER_212_1536 ();
 sg13g2_fill_8 FILLER_212_1544 ();
 sg13g2_fill_8 FILLER_212_1552 ();
 sg13g2_fill_8 FILLER_212_1560 ();
 sg13g2_fill_8 FILLER_212_1568 ();
 sg13g2_fill_8 FILLER_212_1576 ();
 sg13g2_fill_8 FILLER_212_1584 ();
 sg13g2_fill_8 FILLER_213_0 ();
 sg13g2_fill_8 FILLER_213_8 ();
 sg13g2_fill_8 FILLER_213_16 ();
 sg13g2_fill_8 FILLER_213_24 ();
 sg13g2_fill_8 FILLER_213_32 ();
 sg13g2_fill_8 FILLER_213_40 ();
 sg13g2_fill_8 FILLER_213_48 ();
 sg13g2_fill_8 FILLER_213_56 ();
 sg13g2_fill_8 FILLER_213_64 ();
 sg13g2_fill_8 FILLER_213_72 ();
 sg13g2_fill_8 FILLER_213_80 ();
 sg13g2_fill_8 FILLER_213_88 ();
 sg13g2_fill_8 FILLER_213_96 ();
 sg13g2_fill_8 FILLER_213_104 ();
 sg13g2_fill_8 FILLER_213_112 ();
 sg13g2_fill_8 FILLER_213_120 ();
 sg13g2_fill_8 FILLER_213_128 ();
 sg13g2_fill_8 FILLER_213_136 ();
 sg13g2_fill_8 FILLER_213_144 ();
 sg13g2_fill_8 FILLER_213_152 ();
 sg13g2_fill_8 FILLER_213_160 ();
 sg13g2_fill_8 FILLER_213_168 ();
 sg13g2_fill_8 FILLER_213_176 ();
 sg13g2_fill_8 FILLER_213_184 ();
 sg13g2_fill_8 FILLER_213_192 ();
 sg13g2_fill_8 FILLER_213_200 ();
 sg13g2_fill_8 FILLER_213_208 ();
 sg13g2_fill_8 FILLER_213_216 ();
 sg13g2_fill_8 FILLER_213_224 ();
 sg13g2_fill_8 FILLER_213_232 ();
 sg13g2_fill_8 FILLER_213_240 ();
 sg13g2_fill_8 FILLER_213_248 ();
 sg13g2_fill_8 FILLER_213_256 ();
 sg13g2_fill_8 FILLER_213_264 ();
 sg13g2_fill_8 FILLER_213_272 ();
 sg13g2_fill_8 FILLER_213_280 ();
 sg13g2_fill_8 FILLER_213_288 ();
 sg13g2_fill_8 FILLER_213_296 ();
 sg13g2_fill_8 FILLER_213_304 ();
 sg13g2_fill_8 FILLER_213_312 ();
 sg13g2_fill_8 FILLER_213_320 ();
 sg13g2_fill_8 FILLER_213_328 ();
 sg13g2_fill_8 FILLER_213_336 ();
 sg13g2_fill_8 FILLER_213_344 ();
 sg13g2_fill_8 FILLER_213_352 ();
 sg13g2_fill_8 FILLER_213_360 ();
 sg13g2_fill_8 FILLER_213_368 ();
 sg13g2_fill_8 FILLER_213_376 ();
 sg13g2_fill_8 FILLER_213_384 ();
 sg13g2_fill_8 FILLER_213_392 ();
 sg13g2_fill_8 FILLER_213_400 ();
 sg13g2_fill_8 FILLER_213_408 ();
 sg13g2_fill_8 FILLER_213_416 ();
 sg13g2_fill_8 FILLER_213_424 ();
 sg13g2_fill_8 FILLER_213_432 ();
 sg13g2_fill_8 FILLER_213_440 ();
 sg13g2_fill_8 FILLER_213_448 ();
 sg13g2_fill_8 FILLER_213_456 ();
 sg13g2_fill_8 FILLER_213_464 ();
 sg13g2_fill_8 FILLER_213_472 ();
 sg13g2_fill_8 FILLER_213_480 ();
 sg13g2_fill_8 FILLER_213_488 ();
 sg13g2_fill_8 FILLER_213_496 ();
 sg13g2_fill_8 FILLER_213_504 ();
 sg13g2_fill_8 FILLER_213_512 ();
 sg13g2_fill_8 FILLER_213_520 ();
 sg13g2_fill_8 FILLER_213_528 ();
 sg13g2_fill_8 FILLER_213_536 ();
 sg13g2_fill_8 FILLER_213_544 ();
 sg13g2_fill_8 FILLER_213_552 ();
 sg13g2_fill_8 FILLER_213_560 ();
 sg13g2_fill_8 FILLER_213_568 ();
 sg13g2_fill_8 FILLER_213_576 ();
 sg13g2_fill_8 FILLER_213_584 ();
 sg13g2_fill_8 FILLER_213_592 ();
 sg13g2_fill_8 FILLER_213_600 ();
 sg13g2_fill_8 FILLER_213_608 ();
 sg13g2_fill_8 FILLER_213_616 ();
 sg13g2_fill_8 FILLER_213_624 ();
 sg13g2_fill_8 FILLER_213_632 ();
 sg13g2_fill_8 FILLER_213_640 ();
 sg13g2_fill_8 FILLER_213_648 ();
 sg13g2_fill_8 FILLER_213_656 ();
 sg13g2_fill_8 FILLER_213_664 ();
 sg13g2_fill_8 FILLER_213_672 ();
 sg13g2_fill_8 FILLER_213_680 ();
 sg13g2_fill_8 FILLER_213_688 ();
 sg13g2_fill_8 FILLER_213_696 ();
 sg13g2_fill_8 FILLER_213_704 ();
 sg13g2_fill_8 FILLER_213_712 ();
 sg13g2_fill_8 FILLER_213_720 ();
 sg13g2_fill_8 FILLER_213_728 ();
 sg13g2_fill_8 FILLER_213_736 ();
 sg13g2_fill_8 FILLER_213_744 ();
 sg13g2_fill_8 FILLER_213_752 ();
 sg13g2_fill_8 FILLER_213_760 ();
 sg13g2_fill_8 FILLER_213_768 ();
 sg13g2_fill_8 FILLER_213_776 ();
 sg13g2_fill_8 FILLER_213_784 ();
 sg13g2_fill_8 FILLER_213_792 ();
 sg13g2_fill_8 FILLER_213_800 ();
 sg13g2_fill_8 FILLER_213_808 ();
 sg13g2_fill_8 FILLER_213_816 ();
 sg13g2_fill_8 FILLER_213_824 ();
 sg13g2_fill_8 FILLER_213_832 ();
 sg13g2_fill_8 FILLER_213_840 ();
 sg13g2_fill_8 FILLER_213_848 ();
 sg13g2_fill_8 FILLER_213_856 ();
 sg13g2_fill_8 FILLER_213_864 ();
 sg13g2_fill_8 FILLER_213_872 ();
 sg13g2_fill_8 FILLER_213_880 ();
 sg13g2_fill_8 FILLER_213_888 ();
 sg13g2_fill_8 FILLER_213_896 ();
 sg13g2_fill_8 FILLER_213_904 ();
 sg13g2_fill_8 FILLER_213_912 ();
 sg13g2_fill_8 FILLER_213_920 ();
 sg13g2_fill_8 FILLER_213_928 ();
 sg13g2_fill_8 FILLER_213_936 ();
 sg13g2_fill_8 FILLER_213_944 ();
 sg13g2_fill_8 FILLER_213_952 ();
 sg13g2_fill_8 FILLER_213_960 ();
 sg13g2_fill_8 FILLER_213_968 ();
 sg13g2_fill_8 FILLER_213_976 ();
 sg13g2_fill_8 FILLER_213_984 ();
 sg13g2_fill_8 FILLER_213_992 ();
 sg13g2_fill_8 FILLER_213_1000 ();
 sg13g2_fill_8 FILLER_213_1008 ();
 sg13g2_fill_8 FILLER_213_1016 ();
 sg13g2_fill_8 FILLER_213_1024 ();
 sg13g2_fill_8 FILLER_213_1032 ();
 sg13g2_fill_8 FILLER_213_1040 ();
 sg13g2_fill_8 FILLER_213_1048 ();
 sg13g2_fill_8 FILLER_213_1056 ();
 sg13g2_fill_8 FILLER_213_1064 ();
 sg13g2_fill_8 FILLER_213_1072 ();
 sg13g2_fill_8 FILLER_213_1080 ();
 sg13g2_fill_8 FILLER_213_1088 ();
 sg13g2_fill_8 FILLER_213_1096 ();
 sg13g2_fill_8 FILLER_213_1104 ();
 sg13g2_fill_8 FILLER_213_1112 ();
 sg13g2_fill_8 FILLER_213_1120 ();
 sg13g2_fill_8 FILLER_213_1128 ();
 sg13g2_fill_8 FILLER_213_1136 ();
 sg13g2_fill_8 FILLER_213_1144 ();
 sg13g2_fill_8 FILLER_213_1152 ();
 sg13g2_fill_8 FILLER_213_1160 ();
 sg13g2_fill_8 FILLER_213_1168 ();
 sg13g2_fill_8 FILLER_213_1176 ();
 sg13g2_fill_4 FILLER_213_1184 ();
 sg13g2_fill_2 FILLER_213_1188 ();
 sg13g2_fill_4 FILLER_213_1211 ();
 sg13g2_fill_2 FILLER_213_1215 ();
 sg13g2_fill_1 FILLER_213_1235 ();
 sg13g2_fill_1 FILLER_213_1240 ();
 sg13g2_fill_1 FILLER_213_1245 ();
 sg13g2_fill_2 FILLER_213_1260 ();
 sg13g2_fill_8 FILLER_213_1267 ();
 sg13g2_fill_8 FILLER_213_1275 ();
 sg13g2_fill_8 FILLER_213_1283 ();
 sg13g2_fill_8 FILLER_213_1291 ();
 sg13g2_fill_8 FILLER_213_1299 ();
 sg13g2_fill_8 FILLER_213_1307 ();
 sg13g2_fill_8 FILLER_213_1315 ();
 sg13g2_fill_8 FILLER_213_1323 ();
 sg13g2_fill_8 FILLER_213_1331 ();
 sg13g2_fill_8 FILLER_213_1339 ();
 sg13g2_fill_8 FILLER_213_1347 ();
 sg13g2_fill_8 FILLER_213_1355 ();
 sg13g2_fill_8 FILLER_213_1363 ();
 sg13g2_fill_8 FILLER_213_1371 ();
 sg13g2_fill_8 FILLER_213_1379 ();
 sg13g2_fill_8 FILLER_213_1387 ();
 sg13g2_fill_8 FILLER_213_1395 ();
 sg13g2_fill_8 FILLER_213_1403 ();
 sg13g2_fill_8 FILLER_213_1411 ();
 sg13g2_fill_8 FILLER_213_1419 ();
 sg13g2_fill_8 FILLER_213_1427 ();
 sg13g2_fill_8 FILLER_213_1435 ();
 sg13g2_fill_8 FILLER_213_1443 ();
 sg13g2_fill_8 FILLER_213_1451 ();
 sg13g2_fill_8 FILLER_213_1459 ();
 sg13g2_fill_8 FILLER_213_1467 ();
 sg13g2_fill_8 FILLER_213_1475 ();
 sg13g2_fill_8 FILLER_213_1483 ();
 sg13g2_fill_8 FILLER_213_1491 ();
 sg13g2_fill_8 FILLER_213_1499 ();
 sg13g2_fill_8 FILLER_213_1507 ();
 sg13g2_fill_8 FILLER_213_1515 ();
 sg13g2_fill_8 FILLER_213_1523 ();
 sg13g2_fill_8 FILLER_213_1531 ();
 sg13g2_fill_8 FILLER_213_1539 ();
 sg13g2_fill_8 FILLER_213_1547 ();
 sg13g2_fill_8 FILLER_213_1555 ();
 sg13g2_fill_8 FILLER_213_1563 ();
 sg13g2_fill_8 FILLER_213_1571 ();
 sg13g2_fill_8 FILLER_213_1579 ();
 sg13g2_fill_4 FILLER_213_1587 ();
 sg13g2_fill_1 FILLER_213_1591 ();
 sg13g2_fill_8 FILLER_214_0 ();
 sg13g2_fill_8 FILLER_214_8 ();
 sg13g2_fill_8 FILLER_214_16 ();
 sg13g2_fill_8 FILLER_214_24 ();
 sg13g2_fill_8 FILLER_214_32 ();
 sg13g2_fill_8 FILLER_214_40 ();
 sg13g2_fill_8 FILLER_214_48 ();
 sg13g2_fill_8 FILLER_214_56 ();
 sg13g2_fill_8 FILLER_214_64 ();
 sg13g2_fill_8 FILLER_214_72 ();
 sg13g2_fill_8 FILLER_214_80 ();
 sg13g2_fill_8 FILLER_214_88 ();
 sg13g2_fill_8 FILLER_214_96 ();
 sg13g2_fill_8 FILLER_214_104 ();
 sg13g2_fill_8 FILLER_214_112 ();
 sg13g2_fill_8 FILLER_214_120 ();
 sg13g2_fill_8 FILLER_214_128 ();
 sg13g2_fill_8 FILLER_214_136 ();
 sg13g2_fill_8 FILLER_214_144 ();
 sg13g2_fill_8 FILLER_214_152 ();
 sg13g2_fill_8 FILLER_214_160 ();
 sg13g2_fill_8 FILLER_214_168 ();
 sg13g2_fill_8 FILLER_214_176 ();
 sg13g2_fill_8 FILLER_214_184 ();
 sg13g2_fill_8 FILLER_214_192 ();
 sg13g2_fill_8 FILLER_214_200 ();
 sg13g2_fill_8 FILLER_214_208 ();
 sg13g2_fill_8 FILLER_214_216 ();
 sg13g2_fill_8 FILLER_214_224 ();
 sg13g2_fill_8 FILLER_214_232 ();
 sg13g2_fill_8 FILLER_214_240 ();
 sg13g2_fill_8 FILLER_214_248 ();
 sg13g2_fill_8 FILLER_214_256 ();
 sg13g2_fill_8 FILLER_214_264 ();
 sg13g2_fill_8 FILLER_214_272 ();
 sg13g2_fill_8 FILLER_214_280 ();
 sg13g2_fill_8 FILLER_214_288 ();
 sg13g2_fill_8 FILLER_214_296 ();
 sg13g2_fill_8 FILLER_214_304 ();
 sg13g2_fill_8 FILLER_214_312 ();
 sg13g2_fill_8 FILLER_214_320 ();
 sg13g2_fill_8 FILLER_214_328 ();
 sg13g2_fill_8 FILLER_214_336 ();
 sg13g2_fill_8 FILLER_214_344 ();
 sg13g2_fill_8 FILLER_214_352 ();
 sg13g2_fill_8 FILLER_214_360 ();
 sg13g2_fill_8 FILLER_214_368 ();
 sg13g2_fill_8 FILLER_214_376 ();
 sg13g2_fill_8 FILLER_214_384 ();
 sg13g2_fill_8 FILLER_214_392 ();
 sg13g2_fill_8 FILLER_214_400 ();
 sg13g2_fill_8 FILLER_214_408 ();
 sg13g2_fill_8 FILLER_214_416 ();
 sg13g2_fill_8 FILLER_214_424 ();
 sg13g2_fill_8 FILLER_214_432 ();
 sg13g2_fill_8 FILLER_214_440 ();
 sg13g2_fill_8 FILLER_214_448 ();
 sg13g2_fill_8 FILLER_214_456 ();
 sg13g2_fill_8 FILLER_214_464 ();
 sg13g2_fill_8 FILLER_214_472 ();
 sg13g2_fill_8 FILLER_214_480 ();
 sg13g2_fill_8 FILLER_214_488 ();
 sg13g2_fill_8 FILLER_214_496 ();
 sg13g2_fill_8 FILLER_214_504 ();
 sg13g2_fill_8 FILLER_214_512 ();
 sg13g2_fill_8 FILLER_214_520 ();
 sg13g2_fill_8 FILLER_214_528 ();
 sg13g2_fill_8 FILLER_214_536 ();
 sg13g2_fill_8 FILLER_214_544 ();
 sg13g2_fill_8 FILLER_214_552 ();
 sg13g2_fill_8 FILLER_214_560 ();
 sg13g2_fill_8 FILLER_214_568 ();
 sg13g2_fill_8 FILLER_214_576 ();
 sg13g2_fill_8 FILLER_214_584 ();
 sg13g2_fill_8 FILLER_214_592 ();
 sg13g2_fill_8 FILLER_214_600 ();
 sg13g2_fill_8 FILLER_214_608 ();
 sg13g2_fill_8 FILLER_214_616 ();
 sg13g2_fill_8 FILLER_214_624 ();
 sg13g2_fill_8 FILLER_214_632 ();
 sg13g2_fill_8 FILLER_214_640 ();
 sg13g2_fill_8 FILLER_214_648 ();
 sg13g2_fill_8 FILLER_214_656 ();
 sg13g2_fill_8 FILLER_214_664 ();
 sg13g2_fill_8 FILLER_214_672 ();
 sg13g2_fill_8 FILLER_214_680 ();
 sg13g2_fill_8 FILLER_214_688 ();
 sg13g2_fill_8 FILLER_214_696 ();
 sg13g2_fill_8 FILLER_214_704 ();
 sg13g2_fill_8 FILLER_214_712 ();
 sg13g2_fill_8 FILLER_214_720 ();
 sg13g2_fill_8 FILLER_214_728 ();
 sg13g2_fill_8 FILLER_214_736 ();
 sg13g2_fill_8 FILLER_214_744 ();
 sg13g2_fill_8 FILLER_214_752 ();
 sg13g2_fill_8 FILLER_214_760 ();
 sg13g2_fill_8 FILLER_214_768 ();
 sg13g2_fill_8 FILLER_214_776 ();
 sg13g2_fill_8 FILLER_214_784 ();
 sg13g2_fill_8 FILLER_214_792 ();
 sg13g2_fill_8 FILLER_214_800 ();
 sg13g2_fill_8 FILLER_214_808 ();
 sg13g2_fill_8 FILLER_214_816 ();
 sg13g2_fill_8 FILLER_214_824 ();
 sg13g2_fill_8 FILLER_214_832 ();
 sg13g2_fill_8 FILLER_214_840 ();
 sg13g2_fill_8 FILLER_214_848 ();
 sg13g2_fill_8 FILLER_214_856 ();
 sg13g2_fill_8 FILLER_214_864 ();
 sg13g2_fill_8 FILLER_214_872 ();
 sg13g2_fill_8 FILLER_214_880 ();
 sg13g2_fill_8 FILLER_214_888 ();
 sg13g2_fill_8 FILLER_214_896 ();
 sg13g2_fill_8 FILLER_214_904 ();
 sg13g2_fill_8 FILLER_214_912 ();
 sg13g2_fill_8 FILLER_214_920 ();
 sg13g2_fill_8 FILLER_214_928 ();
 sg13g2_fill_8 FILLER_214_936 ();
 sg13g2_fill_8 FILLER_214_944 ();
 sg13g2_fill_8 FILLER_214_952 ();
 sg13g2_fill_8 FILLER_214_960 ();
 sg13g2_fill_8 FILLER_214_968 ();
 sg13g2_fill_8 FILLER_214_976 ();
 sg13g2_fill_8 FILLER_214_984 ();
 sg13g2_fill_8 FILLER_214_992 ();
 sg13g2_fill_8 FILLER_214_1000 ();
 sg13g2_fill_8 FILLER_214_1008 ();
 sg13g2_fill_8 FILLER_214_1016 ();
 sg13g2_fill_8 FILLER_214_1024 ();
 sg13g2_fill_8 FILLER_214_1032 ();
 sg13g2_fill_8 FILLER_214_1040 ();
 sg13g2_fill_8 FILLER_214_1048 ();
 sg13g2_fill_8 FILLER_214_1056 ();
 sg13g2_fill_8 FILLER_214_1064 ();
 sg13g2_fill_8 FILLER_214_1072 ();
 sg13g2_fill_8 FILLER_214_1080 ();
 sg13g2_fill_8 FILLER_214_1088 ();
 sg13g2_fill_8 FILLER_214_1096 ();
 sg13g2_fill_8 FILLER_214_1104 ();
 sg13g2_fill_8 FILLER_214_1112 ();
 sg13g2_fill_8 FILLER_214_1120 ();
 sg13g2_fill_8 FILLER_214_1128 ();
 sg13g2_fill_8 FILLER_214_1136 ();
 sg13g2_fill_8 FILLER_214_1144 ();
 sg13g2_fill_8 FILLER_214_1152 ();
 sg13g2_fill_8 FILLER_214_1160 ();
 sg13g2_fill_8 FILLER_214_1168 ();
 sg13g2_fill_8 FILLER_214_1176 ();
 sg13g2_fill_8 FILLER_214_1184 ();
 sg13g2_fill_2 FILLER_214_1192 ();
 sg13g2_fill_8 FILLER_214_1199 ();
 sg13g2_fill_4 FILLER_214_1207 ();
 sg13g2_fill_1 FILLER_214_1211 ();
 sg13g2_fill_8 FILLER_214_1275 ();
 sg13g2_fill_8 FILLER_214_1283 ();
 sg13g2_fill_8 FILLER_214_1291 ();
 sg13g2_fill_8 FILLER_214_1299 ();
 sg13g2_fill_8 FILLER_214_1307 ();
 sg13g2_fill_8 FILLER_214_1315 ();
 sg13g2_fill_8 FILLER_214_1323 ();
 sg13g2_fill_8 FILLER_214_1331 ();
 sg13g2_fill_8 FILLER_214_1339 ();
 sg13g2_fill_8 FILLER_214_1347 ();
 sg13g2_fill_8 FILLER_214_1355 ();
 sg13g2_fill_8 FILLER_214_1363 ();
 sg13g2_fill_8 FILLER_214_1371 ();
 sg13g2_fill_8 FILLER_214_1379 ();
 sg13g2_fill_8 FILLER_214_1387 ();
 sg13g2_fill_8 FILLER_214_1395 ();
 sg13g2_fill_8 FILLER_214_1403 ();
 sg13g2_fill_8 FILLER_214_1411 ();
 sg13g2_fill_8 FILLER_214_1419 ();
 sg13g2_fill_8 FILLER_214_1427 ();
 sg13g2_fill_8 FILLER_214_1435 ();
 sg13g2_fill_8 FILLER_214_1443 ();
 sg13g2_fill_8 FILLER_214_1451 ();
 sg13g2_fill_8 FILLER_214_1459 ();
 sg13g2_fill_8 FILLER_214_1467 ();
 sg13g2_fill_8 FILLER_214_1475 ();
 sg13g2_fill_8 FILLER_214_1483 ();
 sg13g2_fill_8 FILLER_214_1491 ();
 sg13g2_fill_8 FILLER_214_1499 ();
 sg13g2_fill_8 FILLER_214_1507 ();
 sg13g2_fill_8 FILLER_214_1515 ();
 sg13g2_fill_8 FILLER_214_1523 ();
 sg13g2_fill_8 FILLER_214_1531 ();
 sg13g2_fill_8 FILLER_214_1539 ();
 sg13g2_fill_8 FILLER_214_1547 ();
 sg13g2_fill_8 FILLER_214_1555 ();
 sg13g2_fill_8 FILLER_214_1563 ();
 sg13g2_fill_8 FILLER_214_1571 ();
 sg13g2_fill_8 FILLER_214_1579 ();
 sg13g2_fill_4 FILLER_214_1587 ();
 sg13g2_fill_1 FILLER_214_1591 ();
 sg13g2_fill_8 FILLER_215_0 ();
 sg13g2_fill_8 FILLER_215_8 ();
 sg13g2_fill_8 FILLER_215_16 ();
 sg13g2_fill_8 FILLER_215_24 ();
 sg13g2_fill_8 FILLER_215_32 ();
 sg13g2_fill_8 FILLER_215_40 ();
 sg13g2_fill_8 FILLER_215_48 ();
 sg13g2_fill_8 FILLER_215_56 ();
 sg13g2_fill_8 FILLER_215_64 ();
 sg13g2_fill_8 FILLER_215_72 ();
 sg13g2_fill_8 FILLER_215_80 ();
 sg13g2_fill_8 FILLER_215_88 ();
 sg13g2_fill_8 FILLER_215_96 ();
 sg13g2_fill_8 FILLER_215_104 ();
 sg13g2_fill_8 FILLER_215_112 ();
 sg13g2_fill_8 FILLER_215_120 ();
 sg13g2_fill_8 FILLER_215_128 ();
 sg13g2_fill_8 FILLER_215_136 ();
 sg13g2_fill_8 FILLER_215_144 ();
 sg13g2_fill_8 FILLER_215_152 ();
 sg13g2_fill_8 FILLER_215_160 ();
 sg13g2_fill_8 FILLER_215_168 ();
 sg13g2_fill_8 FILLER_215_176 ();
 sg13g2_fill_8 FILLER_215_184 ();
 sg13g2_fill_8 FILLER_215_192 ();
 sg13g2_fill_8 FILLER_215_200 ();
 sg13g2_fill_8 FILLER_215_208 ();
 sg13g2_fill_8 FILLER_215_216 ();
 sg13g2_fill_8 FILLER_215_224 ();
 sg13g2_fill_8 FILLER_215_232 ();
 sg13g2_fill_8 FILLER_215_240 ();
 sg13g2_fill_8 FILLER_215_248 ();
 sg13g2_fill_8 FILLER_215_256 ();
 sg13g2_fill_8 FILLER_215_264 ();
 sg13g2_fill_8 FILLER_215_272 ();
 sg13g2_fill_8 FILLER_215_280 ();
 sg13g2_fill_8 FILLER_215_288 ();
 sg13g2_fill_8 FILLER_215_296 ();
 sg13g2_fill_8 FILLER_215_304 ();
 sg13g2_fill_8 FILLER_215_312 ();
 sg13g2_fill_8 FILLER_215_320 ();
 sg13g2_fill_8 FILLER_215_328 ();
 sg13g2_fill_8 FILLER_215_336 ();
 sg13g2_fill_8 FILLER_215_344 ();
 sg13g2_fill_8 FILLER_215_352 ();
 sg13g2_fill_8 FILLER_215_360 ();
 sg13g2_fill_8 FILLER_215_368 ();
 sg13g2_fill_8 FILLER_215_376 ();
 sg13g2_fill_8 FILLER_215_384 ();
 sg13g2_fill_8 FILLER_215_392 ();
 sg13g2_fill_8 FILLER_215_400 ();
 sg13g2_fill_8 FILLER_215_408 ();
 sg13g2_fill_8 FILLER_215_416 ();
 sg13g2_fill_8 FILLER_215_424 ();
 sg13g2_fill_8 FILLER_215_432 ();
 sg13g2_fill_8 FILLER_215_440 ();
 sg13g2_fill_8 FILLER_215_448 ();
 sg13g2_fill_8 FILLER_215_456 ();
 sg13g2_fill_8 FILLER_215_464 ();
 sg13g2_fill_8 FILLER_215_472 ();
 sg13g2_fill_8 FILLER_215_480 ();
 sg13g2_fill_8 FILLER_215_488 ();
 sg13g2_fill_8 FILLER_215_496 ();
 sg13g2_fill_8 FILLER_215_504 ();
 sg13g2_fill_8 FILLER_215_512 ();
 sg13g2_fill_8 FILLER_215_520 ();
 sg13g2_fill_8 FILLER_215_528 ();
 sg13g2_fill_8 FILLER_215_536 ();
 sg13g2_fill_8 FILLER_215_544 ();
 sg13g2_fill_8 FILLER_215_552 ();
 sg13g2_fill_8 FILLER_215_560 ();
 sg13g2_fill_8 FILLER_215_568 ();
 sg13g2_fill_8 FILLER_215_576 ();
 sg13g2_fill_8 FILLER_215_584 ();
 sg13g2_fill_8 FILLER_215_592 ();
 sg13g2_fill_8 FILLER_215_600 ();
 sg13g2_fill_8 FILLER_215_608 ();
 sg13g2_fill_8 FILLER_215_616 ();
 sg13g2_fill_8 FILLER_215_624 ();
 sg13g2_fill_8 FILLER_215_632 ();
 sg13g2_fill_8 FILLER_215_640 ();
 sg13g2_fill_8 FILLER_215_648 ();
 sg13g2_fill_8 FILLER_215_656 ();
 sg13g2_fill_8 FILLER_215_664 ();
 sg13g2_fill_8 FILLER_215_672 ();
 sg13g2_fill_8 FILLER_215_680 ();
 sg13g2_fill_8 FILLER_215_688 ();
 sg13g2_fill_8 FILLER_215_696 ();
 sg13g2_fill_8 FILLER_215_704 ();
 sg13g2_fill_8 FILLER_215_712 ();
 sg13g2_fill_8 FILLER_215_720 ();
 sg13g2_fill_8 FILLER_215_728 ();
 sg13g2_fill_8 FILLER_215_736 ();
 sg13g2_fill_8 FILLER_215_744 ();
 sg13g2_fill_8 FILLER_215_752 ();
 sg13g2_fill_8 FILLER_215_760 ();
 sg13g2_fill_8 FILLER_215_768 ();
 sg13g2_fill_8 FILLER_215_776 ();
 sg13g2_fill_8 FILLER_215_784 ();
 sg13g2_fill_8 FILLER_215_792 ();
 sg13g2_fill_8 FILLER_215_800 ();
 sg13g2_fill_8 FILLER_215_808 ();
 sg13g2_fill_8 FILLER_215_816 ();
 sg13g2_fill_8 FILLER_215_824 ();
 sg13g2_fill_8 FILLER_215_832 ();
 sg13g2_fill_8 FILLER_215_840 ();
 sg13g2_fill_8 FILLER_215_848 ();
 sg13g2_fill_8 FILLER_215_856 ();
 sg13g2_fill_8 FILLER_215_864 ();
 sg13g2_fill_8 FILLER_215_872 ();
 sg13g2_fill_8 FILLER_215_880 ();
 sg13g2_fill_8 FILLER_215_888 ();
 sg13g2_fill_8 FILLER_215_896 ();
 sg13g2_fill_8 FILLER_215_904 ();
 sg13g2_fill_8 FILLER_215_912 ();
 sg13g2_fill_8 FILLER_215_920 ();
 sg13g2_fill_8 FILLER_215_928 ();
 sg13g2_fill_8 FILLER_215_936 ();
 sg13g2_fill_8 FILLER_215_944 ();
 sg13g2_fill_8 FILLER_215_952 ();
 sg13g2_fill_8 FILLER_215_960 ();
 sg13g2_fill_8 FILLER_215_968 ();
 sg13g2_fill_8 FILLER_215_976 ();
 sg13g2_fill_8 FILLER_215_984 ();
 sg13g2_fill_8 FILLER_215_992 ();
 sg13g2_fill_8 FILLER_215_1000 ();
 sg13g2_fill_8 FILLER_215_1008 ();
 sg13g2_fill_8 FILLER_215_1016 ();
 sg13g2_fill_8 FILLER_215_1024 ();
 sg13g2_fill_8 FILLER_215_1032 ();
 sg13g2_fill_8 FILLER_215_1040 ();
 sg13g2_fill_8 FILLER_215_1048 ();
 sg13g2_fill_8 FILLER_215_1056 ();
 sg13g2_fill_8 FILLER_215_1064 ();
 sg13g2_fill_8 FILLER_215_1072 ();
 sg13g2_fill_8 FILLER_215_1080 ();
 sg13g2_fill_8 FILLER_215_1088 ();
 sg13g2_fill_8 FILLER_215_1096 ();
 sg13g2_fill_8 FILLER_215_1104 ();
 sg13g2_fill_8 FILLER_215_1112 ();
 sg13g2_fill_8 FILLER_215_1120 ();
 sg13g2_fill_8 FILLER_215_1128 ();
 sg13g2_fill_8 FILLER_215_1136 ();
 sg13g2_fill_8 FILLER_215_1144 ();
 sg13g2_fill_8 FILLER_215_1152 ();
 sg13g2_fill_8 FILLER_215_1160 ();
 sg13g2_fill_8 FILLER_215_1168 ();
 sg13g2_fill_8 FILLER_215_1176 ();
 sg13g2_fill_8 FILLER_215_1184 ();
 sg13g2_fill_8 FILLER_215_1192 ();
 sg13g2_fill_8 FILLER_215_1200 ();
 sg13g2_fill_8 FILLER_215_1208 ();
 sg13g2_fill_8 FILLER_215_1216 ();
 sg13g2_fill_2 FILLER_215_1224 ();
 sg13g2_fill_1 FILLER_215_1226 ();
 sg13g2_fill_8 FILLER_215_1235 ();
 sg13g2_fill_2 FILLER_215_1243 ();
 sg13g2_fill_1 FILLER_215_1245 ();
 sg13g2_fill_8 FILLER_215_1264 ();
 sg13g2_fill_8 FILLER_215_1272 ();
 sg13g2_fill_8 FILLER_215_1280 ();
 sg13g2_fill_8 FILLER_215_1288 ();
 sg13g2_fill_8 FILLER_215_1296 ();
 sg13g2_fill_8 FILLER_215_1304 ();
 sg13g2_fill_8 FILLER_215_1312 ();
 sg13g2_fill_8 FILLER_215_1320 ();
 sg13g2_fill_8 FILLER_215_1328 ();
 sg13g2_fill_8 FILLER_215_1336 ();
 sg13g2_fill_8 FILLER_215_1344 ();
 sg13g2_fill_8 FILLER_215_1352 ();
 sg13g2_fill_8 FILLER_215_1360 ();
 sg13g2_fill_8 FILLER_215_1368 ();
 sg13g2_fill_8 FILLER_215_1376 ();
 sg13g2_fill_8 FILLER_215_1384 ();
 sg13g2_fill_8 FILLER_215_1392 ();
 sg13g2_fill_8 FILLER_215_1400 ();
 sg13g2_fill_8 FILLER_215_1408 ();
 sg13g2_fill_8 FILLER_215_1416 ();
 sg13g2_fill_8 FILLER_215_1424 ();
 sg13g2_fill_8 FILLER_215_1432 ();
 sg13g2_fill_8 FILLER_215_1440 ();
 sg13g2_fill_8 FILLER_215_1448 ();
 sg13g2_fill_8 FILLER_215_1456 ();
 sg13g2_fill_8 FILLER_215_1464 ();
 sg13g2_fill_8 FILLER_215_1472 ();
 sg13g2_fill_8 FILLER_215_1480 ();
 sg13g2_fill_8 FILLER_215_1488 ();
 sg13g2_fill_8 FILLER_215_1496 ();
 sg13g2_fill_8 FILLER_215_1504 ();
 sg13g2_fill_8 FILLER_215_1512 ();
 sg13g2_fill_8 FILLER_215_1520 ();
 sg13g2_fill_8 FILLER_215_1528 ();
 sg13g2_fill_8 FILLER_215_1536 ();
 sg13g2_fill_8 FILLER_215_1544 ();
 sg13g2_fill_8 FILLER_215_1552 ();
 sg13g2_fill_8 FILLER_215_1560 ();
 sg13g2_fill_8 FILLER_215_1568 ();
 sg13g2_fill_8 FILLER_215_1576 ();
 sg13g2_fill_8 FILLER_215_1584 ();
 sg13g2_fill_8 FILLER_216_0 ();
 sg13g2_fill_8 FILLER_216_8 ();
 sg13g2_fill_8 FILLER_216_16 ();
 sg13g2_fill_8 FILLER_216_24 ();
 sg13g2_fill_8 FILLER_216_32 ();
 sg13g2_fill_8 FILLER_216_40 ();
 sg13g2_fill_8 FILLER_216_48 ();
 sg13g2_fill_8 FILLER_216_56 ();
 sg13g2_fill_8 FILLER_216_64 ();
 sg13g2_fill_8 FILLER_216_72 ();
 sg13g2_fill_8 FILLER_216_80 ();
 sg13g2_fill_8 FILLER_216_88 ();
 sg13g2_fill_8 FILLER_216_96 ();
 sg13g2_fill_8 FILLER_216_104 ();
 sg13g2_fill_8 FILLER_216_112 ();
 sg13g2_fill_8 FILLER_216_120 ();
 sg13g2_fill_8 FILLER_216_128 ();
 sg13g2_fill_8 FILLER_216_136 ();
 sg13g2_fill_8 FILLER_216_144 ();
 sg13g2_fill_8 FILLER_216_152 ();
 sg13g2_fill_8 FILLER_216_160 ();
 sg13g2_fill_8 FILLER_216_168 ();
 sg13g2_fill_8 FILLER_216_176 ();
 sg13g2_fill_8 FILLER_216_184 ();
 sg13g2_fill_8 FILLER_216_192 ();
 sg13g2_fill_8 FILLER_216_200 ();
 sg13g2_fill_8 FILLER_216_208 ();
 sg13g2_fill_8 FILLER_216_216 ();
 sg13g2_fill_8 FILLER_216_224 ();
 sg13g2_fill_8 FILLER_216_232 ();
 sg13g2_fill_8 FILLER_216_240 ();
 sg13g2_fill_8 FILLER_216_248 ();
 sg13g2_fill_8 FILLER_216_256 ();
 sg13g2_fill_8 FILLER_216_264 ();
 sg13g2_fill_8 FILLER_216_272 ();
 sg13g2_fill_8 FILLER_216_280 ();
 sg13g2_fill_8 FILLER_216_288 ();
 sg13g2_fill_8 FILLER_216_296 ();
 sg13g2_fill_8 FILLER_216_304 ();
 sg13g2_fill_8 FILLER_216_312 ();
 sg13g2_fill_8 FILLER_216_320 ();
 sg13g2_fill_8 FILLER_216_328 ();
 sg13g2_fill_8 FILLER_216_336 ();
 sg13g2_fill_8 FILLER_216_344 ();
 sg13g2_fill_8 FILLER_216_352 ();
 sg13g2_fill_8 FILLER_216_360 ();
 sg13g2_fill_8 FILLER_216_368 ();
 sg13g2_fill_8 FILLER_216_376 ();
 sg13g2_fill_8 FILLER_216_384 ();
 sg13g2_fill_8 FILLER_216_392 ();
 sg13g2_fill_8 FILLER_216_400 ();
 sg13g2_fill_8 FILLER_216_408 ();
 sg13g2_fill_8 FILLER_216_416 ();
 sg13g2_fill_8 FILLER_216_424 ();
 sg13g2_fill_8 FILLER_216_432 ();
 sg13g2_fill_8 FILLER_216_440 ();
 sg13g2_fill_8 FILLER_216_448 ();
 sg13g2_fill_8 FILLER_216_456 ();
 sg13g2_fill_8 FILLER_216_464 ();
 sg13g2_fill_8 FILLER_216_472 ();
 sg13g2_fill_8 FILLER_216_480 ();
 sg13g2_fill_8 FILLER_216_488 ();
 sg13g2_fill_8 FILLER_216_496 ();
 sg13g2_fill_8 FILLER_216_504 ();
 sg13g2_fill_8 FILLER_216_512 ();
 sg13g2_fill_8 FILLER_216_520 ();
 sg13g2_fill_8 FILLER_216_528 ();
 sg13g2_fill_8 FILLER_216_536 ();
 sg13g2_fill_8 FILLER_216_544 ();
 sg13g2_fill_8 FILLER_216_552 ();
 sg13g2_fill_8 FILLER_216_560 ();
 sg13g2_fill_8 FILLER_216_568 ();
 sg13g2_fill_8 FILLER_216_576 ();
 sg13g2_fill_8 FILLER_216_584 ();
 sg13g2_fill_8 FILLER_216_592 ();
 sg13g2_fill_8 FILLER_216_600 ();
 sg13g2_fill_8 FILLER_216_608 ();
 sg13g2_fill_8 FILLER_216_616 ();
 sg13g2_fill_8 FILLER_216_624 ();
 sg13g2_fill_8 FILLER_216_632 ();
 sg13g2_fill_8 FILLER_216_640 ();
 sg13g2_fill_8 FILLER_216_648 ();
 sg13g2_fill_8 FILLER_216_656 ();
 sg13g2_fill_8 FILLER_216_664 ();
 sg13g2_fill_8 FILLER_216_672 ();
 sg13g2_fill_8 FILLER_216_680 ();
 sg13g2_fill_8 FILLER_216_688 ();
 sg13g2_fill_8 FILLER_216_696 ();
 sg13g2_fill_8 FILLER_216_704 ();
 sg13g2_fill_8 FILLER_216_712 ();
 sg13g2_fill_8 FILLER_216_720 ();
 sg13g2_fill_8 FILLER_216_728 ();
 sg13g2_fill_8 FILLER_216_736 ();
 sg13g2_fill_8 FILLER_216_744 ();
 sg13g2_fill_8 FILLER_216_752 ();
 sg13g2_fill_8 FILLER_216_760 ();
 sg13g2_fill_8 FILLER_216_768 ();
 sg13g2_fill_8 FILLER_216_776 ();
 sg13g2_fill_8 FILLER_216_784 ();
 sg13g2_fill_8 FILLER_216_792 ();
 sg13g2_fill_8 FILLER_216_800 ();
 sg13g2_fill_8 FILLER_216_808 ();
 sg13g2_fill_8 FILLER_216_816 ();
 sg13g2_fill_8 FILLER_216_824 ();
 sg13g2_fill_8 FILLER_216_832 ();
 sg13g2_fill_8 FILLER_216_840 ();
 sg13g2_fill_8 FILLER_216_848 ();
 sg13g2_fill_8 FILLER_216_856 ();
 sg13g2_fill_8 FILLER_216_864 ();
 sg13g2_fill_8 FILLER_216_872 ();
 sg13g2_fill_8 FILLER_216_880 ();
 sg13g2_fill_8 FILLER_216_888 ();
 sg13g2_fill_8 FILLER_216_896 ();
 sg13g2_fill_8 FILLER_216_904 ();
 sg13g2_fill_8 FILLER_216_912 ();
 sg13g2_fill_8 FILLER_216_920 ();
 sg13g2_fill_8 FILLER_216_928 ();
 sg13g2_fill_8 FILLER_216_936 ();
 sg13g2_fill_8 FILLER_216_944 ();
 sg13g2_fill_8 FILLER_216_952 ();
 sg13g2_fill_8 FILLER_216_960 ();
 sg13g2_fill_8 FILLER_216_968 ();
 sg13g2_fill_8 FILLER_216_976 ();
 sg13g2_fill_8 FILLER_216_984 ();
 sg13g2_fill_8 FILLER_216_992 ();
 sg13g2_fill_8 FILLER_216_1000 ();
 sg13g2_fill_8 FILLER_216_1008 ();
 sg13g2_fill_8 FILLER_216_1016 ();
 sg13g2_fill_8 FILLER_216_1024 ();
 sg13g2_fill_8 FILLER_216_1032 ();
 sg13g2_fill_8 FILLER_216_1040 ();
 sg13g2_fill_8 FILLER_216_1048 ();
 sg13g2_fill_8 FILLER_216_1056 ();
 sg13g2_fill_8 FILLER_216_1064 ();
 sg13g2_fill_8 FILLER_216_1072 ();
 sg13g2_fill_8 FILLER_216_1080 ();
 sg13g2_fill_8 FILLER_216_1088 ();
 sg13g2_fill_8 FILLER_216_1096 ();
 sg13g2_fill_8 FILLER_216_1104 ();
 sg13g2_fill_8 FILLER_216_1112 ();
 sg13g2_fill_8 FILLER_216_1120 ();
 sg13g2_fill_8 FILLER_216_1128 ();
 sg13g2_fill_8 FILLER_216_1136 ();
 sg13g2_fill_8 FILLER_216_1144 ();
 sg13g2_fill_8 FILLER_216_1152 ();
 sg13g2_fill_8 FILLER_216_1160 ();
 sg13g2_fill_8 FILLER_216_1168 ();
 sg13g2_fill_8 FILLER_216_1176 ();
 sg13g2_fill_8 FILLER_216_1184 ();
 sg13g2_fill_8 FILLER_216_1192 ();
 sg13g2_fill_8 FILLER_216_1200 ();
 sg13g2_fill_8 FILLER_216_1208 ();
 sg13g2_fill_8 FILLER_216_1216 ();
 sg13g2_fill_8 FILLER_216_1224 ();
 sg13g2_fill_8 FILLER_216_1232 ();
 sg13g2_fill_8 FILLER_216_1240 ();
 sg13g2_fill_4 FILLER_216_1248 ();
 sg13g2_fill_8 FILLER_216_1255 ();
 sg13g2_fill_8 FILLER_216_1263 ();
 sg13g2_fill_8 FILLER_216_1271 ();
 sg13g2_fill_8 FILLER_216_1279 ();
 sg13g2_fill_8 FILLER_216_1287 ();
 sg13g2_fill_8 FILLER_216_1295 ();
 sg13g2_fill_8 FILLER_216_1303 ();
 sg13g2_fill_8 FILLER_216_1311 ();
 sg13g2_fill_8 FILLER_216_1319 ();
 sg13g2_fill_8 FILLER_216_1327 ();
 sg13g2_fill_8 FILLER_216_1335 ();
 sg13g2_fill_8 FILLER_216_1343 ();
 sg13g2_fill_8 FILLER_216_1351 ();
 sg13g2_fill_8 FILLER_216_1359 ();
 sg13g2_fill_8 FILLER_216_1367 ();
 sg13g2_fill_8 FILLER_216_1375 ();
 sg13g2_fill_8 FILLER_216_1383 ();
 sg13g2_fill_8 FILLER_216_1391 ();
 sg13g2_fill_8 FILLER_216_1399 ();
 sg13g2_fill_8 FILLER_216_1407 ();
 sg13g2_fill_8 FILLER_216_1415 ();
 sg13g2_fill_8 FILLER_216_1423 ();
 sg13g2_fill_8 FILLER_216_1431 ();
 sg13g2_fill_8 FILLER_216_1439 ();
 sg13g2_fill_8 FILLER_216_1447 ();
 sg13g2_fill_8 FILLER_216_1455 ();
 sg13g2_fill_8 FILLER_216_1463 ();
 sg13g2_fill_8 FILLER_216_1471 ();
 sg13g2_fill_8 FILLER_216_1479 ();
 sg13g2_fill_8 FILLER_216_1487 ();
 sg13g2_fill_8 FILLER_216_1495 ();
 sg13g2_fill_8 FILLER_216_1503 ();
 sg13g2_fill_8 FILLER_216_1511 ();
 sg13g2_fill_8 FILLER_216_1519 ();
 sg13g2_fill_8 FILLER_216_1527 ();
 sg13g2_fill_8 FILLER_216_1535 ();
 sg13g2_fill_8 FILLER_216_1543 ();
 sg13g2_fill_8 FILLER_216_1551 ();
 sg13g2_fill_8 FILLER_216_1559 ();
 sg13g2_fill_8 FILLER_216_1567 ();
 sg13g2_fill_8 FILLER_216_1575 ();
 sg13g2_fill_8 FILLER_216_1583 ();
 sg13g2_fill_1 FILLER_216_1591 ();
 sg13g2_fill_8 FILLER_217_0 ();
 sg13g2_fill_8 FILLER_217_8 ();
 sg13g2_fill_8 FILLER_217_16 ();
 sg13g2_fill_8 FILLER_217_24 ();
 sg13g2_fill_8 FILLER_217_32 ();
 sg13g2_fill_8 FILLER_217_40 ();
 sg13g2_fill_8 FILLER_217_48 ();
 sg13g2_fill_8 FILLER_217_56 ();
 sg13g2_fill_8 FILLER_217_64 ();
 sg13g2_fill_8 FILLER_217_72 ();
 sg13g2_fill_8 FILLER_217_80 ();
 sg13g2_fill_8 FILLER_217_88 ();
 sg13g2_fill_8 FILLER_217_96 ();
 sg13g2_fill_8 FILLER_217_104 ();
 sg13g2_fill_8 FILLER_217_112 ();
 sg13g2_fill_8 FILLER_217_120 ();
 sg13g2_fill_8 FILLER_217_128 ();
 sg13g2_fill_8 FILLER_217_136 ();
 sg13g2_fill_8 FILLER_217_144 ();
 sg13g2_fill_8 FILLER_217_152 ();
 sg13g2_fill_8 FILLER_217_160 ();
 sg13g2_fill_8 FILLER_217_168 ();
 sg13g2_fill_8 FILLER_217_176 ();
 sg13g2_fill_8 FILLER_217_184 ();
 sg13g2_fill_8 FILLER_217_192 ();
 sg13g2_fill_8 FILLER_217_200 ();
 sg13g2_fill_8 FILLER_217_208 ();
 sg13g2_fill_8 FILLER_217_216 ();
 sg13g2_fill_8 FILLER_217_224 ();
 sg13g2_fill_8 FILLER_217_232 ();
 sg13g2_fill_8 FILLER_217_240 ();
 sg13g2_fill_8 FILLER_217_248 ();
 sg13g2_fill_8 FILLER_217_256 ();
 sg13g2_fill_8 FILLER_217_264 ();
 sg13g2_fill_8 FILLER_217_272 ();
 sg13g2_fill_8 FILLER_217_280 ();
 sg13g2_fill_8 FILLER_217_288 ();
 sg13g2_fill_8 FILLER_217_296 ();
 sg13g2_fill_8 FILLER_217_304 ();
 sg13g2_fill_8 FILLER_217_312 ();
 sg13g2_fill_8 FILLER_217_320 ();
 sg13g2_fill_8 FILLER_217_328 ();
 sg13g2_fill_8 FILLER_217_336 ();
 sg13g2_fill_8 FILLER_217_344 ();
 sg13g2_fill_8 FILLER_217_352 ();
 sg13g2_fill_8 FILLER_217_360 ();
 sg13g2_fill_8 FILLER_217_368 ();
 sg13g2_fill_8 FILLER_217_376 ();
 sg13g2_fill_8 FILLER_217_384 ();
 sg13g2_fill_8 FILLER_217_392 ();
 sg13g2_fill_8 FILLER_217_400 ();
 sg13g2_fill_8 FILLER_217_408 ();
 sg13g2_fill_8 FILLER_217_416 ();
 sg13g2_fill_8 FILLER_217_424 ();
 sg13g2_fill_8 FILLER_217_432 ();
 sg13g2_fill_8 FILLER_217_440 ();
 sg13g2_fill_8 FILLER_217_448 ();
 sg13g2_fill_8 FILLER_217_456 ();
 sg13g2_fill_8 FILLER_217_464 ();
 sg13g2_fill_8 FILLER_217_472 ();
 sg13g2_fill_8 FILLER_217_480 ();
 sg13g2_fill_8 FILLER_217_488 ();
 sg13g2_fill_8 FILLER_217_496 ();
 sg13g2_fill_8 FILLER_217_504 ();
 sg13g2_fill_8 FILLER_217_512 ();
 sg13g2_fill_8 FILLER_217_520 ();
 sg13g2_fill_8 FILLER_217_528 ();
 sg13g2_fill_8 FILLER_217_536 ();
 sg13g2_fill_8 FILLER_217_544 ();
 sg13g2_fill_8 FILLER_217_552 ();
 sg13g2_fill_8 FILLER_217_560 ();
 sg13g2_fill_8 FILLER_217_568 ();
 sg13g2_fill_8 FILLER_217_576 ();
 sg13g2_fill_8 FILLER_217_584 ();
 sg13g2_fill_8 FILLER_217_592 ();
 sg13g2_fill_8 FILLER_217_600 ();
 sg13g2_fill_8 FILLER_217_608 ();
 sg13g2_fill_8 FILLER_217_616 ();
 sg13g2_fill_8 FILLER_217_624 ();
 sg13g2_fill_8 FILLER_217_632 ();
 sg13g2_fill_8 FILLER_217_640 ();
 sg13g2_fill_8 FILLER_217_648 ();
 sg13g2_fill_8 FILLER_217_656 ();
 sg13g2_fill_8 FILLER_217_664 ();
 sg13g2_fill_8 FILLER_217_672 ();
 sg13g2_fill_8 FILLER_217_680 ();
 sg13g2_fill_8 FILLER_217_688 ();
 sg13g2_fill_8 FILLER_217_696 ();
 sg13g2_fill_8 FILLER_217_704 ();
 sg13g2_fill_8 FILLER_217_712 ();
 sg13g2_fill_8 FILLER_217_720 ();
 sg13g2_fill_8 FILLER_217_728 ();
 sg13g2_fill_8 FILLER_217_736 ();
 sg13g2_fill_8 FILLER_217_744 ();
 sg13g2_fill_8 FILLER_217_752 ();
 sg13g2_fill_8 FILLER_217_760 ();
 sg13g2_fill_8 FILLER_217_768 ();
 sg13g2_fill_8 FILLER_217_776 ();
 sg13g2_fill_8 FILLER_217_784 ();
 sg13g2_fill_8 FILLER_217_792 ();
 sg13g2_fill_8 FILLER_217_800 ();
 sg13g2_fill_8 FILLER_217_808 ();
 sg13g2_fill_8 FILLER_217_816 ();
 sg13g2_fill_8 FILLER_217_824 ();
 sg13g2_fill_8 FILLER_217_832 ();
 sg13g2_fill_8 FILLER_217_840 ();
 sg13g2_fill_8 FILLER_217_848 ();
 sg13g2_fill_8 FILLER_217_856 ();
 sg13g2_fill_8 FILLER_217_864 ();
 sg13g2_fill_8 FILLER_217_872 ();
 sg13g2_fill_8 FILLER_217_880 ();
 sg13g2_fill_8 FILLER_217_888 ();
 sg13g2_fill_8 FILLER_217_896 ();
 sg13g2_fill_8 FILLER_217_904 ();
 sg13g2_fill_8 FILLER_217_912 ();
 sg13g2_fill_8 FILLER_217_920 ();
 sg13g2_fill_8 FILLER_217_928 ();
 sg13g2_fill_8 FILLER_217_936 ();
 sg13g2_fill_8 FILLER_217_944 ();
 sg13g2_fill_8 FILLER_217_952 ();
 sg13g2_fill_8 FILLER_217_960 ();
 sg13g2_fill_8 FILLER_217_968 ();
 sg13g2_fill_8 FILLER_217_976 ();
 sg13g2_fill_8 FILLER_217_984 ();
 sg13g2_fill_8 FILLER_217_992 ();
 sg13g2_fill_8 FILLER_217_1000 ();
 sg13g2_fill_8 FILLER_217_1008 ();
 sg13g2_fill_8 FILLER_217_1016 ();
 sg13g2_fill_8 FILLER_217_1024 ();
 sg13g2_fill_8 FILLER_217_1032 ();
 sg13g2_fill_8 FILLER_217_1040 ();
 sg13g2_fill_8 FILLER_217_1048 ();
 sg13g2_fill_8 FILLER_217_1056 ();
 sg13g2_fill_8 FILLER_217_1064 ();
 sg13g2_fill_8 FILLER_217_1072 ();
 sg13g2_fill_8 FILLER_217_1080 ();
 sg13g2_fill_8 FILLER_217_1088 ();
 sg13g2_fill_8 FILLER_217_1096 ();
 sg13g2_fill_8 FILLER_217_1104 ();
 sg13g2_fill_8 FILLER_217_1112 ();
 sg13g2_fill_8 FILLER_217_1120 ();
 sg13g2_fill_8 FILLER_217_1128 ();
 sg13g2_fill_8 FILLER_217_1136 ();
 sg13g2_fill_8 FILLER_217_1144 ();
 sg13g2_fill_8 FILLER_217_1152 ();
 sg13g2_fill_8 FILLER_217_1160 ();
 sg13g2_fill_8 FILLER_217_1168 ();
 sg13g2_fill_8 FILLER_217_1176 ();
 sg13g2_fill_8 FILLER_217_1184 ();
 sg13g2_fill_8 FILLER_217_1192 ();
 sg13g2_fill_8 FILLER_217_1200 ();
 sg13g2_fill_8 FILLER_217_1208 ();
 sg13g2_fill_8 FILLER_217_1216 ();
 sg13g2_fill_8 FILLER_217_1224 ();
 sg13g2_fill_8 FILLER_217_1232 ();
 sg13g2_fill_8 FILLER_217_1240 ();
 sg13g2_fill_8 FILLER_217_1248 ();
 sg13g2_fill_8 FILLER_217_1256 ();
 sg13g2_fill_8 FILLER_217_1264 ();
 sg13g2_fill_8 FILLER_217_1272 ();
 sg13g2_fill_8 FILLER_217_1280 ();
 sg13g2_fill_8 FILLER_217_1288 ();
 sg13g2_fill_8 FILLER_217_1296 ();
 sg13g2_fill_8 FILLER_217_1304 ();
 sg13g2_fill_8 FILLER_217_1312 ();
 sg13g2_fill_8 FILLER_217_1320 ();
 sg13g2_fill_8 FILLER_217_1328 ();
 sg13g2_fill_8 FILLER_217_1336 ();
 sg13g2_fill_8 FILLER_217_1344 ();
 sg13g2_fill_8 FILLER_217_1352 ();
 sg13g2_fill_8 FILLER_217_1360 ();
 sg13g2_fill_8 FILLER_217_1368 ();
 sg13g2_fill_8 FILLER_217_1376 ();
 sg13g2_fill_8 FILLER_217_1384 ();
 sg13g2_fill_8 FILLER_217_1392 ();
 sg13g2_fill_8 FILLER_217_1400 ();
 sg13g2_fill_8 FILLER_217_1408 ();
 sg13g2_fill_8 FILLER_217_1416 ();
 sg13g2_fill_8 FILLER_217_1424 ();
 sg13g2_fill_8 FILLER_217_1432 ();
 sg13g2_fill_8 FILLER_217_1440 ();
 sg13g2_fill_8 FILLER_217_1448 ();
 sg13g2_fill_8 FILLER_217_1456 ();
 sg13g2_fill_8 FILLER_217_1464 ();
 sg13g2_fill_8 FILLER_217_1472 ();
 sg13g2_fill_8 FILLER_217_1480 ();
 sg13g2_fill_8 FILLER_217_1488 ();
 sg13g2_fill_8 FILLER_217_1496 ();
 sg13g2_fill_8 FILLER_217_1504 ();
 sg13g2_fill_8 FILLER_217_1512 ();
 sg13g2_fill_8 FILLER_217_1520 ();
 sg13g2_fill_8 FILLER_217_1528 ();
 sg13g2_fill_8 FILLER_217_1536 ();
 sg13g2_fill_8 FILLER_217_1544 ();
 sg13g2_fill_8 FILLER_217_1552 ();
 sg13g2_fill_8 FILLER_217_1560 ();
 sg13g2_fill_8 FILLER_217_1568 ();
 sg13g2_fill_8 FILLER_217_1576 ();
 sg13g2_fill_8 FILLER_217_1584 ();
 sg13g2_fill_8 FILLER_218_0 ();
 sg13g2_fill_8 FILLER_218_8 ();
 sg13g2_fill_8 FILLER_218_16 ();
 sg13g2_fill_8 FILLER_218_24 ();
 sg13g2_fill_8 FILLER_218_32 ();
 sg13g2_fill_8 FILLER_218_40 ();
 sg13g2_fill_8 FILLER_218_48 ();
 sg13g2_fill_8 FILLER_218_56 ();
 sg13g2_fill_8 FILLER_218_64 ();
 sg13g2_fill_8 FILLER_218_72 ();
 sg13g2_fill_8 FILLER_218_80 ();
 sg13g2_fill_8 FILLER_218_88 ();
 sg13g2_fill_8 FILLER_218_96 ();
 sg13g2_fill_8 FILLER_218_104 ();
 sg13g2_fill_8 FILLER_218_112 ();
 sg13g2_fill_8 FILLER_218_120 ();
 sg13g2_fill_8 FILLER_218_128 ();
 sg13g2_fill_8 FILLER_218_136 ();
 sg13g2_fill_8 FILLER_218_144 ();
 sg13g2_fill_8 FILLER_218_152 ();
 sg13g2_fill_8 FILLER_218_160 ();
 sg13g2_fill_8 FILLER_218_168 ();
 sg13g2_fill_8 FILLER_218_176 ();
 sg13g2_fill_8 FILLER_218_184 ();
 sg13g2_fill_8 FILLER_218_192 ();
 sg13g2_fill_8 FILLER_218_200 ();
 sg13g2_fill_8 FILLER_218_208 ();
 sg13g2_fill_8 FILLER_218_216 ();
 sg13g2_fill_8 FILLER_218_224 ();
 sg13g2_fill_8 FILLER_218_232 ();
 sg13g2_fill_8 FILLER_218_240 ();
 sg13g2_fill_8 FILLER_218_248 ();
 sg13g2_fill_8 FILLER_218_256 ();
 sg13g2_fill_8 FILLER_218_264 ();
 sg13g2_fill_8 FILLER_218_272 ();
 sg13g2_fill_8 FILLER_218_280 ();
 sg13g2_fill_8 FILLER_218_288 ();
 sg13g2_fill_8 FILLER_218_296 ();
 sg13g2_fill_8 FILLER_218_304 ();
 sg13g2_fill_8 FILLER_218_312 ();
 sg13g2_fill_8 FILLER_218_320 ();
 sg13g2_fill_8 FILLER_218_328 ();
 sg13g2_fill_8 FILLER_218_336 ();
 sg13g2_fill_8 FILLER_218_344 ();
 sg13g2_fill_8 FILLER_218_352 ();
 sg13g2_fill_8 FILLER_218_360 ();
 sg13g2_fill_8 FILLER_218_368 ();
 sg13g2_fill_8 FILLER_218_376 ();
 sg13g2_fill_8 FILLER_218_384 ();
 sg13g2_fill_8 FILLER_218_392 ();
 sg13g2_fill_8 FILLER_218_400 ();
 sg13g2_fill_8 FILLER_218_408 ();
 sg13g2_fill_8 FILLER_218_416 ();
 sg13g2_fill_8 FILLER_218_424 ();
 sg13g2_fill_8 FILLER_218_432 ();
 sg13g2_fill_8 FILLER_218_440 ();
 sg13g2_fill_8 FILLER_218_448 ();
 sg13g2_fill_8 FILLER_218_456 ();
 sg13g2_fill_8 FILLER_218_464 ();
 sg13g2_fill_8 FILLER_218_472 ();
 sg13g2_fill_8 FILLER_218_480 ();
 sg13g2_fill_8 FILLER_218_488 ();
 sg13g2_fill_8 FILLER_218_496 ();
 sg13g2_fill_8 FILLER_218_504 ();
 sg13g2_fill_8 FILLER_218_512 ();
 sg13g2_fill_8 FILLER_218_520 ();
 sg13g2_fill_8 FILLER_218_528 ();
 sg13g2_fill_8 FILLER_218_536 ();
 sg13g2_fill_8 FILLER_218_544 ();
 sg13g2_fill_8 FILLER_218_552 ();
 sg13g2_fill_8 FILLER_218_560 ();
 sg13g2_fill_8 FILLER_218_568 ();
 sg13g2_fill_8 FILLER_218_576 ();
 sg13g2_fill_8 FILLER_218_584 ();
 sg13g2_fill_8 FILLER_218_592 ();
 sg13g2_fill_8 FILLER_218_600 ();
 sg13g2_fill_8 FILLER_218_608 ();
 sg13g2_fill_8 FILLER_218_616 ();
 sg13g2_fill_8 FILLER_218_624 ();
 sg13g2_fill_8 FILLER_218_632 ();
 sg13g2_fill_8 FILLER_218_640 ();
 sg13g2_fill_8 FILLER_218_648 ();
 sg13g2_fill_8 FILLER_218_656 ();
 sg13g2_fill_8 FILLER_218_664 ();
 sg13g2_fill_8 FILLER_218_672 ();
 sg13g2_fill_8 FILLER_218_680 ();
 sg13g2_fill_8 FILLER_218_688 ();
 sg13g2_fill_8 FILLER_218_696 ();
 sg13g2_fill_8 FILLER_218_704 ();
 sg13g2_fill_8 FILLER_218_712 ();
 sg13g2_fill_8 FILLER_218_720 ();
 sg13g2_fill_8 FILLER_218_728 ();
 sg13g2_fill_8 FILLER_218_736 ();
 sg13g2_fill_8 FILLER_218_744 ();
 sg13g2_fill_8 FILLER_218_752 ();
 sg13g2_fill_8 FILLER_218_760 ();
 sg13g2_fill_8 FILLER_218_768 ();
 sg13g2_fill_8 FILLER_218_776 ();
 sg13g2_fill_8 FILLER_218_784 ();
 sg13g2_fill_8 FILLER_218_792 ();
 sg13g2_fill_8 FILLER_218_800 ();
 sg13g2_fill_8 FILLER_218_808 ();
 sg13g2_fill_8 FILLER_218_816 ();
 sg13g2_fill_8 FILLER_218_824 ();
 sg13g2_fill_8 FILLER_218_832 ();
 sg13g2_fill_8 FILLER_218_840 ();
 sg13g2_fill_8 FILLER_218_848 ();
 sg13g2_fill_8 FILLER_218_856 ();
 sg13g2_fill_8 FILLER_218_864 ();
 sg13g2_fill_8 FILLER_218_872 ();
 sg13g2_fill_8 FILLER_218_880 ();
 sg13g2_fill_8 FILLER_218_888 ();
 sg13g2_fill_8 FILLER_218_896 ();
 sg13g2_fill_8 FILLER_218_904 ();
 sg13g2_fill_8 FILLER_218_912 ();
 sg13g2_fill_8 FILLER_218_920 ();
 sg13g2_fill_8 FILLER_218_928 ();
 sg13g2_fill_8 FILLER_218_936 ();
 sg13g2_fill_8 FILLER_218_944 ();
 sg13g2_fill_8 FILLER_218_952 ();
 sg13g2_fill_8 FILLER_218_960 ();
 sg13g2_fill_8 FILLER_218_968 ();
 sg13g2_fill_8 FILLER_218_976 ();
 sg13g2_fill_8 FILLER_218_984 ();
 sg13g2_fill_8 FILLER_218_992 ();
 sg13g2_fill_8 FILLER_218_1000 ();
 sg13g2_fill_8 FILLER_218_1008 ();
 sg13g2_fill_8 FILLER_218_1016 ();
 sg13g2_fill_8 FILLER_218_1024 ();
 sg13g2_fill_8 FILLER_218_1032 ();
 sg13g2_fill_8 FILLER_218_1040 ();
 sg13g2_fill_8 FILLER_218_1048 ();
 sg13g2_fill_8 FILLER_218_1056 ();
 sg13g2_fill_8 FILLER_218_1064 ();
 sg13g2_fill_8 FILLER_218_1072 ();
 sg13g2_fill_8 FILLER_218_1080 ();
 sg13g2_fill_8 FILLER_218_1088 ();
 sg13g2_fill_8 FILLER_218_1096 ();
 sg13g2_fill_8 FILLER_218_1104 ();
 sg13g2_fill_8 FILLER_218_1112 ();
 sg13g2_fill_8 FILLER_218_1120 ();
 sg13g2_fill_8 FILLER_218_1128 ();
 sg13g2_fill_8 FILLER_218_1136 ();
 sg13g2_fill_8 FILLER_218_1144 ();
 sg13g2_fill_8 FILLER_218_1152 ();
 sg13g2_fill_8 FILLER_218_1160 ();
 sg13g2_fill_8 FILLER_218_1168 ();
 sg13g2_fill_8 FILLER_218_1176 ();
 sg13g2_fill_8 FILLER_218_1184 ();
 sg13g2_fill_8 FILLER_218_1192 ();
 sg13g2_fill_8 FILLER_218_1200 ();
 sg13g2_fill_8 FILLER_218_1208 ();
 sg13g2_fill_8 FILLER_218_1216 ();
 sg13g2_fill_8 FILLER_218_1224 ();
 sg13g2_fill_8 FILLER_218_1232 ();
 sg13g2_fill_8 FILLER_218_1240 ();
 sg13g2_fill_8 FILLER_218_1248 ();
 sg13g2_fill_8 FILLER_218_1256 ();
 sg13g2_fill_8 FILLER_218_1264 ();
 sg13g2_fill_8 FILLER_218_1272 ();
 sg13g2_fill_8 FILLER_218_1280 ();
 sg13g2_fill_8 FILLER_218_1288 ();
 sg13g2_fill_8 FILLER_218_1296 ();
 sg13g2_fill_8 FILLER_218_1304 ();
 sg13g2_fill_8 FILLER_218_1312 ();
 sg13g2_fill_8 FILLER_218_1320 ();
 sg13g2_fill_8 FILLER_218_1328 ();
 sg13g2_fill_8 FILLER_218_1336 ();
 sg13g2_fill_8 FILLER_218_1344 ();
 sg13g2_fill_8 FILLER_218_1352 ();
 sg13g2_fill_8 FILLER_218_1360 ();
 sg13g2_fill_8 FILLER_218_1368 ();
 sg13g2_fill_8 FILLER_218_1376 ();
 sg13g2_fill_8 FILLER_218_1384 ();
 sg13g2_fill_8 FILLER_218_1392 ();
 sg13g2_fill_8 FILLER_218_1400 ();
 sg13g2_fill_8 FILLER_218_1408 ();
 sg13g2_fill_8 FILLER_218_1416 ();
 sg13g2_fill_8 FILLER_218_1424 ();
 sg13g2_fill_8 FILLER_218_1432 ();
 sg13g2_fill_8 FILLER_218_1440 ();
 sg13g2_fill_8 FILLER_218_1448 ();
 sg13g2_fill_8 FILLER_218_1456 ();
 sg13g2_fill_8 FILLER_218_1464 ();
 sg13g2_fill_8 FILLER_218_1472 ();
 sg13g2_fill_8 FILLER_218_1480 ();
 sg13g2_fill_8 FILLER_218_1488 ();
 sg13g2_fill_8 FILLER_218_1496 ();
 sg13g2_fill_8 FILLER_218_1504 ();
 sg13g2_fill_8 FILLER_218_1512 ();
 sg13g2_fill_8 FILLER_218_1520 ();
 sg13g2_fill_8 FILLER_218_1528 ();
 sg13g2_fill_8 FILLER_218_1536 ();
 sg13g2_fill_8 FILLER_218_1544 ();
 sg13g2_fill_8 FILLER_218_1552 ();
 sg13g2_fill_8 FILLER_218_1560 ();
 sg13g2_fill_8 FILLER_218_1568 ();
 sg13g2_fill_8 FILLER_218_1576 ();
 sg13g2_fill_8 FILLER_218_1584 ();
 sg13g2_fill_8 FILLER_219_0 ();
 sg13g2_fill_8 FILLER_219_8 ();
 sg13g2_fill_8 FILLER_219_16 ();
 sg13g2_fill_8 FILLER_219_24 ();
 sg13g2_fill_8 FILLER_219_32 ();
 sg13g2_fill_8 FILLER_219_40 ();
 sg13g2_fill_8 FILLER_219_48 ();
 sg13g2_fill_8 FILLER_219_56 ();
 sg13g2_fill_8 FILLER_219_64 ();
 sg13g2_fill_8 FILLER_219_72 ();
 sg13g2_fill_8 FILLER_219_80 ();
 sg13g2_fill_8 FILLER_219_88 ();
 sg13g2_fill_8 FILLER_219_96 ();
 sg13g2_fill_8 FILLER_219_104 ();
 sg13g2_fill_8 FILLER_219_112 ();
 sg13g2_fill_8 FILLER_219_120 ();
 sg13g2_fill_8 FILLER_219_128 ();
 sg13g2_fill_8 FILLER_219_136 ();
 sg13g2_fill_8 FILLER_219_144 ();
 sg13g2_fill_8 FILLER_219_152 ();
 sg13g2_fill_8 FILLER_219_160 ();
 sg13g2_fill_8 FILLER_219_168 ();
 sg13g2_fill_8 FILLER_219_176 ();
 sg13g2_fill_8 FILLER_219_184 ();
 sg13g2_fill_8 FILLER_219_192 ();
 sg13g2_fill_8 FILLER_219_200 ();
 sg13g2_fill_8 FILLER_219_208 ();
 sg13g2_fill_8 FILLER_219_216 ();
 sg13g2_fill_8 FILLER_219_224 ();
 sg13g2_fill_8 FILLER_219_232 ();
 sg13g2_fill_8 FILLER_219_240 ();
 sg13g2_fill_8 FILLER_219_248 ();
 sg13g2_fill_8 FILLER_219_256 ();
 sg13g2_fill_8 FILLER_219_264 ();
 sg13g2_fill_8 FILLER_219_272 ();
 sg13g2_fill_8 FILLER_219_280 ();
 sg13g2_fill_8 FILLER_219_288 ();
 sg13g2_fill_8 FILLER_219_296 ();
 sg13g2_fill_8 FILLER_219_304 ();
 sg13g2_fill_8 FILLER_219_312 ();
 sg13g2_fill_8 FILLER_219_320 ();
 sg13g2_fill_8 FILLER_219_328 ();
 sg13g2_fill_8 FILLER_219_336 ();
 sg13g2_fill_8 FILLER_219_344 ();
 sg13g2_fill_8 FILLER_219_352 ();
 sg13g2_fill_8 FILLER_219_360 ();
 sg13g2_fill_8 FILLER_219_368 ();
 sg13g2_fill_8 FILLER_219_376 ();
 sg13g2_fill_8 FILLER_219_384 ();
 sg13g2_fill_8 FILLER_219_392 ();
 sg13g2_fill_8 FILLER_219_400 ();
 sg13g2_fill_8 FILLER_219_408 ();
 sg13g2_fill_8 FILLER_219_416 ();
 sg13g2_fill_8 FILLER_219_424 ();
 sg13g2_fill_8 FILLER_219_432 ();
 sg13g2_fill_8 FILLER_219_440 ();
 sg13g2_fill_8 FILLER_219_448 ();
 sg13g2_fill_8 FILLER_219_456 ();
 sg13g2_fill_8 FILLER_219_464 ();
 sg13g2_fill_8 FILLER_219_472 ();
 sg13g2_fill_8 FILLER_219_480 ();
 sg13g2_fill_8 FILLER_219_488 ();
 sg13g2_fill_8 FILLER_219_496 ();
 sg13g2_fill_8 FILLER_219_504 ();
 sg13g2_fill_8 FILLER_219_512 ();
 sg13g2_fill_8 FILLER_219_520 ();
 sg13g2_fill_8 FILLER_219_528 ();
 sg13g2_fill_8 FILLER_219_536 ();
 sg13g2_fill_8 FILLER_219_544 ();
 sg13g2_fill_8 FILLER_219_552 ();
 sg13g2_fill_8 FILLER_219_560 ();
 sg13g2_fill_8 FILLER_219_568 ();
 sg13g2_fill_8 FILLER_219_576 ();
 sg13g2_fill_8 FILLER_219_584 ();
 sg13g2_fill_8 FILLER_219_592 ();
 sg13g2_fill_8 FILLER_219_600 ();
 sg13g2_fill_8 FILLER_219_608 ();
 sg13g2_fill_8 FILLER_219_616 ();
 sg13g2_fill_8 FILLER_219_624 ();
 sg13g2_fill_8 FILLER_219_632 ();
 sg13g2_fill_8 FILLER_219_640 ();
 sg13g2_fill_8 FILLER_219_648 ();
 sg13g2_fill_8 FILLER_219_656 ();
 sg13g2_fill_8 FILLER_219_664 ();
 sg13g2_fill_8 FILLER_219_672 ();
 sg13g2_fill_8 FILLER_219_680 ();
 sg13g2_fill_8 FILLER_219_688 ();
 sg13g2_fill_8 FILLER_219_696 ();
 sg13g2_fill_8 FILLER_219_704 ();
 sg13g2_fill_8 FILLER_219_712 ();
 sg13g2_fill_8 FILLER_219_720 ();
 sg13g2_fill_8 FILLER_219_728 ();
 sg13g2_fill_8 FILLER_219_736 ();
 sg13g2_fill_8 FILLER_219_744 ();
 sg13g2_fill_8 FILLER_219_752 ();
 sg13g2_fill_8 FILLER_219_760 ();
 sg13g2_fill_8 FILLER_219_768 ();
 sg13g2_fill_8 FILLER_219_776 ();
 sg13g2_fill_8 FILLER_219_784 ();
 sg13g2_fill_8 FILLER_219_792 ();
 sg13g2_fill_8 FILLER_219_800 ();
 sg13g2_fill_8 FILLER_219_808 ();
 sg13g2_fill_8 FILLER_219_816 ();
 sg13g2_fill_8 FILLER_219_824 ();
 sg13g2_fill_8 FILLER_219_832 ();
 sg13g2_fill_8 FILLER_219_840 ();
 sg13g2_fill_8 FILLER_219_848 ();
 sg13g2_fill_8 FILLER_219_856 ();
 sg13g2_fill_8 FILLER_219_864 ();
 sg13g2_fill_8 FILLER_219_872 ();
 sg13g2_fill_8 FILLER_219_880 ();
 sg13g2_fill_8 FILLER_219_888 ();
 sg13g2_fill_8 FILLER_219_896 ();
 sg13g2_fill_8 FILLER_219_904 ();
 sg13g2_fill_8 FILLER_219_912 ();
 sg13g2_fill_8 FILLER_219_920 ();
 sg13g2_fill_8 FILLER_219_928 ();
 sg13g2_fill_8 FILLER_219_936 ();
 sg13g2_fill_8 FILLER_219_944 ();
 sg13g2_fill_8 FILLER_219_952 ();
 sg13g2_fill_8 FILLER_219_960 ();
 sg13g2_fill_8 FILLER_219_968 ();
 sg13g2_fill_8 FILLER_219_976 ();
 sg13g2_fill_8 FILLER_219_984 ();
 sg13g2_fill_8 FILLER_219_992 ();
 sg13g2_fill_8 FILLER_219_1000 ();
 sg13g2_fill_8 FILLER_219_1008 ();
 sg13g2_fill_8 FILLER_219_1016 ();
 sg13g2_fill_8 FILLER_219_1024 ();
 sg13g2_fill_8 FILLER_219_1032 ();
 sg13g2_fill_8 FILLER_219_1040 ();
 sg13g2_fill_8 FILLER_219_1048 ();
 sg13g2_fill_8 FILLER_219_1056 ();
 sg13g2_fill_8 FILLER_219_1064 ();
 sg13g2_fill_8 FILLER_219_1072 ();
 sg13g2_fill_8 FILLER_219_1080 ();
 sg13g2_fill_8 FILLER_219_1088 ();
 sg13g2_fill_8 FILLER_219_1096 ();
 sg13g2_fill_8 FILLER_219_1104 ();
 sg13g2_fill_8 FILLER_219_1112 ();
 sg13g2_fill_8 FILLER_219_1120 ();
 sg13g2_fill_8 FILLER_219_1128 ();
 sg13g2_fill_8 FILLER_219_1136 ();
 sg13g2_fill_8 FILLER_219_1144 ();
 sg13g2_fill_8 FILLER_219_1152 ();
 sg13g2_fill_8 FILLER_219_1160 ();
 sg13g2_fill_8 FILLER_219_1168 ();
 sg13g2_fill_8 FILLER_219_1176 ();
 sg13g2_fill_8 FILLER_219_1184 ();
 sg13g2_fill_8 FILLER_219_1192 ();
 sg13g2_fill_8 FILLER_219_1200 ();
 sg13g2_fill_8 FILLER_219_1208 ();
 sg13g2_fill_8 FILLER_219_1216 ();
 sg13g2_fill_8 FILLER_219_1224 ();
 sg13g2_fill_8 FILLER_219_1232 ();
 sg13g2_fill_8 FILLER_219_1240 ();
 sg13g2_fill_8 FILLER_219_1248 ();
 sg13g2_fill_8 FILLER_219_1256 ();
 sg13g2_fill_8 FILLER_219_1264 ();
 sg13g2_fill_8 FILLER_219_1272 ();
 sg13g2_fill_8 FILLER_219_1280 ();
 sg13g2_fill_8 FILLER_219_1288 ();
 sg13g2_fill_8 FILLER_219_1296 ();
 sg13g2_fill_8 FILLER_219_1304 ();
 sg13g2_fill_8 FILLER_219_1312 ();
 sg13g2_fill_8 FILLER_219_1320 ();
 sg13g2_fill_8 FILLER_219_1328 ();
 sg13g2_fill_8 FILLER_219_1336 ();
 sg13g2_fill_8 FILLER_219_1344 ();
 sg13g2_fill_8 FILLER_219_1352 ();
 sg13g2_fill_8 FILLER_219_1360 ();
 sg13g2_fill_8 FILLER_219_1368 ();
 sg13g2_fill_8 FILLER_219_1376 ();
 sg13g2_fill_8 FILLER_219_1384 ();
 sg13g2_fill_8 FILLER_219_1392 ();
 sg13g2_fill_8 FILLER_219_1400 ();
 sg13g2_fill_8 FILLER_219_1408 ();
 sg13g2_fill_8 FILLER_219_1416 ();
 sg13g2_fill_8 FILLER_219_1424 ();
 sg13g2_fill_8 FILLER_219_1432 ();
 sg13g2_fill_8 FILLER_219_1440 ();
 sg13g2_fill_8 FILLER_219_1448 ();
 sg13g2_fill_8 FILLER_219_1456 ();
 sg13g2_fill_8 FILLER_219_1464 ();
 sg13g2_fill_8 FILLER_219_1472 ();
 sg13g2_fill_8 FILLER_219_1480 ();
 sg13g2_fill_8 FILLER_219_1488 ();
 sg13g2_fill_8 FILLER_219_1496 ();
 sg13g2_fill_8 FILLER_219_1504 ();
 sg13g2_fill_8 FILLER_219_1512 ();
 sg13g2_fill_8 FILLER_219_1520 ();
 sg13g2_fill_8 FILLER_219_1528 ();
 sg13g2_fill_8 FILLER_219_1536 ();
 sg13g2_fill_8 FILLER_219_1544 ();
 sg13g2_fill_8 FILLER_219_1552 ();
 sg13g2_fill_8 FILLER_219_1560 ();
 sg13g2_fill_8 FILLER_219_1568 ();
 sg13g2_fill_8 FILLER_219_1576 ();
 sg13g2_fill_8 FILLER_219_1584 ();
 sg13g2_fill_8 FILLER_220_0 ();
 sg13g2_fill_8 FILLER_220_8 ();
 sg13g2_fill_8 FILLER_220_16 ();
 sg13g2_fill_8 FILLER_220_24 ();
 sg13g2_fill_8 FILLER_220_32 ();
 sg13g2_fill_8 FILLER_220_40 ();
 sg13g2_fill_8 FILLER_220_48 ();
 sg13g2_fill_8 FILLER_220_56 ();
 sg13g2_fill_8 FILLER_220_64 ();
 sg13g2_fill_8 FILLER_220_72 ();
 sg13g2_fill_8 FILLER_220_80 ();
 sg13g2_fill_8 FILLER_220_88 ();
 sg13g2_fill_8 FILLER_220_96 ();
 sg13g2_fill_8 FILLER_220_104 ();
 sg13g2_fill_8 FILLER_220_112 ();
 sg13g2_fill_8 FILLER_220_120 ();
 sg13g2_fill_8 FILLER_220_128 ();
 sg13g2_fill_8 FILLER_220_136 ();
 sg13g2_fill_8 FILLER_220_144 ();
 sg13g2_fill_8 FILLER_220_152 ();
 sg13g2_fill_8 FILLER_220_160 ();
 sg13g2_fill_8 FILLER_220_168 ();
 sg13g2_fill_8 FILLER_220_176 ();
 sg13g2_fill_8 FILLER_220_184 ();
 sg13g2_fill_8 FILLER_220_192 ();
 sg13g2_fill_8 FILLER_220_200 ();
 sg13g2_fill_8 FILLER_220_208 ();
 sg13g2_fill_8 FILLER_220_216 ();
 sg13g2_fill_8 FILLER_220_224 ();
 sg13g2_fill_8 FILLER_220_232 ();
 sg13g2_fill_8 FILLER_220_240 ();
 sg13g2_fill_8 FILLER_220_248 ();
 sg13g2_fill_8 FILLER_220_256 ();
 sg13g2_fill_8 FILLER_220_264 ();
 sg13g2_fill_8 FILLER_220_272 ();
 sg13g2_fill_8 FILLER_220_280 ();
 sg13g2_fill_8 FILLER_220_288 ();
 sg13g2_fill_8 FILLER_220_296 ();
 sg13g2_fill_8 FILLER_220_304 ();
 sg13g2_fill_8 FILLER_220_312 ();
 sg13g2_fill_8 FILLER_220_320 ();
 sg13g2_fill_8 FILLER_220_328 ();
 sg13g2_fill_8 FILLER_220_336 ();
 sg13g2_fill_8 FILLER_220_344 ();
 sg13g2_fill_8 FILLER_220_352 ();
 sg13g2_fill_8 FILLER_220_360 ();
 sg13g2_fill_8 FILLER_220_368 ();
 sg13g2_fill_8 FILLER_220_376 ();
 sg13g2_fill_8 FILLER_220_384 ();
 sg13g2_fill_8 FILLER_220_392 ();
 sg13g2_fill_8 FILLER_220_400 ();
 sg13g2_fill_8 FILLER_220_408 ();
 sg13g2_fill_8 FILLER_220_416 ();
 sg13g2_fill_8 FILLER_220_424 ();
 sg13g2_fill_8 FILLER_220_432 ();
 sg13g2_fill_8 FILLER_220_440 ();
 sg13g2_fill_8 FILLER_220_448 ();
 sg13g2_fill_8 FILLER_220_456 ();
 sg13g2_fill_8 FILLER_220_464 ();
 sg13g2_fill_8 FILLER_220_472 ();
 sg13g2_fill_8 FILLER_220_480 ();
 sg13g2_fill_8 FILLER_220_488 ();
 sg13g2_fill_8 FILLER_220_496 ();
 sg13g2_fill_8 FILLER_220_504 ();
 sg13g2_fill_8 FILLER_220_512 ();
 sg13g2_fill_8 FILLER_220_520 ();
 sg13g2_fill_8 FILLER_220_528 ();
 sg13g2_fill_8 FILLER_220_536 ();
 sg13g2_fill_8 FILLER_220_544 ();
 sg13g2_fill_8 FILLER_220_552 ();
 sg13g2_fill_8 FILLER_220_560 ();
 sg13g2_fill_8 FILLER_220_568 ();
 sg13g2_fill_8 FILLER_220_576 ();
 sg13g2_fill_8 FILLER_220_584 ();
 sg13g2_fill_8 FILLER_220_592 ();
 sg13g2_fill_8 FILLER_220_600 ();
 sg13g2_fill_8 FILLER_220_608 ();
 sg13g2_fill_8 FILLER_220_616 ();
 sg13g2_fill_8 FILLER_220_624 ();
 sg13g2_fill_8 FILLER_220_632 ();
 sg13g2_fill_8 FILLER_220_640 ();
 sg13g2_fill_8 FILLER_220_648 ();
 sg13g2_fill_8 FILLER_220_656 ();
 sg13g2_fill_8 FILLER_220_664 ();
 sg13g2_fill_8 FILLER_220_672 ();
 sg13g2_fill_8 FILLER_220_680 ();
 sg13g2_fill_8 FILLER_220_688 ();
 sg13g2_fill_8 FILLER_220_696 ();
 sg13g2_fill_8 FILLER_220_704 ();
 sg13g2_fill_8 FILLER_220_712 ();
 sg13g2_fill_8 FILLER_220_720 ();
 sg13g2_fill_8 FILLER_220_728 ();
 sg13g2_fill_8 FILLER_220_736 ();
 sg13g2_fill_8 FILLER_220_744 ();
 sg13g2_fill_8 FILLER_220_752 ();
 sg13g2_fill_8 FILLER_220_760 ();
 sg13g2_fill_8 FILLER_220_768 ();
 sg13g2_fill_8 FILLER_220_776 ();
 sg13g2_fill_8 FILLER_220_784 ();
 sg13g2_fill_8 FILLER_220_792 ();
 sg13g2_fill_8 FILLER_220_800 ();
 sg13g2_fill_8 FILLER_220_808 ();
 sg13g2_fill_8 FILLER_220_816 ();
 sg13g2_fill_8 FILLER_220_824 ();
 sg13g2_fill_8 FILLER_220_832 ();
 sg13g2_fill_8 FILLER_220_840 ();
 sg13g2_fill_8 FILLER_220_848 ();
 sg13g2_fill_8 FILLER_220_856 ();
 sg13g2_fill_8 FILLER_220_864 ();
 sg13g2_fill_8 FILLER_220_872 ();
 sg13g2_fill_8 FILLER_220_880 ();
 sg13g2_fill_8 FILLER_220_888 ();
 sg13g2_fill_8 FILLER_220_896 ();
 sg13g2_fill_8 FILLER_220_904 ();
 sg13g2_fill_8 FILLER_220_912 ();
 sg13g2_fill_8 FILLER_220_920 ();
 sg13g2_fill_8 FILLER_220_928 ();
 sg13g2_fill_8 FILLER_220_936 ();
 sg13g2_fill_8 FILLER_220_944 ();
 sg13g2_fill_8 FILLER_220_952 ();
 sg13g2_fill_8 FILLER_220_960 ();
 sg13g2_fill_8 FILLER_220_968 ();
 sg13g2_fill_8 FILLER_220_976 ();
 sg13g2_fill_8 FILLER_220_984 ();
 sg13g2_fill_8 FILLER_220_992 ();
 sg13g2_fill_8 FILLER_220_1000 ();
 sg13g2_fill_8 FILLER_220_1008 ();
 sg13g2_fill_8 FILLER_220_1016 ();
 sg13g2_fill_8 FILLER_220_1024 ();
 sg13g2_fill_8 FILLER_220_1032 ();
 sg13g2_fill_8 FILLER_220_1040 ();
 sg13g2_fill_8 FILLER_220_1048 ();
 sg13g2_fill_8 FILLER_220_1056 ();
 sg13g2_fill_8 FILLER_220_1064 ();
 sg13g2_fill_8 FILLER_220_1072 ();
 sg13g2_fill_8 FILLER_220_1080 ();
 sg13g2_fill_8 FILLER_220_1088 ();
 sg13g2_fill_8 FILLER_220_1096 ();
 sg13g2_fill_8 FILLER_220_1104 ();
 sg13g2_fill_8 FILLER_220_1112 ();
 sg13g2_fill_8 FILLER_220_1120 ();
 sg13g2_fill_8 FILLER_220_1128 ();
 sg13g2_fill_8 FILLER_220_1136 ();
 sg13g2_fill_8 FILLER_220_1144 ();
 sg13g2_fill_8 FILLER_220_1152 ();
 sg13g2_fill_8 FILLER_220_1160 ();
 sg13g2_fill_8 FILLER_220_1168 ();
 sg13g2_fill_8 FILLER_220_1176 ();
 sg13g2_fill_8 FILLER_220_1184 ();
 sg13g2_fill_8 FILLER_220_1192 ();
 sg13g2_fill_8 FILLER_220_1200 ();
 sg13g2_fill_8 FILLER_220_1208 ();
 sg13g2_fill_8 FILLER_220_1216 ();
 sg13g2_fill_8 FILLER_220_1224 ();
 sg13g2_fill_8 FILLER_220_1232 ();
 sg13g2_fill_8 FILLER_220_1240 ();
 sg13g2_fill_8 FILLER_220_1248 ();
 sg13g2_fill_8 FILLER_220_1256 ();
 sg13g2_fill_8 FILLER_220_1264 ();
 sg13g2_fill_8 FILLER_220_1272 ();
 sg13g2_fill_8 FILLER_220_1280 ();
 sg13g2_fill_8 FILLER_220_1288 ();
 sg13g2_fill_8 FILLER_220_1296 ();
 sg13g2_fill_8 FILLER_220_1304 ();
 sg13g2_fill_8 FILLER_220_1312 ();
 sg13g2_fill_8 FILLER_220_1320 ();
 sg13g2_fill_8 FILLER_220_1328 ();
 sg13g2_fill_8 FILLER_220_1336 ();
 sg13g2_fill_8 FILLER_220_1344 ();
 sg13g2_fill_8 FILLER_220_1352 ();
 sg13g2_fill_8 FILLER_220_1360 ();
 sg13g2_fill_8 FILLER_220_1368 ();
 sg13g2_fill_8 FILLER_220_1376 ();
 sg13g2_fill_8 FILLER_220_1384 ();
 sg13g2_fill_8 FILLER_220_1392 ();
 sg13g2_fill_8 FILLER_220_1400 ();
 sg13g2_fill_8 FILLER_220_1408 ();
 sg13g2_fill_8 FILLER_220_1416 ();
 sg13g2_fill_8 FILLER_220_1424 ();
 sg13g2_fill_8 FILLER_220_1432 ();
 sg13g2_fill_8 FILLER_220_1440 ();
 sg13g2_fill_8 FILLER_220_1448 ();
 sg13g2_fill_8 FILLER_220_1456 ();
 sg13g2_fill_8 FILLER_220_1464 ();
 sg13g2_fill_8 FILLER_220_1472 ();
 sg13g2_fill_8 FILLER_220_1480 ();
 sg13g2_fill_8 FILLER_220_1488 ();
 sg13g2_fill_8 FILLER_220_1496 ();
 sg13g2_fill_8 FILLER_220_1504 ();
 sg13g2_fill_8 FILLER_220_1512 ();
 sg13g2_fill_8 FILLER_220_1520 ();
 sg13g2_fill_8 FILLER_220_1528 ();
 sg13g2_fill_8 FILLER_220_1536 ();
 sg13g2_fill_8 FILLER_220_1544 ();
 sg13g2_fill_8 FILLER_220_1552 ();
 sg13g2_fill_8 FILLER_220_1560 ();
 sg13g2_fill_8 FILLER_220_1568 ();
 sg13g2_fill_8 FILLER_220_1576 ();
 sg13g2_fill_8 FILLER_220_1584 ();
 sg13g2_fill_8 FILLER_221_0 ();
 sg13g2_fill_8 FILLER_221_8 ();
 sg13g2_fill_8 FILLER_221_16 ();
 sg13g2_fill_8 FILLER_221_24 ();
 sg13g2_fill_8 FILLER_221_32 ();
 sg13g2_fill_8 FILLER_221_40 ();
 sg13g2_fill_8 FILLER_221_48 ();
 sg13g2_fill_8 FILLER_221_56 ();
 sg13g2_fill_8 FILLER_221_64 ();
 sg13g2_fill_8 FILLER_221_72 ();
 sg13g2_fill_8 FILLER_221_80 ();
 sg13g2_fill_8 FILLER_221_88 ();
 sg13g2_fill_8 FILLER_221_96 ();
 sg13g2_fill_8 FILLER_221_104 ();
 sg13g2_fill_8 FILLER_221_112 ();
 sg13g2_fill_8 FILLER_221_120 ();
 sg13g2_fill_8 FILLER_221_128 ();
 sg13g2_fill_8 FILLER_221_136 ();
 sg13g2_fill_8 FILLER_221_144 ();
 sg13g2_fill_8 FILLER_221_152 ();
 sg13g2_fill_8 FILLER_221_160 ();
 sg13g2_fill_8 FILLER_221_168 ();
 sg13g2_fill_8 FILLER_221_176 ();
 sg13g2_fill_8 FILLER_221_184 ();
 sg13g2_fill_8 FILLER_221_192 ();
 sg13g2_fill_8 FILLER_221_200 ();
 sg13g2_fill_8 FILLER_221_208 ();
 sg13g2_fill_8 FILLER_221_216 ();
 sg13g2_fill_8 FILLER_221_224 ();
 sg13g2_fill_8 FILLER_221_232 ();
 sg13g2_fill_8 FILLER_221_240 ();
 sg13g2_fill_8 FILLER_221_248 ();
 sg13g2_fill_8 FILLER_221_256 ();
 sg13g2_fill_8 FILLER_221_264 ();
 sg13g2_fill_8 FILLER_221_272 ();
 sg13g2_fill_8 FILLER_221_280 ();
 sg13g2_fill_8 FILLER_221_288 ();
 sg13g2_fill_8 FILLER_221_296 ();
 sg13g2_fill_8 FILLER_221_304 ();
 sg13g2_fill_8 FILLER_221_312 ();
 sg13g2_fill_8 FILLER_221_320 ();
 sg13g2_fill_8 FILLER_221_328 ();
 sg13g2_fill_8 FILLER_221_336 ();
 sg13g2_fill_8 FILLER_221_344 ();
 sg13g2_fill_8 FILLER_221_352 ();
 sg13g2_fill_8 FILLER_221_360 ();
 sg13g2_fill_8 FILLER_221_368 ();
 sg13g2_fill_8 FILLER_221_376 ();
 sg13g2_fill_8 FILLER_221_384 ();
 sg13g2_fill_8 FILLER_221_392 ();
 sg13g2_fill_8 FILLER_221_400 ();
 sg13g2_fill_8 FILLER_221_408 ();
 sg13g2_fill_8 FILLER_221_416 ();
 sg13g2_fill_8 FILLER_221_424 ();
 sg13g2_fill_8 FILLER_221_432 ();
 sg13g2_fill_8 FILLER_221_440 ();
 sg13g2_fill_8 FILLER_221_448 ();
 sg13g2_fill_8 FILLER_221_456 ();
 sg13g2_fill_8 FILLER_221_464 ();
 sg13g2_fill_8 FILLER_221_472 ();
 sg13g2_fill_8 FILLER_221_480 ();
 sg13g2_fill_8 FILLER_221_488 ();
 sg13g2_fill_8 FILLER_221_496 ();
 sg13g2_fill_8 FILLER_221_504 ();
 sg13g2_fill_8 FILLER_221_512 ();
 sg13g2_fill_8 FILLER_221_520 ();
 sg13g2_fill_8 FILLER_221_528 ();
 sg13g2_fill_8 FILLER_221_536 ();
 sg13g2_fill_8 FILLER_221_544 ();
 sg13g2_fill_8 FILLER_221_552 ();
 sg13g2_fill_8 FILLER_221_560 ();
 sg13g2_fill_8 FILLER_221_568 ();
 sg13g2_fill_8 FILLER_221_576 ();
 sg13g2_fill_8 FILLER_221_584 ();
 sg13g2_fill_8 FILLER_221_592 ();
 sg13g2_fill_8 FILLER_221_600 ();
 sg13g2_fill_8 FILLER_221_608 ();
 sg13g2_fill_8 FILLER_221_616 ();
 sg13g2_fill_8 FILLER_221_624 ();
 sg13g2_fill_8 FILLER_221_632 ();
 sg13g2_fill_8 FILLER_221_640 ();
 sg13g2_fill_8 FILLER_221_648 ();
 sg13g2_fill_8 FILLER_221_656 ();
 sg13g2_fill_8 FILLER_221_664 ();
 sg13g2_fill_8 FILLER_221_672 ();
 sg13g2_fill_8 FILLER_221_680 ();
 sg13g2_fill_8 FILLER_221_688 ();
 sg13g2_fill_8 FILLER_221_696 ();
 sg13g2_fill_8 FILLER_221_704 ();
 sg13g2_fill_8 FILLER_221_712 ();
 sg13g2_fill_8 FILLER_221_720 ();
 sg13g2_fill_8 FILLER_221_728 ();
 sg13g2_fill_8 FILLER_221_736 ();
 sg13g2_fill_8 FILLER_221_744 ();
 sg13g2_fill_8 FILLER_221_752 ();
 sg13g2_fill_8 FILLER_221_760 ();
 sg13g2_fill_8 FILLER_221_768 ();
 sg13g2_fill_8 FILLER_221_776 ();
 sg13g2_fill_8 FILLER_221_784 ();
 sg13g2_fill_8 FILLER_221_792 ();
 sg13g2_fill_8 FILLER_221_800 ();
 sg13g2_fill_8 FILLER_221_808 ();
 sg13g2_fill_8 FILLER_221_816 ();
 sg13g2_fill_8 FILLER_221_824 ();
 sg13g2_fill_8 FILLER_221_832 ();
 sg13g2_fill_8 FILLER_221_840 ();
 sg13g2_fill_8 FILLER_221_848 ();
 sg13g2_fill_8 FILLER_221_856 ();
 sg13g2_fill_8 FILLER_221_864 ();
 sg13g2_fill_8 FILLER_221_872 ();
 sg13g2_fill_8 FILLER_221_880 ();
 sg13g2_fill_8 FILLER_221_888 ();
 sg13g2_fill_8 FILLER_221_896 ();
 sg13g2_fill_8 FILLER_221_904 ();
 sg13g2_fill_8 FILLER_221_912 ();
 sg13g2_fill_8 FILLER_221_920 ();
 sg13g2_fill_8 FILLER_221_928 ();
 sg13g2_fill_8 FILLER_221_936 ();
 sg13g2_fill_8 FILLER_221_944 ();
 sg13g2_fill_8 FILLER_221_952 ();
 sg13g2_fill_8 FILLER_221_960 ();
 sg13g2_fill_8 FILLER_221_968 ();
 sg13g2_fill_8 FILLER_221_976 ();
 sg13g2_fill_8 FILLER_221_984 ();
 sg13g2_fill_8 FILLER_221_992 ();
 sg13g2_fill_8 FILLER_221_1000 ();
 sg13g2_fill_8 FILLER_221_1008 ();
 sg13g2_fill_8 FILLER_221_1016 ();
 sg13g2_fill_8 FILLER_221_1024 ();
 sg13g2_fill_8 FILLER_221_1032 ();
 sg13g2_fill_8 FILLER_221_1040 ();
 sg13g2_fill_8 FILLER_221_1048 ();
 sg13g2_fill_8 FILLER_221_1056 ();
 sg13g2_fill_8 FILLER_221_1064 ();
 sg13g2_fill_8 FILLER_221_1072 ();
 sg13g2_fill_8 FILLER_221_1080 ();
 sg13g2_fill_8 FILLER_221_1088 ();
 sg13g2_fill_8 FILLER_221_1096 ();
 sg13g2_fill_8 FILLER_221_1104 ();
 sg13g2_fill_8 FILLER_221_1112 ();
 sg13g2_fill_8 FILLER_221_1120 ();
 sg13g2_fill_8 FILLER_221_1128 ();
 sg13g2_fill_8 FILLER_221_1136 ();
 sg13g2_fill_8 FILLER_221_1144 ();
 sg13g2_fill_8 FILLER_221_1152 ();
 sg13g2_fill_8 FILLER_221_1160 ();
 sg13g2_fill_8 FILLER_221_1168 ();
 sg13g2_fill_8 FILLER_221_1176 ();
 sg13g2_fill_8 FILLER_221_1184 ();
 sg13g2_fill_8 FILLER_221_1192 ();
 sg13g2_fill_8 FILLER_221_1200 ();
 sg13g2_fill_8 FILLER_221_1208 ();
 sg13g2_fill_8 FILLER_221_1216 ();
 sg13g2_fill_8 FILLER_221_1224 ();
 sg13g2_fill_8 FILLER_221_1232 ();
 sg13g2_fill_8 FILLER_221_1240 ();
 sg13g2_fill_8 FILLER_221_1248 ();
 sg13g2_fill_8 FILLER_221_1256 ();
 sg13g2_fill_8 FILLER_221_1264 ();
 sg13g2_fill_8 FILLER_221_1272 ();
 sg13g2_fill_8 FILLER_221_1280 ();
 sg13g2_fill_8 FILLER_221_1288 ();
 sg13g2_fill_8 FILLER_221_1296 ();
 sg13g2_fill_8 FILLER_221_1304 ();
 sg13g2_fill_8 FILLER_221_1312 ();
 sg13g2_fill_8 FILLER_221_1320 ();
 sg13g2_fill_8 FILLER_221_1328 ();
 sg13g2_fill_8 FILLER_221_1336 ();
 sg13g2_fill_8 FILLER_221_1344 ();
 sg13g2_fill_8 FILLER_221_1352 ();
 sg13g2_fill_8 FILLER_221_1360 ();
 sg13g2_fill_8 FILLER_221_1368 ();
 sg13g2_fill_8 FILLER_221_1376 ();
 sg13g2_fill_8 FILLER_221_1384 ();
 sg13g2_fill_8 FILLER_221_1392 ();
 sg13g2_fill_8 FILLER_221_1400 ();
 sg13g2_fill_8 FILLER_221_1408 ();
 sg13g2_fill_8 FILLER_221_1416 ();
 sg13g2_fill_8 FILLER_221_1424 ();
 sg13g2_fill_8 FILLER_221_1432 ();
 sg13g2_fill_8 FILLER_221_1440 ();
 sg13g2_fill_8 FILLER_221_1448 ();
 sg13g2_fill_8 FILLER_221_1456 ();
 sg13g2_fill_8 FILLER_221_1464 ();
 sg13g2_fill_8 FILLER_221_1472 ();
 sg13g2_fill_8 FILLER_221_1480 ();
 sg13g2_fill_8 FILLER_221_1488 ();
 sg13g2_fill_8 FILLER_221_1496 ();
 sg13g2_fill_8 FILLER_221_1504 ();
 sg13g2_fill_8 FILLER_221_1512 ();
 sg13g2_fill_8 FILLER_221_1520 ();
 sg13g2_fill_8 FILLER_221_1528 ();
 sg13g2_fill_8 FILLER_221_1536 ();
 sg13g2_fill_8 FILLER_221_1544 ();
 sg13g2_fill_8 FILLER_221_1552 ();
 sg13g2_fill_8 FILLER_221_1560 ();
 sg13g2_fill_8 FILLER_221_1568 ();
 sg13g2_fill_8 FILLER_221_1576 ();
 sg13g2_fill_8 FILLER_221_1584 ();
 sg13g2_fill_8 FILLER_222_0 ();
 sg13g2_fill_8 FILLER_222_8 ();
 sg13g2_fill_8 FILLER_222_16 ();
 sg13g2_fill_8 FILLER_222_24 ();
 sg13g2_fill_8 FILLER_222_32 ();
 sg13g2_fill_8 FILLER_222_40 ();
 sg13g2_fill_8 FILLER_222_48 ();
 sg13g2_fill_8 FILLER_222_56 ();
 sg13g2_fill_8 FILLER_222_64 ();
 sg13g2_fill_8 FILLER_222_72 ();
 sg13g2_fill_8 FILLER_222_80 ();
 sg13g2_fill_8 FILLER_222_88 ();
 sg13g2_fill_8 FILLER_222_96 ();
 sg13g2_fill_8 FILLER_222_104 ();
 sg13g2_fill_8 FILLER_222_112 ();
 sg13g2_fill_8 FILLER_222_120 ();
 sg13g2_fill_8 FILLER_222_128 ();
 sg13g2_fill_8 FILLER_222_136 ();
 sg13g2_fill_8 FILLER_222_144 ();
 sg13g2_fill_8 FILLER_222_152 ();
 sg13g2_fill_8 FILLER_222_160 ();
 sg13g2_fill_8 FILLER_222_168 ();
 sg13g2_fill_8 FILLER_222_176 ();
 sg13g2_fill_8 FILLER_222_184 ();
 sg13g2_fill_8 FILLER_222_192 ();
 sg13g2_fill_8 FILLER_222_200 ();
 sg13g2_fill_8 FILLER_222_208 ();
 sg13g2_fill_8 FILLER_222_216 ();
 sg13g2_fill_8 FILLER_222_224 ();
 sg13g2_fill_8 FILLER_222_232 ();
 sg13g2_fill_8 FILLER_222_240 ();
 sg13g2_fill_8 FILLER_222_248 ();
 sg13g2_fill_8 FILLER_222_256 ();
 sg13g2_fill_8 FILLER_222_264 ();
 sg13g2_fill_8 FILLER_222_272 ();
 sg13g2_fill_8 FILLER_222_280 ();
 sg13g2_fill_8 FILLER_222_288 ();
 sg13g2_fill_8 FILLER_222_296 ();
 sg13g2_fill_8 FILLER_222_304 ();
 sg13g2_fill_8 FILLER_222_312 ();
 sg13g2_fill_8 FILLER_222_320 ();
 sg13g2_fill_8 FILLER_222_328 ();
 sg13g2_fill_8 FILLER_222_336 ();
 sg13g2_fill_8 FILLER_222_344 ();
 sg13g2_fill_8 FILLER_222_352 ();
 sg13g2_fill_8 FILLER_222_360 ();
 sg13g2_fill_8 FILLER_222_368 ();
 sg13g2_fill_8 FILLER_222_376 ();
 sg13g2_fill_8 FILLER_222_384 ();
 sg13g2_fill_8 FILLER_222_392 ();
 sg13g2_fill_8 FILLER_222_400 ();
 sg13g2_fill_8 FILLER_222_408 ();
 sg13g2_fill_8 FILLER_222_416 ();
 sg13g2_fill_8 FILLER_222_424 ();
 sg13g2_fill_8 FILLER_222_432 ();
 sg13g2_fill_8 FILLER_222_440 ();
 sg13g2_fill_8 FILLER_222_448 ();
 sg13g2_fill_8 FILLER_222_456 ();
 sg13g2_fill_8 FILLER_222_464 ();
 sg13g2_fill_8 FILLER_222_472 ();
 sg13g2_fill_8 FILLER_222_480 ();
 sg13g2_fill_8 FILLER_222_488 ();
 sg13g2_fill_8 FILLER_222_496 ();
 sg13g2_fill_8 FILLER_222_504 ();
 sg13g2_fill_8 FILLER_222_512 ();
 sg13g2_fill_8 FILLER_222_520 ();
 sg13g2_fill_8 FILLER_222_528 ();
 sg13g2_fill_8 FILLER_222_536 ();
 sg13g2_fill_8 FILLER_222_544 ();
 sg13g2_fill_8 FILLER_222_552 ();
 sg13g2_fill_8 FILLER_222_560 ();
 sg13g2_fill_8 FILLER_222_568 ();
 sg13g2_fill_8 FILLER_222_576 ();
 sg13g2_fill_8 FILLER_222_584 ();
 sg13g2_fill_8 FILLER_222_592 ();
 sg13g2_fill_8 FILLER_222_600 ();
 sg13g2_fill_8 FILLER_222_608 ();
 sg13g2_fill_8 FILLER_222_616 ();
 sg13g2_fill_8 FILLER_222_624 ();
 sg13g2_fill_8 FILLER_222_632 ();
 sg13g2_fill_8 FILLER_222_640 ();
 sg13g2_fill_8 FILLER_222_648 ();
 sg13g2_fill_8 FILLER_222_656 ();
 sg13g2_fill_8 FILLER_222_664 ();
 sg13g2_fill_8 FILLER_222_672 ();
 sg13g2_fill_8 FILLER_222_680 ();
 sg13g2_fill_8 FILLER_222_688 ();
 sg13g2_fill_8 FILLER_222_696 ();
 sg13g2_fill_8 FILLER_222_704 ();
 sg13g2_fill_8 FILLER_222_712 ();
 sg13g2_fill_8 FILLER_222_720 ();
 sg13g2_fill_8 FILLER_222_728 ();
 sg13g2_fill_8 FILLER_222_736 ();
 sg13g2_fill_8 FILLER_222_744 ();
 sg13g2_fill_8 FILLER_222_752 ();
 sg13g2_fill_8 FILLER_222_760 ();
 sg13g2_fill_8 FILLER_222_768 ();
 sg13g2_fill_8 FILLER_222_776 ();
 sg13g2_fill_8 FILLER_222_784 ();
 sg13g2_fill_8 FILLER_222_792 ();
 sg13g2_fill_8 FILLER_222_800 ();
 sg13g2_fill_8 FILLER_222_808 ();
 sg13g2_fill_8 FILLER_222_816 ();
 sg13g2_fill_8 FILLER_222_824 ();
 sg13g2_fill_8 FILLER_222_832 ();
 sg13g2_fill_8 FILLER_222_840 ();
 sg13g2_fill_8 FILLER_222_848 ();
 sg13g2_fill_8 FILLER_222_856 ();
 sg13g2_fill_8 FILLER_222_864 ();
 sg13g2_fill_8 FILLER_222_872 ();
 sg13g2_fill_8 FILLER_222_880 ();
 sg13g2_fill_8 FILLER_222_888 ();
 sg13g2_fill_8 FILLER_222_896 ();
 sg13g2_fill_8 FILLER_222_904 ();
 sg13g2_fill_8 FILLER_222_912 ();
 sg13g2_fill_8 FILLER_222_920 ();
 sg13g2_fill_8 FILLER_222_928 ();
 sg13g2_fill_8 FILLER_222_936 ();
 sg13g2_fill_8 FILLER_222_944 ();
 sg13g2_fill_8 FILLER_222_952 ();
 sg13g2_fill_8 FILLER_222_960 ();
 sg13g2_fill_8 FILLER_222_968 ();
 sg13g2_fill_8 FILLER_222_976 ();
 sg13g2_fill_8 FILLER_222_984 ();
 sg13g2_fill_8 FILLER_222_992 ();
 sg13g2_fill_8 FILLER_222_1000 ();
 sg13g2_fill_8 FILLER_222_1008 ();
 sg13g2_fill_8 FILLER_222_1016 ();
 sg13g2_fill_8 FILLER_222_1024 ();
 sg13g2_fill_8 FILLER_222_1032 ();
 sg13g2_fill_8 FILLER_222_1040 ();
 sg13g2_fill_8 FILLER_222_1048 ();
 sg13g2_fill_8 FILLER_222_1056 ();
 sg13g2_fill_8 FILLER_222_1064 ();
 sg13g2_fill_8 FILLER_222_1072 ();
 sg13g2_fill_8 FILLER_222_1080 ();
 sg13g2_fill_8 FILLER_222_1088 ();
 sg13g2_fill_8 FILLER_222_1096 ();
 sg13g2_fill_8 FILLER_222_1104 ();
 sg13g2_fill_8 FILLER_222_1112 ();
 sg13g2_fill_8 FILLER_222_1120 ();
 sg13g2_fill_8 FILLER_222_1128 ();
 sg13g2_fill_8 FILLER_222_1136 ();
 sg13g2_fill_8 FILLER_222_1144 ();
 sg13g2_fill_8 FILLER_222_1152 ();
 sg13g2_fill_8 FILLER_222_1160 ();
 sg13g2_fill_8 FILLER_222_1168 ();
 sg13g2_fill_8 FILLER_222_1176 ();
 sg13g2_fill_8 FILLER_222_1184 ();
 sg13g2_fill_8 FILLER_222_1192 ();
 sg13g2_fill_8 FILLER_222_1200 ();
 sg13g2_fill_8 FILLER_222_1208 ();
 sg13g2_fill_8 FILLER_222_1216 ();
 sg13g2_fill_8 FILLER_222_1224 ();
 sg13g2_fill_8 FILLER_222_1232 ();
 sg13g2_fill_8 FILLER_222_1240 ();
 sg13g2_fill_8 FILLER_222_1248 ();
 sg13g2_fill_8 FILLER_222_1256 ();
 sg13g2_fill_8 FILLER_222_1264 ();
 sg13g2_fill_8 FILLER_222_1272 ();
 sg13g2_fill_8 FILLER_222_1280 ();
 sg13g2_fill_8 FILLER_222_1288 ();
 sg13g2_fill_8 FILLER_222_1296 ();
 sg13g2_fill_8 FILLER_222_1304 ();
 sg13g2_fill_8 FILLER_222_1312 ();
 sg13g2_fill_8 FILLER_222_1320 ();
 sg13g2_fill_8 FILLER_222_1328 ();
 sg13g2_fill_8 FILLER_222_1336 ();
 sg13g2_fill_8 FILLER_222_1344 ();
 sg13g2_fill_8 FILLER_222_1352 ();
 sg13g2_fill_8 FILLER_222_1360 ();
 sg13g2_fill_8 FILLER_222_1368 ();
 sg13g2_fill_8 FILLER_222_1376 ();
 sg13g2_fill_8 FILLER_222_1384 ();
 sg13g2_fill_8 FILLER_222_1392 ();
 sg13g2_fill_8 FILLER_222_1400 ();
 sg13g2_fill_8 FILLER_222_1408 ();
 sg13g2_fill_8 FILLER_222_1416 ();
 sg13g2_fill_8 FILLER_222_1424 ();
 sg13g2_fill_8 FILLER_222_1432 ();
 sg13g2_fill_8 FILLER_222_1440 ();
 sg13g2_fill_8 FILLER_222_1448 ();
 sg13g2_fill_8 FILLER_222_1456 ();
 sg13g2_fill_8 FILLER_222_1464 ();
 sg13g2_fill_8 FILLER_222_1472 ();
 sg13g2_fill_8 FILLER_222_1480 ();
 sg13g2_fill_8 FILLER_222_1488 ();
 sg13g2_fill_8 FILLER_222_1496 ();
 sg13g2_fill_8 FILLER_222_1504 ();
 sg13g2_fill_8 FILLER_222_1512 ();
 sg13g2_fill_8 FILLER_222_1520 ();
 sg13g2_fill_8 FILLER_222_1528 ();
 sg13g2_fill_8 FILLER_222_1536 ();
 sg13g2_fill_8 FILLER_222_1544 ();
 sg13g2_fill_8 FILLER_222_1552 ();
 sg13g2_fill_8 FILLER_222_1560 ();
 sg13g2_fill_8 FILLER_222_1568 ();
 sg13g2_fill_8 FILLER_222_1576 ();
 sg13g2_fill_8 FILLER_222_1584 ();
 sg13g2_fill_8 FILLER_223_0 ();
 sg13g2_fill_8 FILLER_223_8 ();
 sg13g2_fill_8 FILLER_223_16 ();
 sg13g2_fill_8 FILLER_223_24 ();
 sg13g2_fill_8 FILLER_223_32 ();
 sg13g2_fill_8 FILLER_223_40 ();
 sg13g2_fill_8 FILLER_223_48 ();
 sg13g2_fill_8 FILLER_223_56 ();
 sg13g2_fill_8 FILLER_223_64 ();
 sg13g2_fill_8 FILLER_223_72 ();
 sg13g2_fill_8 FILLER_223_80 ();
 sg13g2_fill_8 FILLER_223_88 ();
 sg13g2_fill_8 FILLER_223_96 ();
 sg13g2_fill_8 FILLER_223_104 ();
 sg13g2_fill_8 FILLER_223_112 ();
 sg13g2_fill_8 FILLER_223_120 ();
 sg13g2_fill_8 FILLER_223_128 ();
 sg13g2_fill_8 FILLER_223_136 ();
 sg13g2_fill_8 FILLER_223_144 ();
 sg13g2_fill_8 FILLER_223_152 ();
 sg13g2_fill_8 FILLER_223_160 ();
 sg13g2_fill_8 FILLER_223_168 ();
 sg13g2_fill_8 FILLER_223_176 ();
 sg13g2_fill_8 FILLER_223_184 ();
 sg13g2_fill_8 FILLER_223_192 ();
 sg13g2_fill_8 FILLER_223_200 ();
 sg13g2_fill_8 FILLER_223_208 ();
 sg13g2_fill_8 FILLER_223_216 ();
 sg13g2_fill_8 FILLER_223_224 ();
 sg13g2_fill_8 FILLER_223_232 ();
 sg13g2_fill_8 FILLER_223_240 ();
 sg13g2_fill_8 FILLER_223_248 ();
 sg13g2_fill_8 FILLER_223_256 ();
 sg13g2_fill_8 FILLER_223_264 ();
 sg13g2_fill_8 FILLER_223_272 ();
 sg13g2_fill_8 FILLER_223_280 ();
 sg13g2_fill_8 FILLER_223_288 ();
 sg13g2_fill_8 FILLER_223_296 ();
 sg13g2_fill_8 FILLER_223_304 ();
 sg13g2_fill_8 FILLER_223_312 ();
 sg13g2_fill_8 FILLER_223_320 ();
 sg13g2_fill_8 FILLER_223_328 ();
 sg13g2_fill_8 FILLER_223_336 ();
 sg13g2_fill_8 FILLER_223_344 ();
 sg13g2_fill_8 FILLER_223_352 ();
 sg13g2_fill_8 FILLER_223_360 ();
 sg13g2_fill_8 FILLER_223_368 ();
 sg13g2_fill_8 FILLER_223_376 ();
 sg13g2_fill_8 FILLER_223_384 ();
 sg13g2_fill_8 FILLER_223_392 ();
 sg13g2_fill_8 FILLER_223_400 ();
 sg13g2_fill_8 FILLER_223_408 ();
 sg13g2_fill_8 FILLER_223_416 ();
 sg13g2_fill_8 FILLER_223_424 ();
 sg13g2_fill_8 FILLER_223_432 ();
 sg13g2_fill_8 FILLER_223_440 ();
 sg13g2_fill_8 FILLER_223_448 ();
 sg13g2_fill_8 FILLER_223_456 ();
 sg13g2_fill_8 FILLER_223_464 ();
 sg13g2_fill_8 FILLER_223_472 ();
 sg13g2_fill_8 FILLER_223_480 ();
 sg13g2_fill_8 FILLER_223_488 ();
 sg13g2_fill_8 FILLER_223_496 ();
 sg13g2_fill_8 FILLER_223_504 ();
 sg13g2_fill_8 FILLER_223_512 ();
 sg13g2_fill_8 FILLER_223_520 ();
 sg13g2_fill_8 FILLER_223_528 ();
 sg13g2_fill_8 FILLER_223_536 ();
 sg13g2_fill_8 FILLER_223_544 ();
 sg13g2_fill_8 FILLER_223_552 ();
 sg13g2_fill_8 FILLER_223_560 ();
 sg13g2_fill_8 FILLER_223_568 ();
 sg13g2_fill_8 FILLER_223_576 ();
 sg13g2_fill_8 FILLER_223_584 ();
 sg13g2_fill_8 FILLER_223_592 ();
 sg13g2_fill_8 FILLER_223_600 ();
 sg13g2_fill_8 FILLER_223_608 ();
 sg13g2_fill_8 FILLER_223_616 ();
 sg13g2_fill_8 FILLER_223_624 ();
 sg13g2_fill_8 FILLER_223_632 ();
 sg13g2_fill_8 FILLER_223_640 ();
 sg13g2_fill_8 FILLER_223_648 ();
 sg13g2_fill_8 FILLER_223_656 ();
 sg13g2_fill_8 FILLER_223_664 ();
 sg13g2_fill_8 FILLER_223_672 ();
 sg13g2_fill_8 FILLER_223_680 ();
 sg13g2_fill_8 FILLER_223_688 ();
 sg13g2_fill_8 FILLER_223_696 ();
 sg13g2_fill_8 FILLER_223_704 ();
 sg13g2_fill_8 FILLER_223_712 ();
 sg13g2_fill_8 FILLER_223_720 ();
 sg13g2_fill_8 FILLER_223_728 ();
 sg13g2_fill_8 FILLER_223_736 ();
 sg13g2_fill_8 FILLER_223_744 ();
 sg13g2_fill_8 FILLER_223_752 ();
 sg13g2_fill_8 FILLER_223_760 ();
 sg13g2_fill_8 FILLER_223_768 ();
 sg13g2_fill_8 FILLER_223_776 ();
 sg13g2_fill_8 FILLER_223_784 ();
 sg13g2_fill_8 FILLER_223_792 ();
 sg13g2_fill_8 FILLER_223_800 ();
 sg13g2_fill_8 FILLER_223_808 ();
 sg13g2_fill_8 FILLER_223_816 ();
 sg13g2_fill_8 FILLER_223_824 ();
 sg13g2_fill_8 FILLER_223_832 ();
 sg13g2_fill_8 FILLER_223_840 ();
 sg13g2_fill_8 FILLER_223_848 ();
 sg13g2_fill_8 FILLER_223_856 ();
 sg13g2_fill_8 FILLER_223_864 ();
 sg13g2_fill_8 FILLER_223_872 ();
 sg13g2_fill_8 FILLER_223_880 ();
 sg13g2_fill_8 FILLER_223_888 ();
 sg13g2_fill_8 FILLER_223_896 ();
 sg13g2_fill_8 FILLER_223_904 ();
 sg13g2_fill_8 FILLER_223_912 ();
 sg13g2_fill_8 FILLER_223_920 ();
 sg13g2_fill_8 FILLER_223_928 ();
 sg13g2_fill_8 FILLER_223_936 ();
 sg13g2_fill_8 FILLER_223_944 ();
 sg13g2_fill_8 FILLER_223_952 ();
 sg13g2_fill_8 FILLER_223_960 ();
 sg13g2_fill_8 FILLER_223_968 ();
 sg13g2_fill_8 FILLER_223_976 ();
 sg13g2_fill_8 FILLER_223_984 ();
 sg13g2_fill_8 FILLER_223_992 ();
 sg13g2_fill_8 FILLER_223_1000 ();
 sg13g2_fill_8 FILLER_223_1008 ();
 sg13g2_fill_8 FILLER_223_1016 ();
 sg13g2_fill_8 FILLER_223_1024 ();
 sg13g2_fill_8 FILLER_223_1032 ();
 sg13g2_fill_8 FILLER_223_1040 ();
 sg13g2_fill_8 FILLER_223_1048 ();
 sg13g2_fill_8 FILLER_223_1056 ();
 sg13g2_fill_8 FILLER_223_1064 ();
 sg13g2_fill_8 FILLER_223_1072 ();
 sg13g2_fill_8 FILLER_223_1080 ();
 sg13g2_fill_8 FILLER_223_1088 ();
 sg13g2_fill_8 FILLER_223_1096 ();
 sg13g2_fill_8 FILLER_223_1104 ();
 sg13g2_fill_8 FILLER_223_1112 ();
 sg13g2_fill_8 FILLER_223_1120 ();
 sg13g2_fill_8 FILLER_223_1128 ();
 sg13g2_fill_8 FILLER_223_1136 ();
 sg13g2_fill_8 FILLER_223_1144 ();
 sg13g2_fill_8 FILLER_223_1152 ();
 sg13g2_fill_8 FILLER_223_1160 ();
 sg13g2_fill_8 FILLER_223_1168 ();
 sg13g2_fill_8 FILLER_223_1176 ();
 sg13g2_fill_8 FILLER_223_1184 ();
 sg13g2_fill_8 FILLER_223_1192 ();
 sg13g2_fill_8 FILLER_223_1200 ();
 sg13g2_fill_8 FILLER_223_1208 ();
 sg13g2_fill_8 FILLER_223_1216 ();
 sg13g2_fill_8 FILLER_223_1224 ();
 sg13g2_fill_8 FILLER_223_1232 ();
 sg13g2_fill_8 FILLER_223_1240 ();
 sg13g2_fill_8 FILLER_223_1248 ();
 sg13g2_fill_8 FILLER_223_1256 ();
 sg13g2_fill_8 FILLER_223_1264 ();
 sg13g2_fill_8 FILLER_223_1272 ();
 sg13g2_fill_8 FILLER_223_1280 ();
 sg13g2_fill_8 FILLER_223_1288 ();
 sg13g2_fill_8 FILLER_223_1296 ();
 sg13g2_fill_8 FILLER_223_1304 ();
 sg13g2_fill_8 FILLER_223_1312 ();
 sg13g2_fill_8 FILLER_223_1320 ();
 sg13g2_fill_8 FILLER_223_1328 ();
 sg13g2_fill_8 FILLER_223_1336 ();
 sg13g2_fill_8 FILLER_223_1344 ();
 sg13g2_fill_8 FILLER_223_1352 ();
 sg13g2_fill_8 FILLER_223_1360 ();
 sg13g2_fill_8 FILLER_223_1368 ();
 sg13g2_fill_8 FILLER_223_1376 ();
 sg13g2_fill_8 FILLER_223_1384 ();
 sg13g2_fill_8 FILLER_223_1392 ();
 sg13g2_fill_8 FILLER_223_1400 ();
 sg13g2_fill_8 FILLER_223_1408 ();
 sg13g2_fill_8 FILLER_223_1416 ();
 sg13g2_fill_8 FILLER_223_1424 ();
 sg13g2_fill_8 FILLER_223_1432 ();
 sg13g2_fill_8 FILLER_223_1440 ();
 sg13g2_fill_8 FILLER_223_1448 ();
 sg13g2_fill_8 FILLER_223_1456 ();
 sg13g2_fill_8 FILLER_223_1464 ();
 sg13g2_fill_8 FILLER_223_1472 ();
 sg13g2_fill_8 FILLER_223_1480 ();
 sg13g2_fill_8 FILLER_223_1488 ();
 sg13g2_fill_8 FILLER_223_1496 ();
 sg13g2_fill_8 FILLER_223_1504 ();
 sg13g2_fill_8 FILLER_223_1512 ();
 sg13g2_fill_8 FILLER_223_1520 ();
 sg13g2_fill_8 FILLER_223_1528 ();
 sg13g2_fill_8 FILLER_223_1536 ();
 sg13g2_fill_8 FILLER_223_1544 ();
 sg13g2_fill_8 FILLER_223_1552 ();
 sg13g2_fill_8 FILLER_223_1560 ();
 sg13g2_fill_8 FILLER_223_1568 ();
 sg13g2_fill_8 FILLER_223_1576 ();
 sg13g2_fill_8 FILLER_223_1584 ();
 sg13g2_fill_8 FILLER_224_0 ();
 sg13g2_fill_8 FILLER_224_8 ();
 sg13g2_fill_8 FILLER_224_16 ();
 sg13g2_fill_8 FILLER_224_24 ();
 sg13g2_fill_8 FILLER_224_32 ();
 sg13g2_fill_8 FILLER_224_40 ();
 sg13g2_fill_8 FILLER_224_48 ();
 sg13g2_fill_8 FILLER_224_56 ();
 sg13g2_fill_8 FILLER_224_64 ();
 sg13g2_fill_8 FILLER_224_72 ();
 sg13g2_fill_8 FILLER_224_80 ();
 sg13g2_fill_8 FILLER_224_88 ();
 sg13g2_fill_8 FILLER_224_96 ();
 sg13g2_fill_8 FILLER_224_104 ();
 sg13g2_fill_8 FILLER_224_112 ();
 sg13g2_fill_8 FILLER_224_120 ();
 sg13g2_fill_8 FILLER_224_128 ();
 sg13g2_fill_8 FILLER_224_136 ();
 sg13g2_fill_8 FILLER_224_144 ();
 sg13g2_fill_8 FILLER_224_152 ();
 sg13g2_fill_8 FILLER_224_160 ();
 sg13g2_fill_8 FILLER_224_168 ();
 sg13g2_fill_8 FILLER_224_176 ();
 sg13g2_fill_8 FILLER_224_184 ();
 sg13g2_fill_8 FILLER_224_192 ();
 sg13g2_fill_8 FILLER_224_200 ();
 sg13g2_fill_8 FILLER_224_208 ();
 sg13g2_fill_8 FILLER_224_216 ();
 sg13g2_fill_8 FILLER_224_224 ();
 sg13g2_fill_8 FILLER_224_232 ();
 sg13g2_fill_8 FILLER_224_240 ();
 sg13g2_fill_8 FILLER_224_248 ();
 sg13g2_fill_8 FILLER_224_256 ();
 sg13g2_fill_8 FILLER_224_264 ();
 sg13g2_fill_8 FILLER_224_272 ();
 sg13g2_fill_8 FILLER_224_280 ();
 sg13g2_fill_8 FILLER_224_288 ();
 sg13g2_fill_8 FILLER_224_296 ();
 sg13g2_fill_8 FILLER_224_304 ();
 sg13g2_fill_8 FILLER_224_312 ();
 sg13g2_fill_8 FILLER_224_320 ();
 sg13g2_fill_8 FILLER_224_328 ();
 sg13g2_fill_8 FILLER_224_336 ();
 sg13g2_fill_8 FILLER_224_344 ();
 sg13g2_fill_8 FILLER_224_352 ();
 sg13g2_fill_8 FILLER_224_360 ();
 sg13g2_fill_8 FILLER_224_368 ();
 sg13g2_fill_8 FILLER_224_376 ();
 sg13g2_fill_8 FILLER_224_384 ();
 sg13g2_fill_8 FILLER_224_392 ();
 sg13g2_fill_8 FILLER_224_400 ();
 sg13g2_fill_8 FILLER_224_408 ();
 sg13g2_fill_8 FILLER_224_416 ();
 sg13g2_fill_8 FILLER_224_424 ();
 sg13g2_fill_8 FILLER_224_432 ();
 sg13g2_fill_8 FILLER_224_440 ();
 sg13g2_fill_8 FILLER_224_448 ();
 sg13g2_fill_8 FILLER_224_456 ();
 sg13g2_fill_8 FILLER_224_464 ();
 sg13g2_fill_8 FILLER_224_472 ();
 sg13g2_fill_8 FILLER_224_480 ();
 sg13g2_fill_8 FILLER_224_488 ();
 sg13g2_fill_8 FILLER_224_496 ();
 sg13g2_fill_8 FILLER_224_504 ();
 sg13g2_fill_8 FILLER_224_512 ();
 sg13g2_fill_8 FILLER_224_520 ();
 sg13g2_fill_8 FILLER_224_528 ();
 sg13g2_fill_8 FILLER_224_536 ();
 sg13g2_fill_8 FILLER_224_544 ();
 sg13g2_fill_8 FILLER_224_552 ();
 sg13g2_fill_8 FILLER_224_560 ();
 sg13g2_fill_8 FILLER_224_568 ();
 sg13g2_fill_8 FILLER_224_576 ();
 sg13g2_fill_8 FILLER_224_584 ();
 sg13g2_fill_8 FILLER_224_592 ();
 sg13g2_fill_8 FILLER_224_600 ();
 sg13g2_fill_8 FILLER_224_608 ();
 sg13g2_fill_8 FILLER_224_616 ();
 sg13g2_fill_8 FILLER_224_624 ();
 sg13g2_fill_8 FILLER_224_632 ();
 sg13g2_fill_8 FILLER_224_640 ();
 sg13g2_fill_8 FILLER_224_648 ();
 sg13g2_fill_8 FILLER_224_656 ();
 sg13g2_fill_8 FILLER_224_664 ();
 sg13g2_fill_8 FILLER_224_672 ();
 sg13g2_fill_8 FILLER_224_680 ();
 sg13g2_fill_8 FILLER_224_688 ();
 sg13g2_fill_8 FILLER_224_696 ();
 sg13g2_fill_8 FILLER_224_704 ();
 sg13g2_fill_8 FILLER_224_712 ();
 sg13g2_fill_8 FILLER_224_720 ();
 sg13g2_fill_8 FILLER_224_728 ();
 sg13g2_fill_8 FILLER_224_736 ();
 sg13g2_fill_8 FILLER_224_744 ();
 sg13g2_fill_8 FILLER_224_752 ();
 sg13g2_fill_8 FILLER_224_760 ();
 sg13g2_fill_8 FILLER_224_768 ();
 sg13g2_fill_8 FILLER_224_776 ();
 sg13g2_fill_8 FILLER_224_784 ();
 sg13g2_fill_8 FILLER_224_792 ();
 sg13g2_fill_8 FILLER_224_800 ();
 sg13g2_fill_8 FILLER_224_808 ();
 sg13g2_fill_8 FILLER_224_816 ();
 sg13g2_fill_8 FILLER_224_824 ();
 sg13g2_fill_8 FILLER_224_832 ();
 sg13g2_fill_8 FILLER_224_840 ();
 sg13g2_fill_8 FILLER_224_848 ();
 sg13g2_fill_8 FILLER_224_856 ();
 sg13g2_fill_8 FILLER_224_864 ();
 sg13g2_fill_8 FILLER_224_872 ();
 sg13g2_fill_8 FILLER_224_880 ();
 sg13g2_fill_8 FILLER_224_888 ();
 sg13g2_fill_8 FILLER_224_896 ();
 sg13g2_fill_8 FILLER_224_904 ();
 sg13g2_fill_8 FILLER_224_912 ();
 sg13g2_fill_8 FILLER_224_920 ();
 sg13g2_fill_8 FILLER_224_928 ();
 sg13g2_fill_8 FILLER_224_936 ();
 sg13g2_fill_8 FILLER_224_944 ();
 sg13g2_fill_8 FILLER_224_952 ();
 sg13g2_fill_8 FILLER_224_960 ();
 sg13g2_fill_8 FILLER_224_968 ();
 sg13g2_fill_8 FILLER_224_976 ();
 sg13g2_fill_8 FILLER_224_984 ();
 sg13g2_fill_8 FILLER_224_992 ();
 sg13g2_fill_8 FILLER_224_1000 ();
 sg13g2_fill_8 FILLER_224_1008 ();
 sg13g2_fill_8 FILLER_224_1016 ();
 sg13g2_fill_8 FILLER_224_1024 ();
 sg13g2_fill_8 FILLER_224_1032 ();
 sg13g2_fill_8 FILLER_224_1040 ();
 sg13g2_fill_8 FILLER_224_1048 ();
 sg13g2_fill_8 FILLER_224_1056 ();
 sg13g2_fill_8 FILLER_224_1064 ();
 sg13g2_fill_8 FILLER_224_1072 ();
 sg13g2_fill_8 FILLER_224_1080 ();
 sg13g2_fill_8 FILLER_224_1088 ();
 sg13g2_fill_8 FILLER_224_1096 ();
 sg13g2_fill_8 FILLER_224_1104 ();
 sg13g2_fill_8 FILLER_224_1112 ();
 sg13g2_fill_8 FILLER_224_1120 ();
 sg13g2_fill_8 FILLER_224_1128 ();
 sg13g2_fill_8 FILLER_224_1136 ();
 sg13g2_fill_8 FILLER_224_1144 ();
 sg13g2_fill_8 FILLER_224_1152 ();
 sg13g2_fill_8 FILLER_224_1160 ();
 sg13g2_fill_8 FILLER_224_1168 ();
 sg13g2_fill_8 FILLER_224_1176 ();
 sg13g2_fill_8 FILLER_224_1184 ();
 sg13g2_fill_8 FILLER_224_1192 ();
 sg13g2_fill_8 FILLER_224_1200 ();
 sg13g2_fill_8 FILLER_224_1208 ();
 sg13g2_fill_8 FILLER_224_1216 ();
 sg13g2_fill_8 FILLER_224_1224 ();
 sg13g2_fill_8 FILLER_224_1232 ();
 sg13g2_fill_8 FILLER_224_1240 ();
 sg13g2_fill_8 FILLER_224_1248 ();
 sg13g2_fill_8 FILLER_224_1256 ();
 sg13g2_fill_8 FILLER_224_1264 ();
 sg13g2_fill_8 FILLER_224_1272 ();
 sg13g2_fill_8 FILLER_224_1280 ();
 sg13g2_fill_8 FILLER_224_1288 ();
 sg13g2_fill_8 FILLER_224_1296 ();
 sg13g2_fill_8 FILLER_224_1304 ();
 sg13g2_fill_8 FILLER_224_1312 ();
 sg13g2_fill_8 FILLER_224_1320 ();
 sg13g2_fill_8 FILLER_224_1328 ();
 sg13g2_fill_8 FILLER_224_1336 ();
 sg13g2_fill_8 FILLER_224_1344 ();
 sg13g2_fill_8 FILLER_224_1352 ();
 sg13g2_fill_8 FILLER_224_1360 ();
 sg13g2_fill_8 FILLER_224_1368 ();
 sg13g2_fill_8 FILLER_224_1376 ();
 sg13g2_fill_8 FILLER_224_1384 ();
 sg13g2_fill_8 FILLER_224_1392 ();
 sg13g2_fill_8 FILLER_224_1400 ();
 sg13g2_fill_8 FILLER_224_1408 ();
 sg13g2_fill_8 FILLER_224_1416 ();
 sg13g2_fill_8 FILLER_224_1424 ();
 sg13g2_fill_8 FILLER_224_1432 ();
 sg13g2_fill_8 FILLER_224_1440 ();
 sg13g2_fill_8 FILLER_224_1448 ();
 sg13g2_fill_8 FILLER_224_1456 ();
 sg13g2_fill_8 FILLER_224_1464 ();
 sg13g2_fill_8 FILLER_224_1472 ();
 sg13g2_fill_8 FILLER_224_1480 ();
 sg13g2_fill_8 FILLER_224_1488 ();
 sg13g2_fill_8 FILLER_224_1496 ();
 sg13g2_fill_8 FILLER_224_1504 ();
 sg13g2_fill_8 FILLER_224_1512 ();
 sg13g2_fill_8 FILLER_224_1520 ();
 sg13g2_fill_8 FILLER_224_1528 ();
 sg13g2_fill_8 FILLER_224_1536 ();
 sg13g2_fill_8 FILLER_224_1544 ();
 sg13g2_fill_8 FILLER_224_1552 ();
 sg13g2_fill_8 FILLER_224_1560 ();
 sg13g2_fill_8 FILLER_224_1568 ();
 sg13g2_fill_8 FILLER_224_1576 ();
 sg13g2_fill_8 FILLER_224_1584 ();
 sg13g2_fill_8 FILLER_225_0 ();
 sg13g2_fill_8 FILLER_225_8 ();
 sg13g2_fill_8 FILLER_225_16 ();
 sg13g2_fill_8 FILLER_225_24 ();
 sg13g2_fill_8 FILLER_225_32 ();
 sg13g2_fill_8 FILLER_225_40 ();
 sg13g2_fill_8 FILLER_225_48 ();
 sg13g2_fill_8 FILLER_225_56 ();
 sg13g2_fill_8 FILLER_225_64 ();
 sg13g2_fill_8 FILLER_225_72 ();
 sg13g2_fill_8 FILLER_225_80 ();
 sg13g2_fill_8 FILLER_225_88 ();
 sg13g2_fill_8 FILLER_225_96 ();
 sg13g2_fill_8 FILLER_225_104 ();
 sg13g2_fill_8 FILLER_225_112 ();
 sg13g2_fill_8 FILLER_225_120 ();
 sg13g2_fill_8 FILLER_225_128 ();
 sg13g2_fill_8 FILLER_225_136 ();
 sg13g2_fill_8 FILLER_225_144 ();
 sg13g2_fill_8 FILLER_225_152 ();
 sg13g2_fill_8 FILLER_225_160 ();
 sg13g2_fill_8 FILLER_225_168 ();
 sg13g2_fill_8 FILLER_225_176 ();
 sg13g2_fill_8 FILLER_225_184 ();
 sg13g2_fill_8 FILLER_225_192 ();
 sg13g2_fill_8 FILLER_225_200 ();
 sg13g2_fill_8 FILLER_225_208 ();
 sg13g2_fill_8 FILLER_225_216 ();
 sg13g2_fill_8 FILLER_225_224 ();
 sg13g2_fill_8 FILLER_225_232 ();
 sg13g2_fill_8 FILLER_225_240 ();
 sg13g2_fill_8 FILLER_225_248 ();
 sg13g2_fill_8 FILLER_225_256 ();
 sg13g2_fill_8 FILLER_225_264 ();
 sg13g2_fill_8 FILLER_225_272 ();
 sg13g2_fill_8 FILLER_225_280 ();
 sg13g2_fill_8 FILLER_225_288 ();
 sg13g2_fill_8 FILLER_225_296 ();
 sg13g2_fill_8 FILLER_225_304 ();
 sg13g2_fill_8 FILLER_225_312 ();
 sg13g2_fill_8 FILLER_225_320 ();
 sg13g2_fill_8 FILLER_225_328 ();
 sg13g2_fill_8 FILLER_225_336 ();
 sg13g2_fill_8 FILLER_225_344 ();
 sg13g2_fill_8 FILLER_225_352 ();
 sg13g2_fill_8 FILLER_225_360 ();
 sg13g2_fill_8 FILLER_225_368 ();
 sg13g2_fill_8 FILLER_225_376 ();
 sg13g2_fill_8 FILLER_225_384 ();
 sg13g2_fill_8 FILLER_225_392 ();
 sg13g2_fill_8 FILLER_225_400 ();
 sg13g2_fill_8 FILLER_225_408 ();
 sg13g2_fill_8 FILLER_225_416 ();
 sg13g2_fill_8 FILLER_225_424 ();
 sg13g2_fill_8 FILLER_225_432 ();
 sg13g2_fill_8 FILLER_225_440 ();
 sg13g2_fill_8 FILLER_225_448 ();
 sg13g2_fill_8 FILLER_225_456 ();
 sg13g2_fill_8 FILLER_225_464 ();
 sg13g2_fill_8 FILLER_225_472 ();
 sg13g2_fill_8 FILLER_225_480 ();
 sg13g2_fill_8 FILLER_225_488 ();
 sg13g2_fill_8 FILLER_225_496 ();
 sg13g2_fill_8 FILLER_225_504 ();
 sg13g2_fill_8 FILLER_225_512 ();
 sg13g2_fill_8 FILLER_225_520 ();
 sg13g2_fill_8 FILLER_225_528 ();
 sg13g2_fill_8 FILLER_225_536 ();
 sg13g2_fill_8 FILLER_225_544 ();
 sg13g2_fill_8 FILLER_225_552 ();
 sg13g2_fill_8 FILLER_225_560 ();
 sg13g2_fill_8 FILLER_225_568 ();
 sg13g2_fill_8 FILLER_225_576 ();
 sg13g2_fill_8 FILLER_225_584 ();
 sg13g2_fill_8 FILLER_225_592 ();
 sg13g2_fill_8 FILLER_225_600 ();
 sg13g2_fill_8 FILLER_225_608 ();
 sg13g2_fill_8 FILLER_225_616 ();
 sg13g2_fill_8 FILLER_225_624 ();
 sg13g2_fill_8 FILLER_225_632 ();
 sg13g2_fill_8 FILLER_225_640 ();
 sg13g2_fill_8 FILLER_225_648 ();
 sg13g2_fill_8 FILLER_225_656 ();
 sg13g2_fill_8 FILLER_225_664 ();
 sg13g2_fill_8 FILLER_225_672 ();
 sg13g2_fill_8 FILLER_225_680 ();
 sg13g2_fill_8 FILLER_225_688 ();
 sg13g2_fill_8 FILLER_225_696 ();
 sg13g2_fill_8 FILLER_225_704 ();
 sg13g2_fill_8 FILLER_225_712 ();
 sg13g2_fill_8 FILLER_225_720 ();
 sg13g2_fill_8 FILLER_225_728 ();
 sg13g2_fill_8 FILLER_225_736 ();
 sg13g2_fill_8 FILLER_225_744 ();
 sg13g2_fill_8 FILLER_225_752 ();
 sg13g2_fill_8 FILLER_225_760 ();
 sg13g2_fill_8 FILLER_225_768 ();
 sg13g2_fill_8 FILLER_225_776 ();
 sg13g2_fill_8 FILLER_225_784 ();
 sg13g2_fill_8 FILLER_225_792 ();
 sg13g2_fill_8 FILLER_225_800 ();
 sg13g2_fill_8 FILLER_225_808 ();
 sg13g2_fill_8 FILLER_225_816 ();
 sg13g2_fill_8 FILLER_225_824 ();
 sg13g2_fill_8 FILLER_225_832 ();
 sg13g2_fill_8 FILLER_225_840 ();
 sg13g2_fill_8 FILLER_225_848 ();
 sg13g2_fill_8 FILLER_225_856 ();
 sg13g2_fill_8 FILLER_225_864 ();
 sg13g2_fill_8 FILLER_225_872 ();
 sg13g2_fill_8 FILLER_225_880 ();
 sg13g2_fill_8 FILLER_225_888 ();
 sg13g2_fill_8 FILLER_225_896 ();
 sg13g2_fill_8 FILLER_225_904 ();
 sg13g2_fill_8 FILLER_225_912 ();
 sg13g2_fill_8 FILLER_225_920 ();
 sg13g2_fill_8 FILLER_225_928 ();
 sg13g2_fill_8 FILLER_225_936 ();
 sg13g2_fill_8 FILLER_225_944 ();
 sg13g2_fill_8 FILLER_225_952 ();
 sg13g2_fill_8 FILLER_225_960 ();
 sg13g2_fill_8 FILLER_225_968 ();
 sg13g2_fill_8 FILLER_225_976 ();
 sg13g2_fill_8 FILLER_225_984 ();
 sg13g2_fill_8 FILLER_225_992 ();
 sg13g2_fill_8 FILLER_225_1000 ();
 sg13g2_fill_8 FILLER_225_1008 ();
 sg13g2_fill_8 FILLER_225_1016 ();
 sg13g2_fill_8 FILLER_225_1024 ();
 sg13g2_fill_8 FILLER_225_1032 ();
 sg13g2_fill_8 FILLER_225_1040 ();
 sg13g2_fill_8 FILLER_225_1048 ();
 sg13g2_fill_8 FILLER_225_1056 ();
 sg13g2_fill_8 FILLER_225_1064 ();
 sg13g2_fill_8 FILLER_225_1072 ();
 sg13g2_fill_8 FILLER_225_1080 ();
 sg13g2_fill_8 FILLER_225_1088 ();
 sg13g2_fill_8 FILLER_225_1096 ();
 sg13g2_fill_8 FILLER_225_1104 ();
 sg13g2_fill_8 FILLER_225_1112 ();
 sg13g2_fill_8 FILLER_225_1120 ();
 sg13g2_fill_8 FILLER_225_1128 ();
 sg13g2_fill_8 FILLER_225_1136 ();
 sg13g2_fill_8 FILLER_225_1144 ();
 sg13g2_fill_8 FILLER_225_1152 ();
 sg13g2_fill_8 FILLER_225_1160 ();
 sg13g2_fill_8 FILLER_225_1168 ();
 sg13g2_fill_8 FILLER_225_1176 ();
 sg13g2_fill_8 FILLER_225_1184 ();
 sg13g2_fill_8 FILLER_225_1192 ();
 sg13g2_fill_8 FILLER_225_1200 ();
 sg13g2_fill_8 FILLER_225_1208 ();
 sg13g2_fill_8 FILLER_225_1216 ();
 sg13g2_fill_8 FILLER_225_1224 ();
 sg13g2_fill_8 FILLER_225_1232 ();
 sg13g2_fill_8 FILLER_225_1240 ();
 sg13g2_fill_8 FILLER_225_1248 ();
 sg13g2_fill_8 FILLER_225_1256 ();
 sg13g2_fill_8 FILLER_225_1264 ();
 sg13g2_fill_8 FILLER_225_1272 ();
 sg13g2_fill_8 FILLER_225_1280 ();
 sg13g2_fill_8 FILLER_225_1288 ();
 sg13g2_fill_8 FILLER_225_1296 ();
 sg13g2_fill_8 FILLER_225_1304 ();
 sg13g2_fill_8 FILLER_225_1312 ();
 sg13g2_fill_8 FILLER_225_1320 ();
 sg13g2_fill_8 FILLER_225_1328 ();
 sg13g2_fill_8 FILLER_225_1336 ();
 sg13g2_fill_8 FILLER_225_1344 ();
 sg13g2_fill_8 FILLER_225_1352 ();
 sg13g2_fill_8 FILLER_225_1360 ();
 sg13g2_fill_8 FILLER_225_1368 ();
 sg13g2_fill_8 FILLER_225_1376 ();
 sg13g2_fill_8 FILLER_225_1384 ();
 sg13g2_fill_8 FILLER_225_1392 ();
 sg13g2_fill_8 FILLER_225_1400 ();
 sg13g2_fill_8 FILLER_225_1408 ();
 sg13g2_fill_8 FILLER_225_1416 ();
 sg13g2_fill_8 FILLER_225_1424 ();
 sg13g2_fill_8 FILLER_225_1432 ();
 sg13g2_fill_8 FILLER_225_1440 ();
 sg13g2_fill_8 FILLER_225_1448 ();
 sg13g2_fill_8 FILLER_225_1456 ();
 sg13g2_fill_8 FILLER_225_1464 ();
 sg13g2_fill_8 FILLER_225_1472 ();
 sg13g2_fill_8 FILLER_225_1480 ();
 sg13g2_fill_8 FILLER_225_1488 ();
 sg13g2_fill_8 FILLER_225_1496 ();
 sg13g2_fill_8 FILLER_225_1504 ();
 sg13g2_fill_8 FILLER_225_1512 ();
 sg13g2_fill_8 FILLER_225_1520 ();
 sg13g2_fill_8 FILLER_225_1528 ();
 sg13g2_fill_8 FILLER_225_1536 ();
 sg13g2_fill_8 FILLER_225_1544 ();
 sg13g2_fill_8 FILLER_225_1552 ();
 sg13g2_fill_8 FILLER_225_1560 ();
 sg13g2_fill_8 FILLER_225_1568 ();
 sg13g2_fill_8 FILLER_225_1576 ();
 sg13g2_fill_8 FILLER_225_1584 ();
 sg13g2_fill_8 FILLER_226_0 ();
 sg13g2_fill_8 FILLER_226_8 ();
 sg13g2_fill_8 FILLER_226_16 ();
 sg13g2_fill_8 FILLER_226_24 ();
 sg13g2_fill_8 FILLER_226_32 ();
 sg13g2_fill_8 FILLER_226_40 ();
 sg13g2_fill_8 FILLER_226_48 ();
 sg13g2_fill_8 FILLER_226_56 ();
 sg13g2_fill_8 FILLER_226_64 ();
 sg13g2_fill_8 FILLER_226_72 ();
 sg13g2_fill_8 FILLER_226_80 ();
 sg13g2_fill_8 FILLER_226_88 ();
 sg13g2_fill_8 FILLER_226_96 ();
 sg13g2_fill_8 FILLER_226_104 ();
 sg13g2_fill_8 FILLER_226_112 ();
 sg13g2_fill_8 FILLER_226_120 ();
 sg13g2_fill_8 FILLER_226_128 ();
 sg13g2_fill_8 FILLER_226_136 ();
 sg13g2_fill_8 FILLER_226_144 ();
 sg13g2_fill_8 FILLER_226_152 ();
 sg13g2_fill_8 FILLER_226_160 ();
 sg13g2_fill_8 FILLER_226_168 ();
 sg13g2_fill_8 FILLER_226_176 ();
 sg13g2_fill_8 FILLER_226_184 ();
 sg13g2_fill_8 FILLER_226_192 ();
 sg13g2_fill_8 FILLER_226_200 ();
 sg13g2_fill_8 FILLER_226_208 ();
 sg13g2_fill_8 FILLER_226_216 ();
 sg13g2_fill_8 FILLER_226_224 ();
 sg13g2_fill_8 FILLER_226_232 ();
 sg13g2_fill_8 FILLER_226_240 ();
 sg13g2_fill_8 FILLER_226_248 ();
 sg13g2_fill_8 FILLER_226_256 ();
 sg13g2_fill_8 FILLER_226_264 ();
 sg13g2_fill_8 FILLER_226_272 ();
 sg13g2_fill_8 FILLER_226_280 ();
 sg13g2_fill_8 FILLER_226_288 ();
 sg13g2_fill_8 FILLER_226_296 ();
 sg13g2_fill_8 FILLER_226_304 ();
 sg13g2_fill_8 FILLER_226_312 ();
 sg13g2_fill_8 FILLER_226_320 ();
 sg13g2_fill_8 FILLER_226_328 ();
 sg13g2_fill_8 FILLER_226_336 ();
 sg13g2_fill_8 FILLER_226_344 ();
 sg13g2_fill_8 FILLER_226_352 ();
 sg13g2_fill_8 FILLER_226_360 ();
 sg13g2_fill_8 FILLER_226_368 ();
 sg13g2_fill_8 FILLER_226_376 ();
 sg13g2_fill_8 FILLER_226_384 ();
 sg13g2_fill_8 FILLER_226_392 ();
 sg13g2_fill_8 FILLER_226_400 ();
 sg13g2_fill_8 FILLER_226_408 ();
 sg13g2_fill_8 FILLER_226_416 ();
 sg13g2_fill_8 FILLER_226_424 ();
 sg13g2_fill_8 FILLER_226_432 ();
 sg13g2_fill_8 FILLER_226_440 ();
 sg13g2_fill_8 FILLER_226_448 ();
 sg13g2_fill_8 FILLER_226_456 ();
 sg13g2_fill_8 FILLER_226_464 ();
 sg13g2_fill_8 FILLER_226_472 ();
 sg13g2_fill_8 FILLER_226_480 ();
 sg13g2_fill_8 FILLER_226_488 ();
 sg13g2_fill_8 FILLER_226_496 ();
 sg13g2_fill_8 FILLER_226_504 ();
 sg13g2_fill_8 FILLER_226_512 ();
 sg13g2_fill_8 FILLER_226_520 ();
 sg13g2_fill_8 FILLER_226_528 ();
 sg13g2_fill_8 FILLER_226_536 ();
 sg13g2_fill_8 FILLER_226_544 ();
 sg13g2_fill_8 FILLER_226_552 ();
 sg13g2_fill_8 FILLER_226_560 ();
 sg13g2_fill_8 FILLER_226_568 ();
 sg13g2_fill_8 FILLER_226_576 ();
 sg13g2_fill_8 FILLER_226_584 ();
 sg13g2_fill_8 FILLER_226_592 ();
 sg13g2_fill_8 FILLER_226_600 ();
 sg13g2_fill_8 FILLER_226_608 ();
 sg13g2_fill_8 FILLER_226_616 ();
 sg13g2_fill_8 FILLER_226_624 ();
 sg13g2_fill_8 FILLER_226_632 ();
 sg13g2_fill_8 FILLER_226_640 ();
 sg13g2_fill_8 FILLER_226_648 ();
 sg13g2_fill_8 FILLER_226_656 ();
 sg13g2_fill_8 FILLER_226_664 ();
 sg13g2_fill_8 FILLER_226_672 ();
 sg13g2_fill_8 FILLER_226_680 ();
 sg13g2_fill_8 FILLER_226_688 ();
 sg13g2_fill_8 FILLER_226_696 ();
 sg13g2_fill_8 FILLER_226_704 ();
 sg13g2_fill_8 FILLER_226_712 ();
 sg13g2_fill_8 FILLER_226_720 ();
 sg13g2_fill_8 FILLER_226_728 ();
 sg13g2_fill_8 FILLER_226_736 ();
 sg13g2_fill_8 FILLER_226_744 ();
 sg13g2_fill_8 FILLER_226_752 ();
 sg13g2_fill_8 FILLER_226_760 ();
 sg13g2_fill_8 FILLER_226_768 ();
 sg13g2_fill_8 FILLER_226_776 ();
 sg13g2_fill_8 FILLER_226_784 ();
 sg13g2_fill_8 FILLER_226_792 ();
 sg13g2_fill_8 FILLER_226_800 ();
 sg13g2_fill_8 FILLER_226_808 ();
 sg13g2_fill_8 FILLER_226_816 ();
 sg13g2_fill_8 FILLER_226_824 ();
 sg13g2_fill_8 FILLER_226_832 ();
 sg13g2_fill_8 FILLER_226_840 ();
 sg13g2_fill_8 FILLER_226_848 ();
 sg13g2_fill_8 FILLER_226_856 ();
 sg13g2_fill_8 FILLER_226_864 ();
 sg13g2_fill_8 FILLER_226_872 ();
 sg13g2_fill_8 FILLER_226_880 ();
 sg13g2_fill_8 FILLER_226_888 ();
 sg13g2_fill_8 FILLER_226_896 ();
 sg13g2_fill_8 FILLER_226_904 ();
 sg13g2_fill_8 FILLER_226_912 ();
 sg13g2_fill_8 FILLER_226_920 ();
 sg13g2_fill_8 FILLER_226_928 ();
 sg13g2_fill_8 FILLER_226_936 ();
 sg13g2_fill_8 FILLER_226_944 ();
 sg13g2_fill_8 FILLER_226_952 ();
 sg13g2_fill_8 FILLER_226_960 ();
 sg13g2_fill_8 FILLER_226_968 ();
 sg13g2_fill_8 FILLER_226_976 ();
 sg13g2_fill_8 FILLER_226_984 ();
 sg13g2_fill_8 FILLER_226_992 ();
 sg13g2_fill_8 FILLER_226_1000 ();
 sg13g2_fill_8 FILLER_226_1008 ();
 sg13g2_fill_8 FILLER_226_1016 ();
 sg13g2_fill_8 FILLER_226_1024 ();
 sg13g2_fill_8 FILLER_226_1032 ();
 sg13g2_fill_8 FILLER_226_1040 ();
 sg13g2_fill_8 FILLER_226_1048 ();
 sg13g2_fill_8 FILLER_226_1056 ();
 sg13g2_fill_8 FILLER_226_1064 ();
 sg13g2_fill_8 FILLER_226_1072 ();
 sg13g2_fill_8 FILLER_226_1080 ();
 sg13g2_fill_8 FILLER_226_1088 ();
 sg13g2_fill_8 FILLER_226_1096 ();
 sg13g2_fill_8 FILLER_226_1104 ();
 sg13g2_fill_8 FILLER_226_1112 ();
 sg13g2_fill_8 FILLER_226_1120 ();
 sg13g2_fill_8 FILLER_226_1128 ();
 sg13g2_fill_8 FILLER_226_1136 ();
 sg13g2_fill_8 FILLER_226_1144 ();
 sg13g2_fill_8 FILLER_226_1152 ();
 sg13g2_fill_8 FILLER_226_1160 ();
 sg13g2_fill_8 FILLER_226_1168 ();
 sg13g2_fill_8 FILLER_226_1176 ();
 sg13g2_fill_8 FILLER_226_1184 ();
 sg13g2_fill_8 FILLER_226_1192 ();
 sg13g2_fill_8 FILLER_226_1200 ();
 sg13g2_fill_8 FILLER_226_1208 ();
 sg13g2_fill_8 FILLER_226_1216 ();
 sg13g2_fill_8 FILLER_226_1224 ();
 sg13g2_fill_8 FILLER_226_1232 ();
 sg13g2_fill_8 FILLER_226_1240 ();
 sg13g2_fill_8 FILLER_226_1248 ();
 sg13g2_fill_8 FILLER_226_1256 ();
 sg13g2_fill_8 FILLER_226_1264 ();
 sg13g2_fill_8 FILLER_226_1272 ();
 sg13g2_fill_8 FILLER_226_1280 ();
 sg13g2_fill_8 FILLER_226_1288 ();
 sg13g2_fill_8 FILLER_226_1296 ();
 sg13g2_fill_8 FILLER_226_1304 ();
 sg13g2_fill_8 FILLER_226_1312 ();
 sg13g2_fill_8 FILLER_226_1320 ();
 sg13g2_fill_8 FILLER_226_1328 ();
 sg13g2_fill_8 FILLER_226_1336 ();
 sg13g2_fill_8 FILLER_226_1344 ();
 sg13g2_fill_8 FILLER_226_1352 ();
 sg13g2_fill_8 FILLER_226_1360 ();
 sg13g2_fill_8 FILLER_226_1368 ();
 sg13g2_fill_8 FILLER_226_1376 ();
 sg13g2_fill_8 FILLER_226_1384 ();
 sg13g2_fill_8 FILLER_226_1392 ();
 sg13g2_fill_8 FILLER_226_1400 ();
 sg13g2_fill_8 FILLER_226_1408 ();
 sg13g2_fill_8 FILLER_226_1416 ();
 sg13g2_fill_8 FILLER_226_1424 ();
 sg13g2_fill_8 FILLER_226_1432 ();
 sg13g2_fill_8 FILLER_226_1440 ();
 sg13g2_fill_8 FILLER_226_1448 ();
 sg13g2_fill_8 FILLER_226_1456 ();
 sg13g2_fill_8 FILLER_226_1464 ();
 sg13g2_fill_8 FILLER_226_1472 ();
 sg13g2_fill_8 FILLER_226_1480 ();
 sg13g2_fill_8 FILLER_226_1488 ();
 sg13g2_fill_8 FILLER_226_1496 ();
 sg13g2_fill_8 FILLER_226_1504 ();
 sg13g2_fill_8 FILLER_226_1512 ();
 sg13g2_fill_8 FILLER_226_1520 ();
 sg13g2_fill_8 FILLER_226_1528 ();
 sg13g2_fill_8 FILLER_226_1536 ();
 sg13g2_fill_8 FILLER_226_1544 ();
 sg13g2_fill_8 FILLER_226_1552 ();
 sg13g2_fill_8 FILLER_226_1560 ();
 sg13g2_fill_8 FILLER_226_1568 ();
 sg13g2_fill_8 FILLER_226_1576 ();
 sg13g2_fill_8 FILLER_226_1584 ();
 sg13g2_fill_8 FILLER_227_0 ();
 sg13g2_fill_8 FILLER_227_8 ();
 sg13g2_fill_8 FILLER_227_16 ();
 sg13g2_fill_8 FILLER_227_24 ();
 sg13g2_fill_8 FILLER_227_32 ();
 sg13g2_fill_8 FILLER_227_40 ();
 sg13g2_fill_8 FILLER_227_48 ();
 sg13g2_fill_8 FILLER_227_56 ();
 sg13g2_fill_8 FILLER_227_64 ();
 sg13g2_fill_8 FILLER_227_72 ();
 sg13g2_fill_8 FILLER_227_80 ();
 sg13g2_fill_8 FILLER_227_88 ();
 sg13g2_fill_8 FILLER_227_96 ();
 sg13g2_fill_8 FILLER_227_104 ();
 sg13g2_fill_8 FILLER_227_112 ();
 sg13g2_fill_8 FILLER_227_120 ();
 sg13g2_fill_8 FILLER_227_128 ();
 sg13g2_fill_8 FILLER_227_136 ();
 sg13g2_fill_8 FILLER_227_144 ();
 sg13g2_fill_8 FILLER_227_152 ();
 sg13g2_fill_8 FILLER_227_160 ();
 sg13g2_fill_8 FILLER_227_168 ();
 sg13g2_fill_8 FILLER_227_176 ();
 sg13g2_fill_8 FILLER_227_184 ();
 sg13g2_fill_8 FILLER_227_192 ();
 sg13g2_fill_8 FILLER_227_200 ();
 sg13g2_fill_8 FILLER_227_208 ();
 sg13g2_fill_8 FILLER_227_216 ();
 sg13g2_fill_8 FILLER_227_224 ();
 sg13g2_fill_8 FILLER_227_232 ();
 sg13g2_fill_8 FILLER_227_240 ();
 sg13g2_fill_8 FILLER_227_248 ();
 sg13g2_fill_8 FILLER_227_256 ();
 sg13g2_fill_8 FILLER_227_264 ();
 sg13g2_fill_8 FILLER_227_272 ();
 sg13g2_fill_8 FILLER_227_280 ();
 sg13g2_fill_8 FILLER_227_288 ();
 sg13g2_fill_8 FILLER_227_296 ();
 sg13g2_fill_8 FILLER_227_304 ();
 sg13g2_fill_8 FILLER_227_312 ();
 sg13g2_fill_8 FILLER_227_320 ();
 sg13g2_fill_8 FILLER_227_328 ();
 sg13g2_fill_8 FILLER_227_336 ();
 sg13g2_fill_8 FILLER_227_344 ();
 sg13g2_fill_8 FILLER_227_352 ();
 sg13g2_fill_8 FILLER_227_360 ();
 sg13g2_fill_8 FILLER_227_368 ();
 sg13g2_fill_8 FILLER_227_376 ();
 sg13g2_fill_8 FILLER_227_384 ();
 sg13g2_fill_8 FILLER_227_392 ();
 sg13g2_fill_8 FILLER_227_400 ();
 sg13g2_fill_8 FILLER_227_408 ();
 sg13g2_fill_8 FILLER_227_416 ();
 sg13g2_fill_8 FILLER_227_424 ();
 sg13g2_fill_8 FILLER_227_432 ();
 sg13g2_fill_8 FILLER_227_440 ();
 sg13g2_fill_8 FILLER_227_448 ();
 sg13g2_fill_8 FILLER_227_456 ();
 sg13g2_fill_8 FILLER_227_464 ();
 sg13g2_fill_8 FILLER_227_472 ();
 sg13g2_fill_8 FILLER_227_480 ();
 sg13g2_fill_8 FILLER_227_488 ();
 sg13g2_fill_8 FILLER_227_496 ();
 sg13g2_fill_8 FILLER_227_504 ();
 sg13g2_fill_8 FILLER_227_512 ();
 sg13g2_fill_8 FILLER_227_520 ();
 sg13g2_fill_8 FILLER_227_528 ();
 sg13g2_fill_8 FILLER_227_536 ();
 sg13g2_fill_8 FILLER_227_544 ();
 sg13g2_fill_8 FILLER_227_552 ();
 sg13g2_fill_8 FILLER_227_560 ();
 sg13g2_fill_8 FILLER_227_568 ();
 sg13g2_fill_8 FILLER_227_576 ();
 sg13g2_fill_8 FILLER_227_584 ();
 sg13g2_fill_8 FILLER_227_592 ();
 sg13g2_fill_8 FILLER_227_600 ();
 sg13g2_fill_8 FILLER_227_608 ();
 sg13g2_fill_8 FILLER_227_616 ();
 sg13g2_fill_8 FILLER_227_624 ();
 sg13g2_fill_8 FILLER_227_632 ();
 sg13g2_fill_8 FILLER_227_640 ();
 sg13g2_fill_8 FILLER_227_648 ();
 sg13g2_fill_8 FILLER_227_656 ();
 sg13g2_fill_8 FILLER_227_664 ();
 sg13g2_fill_8 FILLER_227_672 ();
 sg13g2_fill_8 FILLER_227_680 ();
 sg13g2_fill_8 FILLER_227_688 ();
 sg13g2_fill_8 FILLER_227_696 ();
 sg13g2_fill_8 FILLER_227_704 ();
 sg13g2_fill_8 FILLER_227_712 ();
 sg13g2_fill_8 FILLER_227_720 ();
 sg13g2_fill_8 FILLER_227_728 ();
 sg13g2_fill_8 FILLER_227_736 ();
 sg13g2_fill_8 FILLER_227_744 ();
 sg13g2_fill_8 FILLER_227_752 ();
 sg13g2_fill_8 FILLER_227_760 ();
 sg13g2_fill_8 FILLER_227_768 ();
 sg13g2_fill_8 FILLER_227_776 ();
 sg13g2_fill_8 FILLER_227_784 ();
 sg13g2_fill_8 FILLER_227_792 ();
 sg13g2_fill_8 FILLER_227_800 ();
 sg13g2_fill_8 FILLER_227_808 ();
 sg13g2_fill_8 FILLER_227_816 ();
 sg13g2_fill_8 FILLER_227_824 ();
 sg13g2_fill_8 FILLER_227_832 ();
 sg13g2_fill_8 FILLER_227_840 ();
 sg13g2_fill_8 FILLER_227_848 ();
 sg13g2_fill_8 FILLER_227_856 ();
 sg13g2_fill_8 FILLER_227_864 ();
 sg13g2_fill_8 FILLER_227_872 ();
 sg13g2_fill_8 FILLER_227_880 ();
 sg13g2_fill_8 FILLER_227_888 ();
 sg13g2_fill_8 FILLER_227_896 ();
 sg13g2_fill_8 FILLER_227_904 ();
 sg13g2_fill_8 FILLER_227_912 ();
 sg13g2_fill_8 FILLER_227_920 ();
 sg13g2_fill_8 FILLER_227_928 ();
 sg13g2_fill_8 FILLER_227_936 ();
 sg13g2_fill_8 FILLER_227_944 ();
 sg13g2_fill_8 FILLER_227_952 ();
 sg13g2_fill_8 FILLER_227_960 ();
 sg13g2_fill_8 FILLER_227_968 ();
 sg13g2_fill_8 FILLER_227_976 ();
 sg13g2_fill_8 FILLER_227_984 ();
 sg13g2_fill_8 FILLER_227_992 ();
 sg13g2_fill_8 FILLER_227_1000 ();
 sg13g2_fill_8 FILLER_227_1008 ();
 sg13g2_fill_8 FILLER_227_1016 ();
 sg13g2_fill_8 FILLER_227_1024 ();
 sg13g2_fill_8 FILLER_227_1032 ();
 sg13g2_fill_8 FILLER_227_1040 ();
 sg13g2_fill_8 FILLER_227_1048 ();
 sg13g2_fill_8 FILLER_227_1056 ();
 sg13g2_fill_8 FILLER_227_1064 ();
 sg13g2_fill_8 FILLER_227_1072 ();
 sg13g2_fill_8 FILLER_227_1080 ();
 sg13g2_fill_8 FILLER_227_1088 ();
 sg13g2_fill_8 FILLER_227_1096 ();
 sg13g2_fill_8 FILLER_227_1104 ();
 sg13g2_fill_8 FILLER_227_1112 ();
 sg13g2_fill_8 FILLER_227_1120 ();
 sg13g2_fill_8 FILLER_227_1128 ();
 sg13g2_fill_8 FILLER_227_1136 ();
 sg13g2_fill_8 FILLER_227_1144 ();
 sg13g2_fill_8 FILLER_227_1152 ();
 sg13g2_fill_8 FILLER_227_1160 ();
 sg13g2_fill_8 FILLER_227_1168 ();
 sg13g2_fill_8 FILLER_227_1176 ();
 sg13g2_fill_8 FILLER_227_1184 ();
 sg13g2_fill_8 FILLER_227_1192 ();
 sg13g2_fill_8 FILLER_227_1200 ();
 sg13g2_fill_8 FILLER_227_1208 ();
 sg13g2_fill_8 FILLER_227_1216 ();
 sg13g2_fill_8 FILLER_227_1224 ();
 sg13g2_fill_8 FILLER_227_1232 ();
 sg13g2_fill_8 FILLER_227_1240 ();
 sg13g2_fill_8 FILLER_227_1248 ();
 sg13g2_fill_8 FILLER_227_1256 ();
 sg13g2_fill_8 FILLER_227_1264 ();
 sg13g2_fill_8 FILLER_227_1272 ();
 sg13g2_fill_8 FILLER_227_1280 ();
 sg13g2_fill_8 FILLER_227_1288 ();
 sg13g2_fill_8 FILLER_227_1296 ();
 sg13g2_fill_8 FILLER_227_1304 ();
 sg13g2_fill_8 FILLER_227_1312 ();
 sg13g2_fill_8 FILLER_227_1320 ();
 sg13g2_fill_8 FILLER_227_1328 ();
 sg13g2_fill_8 FILLER_227_1336 ();
 sg13g2_fill_8 FILLER_227_1344 ();
 sg13g2_fill_8 FILLER_227_1352 ();
 sg13g2_fill_8 FILLER_227_1360 ();
 sg13g2_fill_8 FILLER_227_1368 ();
 sg13g2_fill_8 FILLER_227_1376 ();
 sg13g2_fill_8 FILLER_227_1384 ();
 sg13g2_fill_8 FILLER_227_1392 ();
 sg13g2_fill_8 FILLER_227_1400 ();
 sg13g2_fill_8 FILLER_227_1408 ();
 sg13g2_fill_8 FILLER_227_1416 ();
 sg13g2_fill_8 FILLER_227_1424 ();
 sg13g2_fill_8 FILLER_227_1432 ();
 sg13g2_fill_8 FILLER_227_1440 ();
 sg13g2_fill_8 FILLER_227_1448 ();
 sg13g2_fill_8 FILLER_227_1456 ();
 sg13g2_fill_8 FILLER_227_1464 ();
 sg13g2_fill_8 FILLER_227_1472 ();
 sg13g2_fill_8 FILLER_227_1480 ();
 sg13g2_fill_8 FILLER_227_1488 ();
 sg13g2_fill_8 FILLER_227_1496 ();
 sg13g2_fill_8 FILLER_227_1504 ();
 sg13g2_fill_8 FILLER_227_1512 ();
 sg13g2_fill_8 FILLER_227_1520 ();
 sg13g2_fill_8 FILLER_227_1528 ();
 sg13g2_fill_8 FILLER_227_1536 ();
 sg13g2_fill_8 FILLER_227_1544 ();
 sg13g2_fill_8 FILLER_227_1552 ();
 sg13g2_fill_8 FILLER_227_1560 ();
 sg13g2_fill_8 FILLER_227_1568 ();
 sg13g2_fill_8 FILLER_227_1576 ();
 sg13g2_fill_8 FILLER_227_1584 ();
 assign crash_dump_o_64_ = net1;
 assign data_addr_o_0_ = net2;
 assign data_addr_o_1_ = net3;
 assign instr_addr_o_0_ = net4;
 assign instr_addr_o_1_ = net5;
endmodule
