//Latest Update Date: 9th Aug, 2025
//Owner: B Nithin Reddy

//Interface  
interface dff_if;
  
  logic reset;
  logic D;
  logic Q;
  logic clock;
  
endinterface
