VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA croc_chip_via6_7_10000_10000_5_5_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.63 0.5 ;
  ROWCOL 5 5 ;
END croc_chip_via6_7_10000_10000_5_5_1960_1960

VIA croc_chip_via6_7_13330_18000_9_6_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 1.315 0.71 1.315 0.5 ;
  ROWCOL 9 6 ;
END croc_chip_via6_7_13330_18000_9_6_1960_1960

VIA croc_chip_via6_7_13330_10000_5_6_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 1.315 0.5 ;
  ROWCOL 5 6 ;
END croc_chip_via6_7_13330_10000_5_6_1960_1960

VIA croc_chip_via6_7_20000_10000_5_10_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.73 0.5 ;
  ROWCOL 5 10 ;
END croc_chip_via6_7_20000_10000_5_10_1960_1960

VIA croc_chip_via6_7_20000_18000_9_10_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.73 0.71 0.73 0.5 ;
  ROWCOL 9 10 ;
END croc_chip_via6_7_20000_18000_9_10_1960_1960

VIA croc_chip_via6_7_8330_18000_9_4_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.775 0.71 0.775 0.5 ;
  ROWCOL 9 4 ;
END croc_chip_via6_7_8330_18000_9_4_1960_1960

VIA croc_chip_via6_7_8330_10000_5_4_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.775 0.5 ;
  ROWCOL 5 4 ;
END croc_chip_via6_7_8330_10000_5_4_1960_1960

VIA croc_chip_via6_7_6000_10000_5_3_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 0.59 0.5 ;
  ROWCOL 5 3 ;
END croc_chip_via6_7_6000_10000_5_3_1960_1960

VIA croc_chip_via6_7_3330_18000_9_1_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 1.215 0.71 1.215 0.5 ;
  ROWCOL 9 1 ;
END croc_chip_via6_7_3330_18000_9_1_1960_1960

VIA croc_chip_via6_7_3330_10000_5_1_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.63 1.215 0.5 ;
  ROWCOL 5 1 ;
END croc_chip_via6_7_3330_10000_5_1_1960_1960

VIA croc_chip_via3_4_2000_2000_4_4_480_480
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.185 0.05 0.05 0.185 ;
  ROWCOL 4 4 ;
END croc_chip_via3_4_2000_2000_4_4_480_480

VIA croc_chip_via3_4_2000_6000_12_4_480_480
  VIARULE via3Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal3 Via3 Metal4 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.185 0.05 0.05 0.005 ;
  ROWCOL 12 4 ;
END croc_chip_via3_4_2000_6000_12_4_480_480

VIA croc_chip_via4_5_2000_6000_12_4_480_480
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.05 0.005 0.005 0.05 ;
  ROWCOL 12 4 ;
END croc_chip_via4_5_2000_6000_12_4_480_480

VIA croc_chip_via5_6_2000_6000_6_1_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.69 ;
  ROWCOL 6 1 ;
END croc_chip_via5_6_2000_6000_6_1_840_840

VIA croc_chip_via4_5_2810_6000_12_6_480_480
  VIARULE via4Array ;
  CUTSIZE 0.19 0.19 ;
  LAYERS Metal4 Via4 Metal5 ;
  CUTSPACING 0.29 0.29 ;
  ENCLOSURE 0.11 0.265 0.005 0.05 ;
  ROWCOL 12 6 ;
END croc_chip_via4_5_2810_6000_12_6_480_480

VIA croc_chip_via5_6_2810_6000_6_2_840_840
  VIARULE viagen56 ;
  CUTSIZE 0.42 0.42 ;
  LAYERS Metal5 TopVia1 TopMetal1 ;
  CUTSPACING 0.42 0.42 ;
  ENCLOSURE 0.1 0.1 0.42 0.69 ;
  ROWCOL 6 2 ;
END croc_chip_via5_6_2810_6000_6_2_840_840

VIA croc_chip_via6_7_6000_6000_3_3_1960_1960
  VIARULE viagen67 ;
  CUTSIZE 0.9 0.9 ;
  LAYERS TopMetal1 TopVia2 TopMetal2 ;
  CUTSPACING 1.06 1.06 ;
  ENCLOSURE 0.5 0.59 0.59 0.5 ;
  ROWCOL 3 3 ;
END croc_chip_via6_7_6000_6000_3_3_1960_1960

MACRO croc_chip
  FOREIGN croc_chip 0 0 ;
  CLASS BLOCK ;
  SIZE 3470 BY 3470 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1961 0 2031 ;
    END
  END clk_i
  PIN fetch_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 2349 0 2419 ;
    END
  END fetch_en_i
  PIN gpio0_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  593 -70 663 0 ;
    END
  END gpio0_io
  PIN gpio10_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2533 -70 2603 0 ;
    END
  END gpio10_io
  PIN gpio11_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2727 -70 2797 0 ;
    END
  END gpio11_io
  PIN gpio12_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 593 3470 663 ;
    END
  END gpio12_io
  PIN gpio13_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 787 3470 857 ;
    END
  END gpio13_io
  PIN gpio14_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 981 3470 1051 ;
    END
  END gpio14_io
  PIN gpio15_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 1175 3470 1245 ;
    END
  END gpio15_io
  PIN gpio16_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 1369 3470 1439 ;
    END
  END gpio16_io
  PIN gpio17_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 1563 3470 1633 ;
    END
  END gpio17_io
  PIN gpio18_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 1757 3470 1827 ;
    END
  END gpio18_io
  PIN gpio19_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 1951 3470 2021 ;
    END
  END gpio19_io
  PIN gpio1_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  787 -70 857 0 ;
    END
  END gpio1_io
  PIN gpio20_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 2145 3470 2215 ;
    END
  END gpio20_io
  PIN gpio21_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 2339 3470 2409 ;
    END
  END gpio21_io
  PIN gpio22_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 2533 3470 2603 ;
    END
  END gpio22_io
  PIN gpio23_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  3400 2727 3470 2797 ;
    END
  END gpio23_io
  PIN gpio24_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2737 3400 2807 3470 ;
    END
  END gpio24_io
  PIN gpio25_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2543 3400 2613 3470 ;
    END
  END gpio25_io
  PIN gpio26_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2349 3400 2419 3470 ;
    END
  END gpio26_io
  PIN gpio27_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2155 3400 2225 3470 ;
    END
  END gpio27_io
  PIN gpio28_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1961 3400 2031 3470 ;
    END
  END gpio28_io
  PIN gpio29_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1767 3400 1837 3470 ;
    END
  END gpio29_io
  PIN gpio2_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  981 -70 1051 0 ;
    END
  END gpio2_io
  PIN gpio30_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1573 3400 1643 3470 ;
    END
  END gpio30_io
  PIN gpio31_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1379 3400 1449 3470 ;
    END
  END gpio31_io
  PIN gpio3_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1175 -70 1245 0 ;
    END
  END gpio3_io
  PIN gpio4_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1369 -70 1439 0 ;
    END
  END gpio4_io
  PIN gpio5_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1563 -70 1633 0 ;
    END
  END gpio5_io
  PIN gpio6_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1757 -70 1827 0 ;
    END
  END gpio6_io
  PIN gpio7_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1951 -70 2021 0 ;
    END
  END gpio7_io
  PIN gpio8_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2145 -70 2215 0 ;
    END
  END gpio8_io
  PIN gpio9_io
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  2339 -70 2409 0 ;
    END
  END gpio9_io
  PIN jtag_tck_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1379 0 1449 ;
    END
  END jtag_tck_i
  PIN jtag_tdi_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 797 0 867 ;
    END
  END jtag_tdi_i
  PIN jtag_tdo_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 603 0 673 ;
    END
  END jtag_tdo_o
  PIN jtag_tms_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 991 0 1061 ;
    END
  END jtag_tms_i
  PIN jtag_trst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1185 0 1255 ;
    END
  END jtag_trst_ni
  PIN ref_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1767 0 1837 ;
    END
  END ref_clk_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 1573 0 1643 ;
    END
  END rst_ni
  PIN status_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 2155 0 2225 ;
    END
  END status_o
  PIN uart_rx_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 2737 0 2807 ;
    END
  END uart_rx_i
  PIN uart_tx_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  -70 2543 0 2613 ;
    END
  END uart_tx_o
  PIN unused0_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  1185 3400 1255 3470 ;
    END
  END unused0_o
  PIN unused1_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  991 3400 1061 3470 ;
    END
  END unused1_o
  PIN unused2_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  797 3400 867 3470 ;
    END
  END unused2_o
  PIN unused3_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER TopMetal2 ;
        RECT  603 3400 673 3470 ;
    END
  END unused3_o
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER TopMetal2 ;
        RECT  215 3400 285 3470 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  3400 3115 3470 3185 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  3115 -70 3185 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 215 0 285 ;
    END
  END VDD
  PIN VDDIO
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER TopMetal2 ;
        RECT  2931 3400 3001 3470 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  3400 399 3470 469 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  399 -70 469 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 2931 0 3001 ;
    END
  END VDDIO
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal2 ;
        RECT  409 3400 479 3470 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  3400 2921 3470 2991 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  2921 -70 2991 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 409 0 479 ;
    END
  END VSS
  PIN VSSIO
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal2 ;
        RECT  3125 3400 3195 3470 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  3400 205 3470 275 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  205 -70 275 0 ;
    END
    PORT
      LAYER TopMetal2 ;
        RECT  -70 3125 0 3195 ;
    END
  END VSSIO
  OBS
    LAYER Metal1 ;
     RECT  205 -70 275 0 ;
     RECT  399 -70 469 0 ;
     RECT  593 -70 663 0 ;
     RECT  787 -70 857 0 ;
     RECT  981 -70 1051 0 ;
     RECT  1175 -70 1245 0 ;
     RECT  1369 -70 1439 0 ;
     RECT  1563 -70 1633 0 ;
     RECT  1757 -70 1827 0 ;
     RECT  1951 -70 2021 0 ;
     RECT  2145 -70 2215 0 ;
     RECT  2339 -70 2409 0 ;
     RECT  2533 -70 2603 0 ;
     RECT  2727 -70 2797 0 ;
     RECT  2921 -70 2991 0 ;
     RECT  3115 -70 3185 0 ;
     RECT  0 0 3400 180 ;
     RECT  3220 180 3400 205 ;
     RECT  0 180 180 215 ;
     RECT  3220 205 3470 275 ;
     RECT  -70 215 180 285 ;
     RECT  3220 275 3400 399 ;
     RECT  0 285 180 409 ;
     RECT  3220 399 3470 469 ;
     RECT  -70 409 180 479 ;
     RECT  3220 469 3400 593 ;
     RECT  200.16 200.12 3199.68 593.68 ;
     RECT  0 479 180 603 ;
     RECT  3220 593 3470 663 ;
     RECT  -70 603 180 673 ;
     RECT  200.16 593.68 994.56 772.12 ;
     RECT  1392.56 751.54 1392.72 782.36 ;
     RECT  3220 663 3400 787 ;
     RECT  0 673 180 797 ;
     RECT  1392.08 798.58 1392.24 799 ;
     RECT  1392.08 799 1394.16 824.78 ;
     RECT  200.16 772.12 1001.04 827.3 ;
     RECT  1392.08 824.78 1392.24 829.82 ;
     RECT  3220 787 3470 857 ;
     RECT  -70 797 180 867 ;
     RECT  3220 857 3400 981 ;
     RECT  200.16 827.3 994.56 986.36 ;
     RECT  1020.16 622.46 1379.68 986.36 ;
     RECT  1405.44 593.68 3199.68 986.36 ;
     RECT  0 867 180 991 ;
     RECT  200.16 986.36 3199.68 994.36 ;
     RECT  3220 981 3470 1051 ;
     RECT  -70 991 180 1061 ;
     RECT  3220 1051 3400 1175 ;
     RECT  0 1061 180 1185 ;
     RECT  3220 1175 3470 1245 ;
     RECT  -70 1185 180 1255 ;
     RECT  3220 1245 3400 1369 ;
     RECT  0 1255 180 1379 ;
     RECT  3220 1369 3470 1439 ;
     RECT  -70 1379 180 1449 ;
     RECT  3105.12 994.36 3199.68 1474.1 ;
     RECT  1825.44 1026.24 3074.88 1498.04 ;
     RECT  1825.44 1498.04 3075.44 1499.88 ;
     RECT  3088.72 1494.26 3088.88 1500.3 ;
     RECT  3088.72 1521.98 3088.88 1528.44 ;
     RECT  1825.44 1499.88 3074.88 1529.54 ;
     RECT  1825.44 1529.54 3075.44 1537.1 ;
     RECT  1825.44 1537.1 3081.2 1539.78 ;
     RECT  3098.8 1474.1 3199.68 1544.4 ;
     RECT  3220 1439 3400 1563 ;
     RECT  200.16 994.36 1794.72 1566.08 ;
     RECT  0 1449 180 1573 ;
     RECT  3105.12 1544.4 3199.68 1574.9 ;
     RECT  3097.36 1574.9 3199.68 1577.42 ;
     RECT  1825.44 1539.78 3074.88 1577.715 ;
     RECT  1825.44 1577.715 3074.96 1587.5 ;
     RECT  3096.4 1577.42 3199.68 1600.1 ;
     RECT  3089.68 1600.1 3199.68 1631.18 ;
     RECT  3220 1563 3470 1633 ;
     RECT  200.16 1566.08 1801.04 1634.96 ;
     RECT  -70 1573 180 1643 ;
     RECT  200.16 1634.96 1803.92 1645.88 ;
     RECT  1825.44 1587.5 3077.84 1646.46 ;
     RECT  200.16 1645.88 1805.36 1678.38 ;
     RECT  3088.72 1631.18 3199.68 1678.38 ;
     RECT  200.16 1678.38 1801.04 1680.9 ;
     RECT  3089.2 1678.38 3199.68 1691.24 ;
     RECT  1825.44 1646.46 3074.88 1728.62 ;
     RECT  3084.88 1691.24 3199.68 1728.62 ;
     RECT  3220 1633 3400 1757 ;
     RECT  0 1643 180 1767 ;
     RECT  1825.44 1728.62 3199.68 1773.3 ;
     RECT  200.16 1680.9 1794.72 1778.62 ;
     RECT  200.16 1778.62 1795.28 1796.42 ;
     RECT  3084.88 1773.3 3199.68 1804.38 ;
     RECT  3220 1757 3470 1827 ;
     RECT  3088.72 1804.38 3199.68 1833.78 ;
     RECT  200.16 1796.42 1794.72 1834.9 ;
     RECT  -70 1767 180 1837 ;
     RECT  200.16 1834.9 1795.28 1845.98 ;
     RECT  200.16 1845.98 1794.8 1846.4 ;
     RECT  1825.44 1773.3 3074.88 1867.64 ;
     RECT  1825.44 1867.64 3077.84 1920.3 ;
     RECT  3091.6 1833.78 3199.68 1921.4 ;
     RECT  3088.72 1921.4 3199.68 1940.46 ;
     RECT  3091.6 1940.46 3199.68 1942.98 ;
     RECT  3091.6 1942.98 3091.76 1945.5 ;
     RECT  3220 1827 3400 1951 ;
     RECT  0 1837 180 1961 ;
     RECT  200.16 1846.4 1794.72 1992.28 ;
     RECT  1825.44 1920.3 3074.88 1992.8 ;
     RECT  1303.6 1992.28 1794.72 1992.98 ;
     RECT  3105.12 1942.98 3199.68 2007.08 ;
     RECT  1825.44 1992.8 3075.92 2019.68 ;
     RECT  3088.72 1996.58 3088.88 2019.68 ;
     RECT  3220 1951 3470 2021 ;
     RECT  1825.44 2019.68 3088.88 2027.24 ;
     RECT  3098.8 2007.08 3199.68 2027.24 ;
     RECT  -70 1961 180 2031 ;
     RECT  1825.44 2027.24 3199.68 2041.26 ;
     RECT  3097.36 2041.26 3199.68 2048.82 ;
     RECT  3098.8 2048.82 3199.68 2051.34 ;
     RECT  1825.44 2041.26 3084.08 2053.86 ;
     RECT  200.16 1992.28 694.56 2065.86 ;
     RECT  200.16 2065.86 701.04 2088.54 ;
     RECT  720.16 2022.46 1279.84 2088.54 ;
     RECT  1305.12 1992.98 1794.72 2095.72 ;
     RECT  1305.12 2095.72 1795.28 2103.44 ;
     RECT  1305.12 2103.44 1794.72 2122.6 ;
     RECT  1305.12 2122.6 1795.28 2129.32 ;
     RECT  1303.12 2129.32 1795.28 2129.9 ;
     RECT  1303.12 2129.9 1794.72 2132.42 ;
     RECT  1304.56 2132.42 1794.72 2142.08 ;
     RECT  3220 2021 3400 2145 ;
     RECT  0 2031 180 2155 ;
     RECT  1305.12 2142.08 1794.72 2176.74 ;
     RECT  1298.96 2176.74 1794.72 2181.78 ;
     RECT  1298 2181.78 1794.72 2189.34 ;
     RECT  1295.6 2189.34 1794.72 2198.62 ;
     RECT  1295.6 2198.62 1799.6 2199.04 ;
     RECT  1295.6 2199.04 1800.08 2199.2 ;
     RECT  1295.6 2199.2 1794.72 2205.04 ;
     RECT  3220 2145 3470 2215 ;
     RECT  1297.04 2205.04 1794.72 2219.58 ;
     RECT  1294.16 2219.58 1794.72 2222.1 ;
     RECT  -70 2155 180 2225 ;
     RECT  1293.68 2222.1 1794.72 2227.14 ;
     RECT  1290.32 2227.14 1794.72 2239.36 ;
     RECT  1290.32 2239.36 1794.8 2240.78 ;
     RECT  1290.32 2240.78 1794.72 2242 ;
     RECT  1293.68 2242 1794.72 2249.14 ;
     RECT  1296.08 2249.14 1794.72 2255.74 ;
     RECT  1296.08 2255.74 1794.8 2263.42 ;
     RECT  1297.04 2263.42 1794.8 2279.12 ;
     RECT  1825.44 2053.86 3074.88 2279.12 ;
     RECT  3105.12 2051.34 3199.68 2279.12 ;
     RECT  3220 2215 3400 2339 ;
     RECT  0 2225 180 2349 ;
     RECT  1297.04 2279.12 3199.68 2363.22 ;
     RECT  1289.84 2363.22 3199.68 2364.64 ;
     RECT  1297.04 2364.64 3199.68 2366.32 ;
     RECT  200.16 2088.54 1279.84 2370.52 ;
     RECT  200.16 2370.52 702.48 2391.78 ;
     RECT  200.16 2391.78 704.88 2392.2 ;
     RECT  200.16 2392.2 706.32 2393.46 ;
     RECT  200.16 2393.46 707.28 2406.22 ;
     RECT  3220 2339 3470 2409 ;
     RECT  200.16 2406.22 706.8 2416.3 ;
     RECT  -70 2349 180 2419 ;
     RECT  200.16 2416.3 704.88 2423.86 ;
     RECT  200.16 2423.86 702.48 2461.66 ;
     RECT  1297.52 2366.32 3199.68 2461.66 ;
     RECT  717.68 2370.52 1279.84 2479.3 ;
     RECT  200.16 2461.66 702 2481.82 ;
     RECT  200.16 2481.82 701.52 2504.5 ;
     RECT  200.16 2504.5 701.04 2522.14 ;
     RECT  200.16 2522.14 700.56 2529.28 ;
     RECT  3220 2409 3400 2533 ;
     RECT  0 2419 180 2543 ;
     RECT  200.16 2529.28 694.56 2585.3 ;
     RECT  720.16 2479.3 1279.84 2585.3 ;
     RECT  1305.12 2461.66 3199.68 2585.3 ;
     RECT  3220 2533 3470 2603 ;
     RECT  -70 2543 180 2613 ;
     RECT  3220 2603 3400 2727 ;
     RECT  0 2613 180 2737 ;
     RECT  3220 2727 3470 2797 ;
     RECT  -70 2737 180 2807 ;
     RECT  3220 2797 3400 2921 ;
     RECT  0 2807 180 2931 ;
     RECT  3220 2921 3470 2991 ;
     RECT  -70 2931 180 3001 ;
     RECT  200.16 2585.3 3199.68 3044.1 ;
     RECT  1323.76 3044.1 1325.84 3053.74 ;
     RECT  1323.28 3053.74 1325.84 3054.16 ;
     RECT  1338.16 3044.1 1339.28 3054.16 ;
     RECT  2012.56 3044.1 2012.72 3054.16 ;
     RECT  2043.28 3044.1 2043.44 3054.16 ;
     RECT  2055.28 3044.1 2055.44 3054.16 ;
     RECT  2065.36 3053.74 2065.52 3054.16 ;
     RECT  2078.8 3044.1 2081.36 3054.16 ;
     RECT  1323.28 3054.16 1339.28 3054.58 ;
     RECT  2025.52 3053.74 2025.68 3054.58 ;
     RECT  2035.6 3054.16 2043.44 3054.58 ;
     RECT  2055.28 3054.16 2081.36 3054.58 ;
     RECT  1323.28 3054.58 1341.68 3055 ;
     RECT  1401.04 3054.58 1401.2 3055 ;
     RECT  1979.92 3054.16 1980.08 3055 ;
     RECT  200.16 3044.1 1302.8 3055.42 ;
     RECT  1378.48 3054.16 1378.64 3055.42 ;
     RECT  200.16 3055.42 1310 3055.84 ;
     RECT  1378.48 3055.42 1380.08 3055.84 ;
     RECT  1581.04 3055.42 1581.2 3055.84 ;
     RECT  1614.16 3055.42 1614.32 3055.84 ;
     RECT  2002 3054.16 2002.16 3055.84 ;
     RECT  2025.52 3054.58 2081.36 3055.84 ;
     RECT  2092.72 3044.1 3199.68 3055.84 ;
     RECT  1700.08 3055.84 1700.24 3056.26 ;
     RECT  1998.16 3055.84 2002.16 3056.68 ;
     RECT  2012.56 3054.16 2013.2 3056.68 ;
     RECT  200.16 3055.84 1310.48 3057.1 ;
     RECT  1321.36 3055 1341.68 3057.1 ;
     RECT  1632.88 3056.68 1633.04 3057.1 ;
     RECT  1923.28 3055.42 1923.44 3057.94 ;
     RECT  200.16 3057.1 1341.68 3059.1 ;
     RECT  1352.08 3044.1 1353.2 3059.1 ;
     RECT  1363.6 3044.1 1363.76 3059.1 ;
     RECT  1374.64 3055.84 1380.08 3059.1 ;
     RECT  1391.92 3055 1402.64 3059.1 ;
     RECT  1420.72 3055.84 1420.88 3059.1 ;
     RECT  1442.8 3055.84 1442.96 3059.1 ;
     RECT  1467.76 3055.84 1467.92 3059.1 ;
     RECT  1534.96 3055.84 1535.12 3059.1 ;
     RECT  1555.12 3055.84 1555.28 3059.1 ;
     RECT  1566.16 3055.42 1566.32 3059.1 ;
     RECT  1581.04 3055.84 1589.84 3059.1 ;
     RECT  1600.72 3055.84 1600.88 3059.1 ;
     RECT  1614.16 3055.84 1622.96 3059.1 ;
     RECT  1632.88 3057.1 1634.48 3059.1 ;
     RECT  1644.88 3055.42 1645.04 3059.1 ;
     RECT  1694.8 3056.26 1700.24 3059.1 ;
     RECT  1754.8 3055.84 1754.96 3059.1 ;
     RECT  1768.72 3055.84 1777.52 3059.1 ;
     RECT  1788.4 3055.84 1788.56 3059.1 ;
     RECT  1810.96 3055.84 1811.12 3059.1 ;
     RECT  1833.52 3055.84 1833.68 3059.1 ;
     RECT  1855.6 3055.84 1855.76 3059.1 ;
     RECT  1878.16 3055.84 1878.32 3059.1 ;
     RECT  1922.8 3057.94 1924.88 3059.1 ;
     RECT  1942.96 3055.42 1943.12 3059.1 ;
     RECT  1979.92 3055 1988.24 3059.1 ;
     RECT  1998.16 3056.68 2013.2 3059.1 ;
     RECT  2025.52 3055.84 3199.68 3059.1 ;
     RECT  3220 2991 3400 3115 ;
     RECT  0 3001 180 3125 ;
     RECT  3220 3115 3470 3185 ;
     RECT  -70 3125 180 3195 ;
     RECT  200.16 3059.1 3199.68 3198.1 ;
     RECT  0 3195 180 3220 ;
     RECT  3220 3185 3400 3220 ;
     RECT  0 3220 3400 3400 ;
     RECT  215 3400 285 3470 ;
     RECT  409 3400 479 3470 ;
     RECT  603 3400 673 3470 ;
     RECT  797 3400 867 3470 ;
     RECT  991 3400 1061 3470 ;
     RECT  1185 3400 1255 3470 ;
     RECT  1379 3400 1449 3470 ;
     RECT  1573 3400 1643 3470 ;
     RECT  1767 3400 1837 3470 ;
     RECT  1961 3400 2031 3470 ;
     RECT  2155 3400 2225 3470 ;
     RECT  2349 3400 2419 3470 ;
     RECT  2543 3400 2613 3470 ;
     RECT  2737 3400 2807 3470 ;
     RECT  2931 3400 3001 3470 ;
     RECT  3125 3400 3195 3470 ;
    LAYER Metal2 ;
     RECT  -70 215 0 285 ;
     RECT  -70 409 0 479 ;
     RECT  -70 603 0 673 ;
     RECT  -70 797 0 867 ;
     RECT  -70 991 0 1061 ;
     RECT  -70 1185 0 1255 ;
     RECT  -70 1379 0 1449 ;
     RECT  -70 1573 0 1643 ;
     RECT  -70 1767 0 1837 ;
     RECT  -70 1961 0 2031 ;
     RECT  -70 2155 0 2225 ;
     RECT  -70 2349 0 2419 ;
     RECT  -70 2543 0 2613 ;
     RECT  -70 2737 0 2807 ;
     RECT  -70 2931 0 3001 ;
     RECT  -70 3125 0 3195 ;
     RECT  0 0 180 3400 ;
     RECT  180 2448.08 190.46 2448.28 ;
     RECT  180 2843.72 191.14 2843.92 ;
     RECT  190.46 2448.08 191.62 2451.64 ;
     RECT  191.42 2387.6 200.905 2387.8 ;
     RECT  190.94 2773.16 200.905 2773.36 ;
     RECT  200.905 2387.585 201.4 2387.815 ;
     RECT  200.905 2773.145 201.4 2773.375 ;
     RECT  201.4 2386.75 203.9 2387.815 ;
     RECT  201.4 2772.31 203.9 2773.375 ;
     RECT  180 0 205 180 ;
     RECT  203.9 2384.24 208.355 2387.815 ;
     RECT  203.9 2769.8 208.355 2773.375 ;
     RECT  208.355 2384.24 208.805 2386.98 ;
     RECT  208.355 2769.8 208.805 2772.54 ;
     RECT  208.805 2384.24 209.38 2386.96 ;
     RECT  208.805 2769.8 209.38 2770 ;
     RECT  180 3220 215 3400 ;
     RECT  229.34 1745 230.3 1745.2 ;
     RECT  230.3 1744.58 230.78 1745.2 ;
     RECT  230.78 1741.64 231.26 1745.2 ;
     RECT  231.26 1736.6 233.18 1745.2 ;
     RECT  233.18 1735.34 237.98 1745.2 ;
     RECT  237.98 1735.34 243.94 1748.98 ;
     RECT  243.94 1735.34 251.075 1745.215 ;
     RECT  251.075 1735.34 265.06 1744.78 ;
     RECT  205 -70 275 180 ;
     RECT  215 3220 285 3470 ;
     RECT  265.06 1737.44 288.1 1744.78 ;
     RECT  275 0 399 180 ;
     RECT  285 3220 409 3400 ;
     RECT  425.66 2172.14 426.56 2172.34 ;
     RECT  426.56 2171.13 427.58 2172.34 ;
     RECT  180 2577.86 428.26 2578.06 ;
     RECT  429.5 2189.78 430.4 2189.98 ;
     RECT  427.58 2167.1 432.38 2179.9 ;
     RECT  430.4 2189.78 432.38 2190.99 ;
     RECT  432.38 2167.1 438.14 2190.99 ;
     RECT  438.14 2167.1 438.34 2195.02 ;
     RECT  438.34 2167.52 440.54 2195.02 ;
     RECT  440.54 2167.52 441.44 2201.74 ;
     RECT  440.54 2212.04 442.4 2216.86 ;
     RECT  441.44 2167.52 442.46 2201.775 ;
     RECT  442.4 2212.04 443.42 2216.895 ;
     RECT  442.46 2167.52 446.3 2202.16 ;
     RECT  443.42 2212.04 446.3 2217.28 ;
     RECT  446.3 2167.52 448.22 2217.28 ;
     RECT  448.22 2165 450.14 2217.28 ;
     RECT  450.14 2165 450.62 2221.06 ;
     RECT  450.62 2160.38 451.3 2221.9 ;
     RECT  451.3 2165 453.445 2221.9 ;
     RECT  453.445 2165 454.46 2225.26 ;
     RECT  454.46 2165 455.14 2225.68 ;
     RECT  180 635.78 459.94 635.98 ;
     RECT  455.14 2166.68 466.46 2225.68 ;
     RECT  399 -70 469 180 ;
     RECT  466.46 2164.16 470.3 2225.68 ;
     RECT  470.3 2164.16 471.26 2228.2 ;
     RECT  471.26 2164.16 472.22 2229.88 ;
     RECT  472.22 2164.16 472.7 2232.4 ;
     RECT  472.7 2164.16 475.1 2234.08 ;
     RECT  475.1 2157.44 475.3 2239.96 ;
     RECT  475.3 2157.44 478.9 2157.64 ;
     RECT  409 3220 479 3470 ;
     RECT  475.3 2167.1 481.85 2239.96 ;
     RECT  481.85 2167.1 481.92 2240.3 ;
     RECT  201.5 1033.1 482.02 1033.3 ;
     RECT  479.675 2156.6 488.06 2156.8 ;
     RECT  481.92 2167.1 488.06 2240.38 ;
     RECT  488.06 2156.6 489.5 2240.38 ;
     RECT  489.5 2156.6 495.74 2243.74 ;
     RECT  495.74 2156.6 496.7 2248.36 ;
     RECT  496.7 2156.6 501.02 2251.3 ;
     RECT  501.02 2156.6 501.5 2255.5 ;
     RECT  501.5 2156.6 502.4 2258.02 ;
     RECT  502.4 2156.6 503.9 2259.03 ;
     RECT  503.42 2270 503.9 2270.2 ;
     RECT  503.9 2156.6 505.34 2270.2 ;
     RECT  504.38 2117.96 506.24 2121.94 ;
     RECT  506.78 2136.86 507.26 2137.06 ;
     RECT  507.26 2133.08 507.68 2137.06 ;
     RECT  505.34 2156.6 508.22 2278.18 ;
     RECT  507.68 2133.08 509.18 2138.07 ;
     RECT  509.18 2133.08 510.025 2144.62 ;
     RECT  508.22 2156.6 510.025 2285.74 ;
     RECT  510.025 2133.065 510.08 2144.62 ;
     RECT  506.24 2117.96 511.1 2122.95 ;
     RECT  510.08 2133.065 511.1 2145.63 ;
     RECT  510.025 2156.6 511.58 2289.535 ;
     RECT  511.58 2156.6 512.3 2296.24 ;
     RECT  512.3 2156.6 512.54 2297.5 ;
     RECT  511.1 2117.96 513.02 2145.63 ;
     RECT  512.54 2156.6 513.02 2300.02 ;
     RECT  513.02 2117.96 515.36 2300.02 ;
     RECT  515.36 2117.96 516.38 2300.055 ;
     RECT  516.38 2117.96 517.54 2300.44 ;
     RECT  517.54 2165 518.02 2300.44 ;
     RECT  518.02 2167.94 518.78 2300.44 ;
     RECT  517.54 2117.96 519.26 2149.24 ;
     RECT  519.26 2111.66 519.74 2149.24 ;
     RECT  519.74 2108.3 520.9 2149.24 ;
     RECT  521.66 2099.06 522.14 2099.26 ;
     RECT  520.9 2108.3 522.14 2145.88 ;
     RECT  521.66 2088.98 522.56 2089.18 ;
     RECT  522.56 2087.97 522.62 2089.18 ;
     RECT  522.14 2099.06 522.62 2145.88 ;
     RECT  518.78 2167.94 524.06 2306.74 ;
     RECT  524.06 2167.94 524.245 2308 ;
     RECT  524.245 2171.3 525.7 2308 ;
     RECT  522.62 2087.97 526.18 2145.88 ;
     RECT  525.7 2178.02 528.1 2308 ;
     RECT  528.1 2178.02 530.98 2306.74 ;
     RECT  526.18 2087.97 531.26 2143.78 ;
     RECT  530.98 2178.44 532.66 2306.74 ;
     RECT  531.26 2087.72 536.06 2143.78 ;
     RECT  536.06 2084.78 536.96 2143.78 ;
     RECT  532.66 2178.44 537.7 2305.06 ;
     RECT  537.7 2181.8 538.18 2305.06 ;
     RECT  538.18 2183.06 539.14 2305.06 ;
     RECT  536.96 2084.745 541.26 2143.78 ;
     RECT  544.14 2318.72 544.22 2318.92 ;
     RECT  539.14 2186.42 544.7 2305.06 ;
     RECT  541.26 2084.745 545.18 2149.66 ;
     RECT  545.18 2081.42 546.08 2149.66 ;
     RECT  544.22 2318.72 547.1 2319.76 ;
     RECT  547.1 2318.72 548 2330.26 ;
     RECT  544.7 2186.42 548.54 2308.84 ;
     RECT  548 2318.72 548.54 2330.295 ;
     RECT  548.54 2186.42 549.02 2330.295 ;
     RECT  546.08 2080.41 552.3 2149.66 ;
     RECT  549.02 2186.42 553.34 2330.68 ;
     RECT  552.38 2341.82 553.34 2342.02 ;
     RECT  552.3 2076.38 554.5 2149.66 ;
     RECT  553.34 2186.42 562.18 2342.02 ;
     RECT  558.14 2175.5 562.46 2175.7 ;
     RECT  562.18 2186.42 562.46 2248.36 ;
     RECT  562.18 2257.82 563.36 2342.02 ;
     RECT  554.5 2076.46 563.82 2149.66 ;
     RECT  563.82 2073.86 564.595 2149.66 ;
     RECT  562.46 2175.5 566.02 2248.36 ;
     RECT  562.46 2050.34 568.22 2050.54 ;
     RECT  566.02 2175.5 568.22 2240.38 ;
     RECT  568.22 2046.98 569.18 2050.54 ;
     RECT  569.18 2046.98 570.14 2051.38 ;
     RECT  563.36 2257.82 570.62 2342.19 ;
     RECT  564.595 2073.02 572.54 2149.66 ;
     RECT  568.22 2172.56 572.54 2240.38 ;
     RECT  571.58 2000.78 573.385 2001.4 ;
     RECT  570.62 2257.82 573.98 2342.86 ;
     RECT  570.14 2046.98 574.18 2053.48 ;
     RECT  572.54 2073.02 575.42 2240.38 ;
     RECT  573.385 2000.78 576.1 2002.255 ;
     RECT  575.42 2073.02 577.82 2245.42 ;
     RECT  573.98 2257.82 577.82 2343.28 ;
     RECT  574.18 2050.34 578.02 2050.54 ;
     RECT  577.82 2073.02 578.5 2352.94 ;
     RECT  578.5 2167.52 578.72 2352.94 ;
     RECT  578.72 2167.52 579.01 2352.975 ;
     RECT  576.1 2001.19 580.835 2002.255 ;
     RECT  580.835 2001.19 581.285 2001.42 ;
     RECT  578.5 2073.02 586.46 2157.64 ;
     RECT  586.46 2071.76 587.9 2157.64 ;
     RECT  579.01 2167.52 588.38 2352.94 ;
     RECT  587.9 2070.08 590.18 2157.64 ;
     RECT  588.38 2167.1 590.18 2352.94 ;
     RECT  581.285 2001.2 590.3 2001.4 ;
     RECT  590.3 2000.78 590.5 2001.4 ;
     RECT  590.18 2070.08 592.22 2352.94 ;
     RECT  469 0 593 180 ;
     RECT  592.22 2070.08 593.18 2353.36 ;
     RECT  593.18 2070.08 594.62 2356.72 ;
     RECT  594.62 2070.08 595.04 2359.66 ;
     RECT  581.66 2368.7 595.04 2368.9 ;
     RECT  595.04 2070.08 596.06 2368.9 ;
     RECT  479 3220 603 3400 ;
     RECT  596.06 2068.4 604.155 2368.9 ;
     RECT  604.155 2068.9 604.24 2368.9 ;
     RECT  604.24 2069.395 604.9 2368.9 ;
     RECT  604.9 2069.395 605.38 2124.04 ;
     RECT  593 -70 606.38 180 ;
     RECT  606.38 -70 606.82 180.7 ;
     RECT  605.38 2069.395 607.05 2122.95 ;
     RECT  191.62 2451.44 609.22 2451.64 ;
     RECT  607.05 2069.66 618.14 2122.95 ;
     RECT  604.9 2132.66 618.62 2368.9 ;
     RECT  618.14 2069.24 619.1 2122.95 ;
     RECT  618.62 2132.66 619.1 2371.42 ;
     RECT  619.1 2069.24 619.3 2372.68 ;
     RECT  619.3 2069.24 622.18 2371.84 ;
     RECT  586.94 1983.98 622.46 1984.18 ;
     RECT  622.18 2069.24 622.66 2074.48 ;
     RECT  622.18 2084.36 623.62 2371.84 ;
     RECT  623.62 2084.78 624.085 2371.84 ;
     RECT  622.66 2071.76 624.1 2074.48 ;
     RECT  624.085 2085.62 626.5 2371.84 ;
     RECT  626.3 1934.42 626.98 1935.46 ;
     RECT  626.5 2085.62 627.46 2168.31 ;
     RECT  627.46 2085.62 628.9 2108.5 ;
     RECT  624.1 2071.76 629.86 2071.96 ;
     RECT  628.9 2088.98 630.09 2108.5 ;
     RECT  630.09 2108.3 630.34 2108.5 ;
     RECT  626.5 2178.02 630.62 2371.84 ;
     RECT  630.62 2178.02 633.5 2375.62 ;
     RECT  630.09 2088.98 633.7 2099.68 ;
     RECT  627.46 2118.38 635.42 2168.31 ;
     RECT  633.5 2178.02 635.42 2376.04 ;
     RECT  635.42 2118.38 635.9 2376.04 ;
     RECT  428.06 2012.12 636.86 2012.32 ;
     RECT  635.9 2118.38 637.28 2378.56 ;
     RECT  637.28 2118.38 638.665 2379.99 ;
     RECT  637.34 2512.76 638.665 2512.96 ;
     RECT  638.665 2115.425 639.16 2379.99 ;
     RECT  639.16 2114.59 640.22 2379.99 ;
     RECT  640.22 2114.59 640.42 2382.76 ;
     RECT  629.66 1974.32 640.7 1974.52 ;
     RECT  288.1 1737.44 640.9 1744.36 ;
     RECT  640.7 1973.48 640.9 1974.52 ;
     RECT  640.42 2114.59 644.725 2379.99 ;
     RECT  638.665 2512.76 646.115 2516.335 ;
     RECT  644.725 2114.59 646.565 2378.98 ;
     RECT  646.115 2512.76 646.565 2515.5 ;
     RECT  606.82 -70 647.9 180 ;
     RECT  646.565 2512.76 649.06 2512.96 ;
     RECT  590.5 2000.78 649.225 2000.98 ;
     RECT  647.9 -70 654.82 180.7 ;
     RECT  646.565 2114.6 656.165 2378.98 ;
     RECT  649.225 2000.78 656.675 2002.255 ;
     RECT  656.165 2114.6 656.74 2122.36 ;
     RECT  656.675 2000.78 657.7 2002.24 ;
     RECT  656.165 2131.4 659.14 2378.98 ;
     RECT  659.14 2261.18 660.1 2378.98 ;
     RECT  660.1 2292.09 660.38 2378.98 ;
     RECT  660.38 2292.09 661.34 2379.82 ;
     RECT  626.98 1935.26 662.78 1935.46 ;
     RECT  654.82 -70 663 180 ;
     RECT  661.34 2292.09 663.66 2380.24 ;
     RECT  656.74 2120.9 664.62 2122.36 ;
     RECT  659.14 2131.4 664.62 2251.72 ;
     RECT  664.62 2120.9 669.385 2251.72 ;
     RECT  660.1 2261.18 669.385 2282.38 ;
     RECT  640.9 1973.48 669.5 1973.68 ;
     RECT  622.46 1983.14 669.5 1984.18 ;
     RECT  669.385 2120.9 669.5 2282.38 ;
     RECT  663.66 2292.09 669.5 2383.6 ;
     RECT  669.5 2120.9 670.01 2383.6 ;
     RECT  670.01 2120.9 670.08 2383.94 ;
     RECT  603 3220 673 3470 ;
     RECT  669.5 1973.48 675.74 1984.18 ;
     RECT  670.08 2120.9 677.66 2384.02 ;
     RECT  677.66 2116.28 679.78 2384.02 ;
     RECT  675.26 1905.86 680.06 1906.06 ;
     RECT  633.7 2088.98 680.06 2092.12 ;
     RECT  679.78 2220.02 680.26 2384.02 ;
     RECT  679.58 1894.1 681.98 1894.3 ;
     RECT  662.78 1935.26 682.46 1938.4 ;
     RECT  681.98 1894.1 682.94 1896.4 ;
     RECT  680.06 1905.86 682.94 1911.52 ;
     RECT  680.06 2088.98 683.305 2096.32 ;
     RECT  679.78 2116.28 684.81 2210.06 ;
     RECT  684.81 2116.28 688.42 2189.56 ;
     RECT  684.81 2198.18 688.9 2210.06 ;
     RECT  688.9 2201.12 689.66 2210.06 ;
     RECT  680.26 2220.02 689.66 2383.6 ;
     RECT  675.74 1966.34 690.62 1984.18 ;
     RECT  636.86 2012.12 690.62 2012.74 ;
     RECT  689.66 2201.12 690.62 2383.6 ;
     RECT  690.62 2201.12 691.1 2411.74 ;
     RECT  690.62 2012.12 691.58 2019.46 ;
     RECT  691.1 2201.12 691.58 2416.36 ;
     RECT  690.62 1966.34 692.06 1990.06 ;
     RECT  691.58 2201.12 692.06 2422.24 ;
     RECT  692.06 2201.12 692.54 2423.92 ;
     RECT  682.46 1935.26 692.905 1944.28 ;
     RECT  675.26 2437.58 693.02 2437.78 ;
     RECT  678.62 1925.18 693.4 1925.38 ;
     RECT  692.905 1933.985 693.4 1944.28 ;
     RECT  693.02 2437.16 693.5 2437.78 ;
     RECT  691.58 2012.12 693.98 2023.66 ;
     RECT  683.305 2087.705 693.98 2096.32 ;
     RECT  688.42 2116.28 693.98 2187.88 ;
     RECT  692.06 2466.98 693.98 2467.18 ;
     RECT  683.42 2487.14 693.98 2487.34 ;
     RECT  692.06 2497.22 693.98 2497.84 ;
     RECT  692.06 1966.34 694.94 1990.48 ;
     RECT  693.4 1925.18 696.38 1944.28 ;
     RECT  640.9 1737.44 696.745 1743.94 ;
     RECT  693.5 2437.16 696.86 2441.14 ;
     RECT  693.98 2459.84 696.86 2467.18 ;
     RECT  694.94 1966.34 697.34 1991.32 ;
     RECT  693.98 2075.96 698.3 2187.88 ;
     RECT  692.54 2201.12 698.3 2426.44 ;
     RECT  696.86 2435.48 698.3 2441.14 ;
     RECT  693.98 2482.52 698.3 2507.08 ;
     RECT  675.74 2522.42 698.3 2522.62 ;
     RECT  676.22 2534.6 698.3 2534.8 ;
     RECT  662.78 2560.22 698.3 2560.42 ;
     RECT  693.98 2012.12 698.5 2030.8 ;
     RECT  698.5 2030.56 698.78 2030.8 ;
     RECT  693.98 2059.16 698.78 2059.36 ;
     RECT  682.94 1894.1 699.26 1911.52 ;
     RECT  696.38 1922.66 699.26 1944.28 ;
     RECT  672.86 1955 699.26 1955.2 ;
     RECT  697.34 1963.82 699.26 1991.32 ;
     RECT  698.3 2073.4 699.26 2187.88 ;
     RECT  699.26 1894.1 699.74 1944.28 ;
     RECT  699.26 1955 699.74 1991.32 ;
     RECT  698.78 2057.48 699.74 2059.36 ;
     RECT  699.26 2070.88 699.74 2187.88 ;
     RECT  699.74 2046.14 699.98 2046.34 ;
     RECT  699.74 2057.48 699.98 2192.5 ;
     RECT  698.3 2201.12 699.98 2426.86 ;
     RECT  698.3 2435.48 699.98 2448.28 ;
     RECT  696.86 2458.16 699.98 2467.18 ;
     RECT  698.3 2482.52 699.98 2537.74 ;
     RECT  698.3 2553.5 699.98 2573.02 ;
     RECT  698.78 2030.56 700 2035.8 ;
     RECT  699.98 2046.14 700 2469.14 ;
     RECT  699.98 2481.74 700 2539.7 ;
     RECT  699.98 2552.3 700 2574.98 ;
     RECT  700 2030.56 700.72 2580.12 ;
     RECT  700.72 2569.84 700.9 2578.06 ;
     RECT  700.72 2030.6 701.06 2529.72 ;
     RECT  699.74 1894.1 701.18 1991.32 ;
     RECT  657.7 2001.2 701.18 2001.4 ;
     RECT  700.9 2569.84 701.38 2570.04 ;
     RECT  700.72 2542.12 702.34 2542.32 ;
     RECT  699.74 1824.38 703.1 1824.58 ;
     RECT  701.06 2030.6 703.46 2527.2 ;
     RECT  701.18 1894.1 704.06 2001.4 ;
     RECT  696.745 1737.44 704.195 1745.215 ;
     RECT  703.46 2086 704.42 2255.04 ;
     RECT  703.46 2264.92 704.42 2527.2 ;
     RECT  704.195 1737.44 704.645 1744.38 ;
     RECT  704.06 1889.9 705.5 2001.4 ;
     RECT  700.72 2552.66 705.7 2552.86 ;
     RECT  704.645 1737.44 705.865 1744.36 ;
     RECT  704.42 2391.76 706.34 2527.2 ;
     RECT  705.865 1729.865 706.36 1744.36 ;
     RECT  704.42 2264.92 706.82 2381.04 ;
     RECT  706.34 2416.12 706.82 2527.2 ;
     RECT  703.46 2030.6 707.14 2066.5 ;
     RECT  704.42 2086 707.3 2224.8 ;
     RECT  704.42 2234.68 707.3 2255.04 ;
     RECT  706.82 2264.92 707.3 2282.76 ;
     RECT  706.82 2291.38 707.3 2381.04 ;
     RECT  706.34 2391.76 707.3 2406.24 ;
     RECT  703.1 1817.66 707.42 1824.58 ;
     RECT  694.94 1854.62 708.38 1854.82 ;
     RECT  705.5 1884.86 709.82 2001.4 ;
     RECT  708.38 1854.62 710.3 1856.08 ;
     RECT  706.94 1869.74 710.3 1869.94 ;
     RECT  707.3 2088.52 710.66 2108.88 ;
     RECT  706.82 2421.16 710.66 2527.2 ;
     RECT  710.66 2094.4 711.14 2108.88 ;
     RECT  709.82 1882.76 711.46 2001.4 ;
     RECT  707.3 2234.68 711.62 2247.48 ;
     RECT  711.46 1882.76 711.94 1991.32 ;
     RECT  707.3 2141.44 712.1 2146.68 ;
     RECT  706.36 1729.03 712.7 1744.36 ;
     RECT  712.7 1728.62 712.9 1744.36 ;
     RECT  707.3 2277.52 713.06 2280.24 ;
     RECT  712.9 1728.62 713.315 1730.095 ;
     RECT  713.315 1728.62 714.34 1730.08 ;
     RECT  711.14 2094.4 714.5 2106.36 ;
     RECT  707.3 2291.38 717.66 2345.34 ;
     RECT  707.3 2354.38 717.66 2381.04 ;
     RECT  714.5 2094.82 717.86 2106.36 ;
     RECT  710.66 2421.16 717.86 2479.32 ;
     RECT  707.3 2174.2 719.58 2192.04 ;
     RECT  707.3 2204.02 719.58 2204.64 ;
     RECT  707.3 2216.62 719.58 2224.8 ;
     RECT  707.14 2033.08 720.1 2066.5 ;
     RECT  717.86 2421.16 720.26 2476.8 ;
     RECT  719.58 2163.7 720.74 2195.4 ;
     RECT  711.62 2234.68 720.905 2244.96 ;
     RECT  713.06 2280.04 720.905 2280.24 ;
     RECT  717.66 2291.38 721.22 2381.04 ;
     RECT  707.3 2121.28 721.385 2129.04 ;
     RECT  720.905 2261.965 721.4 2262.195 ;
     RECT  712.1 2146.06 721.98 2146.68 ;
     RECT  720.74 2163.7 721.98 2194.98 ;
     RECT  719.58 2204.02 721.98 2224.8 ;
     RECT  720.905 2234.68 721.98 2252.115 ;
     RECT  721.385 2121.28 722.46 2131.155 ;
     RECT  721.98 2141.44 722.46 2146.68 ;
     RECT  717.86 2106.16 722.94 2106.36 ;
     RECT  722.46 2119.6 722.94 2131.155 ;
     RECT  722.46 2141.44 722.94 2150.88 ;
     RECT  721.98 2159.92 722.94 2194.98 ;
     RECT  720.26 2466.52 723.14 2476.8 ;
     RECT  721.98 2204.02 723.42 2252.115 ;
     RECT  721.4 2261.965 723.42 2263.03 ;
     RECT  707.3 2391.76 723.62 2401.2 ;
     RECT  720.905 2280.04 724.38 2282.355 ;
     RECT  721.22 2291.38 724.38 2377.68 ;
     RECT  723.42 2204.02 724.86 2263.03 ;
     RECT  724.38 2278.36 724.86 2377.68 ;
     RECT  717.86 2094.82 725.705 2095.44 ;
     RECT  723.14 2469.04 726.02 2476.8 ;
     RECT  720.26 2421.16 727.94 2456.64 ;
     RECT  722.94 2106.16 729.18 2194.98 ;
     RECT  724.86 2204.02 729.18 2377.68 ;
     RECT  726.02 2469.04 729.86 2472.18 ;
     RECT  729.18 2106.16 733.5 2377.68 ;
     RECT  725.705 2088.085 733.98 2095.44 ;
     RECT  733.5 2105.32 733.98 2377.68 ;
     RECT  733.865 2072.965 734.36 2073.195 ;
     RECT  727.94 2426.2 735.62 2456.64 ;
     RECT  720.1 2033.08 735.9 2063.52 ;
     RECT  733.98 2088.085 737.34 2377.68 ;
     RECT  734.36 2072.965 737.82 2074.03 ;
     RECT  737.82 2072.965 738.3 2076.54 ;
     RECT  737.34 2085.16 738.3 2377.68 ;
     RECT  735.9 2033.08 739.145 2063.94 ;
     RECT  738.3 2072.965 739.145 2377.68 ;
     RECT  714.34 1729.88 741.5 1730.08 ;
     RECT  701.66 1798.34 741.5 1798.54 ;
     RECT  707.42 1817.66 741.5 1832.56 ;
     RECT  710.3 1854.62 741.5 1869.94 ;
     RECT  739.145 2033.08 741.66 2377.68 ;
     RECT  741.5 1729.88 741.7 1731.34 ;
     RECT  741.5 1798.34 741.7 1799.8 ;
     RECT  741.5 1854.62 741.7 1870.36 ;
     RECT  711.94 1882.76 741.7 1990.48 ;
     RECT  741.7 1882.76 752.425 1988.8 ;
     RECT  752.425 1882.76 752.92 1989.655 ;
     RECT  752.92 1882.76 762.62 1990.49 ;
     RECT  711.46 2001.2 762.82 2001.4 ;
     RECT  741.5 1817.66 768.86 1832.98 ;
     RECT  712.9 1743.74 769.06 1743.94 ;
     RECT  741.7 1799.6 783.74 1799.8 ;
     RECT  768.86 1811.78 783.74 1832.98 ;
     RECT  663 0 787 180 ;
     RECT  741.66 2033.08 791.1 2378.1 ;
     RECT  795.26 1706.36 796.22 1710.76 ;
     RECT  673 3220 797 3400 ;
     RECT  796.22 1703.42 797.12 1710.76 ;
     RECT  180 1681.16 797.66 1681.36 ;
     RECT  797.12 1702.41 798.14 1710.76 ;
     RECT  798.14 1702.41 799.04 1717.9 ;
     RECT  799.04 1702.41 799.1 1717.935 ;
     RECT  783.74 1799.6 799.1 1832.98 ;
     RECT  797.66 1681.16 799.58 1688.5 ;
     RECT  799.1 1702.41 799.58 1721.68 ;
     RECT  799.1 1792.88 800.54 1832.98 ;
     RECT  799.1 1665.62 800.96 1669.6 ;
     RECT  800.54 1649.24 801.02 1653.22 ;
     RECT  799.58 1681.16 801.98 1721.68 ;
     RECT  741.7 1731.14 801.98 1731.34 ;
     RECT  801.02 1642.94 802.4 1653.22 ;
     RECT  735.62 2436.28 802.82 2456.64 ;
     RECT  802.4 1642.94 802.88 1654.23 ;
     RECT  802.88 1641.93 802.94 1654.23 ;
     RECT  802.46 1769.78 803.36 1770.82 ;
     RECT  787 -70 803.42 180 ;
     RECT  741.7 1855.04 803.42 1870.36 ;
     RECT  802.94 1635.38 803.84 1654.23 ;
     RECT  800.54 1549.28 803.9 1549.48 ;
     RECT  803.84 1634.37 803.9 1654.23 ;
     RECT  800.96 1664.61 803.9 1669.6 ;
     RECT  801.98 1681.16 803.9 1733.86 ;
     RECT  803.36 1769.78 803.9 1770.855 ;
     RECT  800.54 1787.42 803.9 1832.98 ;
     RECT  803.42 -70 804.1 180.7 ;
     RECT  803.42 1847.06 804.32 1870.36 ;
     RECT  710.66 2489.2 805.22 2527.2 ;
     RECT  803.9 1769.78 805.34 1832.98 ;
     RECT  805.34 1766.84 806.3 1832.98 ;
     RECT  804.32 1846.05 806.3 1870.36 ;
     RECT  803.9 1634.37 806.78 1733.86 ;
     RECT  791.1 2033.08 807.14 2378.52 ;
     RECT  807.74 1619.42 808.22 1619.62 ;
     RECT  808.22 1618.58 808.64 1619.62 ;
     RECT  808.64 1618.58 808.7 1619.655 ;
     RECT  808.22 1755.5 808.7 1755.7 ;
     RECT  806.3 1766.84 808.7 1870.36 ;
     RECT  808.7 1748.78 809.12 1755.7 ;
     RECT  808.7 1615.64 809.18 1619.655 ;
     RECT  809.12 1748.78 809.6 1755.735 ;
     RECT  809.18 1615.22 809.66 1619.655 ;
     RECT  809.6 1747.77 810.14 1755.735 ;
     RECT  810.14 1747.77 810.62 1756.12 ;
     RECT  809.66 1615.22 811.1 1620.04 ;
     RECT  806.78 1630.34 811.1 1733.86 ;
     RECT  810.62 1743.74 811.1 1756.12 ;
     RECT  811.1 1615.22 813.5 1756.12 ;
     RECT  808.7 1766.42 813.5 1870.36 ;
     RECT  807.14 2035.6 814.14 2378.52 ;
     RECT  723.62 2391.76 815.1 2394.06 ;
     RECT  813.5 1615.22 815.9 1870.36 ;
     RECT  814.14 2035.6 817.5 2379.78 ;
     RECT  817.5 2035.6 818.46 2380.62 ;
     RECT  815.9 1612.7 819.26 1870.36 ;
     RECT  819.26 1610.6 820.7 1870.36 ;
     RECT  762.62 1882.76 820.7 1990.9 ;
     RECT  820.7 1610.6 822.14 1871.2 ;
     RECT  820.7 1879.82 822.14 1990.9 ;
     RECT  822.14 1610.6 823.04 1990.9 ;
     RECT  823.04 1608.465 824.06 1990.9 ;
     RECT  818.46 2035.6 824.7 2381.04 ;
     RECT  815.1 2390.5 824.7 2394.06 ;
     RECT  805.22 2489.2 828.26 2524.68 ;
     RECT  797 3220 830.3 3470 ;
     RECT  824.7 2035.6 833.54 2394.06 ;
     RECT  824.06 1608.08 834.62 1990.9 ;
     RECT  833.54 2054.5 839.3 2394.06 ;
     RECT  609.5 1499.3 842.3 1499.5 ;
     RECT  842.3 1499.3 842.5 1499.92 ;
     RECT  839.3 2054.92 842.645 2394.06 ;
     RECT  828.26 2496.76 842.66 2524.68 ;
     RECT  842.66 2516.92 845.54 2524.68 ;
     RECT  842.645 2055.76 846.02 2394.06 ;
     RECT  834.62 1605.56 851.42 1990.9 ;
     RECT  851.42 1604.72 852.86 1990.9 ;
     RECT  729.86 2469.04 854.66 2469.24 ;
     RECT  804.1 -70 857 180 ;
     RECT  833.54 2035.6 858.02 2043.36 ;
     RECT  842.66 2496.76 858.02 2507.04 ;
     RECT  846.02 2056.18 859.69 2394.06 ;
     RECT  859.69 2056.18 865.5 2381.04 ;
     RECT  858.02 2038.12 866.94 2043.36 ;
     RECT  865.5 2051.98 866.94 2381.04 ;
     RECT  830.3 3219.2 867 3470 ;
     RECT  858.02 2496.76 870.98 2496.96 ;
     RECT  866.94 2038.12 873.66 2381.04 ;
     RECT  859.69 2390.5 873.66 2394.06 ;
     RECT  852.86 1600.1 879.74 1990.9 ;
     RECT  803.9 1549.28 883.58 1550.32 ;
     RECT  883.58 1547.18 889.54 1550.32 ;
     RECT  879.74 1597.16 891.74 1990.9 ;
     RECT  889.54 1547.59 893.285 1550.32 ;
     RECT  873.66 2038.12 894.5 2394.06 ;
     RECT  894.5 2038.12 899.78 2043.36 ;
     RECT  891.74 1596.74 901.54 1990.9 ;
     RECT  893.285 1547.6 905.18 1550.32 ;
     RECT  802.82 2441.32 905.54 2456.64 ;
     RECT  903.74 1521.98 905.6 1525.96 ;
     RECT  905.6 1520.97 905.66 1525.96 ;
     RECT  905.18 1537.1 905.66 1537.3 ;
     RECT  905.18 1467.38 906.08 1468.42 ;
     RECT  905.18 1546.76 906.62 1550.32 ;
     RECT  899.9 1566.5 906.62 1566.7 ;
     RECT  906.08 1467.38 907.1 1468.455 ;
     RECT  906.62 1546.76 907.1 1566.7 ;
     RECT  906.62 1509.38 907.52 1509.58 ;
     RECT  907.1 1477.46 907.58 1479.34 ;
     RECT  907.1 1546.34 907.82 1566.7 ;
     RECT  907.58 1477.46 908.48 1486.9 ;
     RECT  842.5 1499.72 908.54 1499.92 ;
     RECT  907.52 1509.38 908.54 1510.59 ;
     RECT  905.66 1520.97 909.02 1537.3 ;
     RECT  907.82 1546.34 909.02 1567.54 ;
     RECT  901.54 1596.74 909.02 1989.64 ;
     RECT  908.48 1477.46 909.5 1487.91 ;
     RECT  908.54 1499.72 909.5 1510.59 ;
     RECT  909.02 1520.97 909.5 1567.54 ;
     RECT  907.1 1467.38 910.46 1468.84 ;
     RECT  909.5 1477.46 910.46 1567.54 ;
     RECT  910.46 1464.44 910.94 1567.54 ;
     RECT  909.02 1596.32 911.62 1989.64 ;
     RECT  910.94 1456.46 912.38 1567.54 ;
     RECT  906.025 1581.185 913.475 1586.455 ;
     RECT  911.62 1597.16 913.54 1989.64 ;
     RECT  913.475 1581.185 913.925 1585.62 ;
     RECT  913.925 1581.185 914.5 1585.6 ;
     RECT  913.54 1598 914.5 1989.64 ;
     RECT  914.5 1598.42 914.98 1989.64 ;
     RECT  912.38 1448.9 915.26 1567.54 ;
     RECT  894.5 2051.98 915.295 2394.06 ;
     RECT  915.295 2051.14 916.86 2394.06 ;
     RECT  916.86 2050.72 918.02 2394.06 ;
     RECT  918.02 2050.72 918.72 2388.6 ;
     RECT  915.26 1441.76 919.58 1567.54 ;
     RECT  917.18 1577.42 919.58 1578.63 ;
     RECT  899.78 2038.12 920.42 2038.32 ;
     RECT  905.54 2443.84 920.42 2456.64 ;
     RECT  918.72 2050.55 920.585 2388.6 ;
     RECT  920.585 2047.765 921.08 2388.6 ;
     RECT  919.58 1441.76 923.42 1578.63 ;
     RECT  921.08 2046.93 923.58 2388.6 ;
     RECT  735.62 2426.2 923.78 2426.4 ;
     RECT  914.98 1600.52 923.9 1989.64 ;
     RECT  923.9 1596.74 924.38 1989.64 ;
     RECT  923.42 1441.76 924.86 1582.24 ;
     RECT  924.38 1595.9 924.86 1989.64 ;
     RECT  923.58 2043.58 925.22 2388.6 ;
     RECT  925.22 2046.52 927.42 2388.6 ;
     RECT  927.42 2046.52 928.82 2390.28 ;
     RECT  928.82 2046.52 929.34 2391.33 ;
     RECT  928.7 1414.46 929.6 1415.5 ;
     RECT  929.34 2046.52 929.82 2391.54 ;
     RECT  929.6 1414.46 930.62 1415.535 ;
     RECT  930.14 1427.48 930.62 1430.62 ;
     RECT  930.62 1414.46 932 1430.62 ;
     RECT  698.5 2012.12 932.26 2019.46 ;
     RECT  932 1414.46 932.54 1430.655 ;
     RECT  934.46 1388.84 935.9 1389.46 ;
     RECT  932.54 1414.46 935.9 1431.04 ;
     RECT  924.86 1441.76 935.9 1989.64 ;
     RECT  935.9 1414.46 936.745 1989.64 ;
     RECT  935.9 1388.84 936.86 1396.18 ;
     RECT  936.745 1412.345 937.24 1989.64 ;
     RECT  936.86 1385.9 937.76 1396.18 ;
     RECT  937.82 1371.2 938.3 1371.4 ;
     RECT  937.24 1411.51 938.78 1989.64 ;
     RECT  938.3 1363.22 939.2 1371.4 ;
     RECT  938.78 1407.74 939.26 1989.64 ;
     RECT  938.78 1346.84 939.74 1350.82 ;
     RECT  939.74 1340.54 940.64 1350.82 ;
     RECT  940.64 1339.53 940.7 1351.83 ;
     RECT  939.2 1362.21 940.7 1371.4 ;
     RECT  937.76 1384.89 940.7 1397.19 ;
     RECT  940.7 1339.53 941.18 1371.4 ;
     RECT  940.7 1327.94 941.6 1328.14 ;
     RECT  940.7 1382.54 941.66 1397.19 ;
     RECT  939.26 1406.9 941.66 1989.64 ;
     RECT  941.6 1327.94 943.1 1329.15 ;
     RECT  941.18 1339.53 943.1 1373.92 ;
     RECT  941.66 1382.54 943.1 1989.64 ;
     RECT  943.1 1325.84 944.54 1329.15 ;
     RECT  943.1 1339.53 944.54 1989.64 ;
     RECT  929.82 2046.52 944.9 2392.38 ;
     RECT  944.54 1325.84 945.5 1989.64 ;
     RECT  845.54 2516.92 948.26 2519.64 ;
     RECT  858.02 2506.84 950.66 2507.04 ;
     RECT  945.5 1325 950.78 1989.64 ;
     RECT  950.78 1323.74 951.68 1989.64 ;
     RECT  951.68 1321.185 952.7 1989.64 ;
     RECT  920.42 2443.84 954.5 2449.08 ;
     RECT  944.9 2046.52 958.34 2391.54 ;
     RECT  958.34 2046.94 961.02 2391.54 ;
     RECT  961.02 2046.94 962.18 2394.48 ;
     RECT  948.26 2516.92 962.66 2517.12 ;
     RECT  962.18 2051.14 963.42 2394.48 ;
     RECT  963.42 2051.14 965.06 2395.74 ;
     RECT  952.7 1320.8 969.02 1989.64 ;
     RECT  965.06 2054.92 971.285 2395.74 ;
     RECT  971.285 2055.76 973.02 2395.74 ;
     RECT  969.02 1319.96 973.34 1989.64 ;
     RECT  973.02 2055.76 973.43 2399.1 ;
     RECT  190.46 761.78 974.3 761.98 ;
     RECT  973.43 2055.76 974.66 2395.74 ;
     RECT  974.66 2058.11 975.125 2395.74 ;
     RECT  975.125 2059.54 978.5 2395.74 ;
     RECT  973.34 1317.44 979.1 1989.64 ;
     RECT  857 0 981 180 ;
     RECT  978.5 2065.67 984.74 2395.74 ;
     RECT  979.1 1317.02 985.76 1989.64 ;
     RECT  984.74 2065.67 986.18 2395.32 ;
     RECT  985.76 1316.85 986.5 1989.64 ;
     RECT  986.18 2065.67 986.645 2394.9 ;
     RECT  986.5 1951.64 986.98 1989.64 ;
     RECT  986.98 1951.64 987.94 1958.98 ;
     RECT  986.645 2065.84 988.1 2394.9 ;
     RECT  988.1 2068.78 989.06 2394.9 ;
     RECT  989.06 2072.14 990.02 2394.9 ;
     RECT  988.7 742.88 990.82 743.08 ;
     RECT  867 3219.2 991 3400 ;
     RECT  990.02 2072.14 993.38 2391.54 ;
     RECT  987.94 1951.64 994.18 1955.62 ;
     RECT  993.38 2077.17 995.685 2391.54 ;
     RECT  994.18 1951.64 996.58 1952.68 ;
     RECT  995.685 2077.18 996.74 2391.54 ;
     RECT  986.5 1316.85 997.76 1940.5 ;
     RECT  974.3 753.38 997.82 761.98 ;
     RECT  992.54 773.54 997.82 773.74 ;
     RECT  992.06 784.46 997.82 784.66 ;
     RECT  991.58 813.02 997.82 813.64 ;
     RECT  987.26 826.46 997.82 826.66 ;
     RECT  978.14 839.06 997.82 839.26 ;
     RECT  993.5 741.62 998.3 741.82 ;
     RECT  997.82 753.38 998.3 793.9 ;
     RECT  997.82 806.3 998.3 813.64 ;
     RECT  981.5 863.84 998.3 864.04 ;
     RECT  986.98 1968.44 998.3 1989.64 ;
     RECT  997.82 826.46 998.78 841.78 ;
     RECT  997.82 928.52 998.78 935.86 ;
     RECT  992.06 960.02 998.78 960.22 ;
     RECT  997.76 1313.625 998.78 1940.5 ;
     RECT  998.3 738.92 999.26 741.82 ;
     RECT  998.3 753.38 999.26 813.64 ;
     RECT  998.78 949.94 999.26 950.14 ;
     RECT  998.78 1313.24 999.46 1940.5 ;
     RECT  999.26 738.92 999.74 813.64 ;
     RECT  998.78 826.46 999.74 847.48 ;
     RECT  998.3 857.36 999.74 864.04 ;
     RECT  998.78 925.4 999.74 935.86 ;
     RECT  999.74 738.92 999.98 816.58 ;
     RECT  999.74 826.46 999.98 871.18 ;
     RECT  973.34 909.62 999.98 909.82 ;
     RECT  999.74 919.7 999.98 935.86 ;
     RECT  999.26 947.42 999.98 950.14 ;
     RECT  998.78 960.02 999.98 976 ;
     RECT  999.98 907.86 1000 935.86 ;
     RECT  999.98 945.66 1000 976 ;
     RECT  1000 907.76 1000.72 981.04 ;
     RECT  1000.72 954.98 1000.9 955.18 ;
     RECT  996.58 1952.06 1000.9 1952.68 ;
     RECT  999.98 738.92 1001.06 871.18 ;
     RECT  1000.72 978.92 1001.38 981.04 ;
     RECT  1001.06 741.02 1001.66 871.18 ;
     RECT  999.46 1313.24 1001.66 1940.08 ;
     RECT  996.74 2077.18 1002.02 2391.12 ;
     RECT  1002.02 2082.22 1002.405 2391.12 ;
     RECT  1002.405 2103.47 1002.485 2391.12 ;
     RECT  1001.66 741.02 1002.5 874.96 ;
     RECT  1002.485 2104.9 1002.965 2391.12 ;
     RECT  1002.5 819.56 1002.98 874.96 ;
     RECT  1001.66 1309.88 1003.3 1940.08 ;
     RECT  1002.5 741.02 1003.46 809.68 ;
     RECT  1002.98 824.6 1003.46 874.96 ;
     RECT  1000.9 1952.48 1003.78 1952.68 ;
     RECT  1000.72 914.24 1004.26 929.14 ;
     RECT  1002.405 2082.22 1005.365 2093.09 ;
     RECT  1001.38 978.92 1005.7 979.12 ;
     RECT  1003.3 1309.88 1005.7 1937.98 ;
     RECT  1003.46 837.2 1006.82 874.96 ;
     RECT  1003.46 761.6 1007.3 809.68 ;
     RECT  1002.965 2104.9 1007.3 2388.6 ;
     RECT  1005.365 2082.22 1007.78 2091.66 ;
     RECT  1007.78 2091.46 1008.74 2091.66 ;
     RECT  1007.3 2104.9 1008.74 2115.18 ;
     RECT  1008.74 2104.9 1009.22 2105.1 ;
     RECT  1008.74 2114.56 1009.22 2114.76 ;
     RECT  1004.26 914.24 1009.54 917.38 ;
     RECT  998.3 1968.44 1010.02 1990.06 ;
     RECT  1007.3 2125.06 1011.42 2388.6 ;
     RECT  1006.82 844.76 1012.42 874.96 ;
     RECT  1004.26 928.94 1013.86 929.14 ;
     RECT  1003.46 824.6 1014.3 824.8 ;
     RECT  1007.3 761.6 1014.5 807.16 ;
     RECT  1014.3 824.6 1014.5 825.22 ;
     RECT  1009.54 914.24 1016.26 914.44 ;
     RECT  1011.42 2125.06 1016.42 2392.38 ;
     RECT  1016.42 2125.06 1020.74 2391.54 ;
     RECT  1020.74 2125.06 1020.98 2390.7 ;
     RECT  1005.7 1309.88 1022.3 1937.56 ;
     RECT  1022.3 1308.62 1027.1 1937.56 ;
     RECT  1020.98 2125.06 1027.94 2388.6 ;
     RECT  1027.1 1306.1 1028 1937.56 ;
     RECT  1003.46 741.02 1028.9 751.72 ;
     RECT  1028 1306.065 1029.02 1937.56 ;
     RECT  1029.02 1303.16 1029.5 1937.56 ;
     RECT  1027.94 2125.06 1031.78 2384.82 ;
     RECT  1029.5 1302.74 1032.1 1937.56 ;
     RECT  1032.1 1302.74 1032.38 1609.54 ;
     RECT  1032.38 1301.06 1033.06 1609.54 ;
     RECT  1012.42 844.76 1033.22 862.6 ;
     RECT  1031.78 2125.06 1033.7 2383.99 ;
     RECT  1028.9 741.02 1036.1 746.68 ;
     RECT  1014.5 761.6 1036.38 806.74 ;
     RECT  1036.38 760.76 1036.86 806.74 ;
     RECT  1014.5 825.02 1036.86 825.22 ;
     RECT  1036.86 760.76 1037.28 825.22 ;
     RECT  1037.28 760.725 1038.3 825.22 ;
     RECT  1033.06 1301.06 1040.26 1601.31 ;
     RECT  1010.02 1976.42 1040.26 1990.06 ;
     RECT  1033.7 2126.74 1041.285 2383.99 ;
     RECT  1032.1 1618.58 1042.46 1937.56 ;
     RECT  1040.26 1301.73 1042.94 1601.31 ;
     RECT  1042.46 1615.64 1042.94 1937.56 ;
     RECT  1038.3 760.34 1043.58 829 ;
     RECT  1042.94 1301.73 1043.9 1937.56 ;
     RECT  1043.58 760.34 1044.06 836.14 ;
     RECT  1033.22 844.76 1044.06 859.66 ;
     RECT  1040.26 1976.42 1044.1 1986.7 ;
     RECT  1043.9 1301.73 1044.565 1939.24 ;
     RECT  1044.565 1302.32 1045.54 1939.24 ;
     RECT  1045.54 1608.08 1046.02 1939.24 ;
     RECT  1046.02 1611.86 1046.26 1939.24 ;
     RECT  954.5 2443.84 1046.66 2446.56 ;
     RECT  1045.54 1302.32 1047.46 1598.2 ;
     RECT  1036.1 741.44 1048.38 746.68 ;
     RECT  1044.06 760.34 1048.38 863.44 ;
     RECT  1048.38 741.44 1049.54 863.44 ;
     RECT  1047.46 1302.32 1050.82 1597.78 ;
     RECT  981 -70 1051 180 ;
     RECT  1041.285 2126.74 1051.46 2380.62 ;
     RECT  1051.46 2130.52 1051.925 2380.62 ;
     RECT  1049.54 752.78 1053.18 863.44 ;
     RECT  1012.42 874.76 1053.18 874.96 ;
     RECT  1049.54 741.44 1058.94 744.16 ;
     RECT  1053.18 752.78 1058.94 878.14 ;
     RECT  1050.82 1302.74 1059.74 1597.78 ;
     RECT  1059.74 1302.32 1060.22 1597.78 ;
     RECT  991 3219.2 1061 3470 ;
     RECT  1058.94 741.44 1061.34 878.14 ;
     RECT  1051.925 2130.94 1061.82 2380.62 ;
     RECT  1045.82 1960.46 1062.14 1960.66 ;
     RECT  1061.34 741.44 1062.5 881.5 ;
     RECT  1060.22 1301.06 1063.1 1597.78 ;
     RECT  1046.26 1612.28 1064.74 1939.24 ;
     RECT  1044.1 1976.84 1065.5 1986.7 ;
     RECT  1062.5 743.96 1065.6 881.5 ;
     RECT  1062.3 892.64 1066.14 892.84 ;
     RECT  1063.1 1298.12 1066.46 1597.78 ;
     RECT  1061.82 2130.1 1066.62 2380.62 ;
     RECT  1066.46 1296.86 1068.38 1597.78 ;
     RECT  1068.38 1296.86 1069.34 1598.2 ;
     RECT  1069.34 1295.18 1070.24 1598.2 ;
     RECT  1062.14 1953.32 1070.3 1960.66 ;
     RECT  1066.14 891.8 1072.38 892.84 ;
     RECT  1064.74 1621.94 1072.7 1939.24 ;
     RECT  1070.3 1948.7 1072.7 1960.66 ;
     RECT  1070.24 1294.17 1073.18 1598.2 ;
     RECT  1065.6 743.96 1073.34 882.09 ;
     RECT  1072.38 891.8 1073.34 893.26 ;
     RECT  1073.18 1290.56 1074.14 1599.88 ;
     RECT  1066.62 2130.1 1074.5 2381.04 ;
     RECT  1074.14 1290.56 1075.1 1600.72 ;
     RECT  1064.74 1612.28 1075.1 1612.9 ;
     RECT  1073.34 743.96 1078.08 893.26 ;
     RECT  1072.7 1621.94 1078.66 1961.5 ;
     RECT  1075.1 1290.56 1079.9 1601.56 ;
     RECT  1075.1 1611.44 1079.9 1612.9 ;
     RECT  1079.9 1290.56 1080.86 1612.9 ;
     RECT  1078.66 1621.94 1080.86 1701.1 ;
     RECT  1078.08 743.96 1081.44 897.21 ;
     RECT  1078.66 1710.14 1083.74 1961.5 ;
     RECT  1065.5 1970.12 1083.74 1986.7 ;
     RECT  1080.86 1290.56 1085.86 1701.1 ;
     RECT  1074.5 2132.62 1086.78 2381.04 ;
     RECT  1086.78 2130.52 1087.26 2381.04 ;
     RECT  1087.26 2130.1 1087.46 2381.04 ;
     RECT  1085.86 1291.82 1088.3 1701.1 ;
     RECT  1083.74 1710.14 1088.3 1986.7 ;
     RECT  932.26 2012.12 1088.74 2012.74 ;
     RECT  1081.44 741.27 1091.1 897.21 ;
     RECT  1087.46 2132.62 1093.7 2381.04 ;
     RECT  1088.3 1291.82 1094.78 1986.7 ;
     RECT  1091.1 741.27 1095.42 897.46 ;
     RECT  1093.7 2133.46 1095.9 2381.04 ;
     RECT  1094.78 1283.84 1096.7 1986.7 ;
     RECT  1095.42 734.3 1097.34 897.46 ;
     RECT  1097.34 733.04 1098.3 897.46 ;
     RECT  1098.3 732.62 1102.62 897.46 ;
     RECT  1096.7 1283 1104.38 1986.7 ;
     RECT  1102.62 732.62 1109.85 900.82 ;
     RECT  1109.85 732.62 1110.32 901.16 ;
     RECT  1046.66 2443.84 1113.86 2444.04 ;
     RECT  1112.22 2471.56 1118.46 2471.76 ;
     RECT  1104.38 1281.74 1121.065 1986.7 ;
     RECT  1121.065 1276.265 1121.56 1986.7 ;
     RECT  1119.42 2123.8 1123.74 2124 ;
     RECT  1095.9 2133.46 1123.74 2381.46 ;
     RECT  1110.32 732.62 1124.25 900.82 ;
     RECT  1118.46 2466.52 1125.66 2471.76 ;
     RECT  1124.25 732.62 1126.62 901.16 ;
     RECT  1126.62 732.62 1127.975 902.5 ;
     RECT  1088.74 2012.12 1128.58 2012.32 ;
     RECT  1127.975 732.62 1128.755 903.76 ;
     RECT  1121.56 1275.43 1128.965 1986.7 ;
     RECT  1123.74 2123.8 1129.02 2381.46 ;
     RECT  1122.78 2453.92 1129.02 2454.12 ;
     RECT  1128.755 732.62 1129.22 904.6 ;
     RECT  1129.02 2123.8 1129.22 2382.72 ;
     RECT  946.62 2428.72 1130.46 2428.92 ;
     RECT  1129.22 733.46 1130.66 904.6 ;
     RECT  1130.66 737.57 1132.1 904.6 ;
     RECT  1132.1 737.66 1132.58 904.6 ;
     RECT  1132.58 738.08 1133.34 904.6 ;
     RECT  1129.22 2123.8 1134.5 2381.04 ;
     RECT  1129.02 2451.4 1134.78 2454.12 ;
     RECT  1133.34 738.08 1139.58 905.02 ;
     RECT  1128.965 1275.44 1142.02 1986.7 ;
     RECT  1139.58 738.08 1144.1 909.22 ;
     RECT  1142.02 1863.02 1144.7 1986.7 ;
     RECT  1144.1 738.08 1144.86 908.8 ;
     RECT  1142.02 1275.44 1146.82 1854.4 ;
     RECT  1144.7 1863.02 1146.82 1987.12 ;
     RECT  1134.5 2123.8 1147.74 2379.36 ;
     RECT  1146.82 1630.34 1150.94 1854.4 ;
     RECT  1146.82 1863.02 1150.94 1964.86 ;
     RECT  1147.74 2123.8 1151.58 2381.46 ;
     RECT  1151.58 2123.8 1153.5 2382.72 ;
     RECT  1153.5 2123.8 1153.98 2386.5 ;
     RECT  1144.86 737.66 1154.46 908.8 ;
     RECT  1134.78 2451.4 1154.94 2456.64 ;
     RECT  1125.66 2466.52 1154.94 2474.28 ;
     RECT  1146.82 1275.44 1155.26 1619.62 ;
     RECT  1150.94 1630.34 1155.26 1964.86 ;
     RECT  1155.26 1275.44 1155.74 1964.86 ;
     RECT  1146.82 1973.48 1155.74 1987.12 ;
     RECT  1153.98 2123.8 1157.34 2387.34 ;
     RECT  1154.46 737.66 1158.78 909.22 ;
     RECT  1157.34 2123.8 1159.26 2390.28 ;
     RECT  1130.46 2421.16 1159.74 2428.92 ;
     RECT  1158.78 736.82 1162.82 909.22 ;
     RECT  1155.74 1275.44 1164.86 1987.12 ;
     RECT  1164.86 1275.44 1167.26 1987.54 ;
     RECT  1159.26 2123.8 1172.22 2392.38 ;
     RECT  1172.22 2123.8 1172.9 2394.06 ;
     RECT  1162.82 736.82 1173.095 908.38 ;
     RECT  1167.26 1275.44 1173.7 1990.06 ;
     RECT  1172.9 2159.08 1174.14 2394.06 ;
     RECT  1174.14 2159.08 1174.33 2396.16 ;
     RECT  1172.9 2123.8 1174.34 2149.62 ;
     RECT  1174.34 2143.96 1174.82 2149.62 ;
     RECT  1051 0 1175 180 ;
     RECT  1173.7 1282.58 1175.075 1990.06 ;
     RECT  1174.82 2143.96 1175.3 2145 ;
     RECT  1174.33 2159.08 1175.3 2214.72 ;
     RECT  1175.075 1967.58 1175.525 1990.06 ;
     RECT  1175.075 1282.58 1175.62 1958.98 ;
     RECT  1173.095 736.82 1176.06 908.8 ;
     RECT  1175.3 2172.1 1176.26 2202.12 ;
     RECT  1175.62 1282.58 1176.58 1953.02 ;
     RECT  1176.58 1283 1176.88 1953.02 ;
     RECT  1176.26 2201.92 1176.98 2202.12 ;
     RECT  1176.26 2172.1 1177.22 2173.14 ;
     RECT  1176.88 1283 1177.3 1952.68 ;
     RECT  1175.3 2159.08 1178.18 2159.7 ;
     RECT  1176.26 2183.02 1178.18 2190.78 ;
     RECT  1177.3 1952.06 1179.69 1952.68 ;
     RECT  1176.06 735.14 1180.265 908.8 ;
     RECT  1180.265 735.14 1182.78 912.595 ;
     RECT  1177.3 1283 1183.3 1941.76 ;
     RECT  1179.69 1952.48 1183.3 1952.68 ;
     RECT  1061 3219.2 1185 3400 ;
     RECT  1182.78 730.1 1185.66 912.595 ;
     RECT  1185.66 729.68 1187.715 912.595 ;
     RECT  1172.22 2441.32 1188.06 2441.52 ;
     RECT  1154.94 2451.4 1188.06 2474.28 ;
     RECT  1187.715 729.68 1188.165 911.76 ;
     RECT  1175 -70 1188.38 180 ;
     RECT  1036.22 226.7 1188.38 226.9 ;
     RECT  1159.74 2421.16 1188.54 2431.44 ;
     RECT  1188.06 2441.32 1188.54 2474.28 ;
     RECT  1188.38 -70 1188.58 180.7 ;
     RECT  1174.33 2229.64 1190.94 2396.16 ;
     RECT  1188.165 729.68 1192.1 911.74 ;
     RECT  1192.1 729.68 1194.3 900.82 ;
     RECT  1183.3 1283 1194.325 1937.98 ;
     RECT  1194.325 1283 1194.34 1646.08 ;
     RECT  1194.34 1283 1195.06 1645.24 ;
     RECT  1194.325 1656.785 1195.3 1937.98 ;
     RECT  1194.3 729.26 1195.94 900.82 ;
     RECT  1195.06 1283 1198.165 1642.3 ;
     RECT  1195.3 1656.785 1198.595 1937.14 ;
     RECT  1195.94 729.68 1201.7 900.82 ;
     RECT  1198.595 1656.8 1202.5 1937.14 ;
     RECT  1175.3 2214.52 1203.9 2214.72 ;
     RECT  1198.165 1283 1204.42 1641.46 ;
     RECT  1202.5 1660.58 1204.9 1937.14 ;
     RECT  1204.42 1287.2 1206.34 1630.12 ;
     RECT  1201.7 730.1 1206.81 900.82 ;
     RECT  1206.81 730.1 1206.88 901.16 ;
     RECT  1190.94 2229.64 1210.62 2403.72 ;
     RECT  1206.88 730.1 1210.82 901.24 ;
     RECT  1210.82 730.1 1213.7 900.82 ;
     RECT  1213.7 730.1 1213.93 897.04 ;
     RECT  1210.62 2229.64 1214.66 2406.24 ;
     RECT  1206.34 1287.2 1214.98 1627.6 ;
     RECT  1214.98 1288.04 1215.46 1627.6 ;
     RECT  1213.93 730.1 1215.62 896.2 ;
     RECT  1215.62 730.52 1216.1 896.2 ;
     RECT  1204.9 1663.1 1216.62 1937.14 ;
     RECT  1216.62 1658.06 1217.395 1937.14 ;
     RECT  1214.66 2353.96 1218.02 2406.24 ;
     RECT  1203.9 2214.52 1218.3 2216.82 ;
     RECT  1185 3219.2 1218.34 3470 ;
     RECT  1215.46 1290.98 1218.805 1627.6 ;
     RECT  1218.805 1291.82 1220.06 1627.6 ;
     RECT  1216.1 731.36 1220.42 896.2 ;
     RECT  1220.06 1291.82 1220.96 1630.54 ;
     RECT  1220.96 1291.82 1222.18 1631.55 ;
     RECT  1217.395 1657.22 1222.46 1937.14 ;
     RECT  1220.42 731.36 1223.78 893.26 ;
     RECT  1222.18 1298.54 1224.1 1631.55 ;
     RECT  1224.1 1309.29 1224.38 1631.55 ;
     RECT  1204.42 1641.26 1224.38 1641.46 ;
     RECT  1214.66 2229.64 1224.54 2344.5 ;
     RECT  1224.1 1298.54 1224.565 1299.58 ;
     RECT  1224.54 2229.64 1224.74 2348.28 ;
     RECT  1224.38 1309.29 1225.045 1641.46 ;
     RECT  1222.46 1653.44 1227.46 1937.14 ;
     RECT  1224.565 1299.38 1227.94 1299.58 ;
     RECT  1227.46 1653.44 1227.94 1828.78 ;
     RECT  1225.045 1310.3 1228.22 1641.46 ;
     RECT  1228.22 1310.3 1228.42 1643.56 ;
     RECT  1223.78 735.14 1228.58 893.26 ;
     RECT  1178.18 2185.54 1228.86 2185.74 ;
     RECT  1228.42 1313.66 1229.365 1643.56 ;
     RECT  1227.94 1653.44 1229.86 1827.52 ;
     RECT  1188.58 -70 1229.9 180 ;
     RECT  1191.74 716.42 1230.14 716.62 ;
     RECT  1229.9 -70 1230.34 180.7 ;
     RECT  1229.86 1774.82 1231.3 1827.52 ;
     RECT  1229.365 1315.76 1231.58 1643.56 ;
     RECT  1229.86 1653.44 1231.58 1760.32 ;
     RECT  1228.58 736.82 1233.66 893.26 ;
     RECT  1231.3 1774.82 1234.66 1825.42 ;
     RECT  1233.66 736.82 1234.82 893.68 ;
     RECT  1231.58 1315.76 1235.14 1760.32 ;
     RECT  1235.14 1638.32 1235.62 1760.32 ;
     RECT  1234.82 744.8 1236.06 893.68 ;
     RECT  1178.18 2159.08 1236.06 2159.28 ;
     RECT  1234.66 1798.34 1236.1 1825.42 ;
     RECT  1235.14 1315.76 1236.58 1628.44 ;
     RECT  1235.42 1953.32 1237.34 1953.52 ;
     RECT  1236.58 1325 1237.54 1628.44 ;
     RECT  1235.62 1638.32 1237.54 1756.54 ;
     RECT  1236.1 1819.76 1237.54 1825.42 ;
     RECT  1237.54 1325.84 1238.02 1628.44 ;
     RECT  1237.34 1951.64 1238.3 1953.52 ;
     RECT  1237.54 1647.14 1238.5 1756.54 ;
     RECT  1238.02 1325.84 1238.74 1627.6 ;
     RECT  1238.3 1948.28 1239.26 1953.52 ;
     RECT  1239.26 1946.18 1240.7 1953.52 ;
     RECT  1238.5 1653.86 1241.365 1756.54 ;
     RECT  1237.54 1638.32 1241.38 1638.52 ;
     RECT  1227.46 1840.34 1241.66 1937.14 ;
     RECT  1240.7 1946.18 1241.66 1955.62 ;
     RECT  1175.525 1973.48 1241.66 1990.06 ;
     RECT  1218.02 2362.78 1242.02 2406.24 ;
     RECT  1238.74 1328.78 1242.58 1627.6 ;
     RECT  1241.66 1840.34 1242.62 1955.62 ;
     RECT  1241.66 1970.12 1242.62 1990.06 ;
     RECT  1242.58 1339.53 1242.82 1627.6 ;
     RECT  1236.06 744.8 1244.22 894.1 ;
     RECT  1242.58 1328.78 1244.725 1329.82 ;
     RECT  1241.365 1654.28 1244.74 1756.54 ;
     RECT  1230.34 -70 1245 180 ;
     RECT  1242.82 1339.53 1245.205 1623.99 ;
     RECT  1244.74 1657.22 1245.22 1756.54 ;
     RECT  1234.66 1774.82 1245.5 1788.88 ;
     RECT  1236.1 1798.34 1245.5 1807.36 ;
     RECT  1245.22 1657.64 1245.74 1756.54 ;
     RECT  1245.74 1657.64 1246.18 1758.64 ;
     RECT  1245.5 1774.82 1246.46 1807.36 ;
     RECT  1244.22 744.8 1246.62 897.88 ;
     RECT  1246.46 1774.82 1246.66 1807.78 ;
     RECT  1246.62 744.8 1247.52 903.76 ;
     RECT  1246.18 1657.64 1247.62 1756.46 ;
     RECT  1244.725 1329.62 1248.1 1329.82 ;
     RECT  1247.62 1658.06 1248.34 1756.46 ;
     RECT  1245.205 1339.53 1248.565 1622.14 ;
     RECT  1248.34 1659.74 1249.06 1756.46 ;
     RECT  1249.06 1660.58 1250.02 1756.46 ;
     RECT  1250.02 1662.26 1250.25 1756.46 ;
     RECT  1250.25 1662.26 1250.98 1755.28 ;
     RECT  1247.52 744.8 1251.14 904.77 ;
     RECT  1250.98 1664.36 1251.46 1755.28 ;
     RECT  1248.565 1340.54 1251.94 1622.14 ;
     RECT  1251.94 1347.09 1252.885 1622.14 ;
     RECT  1252.885 1347.68 1253.86 1622.14 ;
     RECT  1251.46 1664.36 1253.86 1664.56 ;
     RECT  1218.34 3220 1255 3470 ;
     RECT  1255.1 1763.9 1256.06 1764.52 ;
     RECT  1253.86 1348.1 1256.26 1622.14 ;
     RECT  1256.26 1351.46 1256.74 1622.14 ;
     RECT  1256.06 1763.9 1257.02 1766.2 ;
     RECT  1246.66 1774.82 1257.02 1806.1 ;
     RECT  1251.14 755.72 1258.14 904.77 ;
     RECT  1256.74 1354.385 1259.14 1622.14 ;
     RECT  1251.14 744.8 1259.3 745 ;
     RECT  1258.94 1650.92 1259.9 1651.12 ;
     RECT  1251.46 1675.7 1260.38 1755.28 ;
     RECT  1260.38 1675.28 1260.86 1755.28 ;
     RECT  1257.02 1763.9 1260.86 1806.1 ;
     RECT  1259.14 1354.385 1260.995 1355.45 ;
     RECT  1260.995 1355.22 1261.445 1355.45 ;
     RECT  1259.14 1369.94 1262.02 1622.14 ;
     RECT  1259.9 1650.08 1262.3 1651.12 ;
     RECT  1262.02 1378.34 1262.5 1622.14 ;
     RECT  1262.3 1649.24 1262.78 1651.12 ;
     RECT  1260.38 1660.16 1262.78 1660.78 ;
     RECT  1260.86 1675.28 1262.78 1806.1 ;
     RECT  1262.5 1391.78 1262.98 1622.14 ;
     RECT  1262.78 1645.04 1263.26 1651.12 ;
     RECT  1262.78 1660.16 1263.26 1806.1 ;
     RECT  1262.5 1378.34 1263.46 1382.07 ;
     RECT  1262.98 1391.78 1264.405 1604.5 ;
     RECT  1258.14 755.72 1264.86 905.02 ;
     RECT  1263.46 1380.44 1264.885 1382.07 ;
     RECT  1264.405 1405.22 1264.9 1604.5 ;
     RECT  1264.9 1445.54 1265.365 1604.5 ;
     RECT  1264.86 755.72 1266.5 908.38 ;
     RECT  1237.54 1821.44 1266.62 1825.42 ;
     RECT  1264.405 1391.78 1266.82 1396.18 ;
     RECT  1263.26 1645.04 1267.1 1806.1 ;
     RECT  1266.62 1821.44 1267.1 1831.3 ;
     RECT  1242.62 1840.34 1267.1 1990.06 ;
     RECT  1266.82 1391.78 1267.3 1391.98 ;
     RECT  1265.365 1445.54 1267.3 1603.66 ;
     RECT  1267.3 1448.48 1267.54 1603.66 ;
     RECT  1264.9 1405.22 1267.78 1435.66 ;
     RECT  1267.1 1642.94 1268.06 1806.1 ;
     RECT  1264.885 1380.44 1268.26 1380.64 ;
     RECT  1267.54 1453.94 1268.74 1603.66 ;
     RECT  1268.74 1460.66 1268.98 1599.88 ;
     RECT  1266.5 756.14 1269.86 908.38 ;
     RECT  1268.98 1460.66 1270.18 1596.94 ;
     RECT  1267.78 1412.78 1270.645 1435.66 ;
     RECT  1270.645 1412.78 1271.14 1426 ;
     RECT  1269.98 3059.18 1271.42 3059.38 ;
     RECT  1271.14 1415.7 1271.525 1426 ;
     RECT  1271.525 1415.72 1272.1 1426 ;
     RECT  1270.645 1435.46 1272.1 1435.66 ;
     RECT  1268.06 1641.68 1272.38 1806.1 ;
     RECT  1272.1 1420.34 1272.58 1426 ;
     RECT  1270.18 1461.08 1273.525 1596.94 ;
     RECT  1272.38 1637.48 1273.54 1806.1 ;
     RECT  1269.86 756.56 1273.98 908.38 ;
     RECT  1272.58 1425.8 1274.02 1426 ;
     RECT  1271.42 3056.66 1274.3 3059.8 ;
     RECT  1267.1 1821.44 1274.78 1990.06 ;
     RECT  1273.525 1461.08 1275.46 1593.16 ;
     RECT  1274.78 1821.44 1275.46 1991.32 ;
     RECT  1274.3 3056.66 1275.74 3064 ;
     RECT  1275.46 1461.08 1276.355 1578.895 ;
     RECT  1275.46 1590.44 1276.42 1593.16 ;
     RECT  1276.355 1461.08 1276.805 1578.06 ;
     RECT  1276.42 1592.96 1276.9 1593.16 ;
     RECT  1275.74 3055.82 1279.1 3064.84 ;
     RECT  1276.805 1461.08 1279.3 1575.52 ;
     RECT  1279.1 3055.82 1279.58 3066.52 ;
     RECT  1273.98 756.56 1279.74 909.22 ;
     RECT  1279.58 3048.26 1280.06 3066.52 ;
     RECT  1279.3 1465.28 1280.26 1567.13 ;
     RECT  1275.46 1821.44 1281.5 1990.06 ;
     RECT  1280.06 3047.84 1281.5 3066.52 ;
     RECT  1281.5 1816.4 1282.46 1990.06 ;
     RECT  1281.5 3047.84 1282.94 3067.78 ;
     RECT  1279.74 750.26 1284.06 909.22 ;
     RECT  1284.06 750.26 1284.54 912.16 ;
     RECT  1282.94 3047.84 1284.86 3071.56 ;
     RECT  1284.54 742.7 1285.02 912.16 ;
     RECT  1284.86 3047.84 1285.82 3073.66 ;
     RECT  1280.26 1465.7 1286.98 1567.13 ;
     RECT  1286.98 1479.55 1287.845 1567.13 ;
     RECT  1273.54 1638.74 1288.7 1806.1 ;
     RECT  1282.46 1815.56 1288.7 1990.06 ;
     RECT  1285.82 3047.84 1288.7 3074.5 ;
     RECT  1287.845 1484.18 1288.885 1567.13 ;
     RECT  1288.885 1484.18 1288.9 1505.38 ;
     RECT  1288.7 1638.74 1289 1990.06 ;
     RECT  1289 1638.32 1289.18 1990.06 ;
     RECT  1288.9 1484.6 1289.38 1505.38 ;
     RECT  1288.885 1514.42 1289.38 1567.13 ;
     RECT  1289.18 1638.32 1289.86 1991.32 ;
     RECT  1285.02 736.82 1290.02 912.16 ;
     RECT  1174.34 2123.8 1290.3 2134.08 ;
     RECT  1200.06 2146.48 1290.3 2146.68 ;
     RECT  1236.06 2159.08 1290.3 2166.84 ;
     RECT  1228.86 2185.54 1290.3 2192.04 ;
     RECT  1228.86 2204.86 1290.3 2205.06 ;
     RECT  1218.3 2214.52 1290.3 2217.24 ;
     RECT  1224.74 2229.64 1290.3 2320.56 ;
     RECT  1224.74 2329.18 1290.3 2348.28 ;
     RECT  1242.02 2364.04 1290.3 2406.24 ;
     RECT  1289.38 1524.5 1290.34 1567.13 ;
     RECT  1288.7 3047.84 1290.62 3078.7 ;
     RECT  1290.34 1530.38 1290.725 1532.7 ;
     RECT  1289.38 1486.7 1290.82 1505.38 ;
     RECT  1290.34 1546.76 1290.82 1567.13 ;
     RECT  1290.725 1530.38 1291.3 1532.68 ;
     RECT  1289.38 1514.42 1291.78 1515.04 ;
     RECT  1290.82 1559.78 1292.165 1567.13 ;
     RECT  1290.82 1499.3 1292.26 1505.38 ;
     RECT  1290.82 1546.76 1292.26 1550.32 ;
     RECT  1291.58 2936.12 1292.54 2936.32 ;
     RECT  1290.62 3047.84 1292.54 3079.12 ;
     RECT  1292.54 3045.74 1293.02 3079.12 ;
     RECT  1293.02 3044.06 1293.5 3079.12 ;
     RECT  1290.3 2123.8 1293.66 2217.24 ;
     RECT  1290.3 2227.12 1293.66 2348.28 ;
     RECT  1289.86 1638.32 1293.98 1990.48 ;
     RECT  1293.66 2123.8 1294.62 2348.28 ;
     RECT  1290.3 2358.16 1294.62 2406.24 ;
     RECT  1292.165 1559.78 1294.66 1563.34 ;
     RECT  1294.94 2919.32 1295.9 2919.52 ;
     RECT  1292.54 2928.56 1295.9 2936.32 ;
     RECT  1188.54 2421.16 1296.06 2474.28 ;
     RECT  1292.26 1499.3 1296.1 1499.92 ;
     RECT  1293.98 1637.06 1296.86 1990.48 ;
     RECT  1165.82 2039 1296.86 2039.2 ;
     RECT  1294.62 2123.8 1296.86 2406.24 ;
     RECT  1290.02 737.24 1297.45 912.16 ;
     RECT  1296.86 2121.74 1297.5 2406.24 ;
     RECT  1296.06 2416.12 1297.5 2474.28 ;
     RECT  1281.98 3186.86 1297.82 3187.06 ;
     RECT  1297.82 3033.56 1298.3 3033.76 ;
     RECT  1293.5 3044.06 1298.3 3079.96 ;
     RECT  1298.3 3044.06 1298.5 3081.64 ;
     RECT  1297.82 2100.32 1298.78 2100.52 ;
     RECT  1295.9 2919.32 1298.78 2936.32 ;
     RECT  1297.45 737.24 1298.94 911.74 ;
     RECT  1297.5 2121.74 1298.94 2474.28 ;
     RECT  1262.98 1616.06 1299.26 1622.14 ;
     RECT  1298.3 3032.3 1299.26 3033.76 ;
     RECT  1298.5 3044.06 1299.26 3079.96 ;
     RECT  1298.94 2121.74 1299.74 2476.8 ;
     RECT  1298.94 734.72 1299.84 911.74 ;
     RECT  1296.86 2039 1300.22 2041.72 ;
     RECT  1299.26 1616.06 1300.7 1622.98 ;
     RECT  1299.74 2121.74 1301.18 2476.84 ;
     RECT  1300.7 1614.8 1301.66 1622.98 ;
     RECT  1301.18 2117.12 1301.86 2476.84 ;
     RECT  1301.66 1614.8 1302.14 1624.66 ;
     RECT  1296.86 1635.8 1302.14 1990.48 ;
     RECT  1230.14 716.42 1302.3 723.76 ;
     RECT  1299.84 733.71 1302.3 911.74 ;
     RECT  1302.3 716.42 1302.5 911.74 ;
     RECT  1302.14 1614.8 1302.62 1990.48 ;
     RECT  1301.86 2129.3 1303.3 2150.5 ;
     RECT  1302.62 1614.8 1303.58 1991.32 ;
     RECT  1303.58 1614.8 1304.06 1993 ;
     RECT  1298.78 2919.32 1305.98 2938 ;
     RECT  1302.5 716.42 1306.34 909.64 ;
     RECT  1305.5 2004.98 1306.46 2005.6 ;
     RECT  1305.98 2917.64 1306.94 2938 ;
     RECT  1306.94 2917.22 1307.68 2938 ;
     RECT  1299.26 3032.3 1307.68 3079.96 ;
     RECT  1304.06 1611.44 1307.9 1993 ;
     RECT  1306.46 2004.14 1307.9 2008.12 ;
     RECT  1306.46 1600.52 1308.38 1600.72 ;
     RECT  1307.9 1611.44 1308.38 2008.12 ;
     RECT  1307.68 2917.22 1308.38 3177.88 ;
     RECT  1308.38 1600.52 1309.34 2008.12 ;
     RECT  1301.86 2117.12 1309.82 2117.32 ;
     RECT  1306.34 733.04 1310.66 909.64 ;
     RECT  1309.34 1592.12 1310.78 2008.12 ;
     RECT  1303.3 2131.4 1310.78 2150.5 ;
     RECT  1310.3 1582.46 1311.26 1583.08 ;
     RECT  1310.78 1592.12 1311.26 2009.8 ;
     RECT  1310.78 2131.4 1311.26 2151.76 ;
     RECT  1301.86 2161.64 1311.26 2476.84 ;
     RECT  1311.26 2131.4 1311.74 2476.84 ;
     RECT  1310.66 733.46 1312.1 909.64 ;
     RECT  1311.26 1577 1312.22 2009.8 ;
     RECT  1309.82 2110.82 1312.22 2117.32 ;
     RECT  1311.74 2130.56 1312.22 2476.84 ;
     RECT  1312.1 733.46 1313.06 822.28 ;
     RECT  1312.22 1577 1313.18 2013.58 ;
     RECT  1312.22 2130.14 1313.38 2476.84 ;
     RECT  1313.38 2130.14 1313.66 2454.16 ;
     RECT  1298.78 2100.32 1315.58 2101.36 ;
     RECT  1312.1 831.74 1316.105 909.64 ;
     RECT  1313.18 1577 1316.74 2014 ;
     RECT  1316.74 1577 1317.22 2010.64 ;
     RECT  1315.58 2091.92 1317.5 2101.36 ;
     RECT  1312.22 2109.98 1317.5 2117.32 ;
     RECT  1313.66 2129.3 1318.66 2454.16 ;
     RECT  1317.5 2091.5 1318.94 2117.32 ;
     RECT  1308.38 2915.54 1318.94 3177.88 ;
     RECT  1313.06 737.32 1319.12 822.28 ;
     RECT  1318.94 2083.52 1320.38 2117.32 ;
     RECT  1318.66 2129.3 1320.38 2436.1 ;
     RECT  1318.66 2448.08 1320.58 2454.16 ;
     RECT  1316.105 831.74 1320.74 912.595 ;
     RECT  1320.38 2083.52 1321.06 2436.1 ;
     RECT  1319.12 737.815 1321.93 822.28 ;
     RECT  1318.94 2913.44 1322.78 3177.88 ;
     RECT  1321.93 741.02 1323.14 822.28 ;
     RECT  1320.74 851.06 1323.555 912.595 ;
     RECT  1321.06 2083.52 1323.94 2435.26 ;
     RECT  1323.555 851.06 1324.005 911.76 ;
     RECT  1301.18 2069.66 1324.22 2069.86 ;
     RECT  1322.78 2908.82 1324.42 3177.88 ;
     RECT  1294.66 1559.78 1324.7 1559.98 ;
     RECT  1324.22 2062.52 1324.7 2069.86 ;
     RECT  1323.94 2083.52 1325.18 2432.32 ;
     RECT  1317.22 1577.42 1325.66 2010.64 ;
     RECT  1324.7 2062.52 1325.66 2070.28 ;
     RECT  1325.66 1577.42 1325.86 2012.32 ;
     RECT  1324.7 1558.94 1326.14 1559.98 ;
     RECT  1325.86 1577.42 1326.14 2010.22 ;
     RECT  1325.66 2060 1326.14 2070.28 ;
     RECT  1325.18 2083.1 1326.14 2432.32 ;
     RECT  1324.005 851.06 1326.5 908.8 ;
     RECT  1326.62 2050.34 1327.1 2050.96 ;
     RECT  1326.14 2060 1327.1 2432.32 ;
     RECT  1326.5 865.76 1327.46 908.8 ;
     RECT  1323.14 741.02 1327.94 808 ;
     RECT  1300.22 2033.96 1328.06 2041.72 ;
     RECT  1327.1 2050.34 1328.06 2432.32 ;
     RECT  1323.14 817.04 1328.17 822.28 ;
     RECT  1327.46 866.18 1331.78 908.8 ;
     RECT  1331.78 869.12 1332.26 908.8 ;
     RECT  1328.06 2033.96 1333.54 2432.32 ;
     RECT  1332.26 869.79 1334.66 908.8 ;
     RECT  1326.14 1558.94 1334.78 2010.22 ;
     RECT  1324.42 2913.44 1334.78 3177.88 ;
     RECT  1334.78 1558.94 1334.98 2012.32 ;
     RECT  1334.78 2907.56 1335.74 3177.88 ;
     RECT  1334.66 893.06 1336.58 908.8 ;
     RECT  1336.58 893.9 1337.06 908.8 ;
     RECT  1299.26 1343.48 1337.86 1343.68 ;
     RECT  1327.94 741.44 1338.3 808 ;
     RECT  1320.74 831.74 1338.5 834.46 ;
     RECT  1337.06 896 1340.42 908.8 ;
     RECT  1334.66 869.79 1340.885 882.76 ;
     RECT  1340.42 896 1343.53 904.6 ;
     RECT  1334.98 1558.94 1343.9 2010.64 ;
     RECT  1340.885 871.22 1344.26 882.76 ;
     RECT  1338.3 740.6 1344.74 808 ;
     RECT  1344.26 875 1346.18 882.76 ;
     RECT  1346.18 882.56 1346.66 882.76 ;
     RECT  1343.53 896 1347.14 904.18 ;
     RECT  1347.14 896 1348.38 896.2 ;
     RECT  1333.54 2033.96 1348.42 2426.44 ;
     RECT  1348.38 895.58 1348.58 896.2 ;
     RECT  1344.74 741.44 1349.29 808 ;
     RECT  1348.42 2033.96 1349.38 2399.56 ;
     RECT  1348.42 2408.6 1350.82 2426.44 ;
     RECT  1343.9 1558.94 1352.06 2014.42 ;
     RECT  1349.29 741.86 1352.9 808 ;
     RECT  1349.38 2033.96 1353.7 2394.52 ;
     RECT  1338.5 831.74 1353.86 833.62 ;
     RECT  1352.06 1558.94 1354.94 2014.84 ;
     RECT  1352.9 749 1355.1 808 ;
     RECT  1328.17 817.46 1355.1 822.28 ;
     RECT  1353.7 2380.88 1355.62 2393.68 ;
     RECT  1354.94 1558.94 1356.58 2015.68 ;
     RECT  1353.86 832.16 1357.02 833.62 ;
     RECT  1355.62 2380.88 1357.06 2391.16 ;
     RECT  1335.74 2905.46 1360.22 3177.88 ;
     RECT  1357.06 2380.88 1360.42 2386.54 ;
     RECT  1356.58 1773.14 1361.86 2015.68 ;
     RECT  1356.58 1558.94 1362.34 1764.1 ;
     RECT  1353.7 2033.96 1362.82 2365.96 ;
     RECT  1357.02 832.16 1363.26 839.92 ;
     RECT  1326.5 851.06 1363.26 851.26 ;
     RECT  1362.34 1558.94 1363.3 1763.68 ;
     RECT  1362.82 2346.86 1364.06 2365.96 ;
     RECT  1290.82 1486.7 1364.905 1486.9 ;
     RECT  1363.3 1558.94 1367.14 1759.06 ;
     RECT  1362.82 2033.96 1367.14 2334.46 ;
     RECT  1367.14 1558.94 1368.1 1749.4 ;
     RECT  1245 0 1369 180 ;
     RECT  1368.1 1558.94 1370.98 1748.98 ;
     RECT  1367.14 2033.96 1371.46 2331.52 ;
     RECT  1361.86 1773.14 1372.7 2013.58 ;
     RECT  1371.46 2269.41 1372.9 2331.52 ;
     RECT  1364.905 1486.7 1373.18 1488.175 ;
     RECT  1286.98 1465.7 1373.38 1465.9 ;
     RECT  1372.7 1773.14 1373.66 2015.68 ;
     RECT  1372.9 2314.94 1375.05 2331.52 ;
     RECT  1373.18 1486.28 1375.1 1488.175 ;
     RECT  1360.42 2380.88 1375.1 2381.08 ;
     RECT  1375.1 1486.28 1375.3 1489 ;
     RECT  1370.98 1558.94 1375.3 1748.56 ;
     RECT  1373.66 1773.14 1375.3 2017.36 ;
     RECT  1372.9 2269.41 1375.765 2305.9 ;
     RECT  1355.1 749 1376.22 822.28 ;
     RECT  1363.26 832.16 1376.22 851.26 ;
     RECT  1371.46 2033.96 1376.245 2259.03 ;
     RECT  1376.245 2033.96 1378.18 2258.44 ;
     RECT  1375.05 2315.36 1378.18 2331.52 ;
     RECT  1375.3 1793.3 1378.46 2017.36 ;
     RECT  1378.18 2315.36 1378.66 2315.56 ;
     RECT  1255 3220 1379 3400 ;
     RECT  1375.765 2270.84 1379.14 2305.9 ;
     RECT  1379.14 2271.26 1380.005 2305.9 ;
     RECT  1380.005 2292.68 1380.1 2305.9 ;
     RECT  1378.18 2331.32 1381.06 2331.52 ;
     RECT  1378.46 1793.3 1381.34 2021.14 ;
     RECT  1375.3 1559.78 1381.54 1748.56 ;
     RECT  1381.54 1569.44 1382.3 1748.56 ;
     RECT  1367.14 1758.86 1382.3 1759.06 ;
     RECT  1381.34 1793.3 1382.3 2023.24 ;
     RECT  1382.3 1793.3 1383.26 2023.66 ;
     RECT  1378.18 2033.96 1383.26 2257.6 ;
     RECT  1369 -70 1384.7 180 ;
     RECT  1380.005 2271.26 1385.38 2280.28 ;
     RECT  1376.22 746.06 1385.66 851.26 ;
     RECT  1364.06 2346.86 1387.78 2372.26 ;
     RECT  1385.66 737.84 1388.9 851.26 ;
     RECT  1383.26 1793.3 1389.5 2257.6 ;
     RECT  1382.3 1569.44 1390.46 1759.06 ;
     RECT  1390.46 1569.44 1391.42 1759.9 ;
     RECT  1375.3 1773.14 1391.42 1784.68 ;
     RECT  1391.42 1569.44 1392.1 1784.68 ;
     RECT  1392.1 1574.48 1392.38 1784.68 ;
     RECT  1389.5 1793.3 1392.38 2258.44 ;
     RECT  1392.38 1574.48 1393.34 2258.44 ;
     RECT  1296.1 1499.3 1393.82 1499.5 ;
     RECT  1385.38 2271.26 1394.78 2276.08 ;
     RECT  1393.34 1574.48 1395.26 2262.22 ;
     RECT  1394.78 2271.26 1395.26 2281.96 ;
     RECT  1395.26 1574.48 1395.46 2281.96 ;
     RECT  1393.82 1498.46 1397.18 1499.5 ;
     RECT  1388.9 746.48 1398.62 851.26 ;
     RECT  1398.62 746.48 1399.54 854.38 ;
     RECT  1397.18 1498.46 1399.58 1506.22 ;
     RECT  1399.54 746.48 1400 852.52 ;
     RECT  1400 746.48 1400.26 851.86 ;
     RECT  1400.26 799.4 1400.74 851.86 ;
     RECT  1313.38 2465.72 1400.74 2476.84 ;
     RECT  1400.26 746.48 1401.22 790.96 ;
     RECT  1400.74 799.4 1401.7 812.38 ;
     RECT  1395.46 1576.58 1401.7 2281.96 ;
     RECT  1400.74 823.94 1402.18 851.86 ;
     RECT  1401.7 1577 1403.14 1613.32 ;
     RECT  1403.14 1577.84 1403.62 1613.32 ;
     RECT  1292.26 1549.28 1404.38 1550.32 ;
     RECT  1381.54 1559.78 1404.38 1559.98 ;
     RECT  1399.58 1498.46 1404.86 1513.78 ;
     RECT  1403.62 1584.98 1405.06 1613.32 ;
     RECT  1375.3 1486.7 1405.34 1489 ;
     RECT  1404.86 1498.46 1405.34 1516.72 ;
     RECT  1401.7 1621.94 1405.34 2281.96 ;
     RECT  1401.22 753.38 1407.46 787.18 ;
     RECT  1405.34 1621.94 1407.46 2284.9 ;
     RECT  1402.18 826.46 1408.42 849.34 ;
     RECT  1405.06 1592.54 1408.42 1613.32 ;
     RECT  1401.7 803.78 1408.9 812.38 ;
     RECT  1408.42 1592.54 1408.9 1598.2 ;
     RECT  1408.42 1607.24 1408.9 1613.32 ;
     RECT  1408.42 831.5 1409.86 849.34 ;
     RECT  1291.3 1530.38 1410.14 1530.58 ;
     RECT  1405.34 1486.7 1410.34 1516.72 ;
     RECT  1408.9 1607.24 1410.34 1607.44 ;
     RECT  1407.46 755.9 1410.82 787.18 ;
     RECT  1407.46 1621.94 1411.1 1622.14 ;
     RECT  1407.46 1630.75 1411.1 2284.9 ;
     RECT  1411.1 1621.1 1411.3 1622.14 ;
     RECT  1375.1 2380.88 1411.78 2386.96 ;
     RECT  1411.1 1630.75 1412.06 2285.74 ;
     RECT  1410.34 1486.7 1412.74 1513.78 ;
     RECT  1412.06 1630.75 1413.02 2287.84 ;
     RECT  1413.02 1630.75 1414.46 2289.1 ;
     RECT  1380.1 2297.72 1414.46 2305.9 ;
     RECT  1387.78 2350.64 1417.06 2372.26 ;
     RECT  1410.82 755.9 1417.54 783.82 ;
     RECT  1360.22 2905.04 1419.46 3177.88 ;
     RECT  1419.46 3055.4 1420.9 3177.88 ;
     RECT  1400.74 2466.56 1422.82 2476.84 ;
     RECT  1412.74 1499.3 1423.1 1513.78 ;
     RECT  1411.3 1621.1 1423.58 1621.3 ;
     RECT  1414.46 1630.75 1423.58 2305.9 ;
     RECT  1417.54 766.82 1423.78 783.82 ;
     RECT  1423.1 1499.3 1424.54 1516.72 ;
     RECT  1417.54 755.9 1424.74 756.1 ;
     RECT  1410.14 1530.38 1425.5 1531.84 ;
     RECT  1404.38 1549.28 1425.5 1559.98 ;
     RECT  1423.58 1621.1 1427.305 2305.9 ;
     RECT  1424.54 1498.88 1427.62 1516.72 ;
     RECT  1427.62 1499.3 1427.9 1516.72 ;
     RECT  1408.9 808.82 1430.5 812.38 ;
     RECT  1422.82 2466.56 1430.5 2474.32 ;
     RECT  1427.9 1499.3 1430.78 1518.4 ;
     RECT  1417.06 2351.9 1430.78 2372.26 ;
     RECT  1409.86 834.86 1432.42 849.34 ;
     RECT  1430.78 1499.3 1432.7 1521.34 ;
     RECT  1425.5 1530.38 1432.7 1532.26 ;
     RECT  1427.305 1618.985 1432.7 2305.9 ;
     RECT  1432.7 1618.985 1433.18 2308 ;
     RECT  1422.62 1578.26 1433.66 1578.46 ;
     RECT  1432.7 1499.3 1434.14 1532.26 ;
     RECT  1433.66 1578.26 1434.62 1584.76 ;
     RECT  1434.62 1578.26 1435.58 1589.8 ;
     RECT  1423.78 766.82 1435.78 777.52 ;
     RECT  1320.58 2451.44 1435.78 2454.16 ;
     RECT  1433.18 1618.985 1436.06 2308.84 ;
     RECT  1435.58 1578.26 1437.02 1590.64 ;
     RECT  1433.66 1605.14 1437.98 1605.34 ;
     RECT  1436.06 1618.985 1437.98 2310.94 ;
     RECT  1384.7 -70 1439 183.64 ;
     RECT  1437.02 1578.26 1439.14 1596.1 ;
     RECT  1430.78 2345.18 1439.14 2372.26 ;
     RECT  1412.74 1486.7 1439.42 1489 ;
     RECT  1434.14 1499.3 1439.42 1533.1 ;
     RECT  1439.42 1486.7 1439.62 1533.1 ;
     RECT  1439.62 1486.7 1440.265 1532.68 ;
     RECT  1439.14 1590.44 1440.325 1596.1 ;
     RECT  1437.98 1605.14 1440.325 2310.94 ;
     RECT  1440.325 1590.44 1442.02 2310.94 ;
     RECT  1297.82 3186.86 1442.78 3188.32 ;
     RECT  1442.78 3186.86 1442.98 3192.1 ;
     RECT  1188.38 219.56 1443.46 226.9 ;
     RECT  1442.02 1593.38 1443.74 2310.94 ;
     RECT  997.82 586.64 1443.94 586.84 ;
     RECT  1442.98 3187.28 1443.94 3192.1 ;
     RECT  1443.74 1593.38 1444.7 2315.14 ;
     RECT  1350.82 2415.74 1444.9 2426.44 ;
     RECT  1440.265 1482.905 1447.715 1532.68 ;
     RECT  1447.715 1483.74 1448.165 1532.68 ;
     RECT  1379 3220 1449 3470 ;
     RECT  1444.7 1593.38 1449.02 2317.66 ;
     RECT  1420.9 3055.82 1449.5 3177.88 ;
     RECT  1443.94 3187.28 1450.18 3188.32 ;
     RECT  1425.5 1549.28 1450.46 1560.82 ;
     RECT  1419.46 2905.04 1450.46 3044.1 ;
     RECT  1443.46 219.56 1450.66 219.76 ;
     RECT  1444.9 2426.24 1450.66 2426.44 ;
     RECT  1448.165 1483.76 1452.1 1532.68 ;
     RECT  1306.34 716.42 1453.06 723.76 ;
     RECT  1450.46 2901.68 1453.06 3044.1 ;
     RECT  1449.02 1593.38 1453.34 2318.5 ;
     RECT  1389.02 2329.22 1453.34 2329.42 ;
     RECT  1444.9 2415.74 1453.54 2415.94 ;
     RECT  1450.46 1547.18 1453.76 1560.82 ;
     RECT  1450.18 3187.7 1453.82 3188.32 ;
     RECT  1453.76 1547.18 1454.3 1563.51 ;
     RECT  1452.1 1486.28 1454.78 1532.68 ;
     RECT  1449.5 3053.3 1457.38 3177.88 ;
     RECT  994.46 197.72 1457.86 197.92 ;
     RECT  1439.14 2345.18 1457.86 2352.1 ;
     RECT  1439.14 2362.82 1458.34 2372.26 ;
     RECT  1388.9 737.84 1459.78 738.04 ;
     RECT  1453.06 716.42 1460.74 716.62 ;
     RECT  1454.3 1547.18 1461.5 1569.22 ;
     RECT  1435.78 766.82 1463.62 769.54 ;
     RECT  1458.34 2365.76 1463.62 2372.26 ;
     RECT  1439 0 1464.1 183.64 ;
     RECT  1454.78 1486.28 1464.1 1533.52 ;
     RECT  1453.34 1593.38 1466.3 2329.42 ;
     RECT  1461.5 1543.82 1466.78 1569.64 ;
     RECT  1439.14 1578.26 1466.78 1581.82 ;
     RECT  1466.3 1593.38 1469.18 2330.26 ;
     RECT  1453.82 3187.7 1469.38 3192.1 ;
     RECT  1469.18 1593.38 1471.1 2330.68 ;
     RECT  1464.1 1486.7 1472.06 1533.52 ;
     RECT  1466.78 1543.82 1472.06 1581.82 ;
     RECT  1453.06 2905.04 1472.06 3044.1 ;
     RECT  1432.42 834.86 1472.26 842.2 ;
     RECT  1471.1 1593.38 1474.46 2331.94 ;
     RECT  1472.06 1486.7 1474.94 1581.82 ;
     RECT  1474.94 1486.7 1475.9 1583.08 ;
     RECT  1474.46 1593.38 1475.9 2333.62 ;
     RECT  1469.38 3187.7 1476.1 3188.32 ;
     RECT  1476.1 3187.7 1476.38 3187.9 ;
     RECT  1475.9 2726.96 1476.86 2727.16 ;
     RECT  1476.86 2726.96 1477.06 2741.44 ;
     RECT  1472.54 2685.8 1478.5 2693.14 ;
     RECT  1476.38 3187.28 1479.94 3187.9 ;
     RECT  1475.9 1474.94 1480.22 2334.46 ;
     RECT  1457.86 2345.18 1480.9 2345.38 ;
     RECT  1478.5 2692.94 1480.9 2693.14 ;
     RECT  1457.38 3055.82 1480.9 3177.88 ;
     RECT  1480.22 1472 1482.14 2334.46 ;
     RECT  1477.06 2733.68 1482.34 2741.44 ;
     RECT  1482.14 1471.58 1482.62 2334.46 ;
     RECT  1482.62 1471.58 1484.06 2339.08 ;
     RECT  1484.06 1463.6 1486.94 2339.08 ;
     RECT  1486.94 1463.18 1488.32 2339.08 ;
     RECT  1479.94 3187.7 1488.38 3187.9 ;
     RECT  1482.62 1445.54 1488.86 1445.74 ;
     RECT  1488.38 3187.28 1490.5 3187.9 ;
     RECT  1488.86 1440.92 1490.72 1445.74 ;
     RECT  1463.62 769.34 1491.46 769.54 ;
     RECT  1490.72 1440.92 1491.74 1445.775 ;
     RECT  1472.06 2904.2 1491.74 3044.1 ;
     RECT  1491.74 1440.92 1492.22 1446.16 ;
     RECT  1488.32 1460.49 1492.22 2339.08 ;
     RECT  1490.5 3187.7 1492.7 3187.9 ;
     RECT  1492.22 1440.92 1494.62 2339.08 ;
     RECT  1494.62 1440.5 1497.02 2339.08 ;
     RECT  1484.06 2348.12 1497.02 2348.32 ;
     RECT  1482.34 2738.72 1497.5 2738.92 ;
     RECT  1492.7 3187.7 1497.5 3192.1 ;
     RECT  1497.5 2738.72 1497.7 2739.34 ;
     RECT  1480.9 3056.66 1498.94 3177.88 ;
     RECT  1491.74 2900 1501.54 3044.1 ;
     RECT  1411.78 2380.88 1503.46 2381.08 ;
     RECT  1497.02 1440.5 1505.86 2348.32 ;
     RECT  1464.1 0 1506.14 180 ;
     RECT  1497.5 3187.7 1506.82 3193.36 ;
     RECT  1501.54 2904.2 1507.3 3044.1 ;
     RECT  1498.94 3056.24 1509.5 3177.88 ;
     RECT  1505.86 1440.5 1514.3 2339.08 ;
     RECT  1505.86 2348.12 1514.3 2348.32 ;
     RECT  1514.3 1440.5 1515.94 2348.32 ;
     RECT  1430.5 2474.12 1518.82 2474.32 ;
     RECT  1463.62 2372.06 1519.78 2372.26 ;
     RECT  1435.78 2451.44 1522.18 2451.64 ;
     RECT  1515.94 1440.5 1524.1 2339.08 ;
     RECT  1524.1 1440.5 1524.58 2334.46 ;
     RECT  1506.82 3187.7 1524.86 3187.9 ;
     RECT  1524.86 3187.28 1525.06 3187.9 ;
     RECT  1524.58 1440.5 1526.3 2333.62 ;
     RECT  1525.06 3187.28 1526.5 3187.48 ;
     RECT  1507.3 2904.62 1526.98 3044.1 ;
     RECT  1526.3 1440.08 1527.46 2333.62 ;
     RECT  1526.98 2905.04 1529.86 3044.1 ;
     RECT  1527.46 1440.08 1532.74 2330.68 ;
     RECT  1534.94 3191.9 1536.38 3192.1 ;
     RECT  1532.74 1440.08 1542.14 2329.42 ;
     RECT  1509.5 3055.82 1542.62 3177.88 ;
     RECT  1542.14 1437.98 1543.3 2329.42 ;
     RECT  1542.62 3055.4 1547.14 3177.88 ;
     RECT  1536.38 3187.7 1547.9 3192.1 ;
     RECT  1543.3 1437.98 1550.24 2318.5 ;
     RECT  1547.9 3187.7 1555.78 3193.36 ;
     RECT  1529.86 2906.3 1557.98 3044.1 ;
     RECT  1557.98 2905.88 1559.14 3044.1 ;
     RECT  1506.14 0 1559.42 183.64 ;
     RECT  1550.24 1437.81 1562.3 2318.5 ;
     RECT  1559.42 0 1563 184.06 ;
     RECT  1562.3 1433.78 1564.22 2318.5 ;
     RECT  1564.22 1433.36 1564.7 2318.5 ;
     RECT  1564.7 1432.52 1565.18 2318.5 ;
     RECT  1565.18 1430.42 1565.66 2318.5 ;
     RECT  1565.66 1425.8 1565.86 2318.5 ;
     RECT  1547.14 3055.82 1566.14 3177.88 ;
     RECT  1555.78 3187.7 1571.42 3192.1 ;
     RECT  1565.18 997.82 1572.86 998.02 ;
     RECT  1449 3220 1573 3400 ;
     RECT  1565.86 1425.8 1577.18 2313.88 ;
     RECT  1577.18 1424.12 1578.14 2313.88 ;
     RECT  1578.14 1423.28 1578.86 2313.88 ;
     RECT  1578.86 1422.02 1581.02 2313.88 ;
     RECT  1571.42 3187.28 1581.22 3192.1 ;
     RECT  1570.46 1328.36 1581.5 1328.56 ;
     RECT  1581.02 1417.82 1587.26 2313.88 ;
     RECT  1587.26 1415.72 1587.98 2313.88 ;
     RECT  1587.98 1414.46 1592.26 2313.88 ;
     RECT  1592.26 1414.46 1593.5 1609.96 ;
     RECT  1593.5 1410.68 1596.38 1609.96 ;
     RECT  1596.38 1408.16 1598.3 1609.96 ;
     RECT  1581.22 3187.7 1598.3 3192.1 ;
     RECT  1598.3 1407.74 1601.18 1609.96 ;
     RECT  1598.3 3187.7 1601.18 3193.36 ;
     RECT  1601.18 3187.28 1602.34 3193.36 ;
     RECT  1602.34 3187.28 1603.78 3192.1 ;
     RECT  1601.18 1404.38 1606.46 1609.96 ;
     RECT  1592.26 1618.58 1606.46 2313.88 ;
     RECT  1606.46 1404.38 1606.94 2313.88 ;
     RECT  1606.94 1401.02 1611.26 2313.88 ;
     RECT  1611.26 1396.82 1612.22 2313.88 ;
     RECT  1566.14 3055.4 1614.34 3177.88 ;
     RECT  1612.22 1395.56 1614.62 2313.88 ;
     RECT  1614.62 1393.88 1615.1 2313.88 ;
     RECT  1543.3 2329.22 1618.66 2329.42 ;
     RECT  1339.58 1342.64 1618.94 1342.84 ;
     RECT  1615.1 1393.46 1619.42 2313.88 ;
     RECT  1603.78 3187.7 1620.58 3192.1 ;
     RECT  1620.58 3191.9 1622.02 3192.1 ;
     RECT  1614.34 3055.82 1627.1 3177.88 ;
     RECT  1619.42 1388.84 1629.98 2313.88 ;
     RECT  1629.98 1386.32 1630.46 2313.88 ;
     RECT  1618.94 1342.64 1631.9 1349.98 ;
     RECT  1629.5 3187.28 1632.1 3187.48 ;
     RECT  1563 -70 1633 184.06 ;
     RECT  1630.46 1385.9 1633.34 2313.88 ;
     RECT  1633.34 1385.48 1637.66 2315.98 ;
     RECT  1637.66 1381.7 1639.1 2315.98 ;
     RECT  1639.1 1378.76 1640.54 2315.98 ;
     RECT  1640.54 1378.34 1642.46 2315.98 ;
     RECT  1573 3220 1643 3470 ;
     RECT  1625.66 1188.5 1645.82 1188.7 ;
     RECT  1581.5 1321.22 1647.74 1328.56 ;
     RECT  1631.9 1342.64 1647.74 1357.12 ;
     RECT  1642.46 1378.34 1648.7 2318.08 ;
     RECT  1497.7 2739.14 1648.7 2739.34 ;
     RECT  1644.86 3193.16 1648.7 3193.36 ;
     RECT  1648.7 2739.14 1648.9 2742.7 ;
     RECT  1648.7 3187.7 1648.9 3193.36 ;
     RECT  1648.7 1374.14 1650.34 2318.08 ;
     RECT  1650.34 1374.14 1654.66 2315.98 ;
     RECT  1648.9 3187.7 1654.94 3192.1 ;
     RECT  1654.66 1378.34 1658.02 2315.98 ;
     RECT  1654.94 3187.28 1658.02 3192.1 ;
     RECT  1559.14 2906.3 1660.22 3044.1 ;
     RECT  1515.94 2348.12 1661.86 2348.32 ;
     RECT  1658.02 1381.28 1662.34 2315.98 ;
     RECT  1662.34 1385.06 1662.62 2315.98 ;
     RECT  1660.22 2905.88 1663.3 3044.1 ;
     RECT  1658.02 3187.7 1666.66 3192.1 ;
     RECT  1627.1 3055.4 1667.48 3177.88 ;
     RECT  1663.3 2906.3 1667.62 3044.1 ;
     RECT  1662.62 1385.06 1669.54 2316.4 ;
     RECT  1630.46 609.74 1669.82 609.94 ;
     RECT  1669.54 1388 1672.22 2316.4 ;
     RECT  1666.66 3189.8 1672.7 3192.1 ;
     RECT  1672.22 1388 1672.9 2318.08 ;
     RECT  1672.7 3189.8 1674.14 3192.52 ;
     RECT  1672.9 1392.62 1674.62 2318.08 ;
     RECT  1674.62 1392.62 1675.78 2318.5 ;
     RECT  1675.78 1394.3 1677.5 2318.5 ;
     RECT  1667.62 2906.3 1677.5 2916.16 ;
     RECT  1667.62 2925.32 1677.5 3044.1 ;
     RECT  1677.5 1394.3 1677.98 2319.34 ;
     RECT  1674.14 3189.8 1678.94 3195.46 ;
     RECT  1677.98 1394.3 1679.9 2323.54 ;
     RECT  1679.9 1394.3 1680.1 2323.96 ;
     RECT  1680.1 1398.5 1681.82 2323.96 ;
     RECT  1667.48 3059.1 1682.3 3177.88 ;
     RECT  1681.82 1398.5 1684.7 2325.64 ;
     RECT  1678.94 3187.7 1685.86 3195.46 ;
     RECT  1685.86 3191.06 1686.14 3195.46 ;
     RECT  1684.7 1398.5 1687.3 2330.26 ;
     RECT  1682.3 3057.08 1687.58 3177.88 ;
     RECT  1648.9 2742.5 1688.54 2742.7 ;
     RECT  1677.5 2900 1689.02 3044.1 ;
     RECT  1687.3 1409 1690.94 2330.26 ;
     RECT  1688.54 2742.08 1690.94 2742.7 ;
     RECT  1686.14 3191.06 1693.34 3195.88 ;
     RECT  1690.94 1409 1693.82 2331.52 ;
     RECT  1687.58 3056.66 1694.78 3177.88 ;
     RECT  1689.02 2889.5 1694.98 3044.1 ;
     RECT  1690.94 2739.56 1695.26 2742.7 ;
     RECT  1695.26 2732 1698.14 2742.7 ;
     RECT  1693.34 3191.06 1698.14 3196.3 ;
     RECT  1694.78 3056.24 1698.62 3177.88 ;
     RECT  1698.14 3187.28 1699.3 3196.3 ;
     RECT  1698.14 2732 1700.06 2750.26 ;
     RECT  1698.62 3053.72 1700.54 3177.88 ;
     RECT  1699.3 3191.48 1700.74 3196.3 ;
     RECT  1700.74 3191.48 1701.22 3195.88 ;
     RECT  1700.06 2730.74 1702.66 2750.26 ;
     RECT  1702.825 2349.785 1702.895 2350.015 ;
     RECT  1656.38 800.42 1702.94 800.62 ;
     RECT  1430.5 812.18 1702.94 812.38 ;
     RECT  1693.82 1409 1703.42 2333.2 ;
     RECT  1700.54 3053.3 1703.9 3177.88 ;
     RECT  1702.66 2733.68 1704.1 2750.26 ;
     RECT  1687.3 1398.5 1704.38 1398.7 ;
     RECT  1703.42 1409 1704.38 2333.62 ;
     RECT  1704.38 1398.5 1704.86 2333.62 ;
     RECT  1702.895 2345.18 1704.86 2350.015 ;
     RECT  1694.98 2896.89 1706.005 3044.1 ;
     RECT  1704.86 1398.5 1706.5 2350.015 ;
     RECT  1704.1 2734.52 1706.98 2750.26 ;
     RECT  1706.005 2898.32 1706.98 3044.1 ;
     RECT  1706.98 2734.52 1708.42 2747.32 ;
     RECT  1706.98 2898.32 1709.38 2915.74 ;
     RECT  1706.5 1419.5 1710.275 2350.015 ;
     RECT  1710.275 1419.5 1710.725 2349.18 ;
     RECT  1703.9 3052.88 1711.3 3177.88 ;
     RECT  1710.725 1419.5 1711.78 2345.8 ;
     RECT  1708.42 2734.52 1713.98 2742.7 ;
     RECT  1713.98 2733.68 1714.18 2742.7 ;
     RECT  1711.78 1424.12 1714.66 2345.8 ;
     RECT  1714.18 2734.52 1715.14 2742.7 ;
     RECT  1701.22 3191.48 1715.14 3195.46 ;
     RECT  1715.14 3191.48 1715.42 3193.78 ;
     RECT  1709.38 2901.26 1716.04 2915.74 ;
     RECT  1706.98 2925.32 1716.04 3044.1 ;
     RECT  1715.42 3187.28 1718.02 3193.78 ;
     RECT  1714.66 1427.06 1718.5 2345.8 ;
     RECT  1718.5 1431.68 1719.26 2345.8 ;
     RECT  1718.02 3187.28 1719.46 3192.1 ;
     RECT  1715.14 2734.94 1720.42 2742.7 ;
     RECT  1716.04 2901.26 1720.9 3044.1 ;
     RECT  1711.3 3058.34 1720.9 3177.88 ;
     RECT  1719.26 1431.68 1721.38 2346.22 ;
     RECT  1721.38 1434.2 1723.58 2346.22 ;
     RECT  1719.46 3187.28 1723.78 3187.48 ;
     RECT  1723.58 1434.2 1725.22 2348.32 ;
     RECT  1725.22 1434.2 1727.14 2345.8 ;
     RECT  1715.9 1385.9 1727.9 1386.1 ;
     RECT  1706.5 1398.5 1727.9 1406.26 ;
     RECT  1720.9 2901.26 1727.9 2915.74 ;
     RECT  1727.14 1439.24 1728.1 2345.8 ;
     RECT  1728.1 1439.24 1728.58 1667.08 ;
     RECT  1728.58 1443.86 1730.98 1667.08 ;
     RECT  1727.9 2900.42 1732.22 2915.74 ;
     RECT  1720.9 2925.32 1732.22 3044.1 ;
     RECT  1720.9 3059.1 1732.36 3177.88 ;
     RECT  1728.1 1676.12 1735.3 2345.8 ;
     RECT  1735.3 1676.12 1737.7 2341.18 ;
     RECT  1737.7 1705.52 1739.14 2341.18 ;
     RECT  1727.9 1385.9 1739.9 1406.26 ;
     RECT  1731.26 3187.7 1740.86 3187.9 ;
     RECT  1739.14 1705.52 1741.06 2340.76 ;
     RECT  1730.98 1453.94 1741.34 1667.08 ;
     RECT  1737.7 1676.12 1741.34 1696.06 ;
     RECT  1741.06 1706.36 1742.02 2340.76 ;
     RECT  1740.86 3187.28 1742.3 3187.9 ;
     RECT  1739.9 1385.9 1742.78 1413.82 ;
     RECT  1742.02 1706.36 1742.98 2339.08 ;
     RECT  1742.98 1706.36 1743.46 2338.66 ;
     RECT  1742.3 3187.28 1743.94 3192.1 ;
     RECT  1720.42 2739.56 1745.86 2742.7 ;
     RECT  1743.46 1706.78 1746.34 2338.66 ;
     RECT  1746.34 1706.78 1748.74 2334.46 ;
     RECT  1732.36 3055.82 1756.22 3177.88 ;
     RECT  1633 0 1757 184.06 ;
     RECT  1743.94 3187.7 1757.86 3192.1 ;
     RECT  1741.34 1453.94 1758.62 1696.06 ;
     RECT  1748.74 1706.78 1758.62 2333.2 ;
     RECT  1730.98 1443.86 1762.94 1444.06 ;
     RECT  1758.62 1453.94 1762.94 2333.2 ;
     RECT  1756.22 3052.88 1766.02 3177.88 ;
     RECT  1762.94 1443.86 1766.98 2337.82 ;
     RECT  1643 3220 1767 3400 ;
     RECT  1766.02 3055.82 1768.9 3177.88 ;
     RECT  1766.98 1443.86 1769.86 2335.3 ;
     RECT  1769.86 1443.86 1771.035 2334.04 ;
     RECT  1771.035 1886.54 1771.78 2334.04 ;
     RECT  1771.035 1443.86 1772.74 1876.66 ;
     RECT  1772.74 1443.86 1773.22 1873.3 ;
     RECT  1771.78 1886.96 1773.22 2334.04 ;
     RECT  1757.86 3187.7 1773.98 3187.9 ;
     RECT  1773.98 3187.28 1774.18 3192.1 ;
     RECT  1773.22 1886.96 1775.14 2331.52 ;
     RECT  1775.14 1887.38 1777.06 2331.52 ;
     RECT  1768.9 3056.24 1777.34 3177.88 ;
     RECT  1776.86 1022.6 1777.54 1022.8 ;
     RECT  1774.18 3187.7 1778.02 3192.1 ;
     RECT  1777.06 1887.38 1778.5 2330.68 ;
     RECT  1778.5 1887.38 1778.98 2330.26 ;
     RECT  1778.98 1887.38 1780.42 2326.48 ;
     RECT  1725.02 1370.78 1781.18 1370.98 ;
     RECT  1742.78 1380.86 1781.18 1413.82 ;
     RECT  1780.42 1887.38 1781.38 2325.64 ;
     RECT  1773.5 1431.26 1782.14 1431.46 ;
     RECT  1773.22 1443.86 1783.1 1444.06 ;
     RECT  1782.14 1426.22 1783.58 1431.46 ;
     RECT  1783.1 1441.34 1783.58 1444.06 ;
     RECT  1781.38 1887.38 1783.78 2323.96 ;
     RECT  1783.78 1992.8 1784.26 2323.96 ;
     RECT  1783.78 1906.28 1784.74 1983.76 ;
     RECT  1773.22 1453.94 1785.02 1873.3 ;
     RECT  1783.78 1887.38 1785.02 1895.56 ;
     RECT  1785.02 1453.94 1785.7 1895.56 ;
     RECT  1784.26 1992.8 1785.7 2318.5 ;
     RECT  1783.58 1426.22 1785.98 1444.06 ;
     RECT  1785.7 1453.94 1785.98 1880.02 ;
     RECT  1784.74 1907.96 1786.18 1983.76 ;
     RECT  1781.18 1370.78 1786.46 1413.82 ;
     RECT  1785.98 1426.22 1786.46 1880.02 ;
     RECT  1785.7 1892.84 1786.66 1895.56 ;
     RECT  1786.18 1938.2 1786.66 1983.76 ;
     RECT  1786.18 1907.96 1787.14 1927.9 ;
     RECT  1786.66 1941.14 1787.14 1983.76 ;
     RECT  1785.7 2000.78 1787.14 2318.5 ;
     RECT  1787.14 2000.78 1787.38 2008.12 ;
     RECT  1778.02 3187.7 1787.42 3187.9 ;
     RECT  1787.14 1941.14 1787.62 1971.58 ;
     RECT  1786.66 1895.36 1788.1 1895.56 ;
     RECT  1787.62 1941.14 1788.1 1970.32 ;
     RECT  1787.38 2005.82 1788.1 2008.12 ;
     RECT  1787.14 2016.74 1788.1 2315.14 ;
     RECT  1787.14 1909.64 1788.58 1927.9 ;
     RECT  1788.1 1947.44 1788.58 1970.32 ;
     RECT  1472.26 842 1789.06 842.2 ;
     RECT  1788.58 1947.86 1789.06 1970.32 ;
     RECT  1702.94 800.42 1789.54 812.38 ;
     RECT  1789.06 1947.86 1789.54 1968.64 ;
     RECT  1788.1 2027.66 1789.54 2315.14 ;
     RECT  1788.58 1909.64 1790.98 1918.66 ;
     RECT  1789.54 1947.86 1790.98 1962.76 ;
     RECT  1789.54 2035.22 1790.98 2035.42 ;
     RECT  1790.98 1909.64 1791.46 1916.98 ;
     RECT  1788.58 1927.7 1791.94 1927.9 ;
     RECT  1790.98 1947.86 1791.94 1961.08 ;
     RECT  1789.54 2046.56 1791.94 2315.14 ;
     RECT  1791.94 2046.56 1792.9 2063.14 ;
     RECT  1786.46 1370.78 1793.38 1880.02 ;
     RECT  1791.94 1952.9 1793.38 1961.08 ;
     RECT  1792.9 2053.28 1793.38 2063.14 ;
     RECT  1791.94 2081.84 1793.38 2315.14 ;
     RECT  1793.38 1370.78 1793.86 1760.74 ;
     RECT  1793.38 1772.72 1793.86 1880.02 ;
     RECT  1793.38 2081.84 1793.86 2112.28 ;
     RECT  1793.38 2122.58 1793.86 2141.26 ;
     RECT  1793.38 2149.88 1793.86 2315.14 ;
     RECT  1793.86 2095.7 1794.34 2112.28 ;
     RECT  1793.86 2193.14 1794.34 2315.14 ;
     RECT  1793.86 1772.72 1795.3 1778.8 ;
     RECT  1793.86 1788.68 1795.3 1805.26 ;
     RECT  1793.86 1826.9 1795.3 1846.84 ;
     RECT  1794.34 2095.7 1795.3 2103.88 ;
     RECT  1793.86 2122.58 1795.3 2129.92 ;
     RECT  1787.42 3187.7 1795.58 3192.1 ;
     RECT  1795.58 3187.28 1796.74 3192.1 ;
     RECT  1793.86 1370.78 1797.5 1756.54 ;
     RECT  1795.3 1772.72 1798.18 1775.86 ;
     RECT  1793.38 1952.9 1798.18 1956.04 ;
     RECT  1793.38 2059.16 1798.18 2063.14 ;
     RECT  1795.3 2103.68 1798.18 2103.88 ;
     RECT  1795.3 2122.58 1798.18 2122.78 ;
     RECT  1794.34 2213.3 1798.18 2311.78 ;
     RECT  1795.3 1800.02 1798.66 1805.26 ;
     RECT  1798.18 2220.44 1798.66 2311.78 ;
     RECT  1794.34 2193.14 1799.62 2203 ;
     RECT  1791.46 1913.84 1799.9 1916.98 ;
     RECT  1796.74 3187.7 1799.9 3192.1 ;
     RECT  1797.5 1370.76 1800.1 1756.54 ;
     RECT  1798.66 1800.02 1800.1 1801.06 ;
     RECT  1793.86 1815.98 1800.1 1816.6 ;
     RECT  1798.18 1952.9 1800.1 1954.36 ;
     RECT  1647.74 1321.22 1800.58 1357.12 ;
     RECT  1798.66 2221.28 1800.72 2311.78 ;
     RECT  1798.18 1773.98 1801.54 1775.86 ;
     RECT  1800.72 2231.78 1801.54 2233.24 ;
     RECT  1800.1 1370.76 1803.46 1748.98 ;
     RECT  1803.46 1611.42 1803.94 1748.98 ;
     RECT  1793.86 1856.3 1803.94 1880.02 ;
     RECT  1800.72 2253.62 1804.7 2311.78 ;
     RECT  1803.94 1668.12 1804.9 1748.98 ;
     RECT  1799.9 3187.7 1804.9 3193.36 ;
     RECT  1803.94 1611.42 1807.3 1659.52 ;
     RECT  1804.9 1668.12 1807.3 1746.44 ;
     RECT  1799.9 1912.58 1815.94 1916.98 ;
     RECT  1804.9 3187.7 1819.1 3192.1 ;
     RECT  1819.1 3187.28 1820.74 3192.1 ;
     RECT  1799.62 2193.14 1825.06 2199.64 ;
     RECT  1820.74 3187.7 1825.82 3192.1 ;
     RECT  1795.3 1838.24 1826.02 1846.84 ;
     RECT  1757 -70 1827 184.06 ;
     RECT  1825.82 3187.7 1828.9 3192.52 ;
     RECT  1803.46 1558.5 1835.9 1600.28 ;
     RECT  1807.3 1721.04 1836.1 1746.44 ;
     RECT  1767 3220 1837 3470 ;
     RECT  1828.9 3187.7 1837.34 3192.1 ;
     RECT  1837.34 3187.28 1840.42 3192.1 ;
     RECT  1803.94 1856.3 1840.9 1879.6 ;
     RECT  1840.42 3187.7 1844.54 3192.1 ;
     RECT  1804.7 2253.62 1846.66 2314.72 ;
     RECT  1840.9 1868.9 1849.06 1879.6 ;
     RECT  1844.54 3187.7 1849.06 3192.52 ;
     RECT  1849.06 3187.7 1854.14 3192.1 ;
     RECT  1854.14 3187.28 1857.22 3192.1 ;
     RECT  1840.9 1856.3 1865.38 1857.76 ;
     RECT  1857.22 3187.7 1869.7 3192.1 ;
     RECT  1826.02 1838.24 1871.14 1846.42 ;
     RECT  1869.7 3191.9 1871.14 3192.1 ;
     RECT  1732.22 2900.42 1880.26 3044.1 ;
     RECT  1800.1 1815.98 1888.42 1816.18 ;
     RECT  1795.3 1826.9 1893.22 1827.1 ;
     RECT  1890.14 3187.7 1895.42 3187.9 ;
     RECT  1895.42 3187.28 1897.06 3187.9 ;
     RECT  1777.34 3055.82 1898.3 3177.88 ;
     RECT  1880.26 2906.72 1904.06 3044.1 ;
     RECT  1897.06 3187.7 1905.02 3187.9 ;
     RECT  1846.66 2261.6 1907.62 2314.72 ;
     RECT  1898.3 3055.4 1908.58 3177.88 ;
     RECT  1801.54 1775.66 1911.46 1775.86 ;
     RECT  1905.02 3187.7 1913.86 3192.1 ;
     RECT  1825.06 2193.14 1915.78 2199.22 ;
     RECT  1904.06 2904.62 1917.7 3044.1 ;
     RECT  1913.86 3187.7 1920.86 3187.9 ;
     RECT  1920.86 3187.28 1921.06 3187.9 ;
     RECT  1921.06 3187.28 1922.02 3187.48 ;
     RECT  1917.7 2907.14 1922.5 3044.1 ;
     RECT  1908.58 3056.66 1923.26 3177.88 ;
     RECT  1871.14 1838.66 1923.46 1846.42 ;
     RECT  1849.06 1871.84 1938.34 1879.6 ;
     RECT  1923.26 3055.4 1943.14 3177.88 ;
     RECT  1940.06 3188.54 1943.42 3188.74 ;
     RECT  1922.5 2907.56 1946.78 3044.1 ;
     RECT  1943.42 3188.54 1950.62 3192.1 ;
     RECT  1827 0 1951 184.06 ;
     RECT  1950.62 3187.7 1951.1 3192.1 ;
     RECT  1946.78 2907.56 1953.98 3046.36 ;
     RECT  1953.98 2905.88 1954.94 3046.36 ;
     RECT  1954.94 2904.62 1957.82 3046.36 ;
     RECT  1943.14 3056.24 1957.82 3177.88 ;
     RECT  1951.1 3187.7 1958.3 3193.36 ;
     RECT  1865.38 1856.3 1958.98 1856.5 ;
     RECT  1837 3220 1961 3400 ;
     RECT  1951 -70 1962.34 184.06 ;
     RECT  1958.3 3187.7 1964.74 3195.04 ;
     RECT  1957.82 2904.62 1969.54 3177.88 ;
     RECT  1964.74 3187.7 1970.3 3193.36 ;
     RECT  1970.3 3187.28 1970.5 3193.36 ;
     RECT  1907.62 2292.26 1970.98 2314.72 ;
     RECT  1970.5 3187.28 1971.94 3192.1 ;
     RECT  1971.94 3187.28 1974.34 3187.48 ;
     RECT  1800.72 2221.28 1976.26 2221.9 ;
     RECT  1969.54 2905.88 1976.74 3177.88 ;
     RECT  1938.34 1872.26 1977.7 1879.6 ;
     RECT  1976.26 2221.7 1988.26 2221.9 ;
     RECT  1970.98 2301.5 2008.9 2314.72 ;
     RECT  1976.74 2907.56 2009.38 3177.88 ;
     RECT  1962.34 -70 2021 183.64 ;
     RECT  1798.18 2062.94 2028.58 2063.14 ;
     RECT  2009.38 2907.98 2030.3 3177.88 ;
     RECT  1915.78 2193.14 2030.5 2198.8 ;
     RECT  1961 3220 2031 3470 ;
     RECT  2030.3 2907.56 2040.86 3177.88 ;
     RECT  1800.1 1800.86 2041.06 1801.06 ;
     RECT  1815.94 1912.58 2051.14 1915.72 ;
     RECT  2030.5 2198.6 2051.62 2198.8 ;
     RECT  2051.14 1915.52 2066.98 1915.72 ;
     RECT  2062.46 1792.88 2078.02 1793.08 ;
     RECT  2008.9 2306.54 2079.94 2314.72 ;
     RECT  2040.86 2905.04 2089.06 3177.88 ;
     RECT  2089.06 2915.54 2092.16 3177.88 ;
     RECT  1923.46 1846.22 2092.9 1846.42 ;
     RECT  2092.16 2915.54 2093.38 2936.32 ;
     RECT  2048.06 1781.96 2098.66 1782.16 ;
     RECT  2093.38 2916.38 2099.14 2936.32 ;
     RECT  2099.14 2916.38 2099.62 2924.56 ;
     RECT  2092.16 2944.94 2099.62 2945.14 ;
     RECT  2092.16 3040.7 2099.62 3078.7 ;
     RECT  1810.94 1926.02 2100.1 1926.22 ;
     RECT  2089.06 2905.04 2101.54 2905.24 ;
     RECT  2092.16 3021.38 2105.66 3021.58 ;
     RECT  2099.62 2916.38 2105.86 2916.58 ;
     RECT  2105.66 3020.96 2106.14 3021.58 ;
     RECT  1800.1 1954.16 2106.82 1954.36 ;
     RECT  1977.7 1879.4 2107.3 1879.6 ;
     RECT  2106.14 3018.02 2108.54 3021.58 ;
     RECT  1745.86 2739.56 2109.22 2739.76 ;
     RECT  2108.54 3018.02 2109.22 3022 ;
     RECT  2099.62 3041.12 2109.22 3074.92 ;
     RECT  2077.82 1801.7 2109.5 1801.9 ;
     RECT  2109.5 1801.7 2109.7 1807.36 ;
     RECT  2109.22 3045.32 2110.66 3074.92 ;
     RECT  2099.14 2936.12 2111.14 2936.32 ;
     RECT  2110.66 3049.1 2112.58 3074.92 ;
     RECT  2112.58 3049.1 2115.46 3074.5 ;
     RECT  2115.46 3050.78 2115.94 3074.5 ;
     RECT  2115.94 3051.2 2116.9 3074.5 ;
     RECT  2098.46 1825.22 2117.18 1825.42 ;
     RECT  2109.7 1807.16 2117.38 1807.36 ;
     RECT  1836.1 1721.04 2118.14 1745.6 ;
     RECT  2116.9 3051.2 2118.34 3074.08 ;
     RECT  2117.18 1817.66 2120.26 1825.42 ;
     RECT  2118.34 3051.2 2121.7 3064.84 ;
     RECT  2109.22 3018.02 2122.46 3021.16 ;
     RECT  2121.7 3055.82 2122.66 3064.84 ;
     RECT  2122.66 3055.82 2124.1 3060.22 ;
     RECT  2122.46 3018.02 2126.02 3022 ;
     RECT  2124.1 3055.82 2128.42 3057.28 ;
     RECT  2126.02 3018.02 2129.38 3018.22 ;
     RECT  2128.42 3055.82 2129.86 3056.02 ;
     RECT  2118.14 1721.04 2134.18 1746.04 ;
     RECT  2021 0 2145 183.64 ;
     RECT  2031 3220 2155 3400 ;
     RECT  2145 -70 2156.26 183.64 ;
     RECT  2133.98 1756.34 2160.1 1756.54 ;
     RECT  2120.26 1817.66 2181.5 1817.86 ;
     RECT  2159.9 1778.6 2181.7 1778.8 ;
     RECT  2181.5 1817.66 2181.7 1826.26 ;
     RECT  2120.06 1954.58 2192.26 1954.78 ;
     RECT  2181.7 1826.06 2203.3 1826.26 ;
     RECT  2203.58 1860.5 2213.86 1860.7 ;
     RECT  2156.26 -70 2215 180 ;
     RECT  2213.66 1912.58 2224.9 1912.78 ;
     RECT  2155 3220 2225 3470 ;
     RECT  2224.7 1926.02 2232.1 1926.22 ;
     RECT  2192.06 2027.24 2235.46 2027.44 ;
     RECT  2231.9 1944.08 2249.86 1944.28 ;
     RECT  2235.26 2238.92 2253.22 2239.12 ;
     RECT  2181.5 1796.24 2257.06 1796.44 ;
     RECT  2249.66 2021.36 2260.9 2021.56 ;
     RECT  2256.86 1843.28 2264.26 1843.48 ;
     RECT  2264.06 1886.54 2271.46 1886.74 ;
     RECT  1807.3 1645.44 2282.5 1659.52 ;
     RECT  2271.26 1929.8 2282.5 1930 ;
     RECT  2260.7 2057.9 2282.5 2058.1 ;
     RECT  2282.3 1965.5 2293.06 1965.7 ;
     RECT  2292.86 2020.52 2304.1 2020.72 ;
     RECT  1803.46 1370.76 2314.94 1479.32 ;
     RECT  1803.46 1489.2 2314.94 1548.62 ;
     RECT  2282.3 2077.22 2325.22 2077.42 ;
     RECT  2304.38 2037.74 2329.06 2037.94 ;
     RECT  2325.02 2109.14 2332.7 2109.34 ;
     RECT  2332.7 2109.14 2332.9 2109.76 ;
     RECT  2334.62 1904.58 2335.1 1913.18 ;
     RECT  2334.62 1928.52 2335.1 1928.72 ;
     RECT  2334.62 1892.82 2335.58 1893.02 ;
     RECT  2335.1 1904.58 2335.58 1928.72 ;
     RECT  2335.58 1892.82 2337.02 1928.72 ;
     RECT  2337.02 1886.94 2337.98 1928.72 ;
     RECT  2215 0 2339 180 ;
     RECT  2282.5 1645.44 2340.1 1653.2 ;
     RECT  1807.3 1668.12 2340.1 1683.44 ;
     RECT  2134.18 1721.04 2340.1 1745.6 ;
     RECT  2337.98 1879.8 2340.38 1928.72 ;
     RECT  2340.38 1945.74 2340.86 1947.2 ;
     RECT  2340.38 1965.48 2340.86 1965.68 ;
     RECT  2340.38 1856.7 2341.34 1863.62 ;
     RECT  2340.38 1878.96 2341.34 1935.86 ;
     RECT  2340.86 1945.74 2341.34 1955.18 ;
     RECT  2340.86 1965.48 2341.34 1966.52 ;
     RECT  2341.34 1856.7 2342.24 1866.98 ;
     RECT  2328.86 2144.42 2343.74 2144.62 ;
     RECT  2343.26 1822.26 2345.12 1830.44 ;
     RECT  2345.12 1822.225 2346.14 1830.44 ;
     RECT  2346.14 1821.84 2347.1 1830.44 ;
     RECT  2342.24 1856.7 2347.1 1867.99 ;
     RECT  2343.74 2139.36 2347.1 2144.62 ;
     RECT  2343.26 2174.66 2347.1 2174.86 ;
     RECT  2314.94 1370.76 2347.3 1548.62 ;
     RECT  2347.1 1821.84 2347.58 1833.8 ;
     RECT  2347.1 1849.56 2347.58 1867.99 ;
     RECT  2332.9 2109.56 2347.58 2109.76 ;
     RECT  2347.1 2138.52 2347.58 2144.62 ;
     RECT  2347.1 2174.66 2348.06 2181.56 ;
     RECT  2341.34 1878.96 2348.54 1966.52 ;
     RECT  2343.74 2080.14 2348.54 2086.64 ;
     RECT  2347.58 2101.56 2348.54 2109.76 ;
     RECT  2347.58 2130.54 2348.54 2144.62 ;
     RECT  2225 3220 2349 3400 ;
     RECT  2348.54 1878.96 2349.02 1969.46 ;
     RECT  2348.06 2174.66 2349.02 2184.94 ;
     RECT  2347.58 1821.84 2349.5 1867.99 ;
     RECT  2348.54 2064.18 2349.5 2064.38 ;
     RECT  2348.54 2074.26 2349.5 2086.64 ;
     RECT  2349.5 1821.84 2349.98 1868.66 ;
     RECT  2349.02 1878.96 2349.98 1969.88 ;
     RECT  2349.5 2064.18 2349.98 2086.64 ;
     RECT  2348.54 2101.56 2349.98 2144.62 ;
     RECT  2349.98 2101.14 2350.46 2163.08 ;
     RECT  2349.98 2059.56 2350.88 2086.64 ;
     RECT  2349.02 2174.22 2350.94 2184.94 ;
     RECT  2350.88 2059.56 2351.42 2090.455 ;
     RECT  2349.98 1821.84 2351.9 1969.88 ;
     RECT  2339 -70 2352.38 180 ;
     RECT  2352.38 -70 2352.58 180.7 ;
     RECT  1800.58 1321.22 2352.58 1335.7 ;
     RECT  2351.42 2059.56 2352.86 2090.84 ;
     RECT  2350.46 2100.72 2352.86 2163.08 ;
     RECT  2352.86 2059.56 2354.78 2163.08 ;
     RECT  2350.94 2172.54 2354.78 2184.94 ;
     RECT  2351.9 1814.28 2355.16 1969.88 ;
     RECT  2355.16 1814.28 2355.5 1969.89 ;
     RECT  2355.5 1813.44 2355.74 1969.89 ;
     RECT  2354.78 1980.6 2355.74 1982.48 ;
     RECT  2352.58 1321.22 2355.94 1321.42 ;
     RECT  2355.74 1811.34 2356.22 1982.48 ;
     RECT  2356.22 1811.34 2356.7 1986.68 ;
     RECT  2356.7 1811.34 2357.12 1987.52 ;
     RECT  2357.66 2019.66 2358.14 2025.74 ;
     RECT  2354.78 2059.56 2358.325 2184.94 ;
     RECT  2358.14 2012.1 2358.62 2025.74 ;
     RECT  2358.325 2097.78 2358.62 2184.94 ;
     RECT  2349.5 2196.08 2358.62 2196.28 ;
     RECT  2358.62 2044.02 2359.1 2048.42 ;
     RECT  2358.325 2059.56 2359.1 2086.64 ;
     RECT  2358.62 2004.54 2359.52 2025.74 ;
     RECT  2359.52 2004.54 2360.54 2026.75 ;
     RECT  2360.54 2002.02 2361.02 2026.75 ;
     RECT  2361.02 1999.5 2361.5 2026.75 ;
     RECT  2358.62 2097.78 2361.5 2196.28 ;
     RECT  2357.12 1810.33 2362.46 1987.52 ;
     RECT  2361.5 2097.78 2362.46 2204.66 ;
     RECT  2354.78 2214.96 2362.46 2215.16 ;
     RECT  2362.46 1810.33 2362.94 1988.36 ;
     RECT  2361.5 1998.24 2362.94 2026.75 ;
     RECT  2362.94 1998.24 2363.9 2029.1 ;
     RECT  2362.46 2097.78 2364.38 2218.1 ;
     RECT  2363.42 2226.72 2364.38 2226.92 ;
     RECT  2363.9 1998.24 2365.34 2030.36 ;
     RECT  2364.38 2097.78 2365.82 2226.92 ;
     RECT  2365.34 1998.24 2366.3 2032.88 ;
     RECT  2365.82 2097.78 2366.78 2234.06 ;
     RECT  2362.46 2248.14 2366.78 2248.34 ;
     RECT  2362.94 1810.33 2368.7 1989.62 ;
     RECT  2366.3 1998.24 2368.7 2033.3 ;
     RECT  2368.7 1810.33 2369.66 2034.14 ;
     RECT  2359.1 2044.02 2369.66 2086.64 ;
     RECT  2366.78 2097.78 2370.14 2248.34 ;
     RECT  2369.66 1807.14 2370.56 2086.64 ;
     RECT  2370.56 1802.77 2370.62 2086.64 ;
     RECT  2370.14 2097.78 2371.58 2250.46 ;
     RECT  2370.62 1802.77 2372.06 2087.06 ;
     RECT  2372.06 1802.77 2373.02 2087.48 ;
     RECT  2371.58 2097.36 2373.02 2250.46 ;
     RECT  2373.02 1802.77 2378.005 2250.46 ;
     RECT  2378.005 1802.94 2387.42 2250.46 ;
     RECT  1907.62 2261.6 2387.42 2283.22 ;
     RECT  2387.42 1802.94 2392.22 2283.22 ;
     RECT  2392.22 1800.42 2393.18 2283.22 ;
     RECT  2352.58 -70 2393.9 180 ;
     RECT  2393.9 -70 2394.34 180.7 ;
     RECT  2393.18 1799.16 2400.38 2283.22 ;
     RECT  1970.98 2292.26 2400.38 2292.46 ;
     RECT  2400.38 1799.16 2401.82 2292.46 ;
     RECT  2401.82 1796.22 2402.02 2292.46 ;
     RECT  2402.02 1796.22 2403.46 1796.42 ;
     RECT  2079.94 2311.58 2404.42 2314.72 ;
     RECT  2340.1 1723.56 2404.62 1745.6 ;
     RECT  2404.22 1776.48 2404.7 1776.68 ;
     RECT  2404.62 1723.56 2405.395 1753.58 ;
     RECT  2402.78 1762.62 2405.395 1765.76 ;
     RECT  2405.395 1723.56 2405.66 1765.76 ;
     RECT  2404.7 1776.48 2405.66 1777.52 ;
     RECT  1807.3 1611.42 2406.34 1635.56 ;
     RECT  2340.1 1668.54 2407.78 1683.44 ;
     RECT  2394.34 -70 2409 180 ;
     RECT  2405.66 1723.56 2409.02 1777.52 ;
     RECT  2409.02 1723.56 2409.5 1781.3 ;
     RECT  2409.5 1723.56 2411.9 1781.72 ;
     RECT  2405.18 1795.8 2411.9 1796 ;
     RECT  2411.9 1723.56 2412.38 1796 ;
     RECT  2402.02 1806.3 2412.38 2283.22 ;
     RECT  2347.3 1489.2 2415.94 1548.62 ;
     RECT  2349 3220 2419 3470 ;
     RECT  2407.78 1668.54 2419.1 1668.74 ;
     RECT  2419.1 1668.54 2419.3 1669.16 ;
     RECT  2406.34 1611.42 2420.06 1635.14 ;
     RECT  2340.1 1645.44 2420.06 1652.78 ;
     RECT  2420.06 1611.42 2420.54 1652.78 ;
     RECT  1835.9 1558.5 2420.74 1600.7 ;
     RECT  2419.3 1668.96 2421.5 1669.16 ;
     RECT  2407.78 1683.24 2421.5 1683.44 ;
     RECT  2415.94 1489.2 2421.7 1507.04 ;
     RECT  1807.3 1695.84 2422.46 1711.16 ;
     RECT  2412.38 1723.56 2422.46 2283.22 ;
     RECT  2422.46 1695.84 2423.9 2283.22 ;
     RECT  2421.5 1668.96 2424.86 1683.44 ;
     RECT  2423.9 1693.32 2424.86 2283.22 ;
     RECT  2420.54 1611.42 2434.94 1659.92 ;
     RECT  2424.86 1668.96 2434.94 2283.22 ;
     RECT  2420.74 1590 2439.94 1600.7 ;
     RECT  2347.3 1370.76 2444.26 1479.32 ;
     RECT  2439.94 1590 2452.9 1590.2 ;
     RECT  2415.94 1516.92 2460.1 1548.62 ;
     RECT  2460.1 1516.92 2461.54 1534.76 ;
     RECT  2434.94 1611.42 2462.98 2283.22 ;
     RECT  2462.98 1624.44 2464.9 2283.22 ;
     RECT  2461.54 1519.44 2466.82 1534.76 ;
     RECT  2464.9 1624.44 2468.26 2250.44 ;
     RECT  2468.26 1624.44 2471.14 2249.18 ;
     RECT  2471.14 1625.28 2472.1 2249.18 ;
     RECT  2466.82 1519.44 2477.86 1532.24 ;
     RECT  2444.26 1436.28 2482.18 1479.32 ;
     RECT  2462.98 1611.42 2487.94 1612.88 ;
     RECT  2444.26 1370.76 2489.86 1423.88 ;
     RECT  2489.86 1370.76 2491.78 1406.24 ;
     RECT  2421.7 1489.2 2492.74 1494.44 ;
     RECT  2472.1 1625.28 2493.22 2248.76 ;
     RECT  2493.22 1625.28 2493.7 2237.42 ;
     RECT  2477.86 1522.8 2496.58 1532.24 ;
     RECT  2493.7 1625.28 2502.62 2234.48 ;
     RECT  2493.22 2248.56 2502.82 2248.76 ;
     RECT  2502.62 1625.28 2507.42 2235.32 ;
     RECT  2496.58 1522.8 2508.38 1529.72 ;
     RECT  2507.42 1625.28 2512.7 2237 ;
     RECT  2512.7 1625.28 2520.38 2242.04 ;
     RECT  2520.38 1625.28 2522.78 2242.46 ;
     RECT  2482.18 1441.32 2525.86 1479.32 ;
     RECT  2508.38 1520.72 2530.46 1529.72 ;
     RECT  2460.1 1543.8 2530.46 1548.62 ;
     RECT  2409 0 2533 180 ;
     RECT  2522.78 1625.28 2533.82 2242.88 ;
     RECT  2489.86 1416.12 2534.3 1423.88 ;
     RECT  2533.82 1621.08 2539.945 2242.88 ;
     RECT  2525.86 1474.08 2541.22 1479.32 ;
     RECT  2420.74 1558.5 2541.5 1581.38 ;
     RECT  2530.46 1520.72 2541.7 1548.62 ;
     RECT  2541.02 1590.42 2541.7 1590.62 ;
     RECT  2487.94 1611.42 2542.825 1611.62 ;
     RECT  2539.945 1621.065 2542.825 2242.88 ;
     RECT  2419 3220 2543 3400 ;
     RECT  1800.58 1349.78 2546.98 1357.12 ;
     RECT  2533 -70 2549.42 180 ;
     RECT  2549.42 -70 2549.86 180.7 ;
     RECT  2542.825 1611.42 2550.08 2242.88 ;
     RECT  2492.74 1491.72 2552.06 1494.44 ;
     RECT  2550.08 1611.42 2552.54 2245.99 ;
     RECT  2552.54 1611.42 2553.7 2249.6 ;
     RECT  2541.22 1476.6 2554.66 1479.32 ;
     RECT  2541.7 1520.72 2555.62 1530.16 ;
     RECT  2421.7 1506.84 2555.9 1507.04 ;
     RECT  2555.62 1520.72 2555.9 1529.72 ;
     RECT  2554.66 1479.12 2560.42 1479.32 ;
     RECT  2553.7 1621.92 2567.14 2249.6 ;
     RECT  2567.14 1621.92 2567.65 2249.215 ;
     RECT  2555.9 1506.84 2568.38 1529.72 ;
     RECT  2567.65 1621.92 2579.14 2249.18 ;
     RECT  2579.14 1643.745 2580.035 2249.18 ;
     RECT  2580.035 1644.58 2580.485 2249.18 ;
     RECT  2580.485 1645.44 2580.86 2249.18 ;
     RECT  2579.14 1621.92 2581.06 1635.14 ;
     RECT  2580.86 1645.44 2583.26 2252.96 ;
     RECT  2464.9 2261.6 2583.26 2283.22 ;
     RECT  2568.38 1506.84 2584.9 1531.42 ;
     RECT  2583.26 1645.44 2585.86 2283.22 ;
     RECT  2585.86 1645.44 2587.78 2249.18 ;
     RECT  2552.06 1491.72 2588.06 1494.88 ;
     RECT  2584.9 1506.84 2588.26 1529.72 ;
     RECT  2587.78 1645.86 2590.18 2249.18 ;
     RECT  2590.18 1660.56 2591.605 2249.18 ;
     RECT  2588.06 1490.48 2591.9 1494.88 ;
     RECT  2591.605 1660.56 2594.02 2248.34 ;
     RECT  2594.02 1663.08 2594.5 2248.34 ;
     RECT  2581.06 1629.9 2598.505 1635.14 ;
     RECT  2594.5 1663.5 2600.06 2248.34 ;
     RECT  2600.06 1663.5 2600.74 2249.6 ;
     RECT  2590.18 1645.86 2601.02 1647.74 ;
     RECT  2600.74 1664.34 2601.22 2249.215 ;
     RECT  2601.22 1668.12 2601.25 2249.215 ;
     RECT  2601.02 1645.86 2601.7 1649.42 ;
     RECT  2439.94 1600.5 2602.46 1600.7 ;
     RECT  2525.86 1441.32 2602.66 1464.2 ;
     RECT  2549.86 -70 2603 180 ;
     RECT  2601.7 1645.86 2603.14 1648.16 ;
     RECT  2601.25 1668.12 2604.1 2249.18 ;
     RECT  2598.505 1628.625 2605.955 1635.14 ;
     RECT  2604.1 1669.8 2606.02 2249.18 ;
     RECT  2603.14 1645.86 2606.3 1647.74 ;
     RECT  2605.955 1629.46 2606.405 1635.14 ;
     RECT  2606.3 1644.18 2606.5 1647.74 ;
     RECT  2602.46 1592.52 2608.7 1600.7 ;
     RECT  2553.7 1611.42 2608.7 1611.62 ;
     RECT  2606.405 1629.48 2610.34 1635.14 ;
     RECT  2608.7 1592.52 2610.62 1611.62 ;
     RECT  2610.34 1630.32 2610.62 1635.14 ;
     RECT  2606.5 1644.18 2610.62 1646.06 ;
     RECT  2610.62 1630.32 2610.82 1646.06 ;
     RECT  2606.02 1669.8 2610.82 2047.16 ;
     RECT  2610.62 1591.68 2611.3 1611.62 ;
     RECT  2602.66 1458.96 2611.58 1464.2 ;
     RECT  2591.9 1490.06 2612.54 1494.88 ;
     RECT  2612.54 1483.34 2612.74 1494.88 ;
     RECT  2543 3220 2613 3470 ;
     RECT  2606.02 2055.78 2613.02 2249.18 ;
     RECT  2602.66 1441.32 2613.5 1449.08 ;
     RECT  2611.58 1458.96 2613.5 1469.26 ;
     RECT  2610.82 1644.18 2614.18 1646.06 ;
     RECT  2610.82 1670.64 2614.46 2047.16 ;
     RECT  2613.02 2055.78 2614.46 2249.6 ;
     RECT  2614.46 1670.64 2615.42 2249.6 ;
     RECT  2615.42 1670.64 2617.06 2250.02 ;
     RECT  2617.06 1670.64 2619.94 2244.98 ;
     RECT  2588.26 1506.84 2620.7 1507.04 ;
     RECT  2541.7 1543.8 2620.7 1548.62 ;
     RECT  2541.5 1558.5 2620.7 1581.8 ;
     RECT  2614.18 1645.86 2620.7 1646.06 ;
     RECT  2612.74 1483.34 2620.9 1494.44 ;
     RECT  2620.7 1506.42 2620.9 1507.04 ;
     RECT  2588.26 1521.98 2620.9 1529.72 ;
     RECT  2611.3 1597.14 2620.9 1611.62 ;
     RECT  2613.5 1441.32 2621.18 1469.26 ;
     RECT  2620.9 1483.34 2621.18 1494.02 ;
     RECT  2620.9 1521.98 2624.74 1528.04 ;
     RECT  2619.94 1675.26 2627.14 2244.98 ;
     RECT  2620.7 1645.86 2627.9 1646.9 ;
     RECT  2621.18 1441.32 2628.1 1494.02 ;
     RECT  2627.9 1643.76 2628.38 1652.78 ;
     RECT  2627.14 1675.26 2629.34 2234.49 ;
     RECT  2610.82 1630.32 2630.3 1635.14 ;
     RECT  2628.38 1643.76 2630.3 1656.98 ;
     RECT  2620.9 1597.14 2630.78 1609.52 ;
     RECT  2630.78 1597.14 2631.26 1618.76 ;
     RECT  2630.3 1629.9 2631.26 1656.98 ;
     RECT  2620.7 1543.8 2637.02 1581.8 ;
     RECT  2620.9 1506.42 2637.5 1506.62 ;
     RECT  2637.02 1543.8 2637.5 1583.48 ;
     RECT  2534.3 1416.12 2638.46 1429.36 ;
     RECT  2628.1 1441.32 2638.46 1478.08 ;
     RECT  2637.5 1543.8 2638.94 1584.32 ;
     RECT  2631.26 1597.14 2638.94 1656.98 ;
     RECT  2637.5 1506.42 2639.42 1512.08 ;
     RECT  2629.34 1674.42 2640.005 2234.49 ;
     RECT  2638.46 1416.12 2640.1 1478.08 ;
     RECT  2638.94 1543.8 2640.265 1659.92 ;
     RECT  2640.005 1674.42 2640.565 2231.12 ;
     RECT  2628.1 1491.72 2640.86 1494.02 ;
     RECT  2639.42 1504.74 2640.86 1512.08 ;
     RECT  2624.74 1522.8 2640.86 1528.04 ;
     RECT  2640.265 1543.8 2640.86 1660.34 ;
     RECT  2640.86 1543.8 2641.34 1661.18 ;
     RECT  2640.565 1674.42 2641.34 1727.12 ;
     RECT  2640.1 1445.1 2641.82 1478.08 ;
     RECT  2640.86 1487.94 2641.82 1494.02 ;
     RECT  2641.82 1445.1 2642.3 1494.02 ;
     RECT  2640.86 1504.74 2642.3 1528.04 ;
     RECT  2640.1 1416.12 2642.5 1433.14 ;
     RECT  2642.3 1445.1 2642.5 1528.04 ;
     RECT  2640.565 1735.74 2642.5 2231.12 ;
     RECT  2641.34 1543.8 2646.06 1727.12 ;
     RECT  2646.06 1539.18 2646.835 1727.12 ;
     RECT  2642.5 1445.52 2647.58 1528.04 ;
     RECT  2646.835 1538.34 2647.58 1727.12 ;
     RECT  2647.58 1445.52 2649.7 1727.12 ;
     RECT  2649.7 1474.08 2650.46 1727.12 ;
     RECT  2642.5 1735.74 2650.46 2230.28 ;
     RECT  2642.5 1432.94 2652.86 1433.14 ;
     RECT  2650.46 1474.08 2655.2 2230.28 ;
     RECT  2652.86 1432.52 2656.42 1433.14 ;
     RECT  2655.2 1474.08 2657.18 2230.87 ;
     RECT  2649.7 1445.52 2657.86 1464.2 ;
     RECT  2657.18 1474.08 2657.86 2234.48 ;
     RECT  2657.86 1445.52 2658.34 1449.08 ;
     RECT  2657.86 1474.08 2658.37 2234.095 ;
     RECT  2657.86 1458.96 2658.62 1464.2 ;
     RECT  2658.37 1474.08 2658.62 2234.06 ;
     RECT  2658.62 1458.96 2665.525 2234.06 ;
     RECT  2656.42 1432.52 2666.5 1432.72 ;
     RECT  2665.525 1458.96 2668.7 2229.86 ;
     RECT  2658.34 1445.52 2672.06 1446.56 ;
     RECT  2668.7 1456.02 2672.06 2229.86 ;
     RECT  2672.06 1444.26 2673.92 2229.86 ;
     RECT  2673.92 1444.225 2674.94 2229.86 ;
     RECT  2491.78 1370.76 2677.82 1401.2 ;
     RECT  2642.5 1416.12 2677.82 1423.88 ;
     RECT  2674.94 1443.84 2677.82 2229.86 ;
     RECT  2677.82 1443.84 2681.66 2231.12 ;
     RECT  2681.66 1436.28 2681.86 2231.12 ;
     RECT  2681.86 1436.28 2683.1 2230.7 ;
     RECT  2683.1 1435.86 2683.98 2230.7 ;
     RECT  2683.98 1433.34 2684.755 2230.7 ;
     RECT  2677.82 1370.76 2685.98 1423.88 ;
     RECT  2684.755 1432.5 2685.98 2230.7 ;
     RECT  2685.98 1370.76 2693.86 2230.7 ;
     RECT  2693.86 1380.84 2700.1 2230.7 ;
     RECT  2700.1 1418.64 2701.54 2230.7 ;
     RECT  2700.1 1380.84 2705.86 1407.52 ;
     RECT  2701.54 1422.84 2714.78 2230.7 ;
     RECT  2714.78 1421.16 2721.7 2230.7 ;
     RECT  2721.7 1421.545 2721.92 2230.7 ;
     RECT  2705.86 1380.84 2724.1 1388.6 ;
     RECT  2721.92 1421.545 2726.05 2230.87 ;
     RECT  2603 0 2727 180 ;
     RECT  2705.86 1398.48 2728.7 1407.52 ;
     RECT  2726.05 1421.58 2735.62 2230.87 ;
     RECT  2728.7 1393.04 2735.9 1407.52 ;
     RECT  2735.62 1421.58 2735.9 1993.4 ;
     RECT  2735.62 2003.7 2736.38 2230.87 ;
     RECT  2613 3220 2737 3400 ;
     RECT  2736.38 2003.7 2737.82 2231.12 ;
     RECT  2737.82 2003.7 2738.3 2233.22 ;
     RECT  2735.9 1393.04 2739.46 1993.4 ;
     RECT  2738.3 2003.7 2740.42 2234.48 ;
     RECT  2352.58 1335.5 2740.9 1335.7 ;
     RECT  2546.98 1356.92 2743.78 1357.12 ;
     RECT  2739.46 1988.16 2744.06 1993.4 ;
     RECT  2740.42 2003.7 2744.06 2234.06 ;
     RECT  2744.06 1988.16 2747.9 2234.06 ;
     RECT  2739.46 1393.04 2748.38 1978.28 ;
     RECT  2747.9 1987.74 2748.38 2234.06 ;
     RECT  2748.38 1393.04 2750.5 2234.06 ;
     RECT  2750.5 1393.04 2757.7 2230.28 ;
     RECT  2757.7 1393.04 2760.085 2218.94 ;
     RECT  2760.085 1393.04 2763.46 2218.1 ;
     RECT  2763.46 1393.04 2764.9 2211.8 ;
     RECT  2764.9 2191.44 2765.38 2211.8 ;
     RECT  2764.9 1393.04 2767.78 2182.4 ;
     RECT  2767.78 2175.9 2769.22 2182.4 ;
     RECT  2765.38 2195.22 2769.22 2211.8 ;
     RECT  2769.22 2195.22 2769.7 2210.54 ;
     RECT  2769.7 2195.22 2770.66 2201.3 ;
     RECT  2769.22 2175.9 2772.1 2177.95 ;
     RECT  2767.78 1393.04 2773.06 2167.28 ;
     RECT  2773.06 1393.04 2773.54 2166.45 ;
     RECT  2585.86 2261.6 2774.3 2283.22 ;
     RECT  2402.02 2292.26 2774.3 2292.46 ;
     RECT  2773.54 2165.385 2774.915 2166.45 ;
     RECT  2774.915 2166.22 2775.365 2166.45 ;
     RECT  2772.1 2176.32 2775.445 2177.95 ;
     RECT  2770.66 2195.22 2776.42 2200.895 ;
     RECT  2775.445 2176.32 2778.82 2176.52 ;
     RECT  2776.42 2197.32 2779.1 2200.895 ;
     RECT  2775.365 2166.24 2779.3 2166.44 ;
     RECT  2779.1 2197.32 2779.3 2202.98 ;
     RECT  2757.7 2230.08 2779.3 2230.28 ;
     RECT  1591.58 197.72 2779.78 197.92 ;
     RECT  2779.3 2199.42 2780.26 2202.14 ;
     RECT  2773.54 1393.04 2783.42 2155.94 ;
     RECT  2783.42 1393.04 2785.82 2157.2 ;
     RECT  2785.82 1393.04 2787.74 2158.88 ;
     RECT  2787.74 1393.04 2789.66 2163.08 ;
     RECT  2789.66 1393.04 2791.1 2169.8 ;
     RECT  2404.42 2311.58 2793.5 2311.78 ;
     RECT  2774.3 2261.6 2793.7 2292.46 ;
     RECT  2791.1 1393.04 2794.94 2173.16 ;
     RECT  2794.94 1393.04 2795.9 2174 ;
     RECT  2795.9 1393.04 2796.1 2176.94 ;
     RECT  2796.1 1421.16 2796.38 2176.94 ;
     RECT  2796.38 1421.16 2796.58 2184.08 ;
     RECT  2727 -70 2797 180 ;
     RECT  2796.58 1421.58 2799.74 2184.08 ;
     RECT  2799.74 1421.58 2802.325 2185.34 ;
     RECT  2802.325 1425.15 2804.5 2185.34 ;
     RECT  2804.5 1425.36 2805.02 2185.34 ;
     RECT  2737 3220 2807 3470 ;
     RECT  2805.02 1425.36 2809.54 2192.06 ;
     RECT  2809.54 1427.88 2810.78 2192.06 ;
     RECT  2810.78 1427.88 2815.1 2192.9 ;
     RECT  2793.5 2311.16 2815.3 2311.78 ;
     RECT  2815.1 1427.88 2815.58 2195 ;
     RECT  2815.58 1427.88 2815.78 2196.68 ;
     RECT  2815.78 1427.88 2821.06 2196.26 ;
     RECT  2821.06 1427.88 2823.46 2193.32 ;
     RECT  2823.46 1429.56 2830.66 2193.32 ;
     RECT  2830.66 1438.38 2832.58 2193.32 ;
     RECT  2832.58 1439.64 2835.46 2193.32 ;
     RECT  2830.66 1429.56 2836.42 1429.76 ;
     RECT  2835.46 1440.48 2840.26 2193.32 ;
     RECT  2840.26 1440.48 2841.22 2189.54 ;
     RECT  2841.22 1440.48 2847.46 2186.18 ;
     RECT  2847.46 1458.96 2848.42 2186.18 ;
     RECT  2848.42 1462.57 2852.26 2186.18 ;
     RECT  2852.26 1462.57 2852.725 2185.76 ;
     RECT  2852.725 1462.74 2854.66 2185.76 ;
     RECT  2724.1 1380.84 2857.06 1381.04 ;
     RECT  2847.46 1440.48 2858.02 1449.5 ;
     RECT  2854.66 1465.68 2858.02 2185.76 ;
     RECT  2858.02 1465.68 2860.42 1533.92 ;
     RECT  2860.42 1466.94 2866.94 1533.92 ;
     RECT  2858.02 1542.54 2866.94 2185.76 ;
     RECT  2866.94 1466.94 2871.46 2185.76 ;
     RECT  2858.02 1445.1 2872.9 1449.5 ;
     RECT  2871.46 1486.26 2872.9 2185.76 ;
     RECT  2815.1 2343.5 2876.26 2343.7 ;
     RECT  2796.1 1393.04 2879.62 1407.52 ;
     RECT  2872.9 1486.68 2881.06 2183.66 ;
     RECT  2871.46 1466.94 2882.5 1473.44 ;
     RECT  2872.9 1445.1 2888.06 1445.3 ;
     RECT  2881.06 1486.68 2889.7 2183.24 ;
     RECT  2889.7 1496.76 2890.66 2183.24 ;
     RECT  2693.86 1370.76 2892.1 1370.96 ;
     RECT  2890.66 1499.7 2892.58 2183.24 ;
     RECT  2882.5 1466.94 2894.3 1467.14 ;
     RECT  2894.3 1466.94 2894.5 1467.98 ;
     RECT  2892.58 1503.48 2897.86 2183.24 ;
     RECT  2793.7 2261.6 2901.5 2283.22 ;
     RECT  2793.7 2292.26 2901.5 2292.46 ;
     RECT  2879.42 1382.12 2901.7 1382.32 ;
     RECT  2888.06 1445.1 2901.7 1451.62 ;
     RECT  2894.5 1467.78 2903.14 1467.98 ;
     RECT  2897.86 1503.9 2908.42 2183.24 ;
     RECT  2889.7 1486.68 2912.26 1486.88 ;
     RECT  2901.7 1445.1 2920.42 1445.3 ;
     RECT  2797 0 2921 180 ;
     RECT  2908.42 1504.32 2923.3 2183.24 ;
     RECT  2901.5 1371.62 2928.38 1371.82 ;
     RECT  2928.38 1364.06 2928.58 1371.82 ;
     RECT  2923.3 1504.32 2930.5 2182.4 ;
     RECT  2807 3220 2931 3400 ;
     RECT  2901.5 2261.6 2937.5 2292.46 ;
     RECT  2937.5 2261.6 2937.7 2300.44 ;
     RECT  2930.5 2182.2 2941.06 2182.4 ;
     RECT  2930.5 1504.32 2942.02 2171.48 ;
     RECT  2942.02 1522.785 2943.94 2171.48 ;
     RECT  2942.02 1504.32 2946.34 1513.34 ;
     RECT  2937.7 2292.26 2951.9 2300.44 ;
     RECT  2943.94 1522.785 2953.285 2168.12 ;
     RECT  2953.285 1522.785 2953.475 2169.38 ;
     RECT  2953.475 1523.62 2953.925 2169.38 ;
     RECT  2953.925 1523.64 2954.5 2169.38 ;
     RECT  2954.5 1526.58 2954.78 2169.38 ;
     RECT  2954.78 1526.58 2955.94 2169.8 ;
     RECT  2955.94 1530.78 2960.26 2169.38 ;
     RECT  2960.26 2153.64 2961.22 2168.54 ;
     RECT  2961.22 2154.06 2963.62 2168.54 ;
     RECT  2963.62 2154.48 2965.54 2159.72 ;
     RECT  2965.54 2155.74 2966.02 2159.72 ;
     RECT  2960.26 1530.78 2966.5 2144.6 ;
     RECT  2966.02 2158.68 2967.22 2159.72 ;
     RECT  2967.22 2158.68 2967.94 2158.88 ;
     RECT  2963.62 2168.34 2967.94 2168.54 ;
     RECT  2946.34 1504.32 2968.42 1511.66 ;
     RECT  2966.5 1532.46 2968.9 2144.6 ;
     RECT  2951.9 1439.24 2970.34 1439.44 ;
     RECT  2968.9 2144.4 2970.82 2144.6 ;
     RECT  2968.9 1532.46 2971.3 2125.28 ;
     RECT  2968.42 1507.26 2974.18 1511.66 ;
     RECT  2971.3 1532.46 2976.38 2124.86 ;
     RECT  2976.38 1532.04 2976.58 2124.86 ;
     RECT  2976.58 1532.04 2980.9 2123.6 ;
     RECT  2980.9 1532.04 2981.14 2120.66 ;
     RECT  2981.14 1532.04 2981.86 2117.72 ;
     RECT  2981.86 1532.04 2983.3 2116.04 ;
     RECT  2970.14 1483.34 2984.26 1483.54 ;
     RECT  2983.3 1532.04 2984.74 2113.94 ;
     RECT  2984.74 1532.04 2986.66 2112.68 ;
     RECT  2986.66 1532.04 2988.1 2111 ;
     RECT  2988.1 1532.04 2989.54 2110.58 ;
     RECT  2989.54 2081.82 2990.02 2109.32 ;
     RECT  2990.02 2081.82 2990.74 2108.48 ;
     RECT  2989.54 1532.04 2990.98 2072.78 ;
     RECT  2921 -70 2991 180 ;
     RECT  2990.98 1532.04 2991.46 2072.36 ;
     RECT  2991.46 1532.04 2992.7 2071.94 ;
     RECT  2990.74 2081.82 2994.82 2107.22 ;
     RECT  2992.7 1527.42 2995.3 2071.94 ;
     RECT  2995.3 1527.42 2996.06 2066.06 ;
     RECT  2994.82 2083.08 2996.26 2107.22 ;
     RECT  2996.06 1526.58 2997.02 2066.06 ;
     RECT  2974.18 1507.26 2997.5 1507.46 ;
     RECT  2997.02 1524.06 2997.92 2066.06 ;
     RECT  2997.5 1504.74 2997.98 1507.46 ;
     RECT  2997.98 1504.74 2998.4 1508.3 ;
     RECT  2997.02 1495.92 2999.42 1496.12 ;
     RECT  2998.4 1504.705 2999.42 1508.3 ;
     RECT  2999.42 1495.92 2999.9 1512.5 ;
     RECT  2997.92 1523.05 2999.9 2066.06 ;
     RECT  2996.26 2091.9 3000.58 2107.22 ;
     RECT  2931 3220 3001 3470 ;
     RECT  3000.58 2094 3001.06 2097.56 ;
     RECT  3000.58 2107.02 3001.54 2107.22 ;
     RECT  3001.06 2094.21 3002.02 2097.56 ;
     RECT  2999.9 1495.92 3003.46 2066.06 ;
     RECT  3003.46 1495.92 3003.94 2062.28 ;
     RECT  3003.94 1495.92 3004.9 2058.92 ;
     RECT  3004.9 1495.92 3007.3 2055.98 ;
     RECT  2951.9 2292.26 3013.06 2300.86 ;
     RECT  3007.3 1496.76 3016.7 2049.43 ;
     RECT  2876.06 2401.04 3016.9 2401.24 ;
     RECT  3016.7 1496.76 3017.66 2049.68 ;
     RECT  3013.06 2292.26 3020.26 2300.44 ;
     RECT  3017.66 1492.98 3021.02 2049.68 ;
     RECT  3021.02 1492.14 3023.14 2049.68 ;
     RECT  3023.14 1492.14 3023.9 2046.74 ;
     RECT  3023.9 1491.72 3026.5 2046.74 ;
     RECT  3026.5 1491.72 3026.98 2045.48 ;
     RECT  3026.98 2036.88 3029.38 2045.48 ;
     RECT  3012.86 2343.5 3031.1 2343.7 ;
     RECT  3029.38 2037.72 3031.3 2045.48 ;
     RECT  3020.06 2328.38 3031.3 2328.58 ;
     RECT  3031.3 2037.72 3034.18 2037.92 ;
     RECT  3031.1 2339.72 3038.5 2343.7 ;
     RECT  3016.7 2413.22 3045.7 2413.42 ;
     RECT  3026.98 1491.72 3045.98 2027.84 ;
     RECT  1911.26 2352.74 3052.7 2352.94 ;
     RECT  3038.5 2340.14 3052.9 2343.7 ;
     RECT  3040.7 1476.6 3055.58 1476.8 ;
     RECT  3045.98 1487.94 3060.38 2027.84 ;
     RECT  3060.38 1487.94 3062.3 2029.1 ;
     RECT  3052.7 2352.74 3063.46 2354.62 ;
     RECT  3060.38 2046.12 3063.74 2046.32 ;
     RECT  3055.58 1476.6 3064.22 1479.32 ;
     RECT  3062.3 1487.94 3064.22 2030.36 ;
     RECT  3064.22 1476.6 3065.18 2030.36 ;
     RECT  3065.18 1476.6 3065.66 2031.2 ;
     RECT  3045.5 2422.46 3065.66 2422.66 ;
     RECT  3063.26 2433.8 3065.66 2434 ;
     RECT  3065.66 2422.46 3065.86 2434 ;
     RECT  2928.58 1364.06 3067.1 1364.26 ;
     RECT  3065.66 1476.6 3068.5 2033.72 ;
     RECT  3068.5 1621.5 3068.73 2033.72 ;
     RECT  3068.73 1621.5 3070.41 1852.7 ;
     RECT  3068.5 1476.6 3071.62 1611.62 ;
     RECT  3068.73 1863 3072.1 2033.72 ;
     RECT  3071.62 1611.42 3073.06 1611.62 ;
     RECT  3072.1 1863 3073.06 1889.66 ;
     RECT  3072.1 1898.7 3073.06 2033.72 ;
     RECT  3071.62 1476.6 3073.54 1601.96 ;
     RECT  3070.41 1621.92 3073.54 1852.7 ;
     RECT  3073.06 1863 3073.54 1877.48 ;
     RECT  3073.06 1898.7 3073.54 1937.96 ;
     RECT  3073.06 1947.84 3073.54 1961.06 ;
     RECT  3073.06 1970.52 3073.82 2033.72 ;
     RECT  3063.74 2043.6 3073.82 2046.32 ;
     RECT  3073.54 1621.92 3074.02 1670.84 ;
     RECT  3073.54 1679.88 3074.02 1852.7 ;
     RECT  3073.54 1476.6 3074.5 1595.24 ;
     RECT  3073.54 1863 3074.5 1876.64 ;
     RECT  3073.06 1886.52 3074.5 1889.66 ;
     RECT  3065.86 2426.66 3074.5 2434 ;
     RECT  3074.5 1579.08 3074.98 1595.24 ;
     RECT  3074.5 1886.52 3074.98 1888.82 ;
     RECT  3067.1 1364.06 3077.86 1371.82 ;
     RECT  3074.3 2448.08 3081.5 2448.28 ;
     RECT  3074.5 2426.66 3081.7 2426.86 ;
     RECT  3073.82 1970.52 3083.9 2046.32 ;
     RECT  2815.3 2311.58 3085.06 2311.78 ;
     RECT  3081.5 2448.08 3085.06 2455.42 ;
     RECT  2937.7 2261.6 3087.46 2283.22 ;
     RECT  2879.62 1400.18 3088.42 1407.52 ;
     RECT  3087.46 2264.12 3088.42 2283.22 ;
     RECT  3074.5 1476.6 3088.7 1570.04 ;
     RECT  3074.98 1582.44 3088.7 1595.24 ;
     RECT  3074.02 1623.18 3088.7 1670.84 ;
     RECT  3074.02 1679.88 3088.7 1833.8 ;
     RECT  3074.5 1863.42 3088.7 1876.64 ;
     RECT  3073.54 1899.96 3088.7 1937.96 ;
     RECT  3073.54 1947.84 3088.7 1960.64 ;
     RECT  3083.9 1970.52 3088.7 2053.88 ;
     RECT  3074.98 1887.36 3089.18 1888.82 ;
     RECT  3088.7 1897.44 3089.18 2053.88 ;
     RECT  3088.7 1582.44 3090.14 1602.8 ;
     RECT  3084.86 2512.34 3092.26 2512.54 ;
     RECT  3090.14 1582.44 3092.54 1607.84 ;
     RECT  3074.02 1849.56 3093.02 1852.7 ;
     RECT  3088.7 1862.16 3093.02 1876.64 ;
     RECT  3093.02 1849.56 3093.5 1876.64 ;
     RECT  3089.18 1887.36 3093.5 2053.88 ;
     RECT  3092.54 1582.44 3094.46 1612.88 ;
     RECT  3088.7 1622.76 3094.46 1833.8 ;
     RECT  3093.5 1849.56 3094.46 2053.88 ;
     RECT  3088.7 1469.04 3095.9 1570.04 ;
     RECT  3095.9 1469.04 3096.38 1572.56 ;
     RECT  3094.46 1582.44 3096.38 2053.88 ;
     RECT  3020.26 2292.26 3098.98 2292.46 ;
     RECT  3096.38 1469.04 3099.26 2055.58 ;
     RECT  3092.06 2577.02 3099.46 2577.22 ;
     RECT  3099.26 1467.8 3099.7 2055.58 ;
     RECT  3099.7 1467.8 3099.94 2053.88 ;
     RECT  3099.94 1469.04 3100 2053.88 ;
     RECT  3100 1477.04 3100.42 1484.8 ;
     RECT  3100 2015.06 3100.42 2015.26 ;
     RECT  3100 1496.76 3100.9 1499.48 ;
     RECT  3100 1962.14 3100.9 1980.8 ;
     RECT  3100 2051.16 3100.9 2051.36 ;
     RECT  3100 1514.4 3101.38 1514.6 ;
     RECT  3100.9 1964.24 3101.38 1980.8 ;
     RECT  3088.42 2267.06 3101.38 2283.22 ;
     RECT  3100.9 1499.28 3101.86 1499.48 ;
     RECT  3100 2028.48 3101.86 2028.68 ;
     RECT  3099.26 2666.48 3105.22 2666.68 ;
     RECT  3077.66 1310.3 3107.62 1310.5 ;
     RECT  3100 1941.98 3107.62 1947.22 ;
     RECT  3100 1558.94 3110.98 1559.14 ;
     RECT  3101.38 1964.24 3110.98 1972.42 ;
     RECT  3101.38 2283.02 3110.98 2283.22 ;
     RECT  3110.98 1965.92 3111.46 1972.42 ;
     RECT  3101.38 2267.06 3111.46 2269.78 ;
     RECT  3111.46 2267.06 3111.94 2267.26 ;
     RECT  3111.46 1965.92 3112.42 1969.9 ;
     RECT  3107.62 1947.02 3112.9 1947.22 ;
     RECT  3100 1900.4 3113.38 1900.6 ;
     RECT  3112.42 1969.7 3113.38 1969.9 ;
     RECT  3085.06 2455.22 3114.82 2455.42 ;
     RECT  2991 0 3115 180 ;
     RECT  3107.42 1241 3117.22 1241.2 ;
     RECT  3059.9 1385.9 3117.7 1386.1 ;
     RECT  3105.02 2691.68 3117.7 2691.88 ;
     RECT  3117.5 1376.24 3124.9 1376.44 ;
     RECT  3001 3220 3125 3400 ;
     RECT  3117.02 1216.64 3128.26 1216.84 ;
     RECT  3128.06 1137.68 3131.9 1137.88 ;
     RECT  3131.9 1137.26 3132.1 1137.88 ;
     RECT  3117.5 2718.14 3132.58 2718.34 ;
     RECT  3088.42 1400.18 3137.86 1404.16 ;
     RECT  3124.7 1353.14 3139.3 1353.34 ;
     RECT  3132.1 1137.26 3142.66 1137.46 ;
     RECT  3139.1 1317.86 3146.3 1318.06 ;
     RECT  3146.3 1317.44 3146.5 1318.06 ;
     RECT  3114.62 2464.46 3146.5 2464.66 ;
     RECT  3132.38 2743.34 3146.5 2743.54 ;
     RECT  3142.46 969.68 3149.86 969.88 ;
     RECT  3149.66 884.42 3153.7 884.62 ;
     RECT  3146.5 1317.44 3157.06 1317.64 ;
     RECT  3052.9 2343.5 3160.42 2343.7 ;
     RECT  3063.46 2352.74 3160.7 2352.94 ;
     RECT  3153.5 870.98 3164.26 871.18 ;
     RECT  3146.3 2757.62 3165.7 2757.82 ;
     RECT  3077.86 1364.06 3168.1 1364.26 ;
     RECT  3137.66 1380.02 3170.5 1380.22 ;
     RECT  3156.86 1281.32 3171.46 1281.52 ;
     RECT  3146.3 2473.28 3171.46 2473.48 ;
     RECT  3160.7 2352.74 3175.3 2357.98 ;
     RECT  3169.82 1328.36 3180.86 1328.56 ;
     RECT  3170.3 1360.7 3181.06 1360.9 ;
     RECT  3165.5 2771.9 3182.98 2772.1 ;
     RECT  3115 -70 3185 180 ;
     RECT  3164.06 712.64 3185.86 712.84 ;
     RECT  3171.26 1120.04 3185.86 1120.24 ;
     RECT  3100 1760.12 3193.06 1760.32 ;
     RECT  3169.82 2116.7 3193.06 2116.9 ;
     RECT  3171.26 2534.6 3193.06 2534.8 ;
     RECT  3125 3220 3195 3470 ;
     RECT  3180.86 1328.36 3196.9 1333.6 ;
     RECT  3185.66 673.58 3198.82 673.78 ;
     RECT  3196.9 1328.36 3200.26 1328.56 ;
     RECT  3185.66 1050.74 3203.62 1050.94 ;
     RECT  3192.86 2570.3 3204.1 2570.5 ;
     RECT  3207.26 1579.52 3207.74 1579.72 ;
     RECT  3192.86 2078.9 3207.94 2079.1 ;
     RECT  1669.82 606.8 3217.82 609.94 ;
     RECT  1789.54 800.42 3217.82 803.98 ;
     RECT  3214.46 842 3217.82 842.2 ;
     RECT  1572.86 994.46 3217.82 998.02 ;
     RECT  3203.42 1036.04 3217.82 1036.24 ;
     RECT  1645.82 1188.5 3217.82 1192.06 ;
     RECT  3171.26 1618.16 3217.82 1618.36 ;
     RECT  3192.86 1811.78 3217.82 1811.98 ;
     RECT  3207.74 2005.82 3217.82 2006.02 ;
     RECT  3175.3 2352.74 3217.82 2352.94 ;
     RECT  3175.1 2393.9 3217.82 2394.1 ;
     RECT  3203.9 2587.94 3217.82 2588.14 ;
     RECT  3182.78 2781.98 3217.82 2782.18 ;
     RECT  3185 0 3220 180 ;
     RECT  3217.82 606.375 3220 609.94 ;
     RECT  3198.62 647.96 3220 648.16 ;
     RECT  3217.82 800.375 3220 803.98 ;
     RECT  3217.82 841.875 3220 842.2 ;
     RECT  3217.82 994.375 3220 998.02 ;
     RECT  3217.82 1035.875 3220 1036.24 ;
     RECT  3217.82 1188.375 3220 1192.06 ;
     RECT  3200.06 1216.64 3220 1216.84 ;
     RECT  3214.46 1230.08 3220 1230.28 ;
     RECT  3196.7 1309.04 3220 1309.24 ;
     RECT  3137.86 1403.96 3220 1404.16 ;
     RECT  3196.7 1423.7 3220 1423.9 ;
     RECT  3207.74 1576.58 3220 1579.72 ;
     RECT  3217.82 1617.875 3220 1618.36 ;
     RECT  3217.82 1811.78 3220 1812.075 ;
     RECT  3207.26 1967.6 3220 1967.8 ;
     RECT  3217.82 2005.82 3220 2006.075 ;
     RECT  3207.74 2161.22 3220 2161.42 ;
     RECT  3217.82 2352.375 3220 2352.94 ;
     RECT  3217.82 2393.875 3220 2394.1 ;
     RECT  3217.82 2587.875 3220 2588.14 ;
     RECT  3217.82 2781.875 3220 2782.18 ;
     RECT  3195 3220 3220 3400 ;
     RECT  3220 0 3400 3400 ;
     RECT  3400 205 3470 275 ;
     RECT  3400 399 3470 469 ;
     RECT  3400 593 3470 663 ;
     RECT  3400 787 3470 857 ;
     RECT  3400 981 3470 1051 ;
     RECT  3400 1175 3470 1245 ;
     RECT  3400 1369 3470 1439 ;
     RECT  3400 1563 3470 1633 ;
     RECT  3400 1757 3470 1827 ;
     RECT  3400 1951 3470 2021 ;
     RECT  3400 2145 3470 2215 ;
     RECT  3400 2339 3470 2409 ;
     RECT  3400 2533 3470 2603 ;
     RECT  3400 2727 3470 2797 ;
     RECT  3400 2921 3470 2991 ;
     RECT  3400 3115 3470 3185 ;
    LAYER Metal3 ;
     RECT  205 -70 275 0 ;
     RECT  399 -70 469 0 ;
     RECT  593 -70 663 0 ;
     RECT  787 -70 857 0 ;
     RECT  981 -70 1051 0 ;
     RECT  1175 -70 1245 0 ;
     RECT  1369 -70 1439 0 ;
     RECT  1563 -70 1633 0 ;
     RECT  1757 -70 1827 0 ;
     RECT  1951 -70 2021 0 ;
     RECT  2145 -70 2215 0 ;
     RECT  2339 -70 2409 0 ;
     RECT  2533 -70 2603 0 ;
     RECT  2727 -70 2797 0 ;
     RECT  2921 -70 2991 0 ;
     RECT  3115 -70 3185 0 ;
     RECT  0 0 3400 178 ;
     RECT  0 178 180 180 ;
     RECT  606.225 178 609.775 180 ;
     RECT  647.725 178 654.82 180 ;
     RECT  800.225 178 804.1 180 ;
     RECT  841.725 178 842.225 180 ;
     RECT  994.225 178 998.02 180 ;
     RECT  1035.725 178 1036.42 180 ;
     RECT  1188.225 178 1191.94 180 ;
     RECT  1229.725 178 1230.34 180 ;
     RECT  1382.225 178 1385.86 180 ;
     RECT  1423.725 178 1425.22 180 ;
     RECT  1617.5 178 1618.225 180 ;
     RECT  1770.225 178 1773.775 180 ;
     RECT  1811.725 178 1812.225 180 ;
     RECT  2005.725 178 2006.5 180 ;
     RECT  2199.725 178 2200.42 180 ;
     RECT  2352.225 178 2355.94 180 ;
     RECT  2393.725 178 2394.34 180 ;
     RECT  2546.225 178 2549.86 180 ;
     RECT  2587.725 178 2588.26 180 ;
     RECT  2740.225 178 2743.78 180 ;
     RECT  2779.58 178 2782.225 180 ;
     RECT  3220 178 3400 180 ;
     RECT  1617.5 180 1617.94 181.96 ;
     RECT  1770.62 180 1773.46 181.96 ;
     RECT  2006.06 180 2006.5 181.96 ;
     RECT  2546.54 180 2549.86 181.96 ;
     RECT  1384.7 180 1385.86 183.64 ;
     RECT  1576.22 178 1580.26 183.64 ;
     RECT  2156.06 178 2162.02 183.64 ;
     RECT  1962.14 178 1968.1 184.06 ;
     RECT  1463.9 178 1464.1 197.72 ;
     RECT  994.46 180 998.02 197.92 ;
     RECT  2779.58 180 2779.78 197.92 ;
     RECT  3222 180 3400 205 ;
     RECT  0 180 178 215 ;
     RECT  1457.66 197.72 1464.1 219.56 ;
     RECT  1188.38 180 1191.94 219.76 ;
     RECT  1450.46 219.56 1464.1 226.7 ;
     RECT  1036.22 180 1036.42 226.9 ;
     RECT  3222 205 3470 275 ;
     RECT  -70 215 178 285 ;
     RECT  3222 275 3400 399 ;
     RECT  0 285 178 409 ;
     RECT  3222 399 3470 469 ;
     RECT  -70 409 178 479 ;
     RECT  997.82 197.92 998.02 586.84 ;
     RECT  3222 469 3400 593 ;
     RECT  993 594.8 995 597.4 ;
     RECT  1405 594.8 1407 597.4 ;
     RECT  0 479 178 603 ;
     RECT  3222 593 3470 606.225 ;
     RECT  3220 606.225 3470 609.775 ;
     RECT  -70 603 178 635.78 ;
     RECT  -70 635.78 180.58 636.4 ;
     RECT  -70 636.4 180 639.855 ;
     RECT  3222 609.775 3470 647.725 ;
     RECT  3220 647.725 3470 647.96 ;
     RECT  3219.26 647.96 3470 648.16 ;
     RECT  3220 648.16 3470 648.225 ;
     RECT  3222 648.225 3470 663 ;
     RECT  -70 639.855 178 673 ;
     RECT  3198.62 647.96 3198.82 673.78 ;
     RECT  3185.66 673.58 3185.86 712.84 ;
     RECT  1191.74 219.76 1191.94 716.62 ;
     RECT  1230.14 180 1230.34 723.76 ;
     RECT  1186.14 729.68 1187.3 730.1 ;
     RECT  1302.3 729.26 1302.5 730.1 ;
     RECT  1215.42 730.1 1215.62 730.52 ;
     RECT  1215.42 730.52 1216.1 731.36 ;
     RECT  1302.3 730.1 1305.86 733.04 ;
     RECT  1208.22 731.36 1223.78 733.46 ;
     RECT  1113.66 733.04 1113.86 733.88 ;
     RECT  1182.78 730.1 1195.94 733.88 ;
     RECT  1205.82 733.46 1223.78 733.88 ;
     RECT  1302.3 733.04 1310.18 733.88 ;
     RECT  1182.78 733.88 1223.78 734.3 ;
     RECT  1302.3 733.88 1316.42 734.72 ;
     RECT  1181.34 734.3 1223.78 735.14 ;
     RECT  1181.34 735.14 1228.58 736.82 ;
     RECT  1161.66 736.82 1161.86 737.24 ;
     RECT  1174.14 736.82 1228.58 737.24 ;
     RECT  1098.3 732.62 1098.5 737.66 ;
     RECT  1109.34 733.88 1113.86 737.66 ;
     RECT  1126.62 734.3 1126.82 737.66 ;
     RECT  1289.82 736.82 1290.02 737.66 ;
     RECT  1300.38 734.72 1316.42 737.66 ;
     RECT  1385.66 183.64 1385.86 738.04 ;
     RECT  1095.42 737.66 1126.82 738.08 ;
     RECT  1161.66 737.24 1228.58 738.08 ;
     RECT  1288.86 737.66 1290.02 738.08 ;
     RECT  1300.38 737.66 1318.82 738.08 ;
     RECT  993 597.4 997.6 738.92 ;
     RECT  1095.42 738.08 1131.62 741.02 ;
     RECT  993 738.92 998.5 741.2 ;
     RECT  1288.86 738.08 1318.82 741.44 ;
     RECT  1344.54 740.6 1344.74 741.44 ;
     RECT  1143.42 738.92 1143.62 741.86 ;
     RECT  1161.66 738.08 1231.94 741.86 ;
     RECT  1287.9 741.44 1318.82 741.86 ;
     RECT  1344.06 741.44 1344.74 741.86 ;
     RECT  1081.5 741.44 1081.7 742.28 ;
     RECT  1092.06 741.02 1131.62 742.28 ;
     RECT  1141.98 741.86 1231.94 742.28 ;
     RECT  1337.34 741.86 1344.74 742.28 ;
     RECT  1080.54 742.28 1081.7 742.7 ;
     RECT  1092.06 742.28 1231.94 742.7 ;
     RECT  993 741.2 999.46 742.88 ;
     RECT  988.7 742.88 999.46 743.96 ;
     RECT  1062.3 741.44 1062.5 744.38 ;
     RECT  1080.54 742.7 1231.94 744.38 ;
     RECT  1062.3 744.38 1231.94 744.8 ;
     RECT  1062.3 744.8 1237.22 745.22 ;
     RECT  988.7 743.96 1000.66 745.6 ;
     RECT  1287.9 741.86 1325.54 745.64 ;
     RECT  1336.86 742.28 1344.74 745.64 ;
     RECT  1062.3 745.22 1242.02 746.48 ;
     RECT  1402.4 597.4 1407 746.48 ;
     RECT  1049.34 746.48 1049.54 749 ;
     RECT  1062.3 746.48 1242.5 749 ;
     RECT  1287.9 745.64 1344.74 749 ;
     RECT  1401.02 746.48 1407 749 ;
     RECT  1049.34 749 1242.5 749.42 ;
     RECT  1399.34 749 1407 750.64 ;
     RECT  1049.34 749.42 1246.34 751.52 ;
     RECT  1259.1 751.1 1259.3 751.52 ;
     RECT  1279.74 749 1344.74 751.94 ;
     RECT  1358.46 749 1358.66 751.94 ;
     RECT  1399.58 750.64 1407 753.38 ;
     RECT  1279.74 751.94 1358.66 753.4 ;
     RECT  1425.02 180 1425.22 755.9 ;
     RECT  1049.34 751.52 1259.3 756.98 ;
     RECT  1301.34 753.4 1358.66 756.98 ;
     RECT  1049.34 756.98 1265.06 757.4 ;
     RECT  1279.74 753.4 1291.46 757.4 ;
     RECT  1301.34 756.98 1359.14 758.66 ;
     RECT  1301.34 758.66 1361.06 759.7 ;
     RECT  1049.34 757.4 1291.46 760.76 ;
     RECT  1424.54 755.9 1425.22 763.04 ;
     RECT  1399.58 753.38 1407.46 763.24 ;
     RECT  988.7 745.6 999.46 764.12 ;
     RECT  1046.46 760.76 1291.46 764.54 ;
     RECT  1301.34 759.7 1359.14 764.54 ;
     RECT  1046.46 764.54 1359.14 764.74 ;
     RECT  988.7 764.12 1007.3 765.16 ;
     RECT  1046.46 764.74 1293.38 766 ;
     RECT  1046.46 766 1292.42 767.68 ;
     RECT  1046.46 767.68 1290.98 768.74 ;
     RECT  1036.86 768.74 1290.98 772.3 ;
     RECT  1400.54 763.24 1407.46 776.06 ;
     RECT  1417.34 763.04 1425.22 776.06 ;
     RECT  1304.22 764.74 1359.14 776.3 ;
     RECT  988.7 765.16 999.94 776.72 ;
     RECT  1303.26 776.3 1359.14 777.14 ;
     RECT  1443.26 226.7 1464.1 777.32 ;
     RECT  1039.26 772.3 1290.98 779.66 ;
     RECT  1300.86 777.14 1359.14 779.66 ;
     RECT  1039.26 779.66 1359.14 783.22 ;
     RECT  988.7 776.72 1000.66 783.86 ;
     RECT  3222 663 3400 787 ;
     RECT  1039.26 783.22 1331.78 787.22 ;
     RECT  1033.98 787.22 1331.78 787.42 ;
     RECT  1341.66 783.22 1359.14 790.78 ;
     RECT  1400.54 776.06 1425.22 791.6 ;
     RECT  1389.98 791.6 1425.22 792.04 ;
     RECT  1033.98 787.42 1330.34 795.2 ;
     RECT  0 673 178 797 ;
     RECT  3222 787 3470 800.225 ;
     RECT  1341.66 790.78 1357.22 801.28 ;
     RECT  1341.66 801.28 1344.26 801.7 ;
     RECT  1033.02 795.2 1330.34 802.34 ;
     RECT  1341.66 801.7 1343.78 802.34 ;
     RECT  3220 800.225 3470 803.775 ;
     RECT  1389.98 792.04 1390.18 804.44 ;
     RECT  1400.06 792.04 1425.22 804.44 ;
     RECT  1033.02 802.34 1343.78 805.06 ;
     RECT  1038.78 805.06 1342.34 805.9 ;
     RECT  1038.78 805.9 1330.34 806.32 ;
     RECT  1389.98 804.44 1425.22 808.82 ;
     RECT  1435.58 777.32 1464.1 808.82 ;
     RECT  988.7 783.86 1001.54 809.48 ;
     RECT  1039.74 806.32 1330.34 813.04 ;
     RECT  1040.22 813.04 1330.34 817.66 ;
     RECT  1040.22 817.66 1287.14 818.5 ;
     RECT  1330.14 817.66 1330.34 821.02 ;
     RECT  1299.42 817.66 1319.78 821.44 ;
     RECT  1299.42 821.44 1315.94 824.8 ;
     RECT  988.7 809.48 1007.3 825.22 ;
     RECT  988.7 825.22 1006.82 826.46 ;
     RECT  1040.22 818.5 1285.22 828.38 ;
     RECT  1299.42 824.8 1312.1 828.38 ;
     RECT  -70 797 178 831.725 ;
     RECT  1354.62 801.28 1357.22 831.94 ;
     RECT  -70 831.725 180 832.225 ;
     RECT  1389.98 808.82 1464.1 834.86 ;
     RECT  1356.54 831.94 1357.22 835.72 ;
     RECT  1040.22 828.38 1312.1 836.78 ;
     RECT  987.26 826.46 1006.82 837.4 ;
     RECT  974.3 753.38 974.5 839.06 ;
     RECT  987.26 837.4 1002.5 839.06 ;
     RECT  1357.02 835.72 1357.22 839.92 ;
     RECT  3222 803.775 3470 841.725 ;
     RECT  1789.34 812.18 1789.54 842 ;
     RECT  3220 841.725 3470 842 ;
     RECT  974.3 839.06 1002.5 847.48 ;
     RECT  1040.22 836.78 1312.58 851.06 ;
     RECT  1040.22 851.06 1317.38 852.52 ;
     RECT  1044.54 852.52 1317.38 855.26 ;
     RECT  1044.54 855.26 1326.5 855.88 ;
     RECT  3214.46 842 3470 857 ;
     RECT  1044.54 855.88 1314.5 857.56 ;
     RECT  1050.3 857.56 1314.5 861.76 ;
     RECT  1053.18 861.76 1314.5 863.02 ;
     RECT  1281.66 863.02 1314.5 863.44 ;
     RECT  974.3 847.48 1001.86 863.84 ;
     RECT  1326.3 855.88 1326.5 866.18 ;
     RECT  1341.66 805.9 1342.34 866.18 ;
     RECT  -70 832.225 178 867 ;
     RECT  1319.58 866.18 1342.34 869.32 ;
     RECT  974.3 863.84 1009.06 870.98 ;
     RECT  1020.38 863.42 1020.58 870.98 ;
     RECT  3164.06 712.64 3164.26 871.18 ;
     RECT  1053.18 863.02 1268.42 873.52 ;
     RECT  1061.34 873.52 1268.42 873.74 ;
     RECT  1281.66 863.44 1309.7 873.74 ;
     RECT  1319.58 869.32 1341.86 873.74 ;
     RECT  974.3 870.98 1020.58 874.96 ;
     RECT  1061.34 873.74 1341.86 876.88 ;
     RECT  1061.34 876.88 1337.06 878.14 ;
     RECT  1061.34 878.14 1258.82 881.5 ;
     RECT  1270.62 878.14 1337.06 881.5 ;
     RECT  3153.5 870.98 3153.7 884.42 ;
     RECT  1062.3 881.5 1256.42 884.44 ;
     RECT  3149.66 884.42 3153.7 884.62 ;
     RECT  1072.86 884.44 1256.42 888.22 ;
     RECT  1237.5 888.22 1256.42 888.64 ;
     RECT  1238.94 888.64 1256.42 889.06 ;
     RECT  1072.86 888.22 1227.14 891.58 ;
     RECT  1247.58 889.06 1256.42 892.64 ;
     RECT  1062.3 884.44 1062.5 892.84 ;
     RECT  1247.58 892.64 1258.82 893.06 ;
     RECT  1270.62 881.5 1336.1 893.06 ;
     RECT  1072.86 891.58 1220.42 893.26 ;
     RECT  1077.18 893.26 1217.54 893.68 ;
     RECT  1089.66 893.68 1217.54 895.78 ;
     RECT  1077.18 893.68 1079.3 896.2 ;
     RECT  1105.98 895.78 1217.54 896.2 ;
     RECT  1247.58 893.06 1336.1 896.42 ;
     RECT  1079.1 896.2 1079.3 896.62 ;
     RECT  1094.46 895.78 1094.66 896.62 ;
     RECT  1105.98 896.2 1194.02 896.62 ;
     RECT  1205.34 896.2 1217.54 896.62 ;
     RECT  1205.34 896.62 1211.78 897.04 ;
     RECT  1247.58 896.42 1340.42 897.04 ;
     RECT  1105.98 896.62 1193.54 899.56 ;
     RECT  1105.98 899.56 1190.66 899.98 ;
     RECT  1107.9 899.98 1190.66 900.4 ;
     RECT  1258.62 897.04 1340.42 900.4 ;
     RECT  1109.82 900.4 1190.66 900.82 ;
     RECT  1210.62 897.04 1211.78 900.82 ;
     RECT  1284.06 900.4 1340.42 900.82 ;
     RECT  1210.62 900.82 1210.82 901.24 ;
     RECT  1259.1 900.4 1272.74 903.34 ;
     RECT  1129.5 900.82 1179.62 903.76 ;
     RECT  1247.58 897.04 1248.74 904.18 ;
     RECT  1263.9 903.34 1272.74 904.18 ;
     RECT  1284.06 900.82 1312.1 904.18 ;
     RECT  1247.58 904.18 1247.78 904.6 ;
     RECT  1133.34 903.76 1179.62 905.02 ;
     RECT  1141.5 905.02 1179.62 907.12 ;
     RECT  1323.9 900.82 1340.42 907.12 ;
     RECT  1156.86 907.12 1179.62 907.96 ;
     RECT  1284.06 904.18 1309.7 907.96 ;
     RECT  1141.5 907.12 1144.1 908.38 ;
     RECT  1156.86 907.96 1165.7 908.38 ;
     RECT  1264.86 904.18 1269.86 908.38 ;
     RECT  1284.06 907.96 1308.74 908.38 ;
     RECT  1326.3 907.12 1340.42 908.38 ;
     RECT  1177.02 907.96 1179.62 908.8 ;
     RECT  1340.22 908.38 1340.42 908.8 ;
     RECT  1143.9 908.38 1144.1 909.22 ;
     RECT  1306.14 908.38 1308.74 909.22 ;
     RECT  974.3 874.96 998.5 909.62 ;
     RECT  1308.54 909.22 1308.74 909.64 ;
     RECT  1284.06 908.38 1293.86 911.32 ;
     RECT  1326.3 908.38 1326.5 911.74 ;
     RECT  1284.06 911.32 1284.26 912.16 ;
     RECT  973.34 909.62 998.5 919.7 ;
     RECT  1008.86 874.96 1020.58 919.7 ;
     RECT  3149.66 884.62 3149.86 969.68 ;
     RECT  3142.46 969.68 3149.86 969.88 ;
     RECT  3214.46 857 3400 981 ;
     RECT  0 867 178 991 ;
     RECT  1579.58 183.64 1580.26 994.46 ;
     RECT  1788.86 842 1789.54 994.8 ;
     RECT  1788.86 994.8 1795 997.4 ;
     RECT  3105 994.8 3107 997.4 ;
     RECT  1559.42 178 1559.62 997.82 ;
     RECT  1572.86 994.46 1580.26 997.82 ;
     RECT  1770.62 181.96 1773.22 1019.24 ;
     RECT  1770.62 1019.24 1777.54 1022.8 ;
     RECT  -70 991 178 1025.725 ;
     RECT  -70 1025.725 180 1026.225 ;
     RECT  201.5 1025.96 201.7 1033.3 ;
     RECT  3203.42 1036.04 3203.62 1050.94 ;
     RECT  3214.46 981 3470 1051 ;
     RECT  -70 1026.225 178 1061 ;
     RECT  3185.66 1050.74 3185.86 1120.24 ;
     RECT  3142.46 969.88 3142.66 1137.46 ;
     RECT  3214.46 1051 3400 1175 ;
     RECT  0 1061 178 1185 ;
     RECT  1617.5 181.96 1617.7 1188.5 ;
     RECT  1630.46 609.74 1630.66 1188.5 ;
     RECT  3128.06 1137.68 3128.26 1216.84 ;
     RECT  3214.46 1175 3470 1216.84 ;
     RECT  -70 1185 178 1219.725 ;
     RECT  -70 1219.725 180 1220.225 ;
     RECT  3222 1216.84 3470 1229.725 ;
     RECT  3220 1229.725 3470 1230.08 ;
     RECT  3102.4 997.4 3107 1241 ;
     RECT  3117.02 1216.64 3117.22 1241 ;
     RECT  3102.4 1241 3117.22 1241.2 ;
     RECT  3214.46 1230.08 3470 1245 ;
     RECT  -70 1220.225 178 1255 ;
     RECT  973.34 919.7 1020.58 1274.3 ;
     RECT  1130.3 1275.44 1130.5 1275.86 ;
     RECT  1129.82 1275.86 1130.5 1276.7 ;
     RECT  1144.22 1275.44 1144.42 1276.7 ;
     RECT  1159.58 1276.28 1159.78 1276.7 ;
     RECT  1173.5 1275.44 1173.7 1276.7 ;
     RECT  1129.82 1276.7 1144.42 1279.64 ;
     RECT  1156.22 1276.7 1159.78 1279.64 ;
     RECT  1170.62 1276.7 1173.7 1279.64 ;
     RECT  1124.06 1279.64 1144.42 1280.06 ;
     RECT  1156.22 1279.64 1173.7 1280.06 ;
     RECT  1124.06 1280.06 1173.7 1280.48 ;
     RECT  3171.26 1120.04 3171.46 1281.52 ;
     RECT  1124.06 1280.48 1177.06 1282.58 ;
     RECT  1108.7 1282.58 1177.06 1283 ;
     RECT  1096.7 1283 1096.9 1287.62 ;
     RECT  1192.7 1287.2 1192.9 1287.62 ;
     RECT  1214.78 1287.2 1214.98 1288.04 ;
     RECT  1192.7 1287.62 1196.26 1288.88 ;
     RECT  1206.14 1288.04 1215.46 1288.88 ;
     RECT  1108.7 1283 1180.9 1290.98 ;
     RECT  1073.18 1290.56 1073.38 1291.82 ;
     RECT  1096.7 1287.62 1097.38 1291.82 ;
     RECT  1108.7 1290.98 1182.34 1291.82 ;
     RECT  1096.7 1291.82 1182.34 1293.08 ;
     RECT  1096.7 1293.08 1182.82 1294.76 ;
     RECT  1192.7 1288.88 1215.46 1294.76 ;
     RECT  1073.18 1291.82 1074.34 1295.18 ;
     RECT  1086.62 1291.82 1086.82 1295.18 ;
     RECT  1071.74 1295.18 1086.82 1295.6 ;
     RECT  1096.7 1294.76 1215.46 1295.6 ;
     RECT  1071.74 1295.6 1215.94 1298.12 ;
     RECT  1065.5 1298.12 1218.34 1299.38 ;
     RECT  1049.18 874.76 1049.38 1301.06 ;
     RECT  1063.58 1299.38 1218.34 1301.48 ;
     RECT  1040.06 1301.06 1049.38 1302.32 ;
     RECT  1063.1 1301.48 1218.34 1302.32 ;
     RECT  1033.34 1302.32 1049.38 1302.74 ;
     RECT  1062.14 1302.32 1218.34 1302.74 ;
     RECT  972.86 1274.3 1020.58 1303.16 ;
     RECT  1033.34 1302.74 1051.78 1303.16 ;
     RECT  1062.14 1302.74 1220.26 1305.68 ;
     RECT  3200.06 1216.64 3200.26 1309.04 ;
     RECT  3214.46 1245 3400 1309.24 ;
     RECT  972.86 1303.16 1051.78 1310.3 ;
     RECT  1062.14 1305.68 1224.1 1310.3 ;
     RECT  3102.4 1241.2 3107.62 1310.5 ;
     RECT  972.86 1310.3 1224.1 1313.66 ;
     RECT  972.86 1313.66 1226.5 1314.5 ;
     RECT  3156.86 1281.32 3157.06 1317.64 ;
     RECT  972.86 1314.5 1232.74 1320.38 ;
     RECT  972.38 1320.38 1232.74 1320.8 ;
     RECT  965.66 1320.8 1232.74 1321.22 ;
     RECT  1559.42 997.82 1580.26 1321.22 ;
     RECT  2352.38 180 2355.94 1321.42 ;
     RECT  950.78 1321.22 1232.74 1325 ;
     RECT  944.06 1325 1237.54 1326.46 ;
     RECT  2352.38 1321.42 2352.58 1328.56 ;
     RECT  3196.7 1309.04 3200.26 1328.56 ;
     RECT  944.54 1326.46 1237.54 1328.78 ;
     RECT  944.54 1328.78 1240.42 1332.34 ;
     RECT  3196.7 1328.56 3196.9 1333.6 ;
     RECT  1645.82 1191.86 1646.02 1335.5 ;
     RECT  1656.38 800.42 1656.58 1335.5 ;
     RECT  2740.7 180 2743.78 1335.7 ;
     RECT  1107.26 1332.34 1240.42 1337.18 ;
     RECT  944.54 1332.34 1097.38 1340.12 ;
     RECT  1107.26 1337.18 1242.34 1340.12 ;
     RECT  1788.86 997.4 1797.6 1342.64 ;
     RECT  1339.58 918.02 1339.78 1342.84 ;
     RECT  941.66 1340.12 1097.38 1343.9 ;
     RECT  1107.26 1340.12 1246.66 1343.9 ;
     RECT  1788.86 1342.64 1800.58 1346.3 ;
     RECT  3169.82 1328.36 3170.02 1346.3 ;
     RECT  1559.42 1321.22 1581.7 1346.5 ;
     RECT  3167.9 1346.3 3170.02 1346.5 ;
     RECT  941.66 1343.9 1246.66 1347.26 ;
     RECT  941.66 1347.26 1250.02 1347.68 ;
     RECT  2546.78 181.96 2549.86 1349.98 ;
     RECT  941.66 1347.68 1253.86 1351.46 ;
     RECT  3139.1 1317.86 3139.3 1353.34 ;
     RECT  941.66 1351.46 1256.74 1355.24 ;
     RECT  1617.5 1188.5 1630.66 1356.92 ;
     RECT  2743.58 1335.7 2743.78 1357.12 ;
     RECT  941.66 1355.24 1262.02 1358.6 ;
     RECT  3167.9 1346.5 3168.1 1360.7 ;
     RECT  3180.86 1333.4 3181.06 1360.9 ;
     RECT  940.7 1358.6 1262.02 1362.8 ;
     RECT  3167.9 1360.7 3170.5 1364.26 ;
     RECT  940.22 1362.8 1262.02 1366.36 ;
     RECT  3222 1309.24 3400 1369 ;
     RECT  2891.9 1370.76 2892.1 1371.62 ;
     RECT  2928.38 1364.06 2928.58 1371.82 ;
     RECT  3077.66 1310.3 3077.86 1371.82 ;
     RECT  940.7 1366.36 1262.02 1374.98 ;
     RECT  1770.62 1022.8 1773.22 1375.82 ;
     RECT  1788.86 1346.3 1801.06 1375.82 ;
     RECT  3124.7 1353.14 3124.9 1376.24 ;
     RECT  3117.5 1376.24 3124.9 1376.44 ;
     RECT  940.7 1374.98 1263.46 1378.54 ;
     RECT  1617.5 1356.92 1632.1 1378.76 ;
     RECT  1645.82 1335.5 1656.58 1378.76 ;
     RECT  0 1255 178 1379 ;
     RECT  3170.3 1364.26 3170.5 1380.22 ;
     RECT  1617.5 1378.76 1656.58 1381.7 ;
     RECT  1669.82 606.8 1670.02 1381.7 ;
     RECT  940.7 1378.54 1262.02 1381.9 ;
     RECT  3222 1369 3470 1382.225 ;
     RECT  2891.9 1371.62 2901.7 1382.32 ;
     RECT  3220 1382.225 3470 1382.54 ;
     RECT  940.7 1381.9 1021.06 1385.48 ;
     RECT  1725.02 1370.78 1725.22 1385.9 ;
     RECT  3067.1 1371.62 3067.3 1385.9 ;
     RECT  3117.5 1376.44 3117.7 1386.1 ;
     RECT  938.78 1385.48 1021.06 1388.84 ;
     RECT  2693.66 1373.28 2693.86 1389.26 ;
     RECT  2494.94 1375.8 2495.14 1390.92 ;
     RECT  1715.9 1385.9 1725.22 1390.94 ;
     RECT  1617.5 1381.7 1670.02 1392.62 ;
     RECT  934.46 1388.84 1021.06 1393.04 ;
     RECT  1031.9 1381.9 1262.02 1393.04 ;
     RECT  1617.5 1392.62 1670.5 1393.04 ;
     RECT  2723.9 1388.4 2724.1 1393.04 ;
     RECT  2879.42 1382.12 2879.62 1393.24 ;
     RECT  2490.14 1390.92 2495.14 1393.44 ;
     RECT  1617.5 1393.04 1673.38 1393.88 ;
     RECT  1616.54 1393.88 1673.86 1395.56 ;
     RECT  1770.62 1375.82 1801.06 1396.18 ;
     RECT  1613.18 1395.56 1673.86 1396.82 ;
     RECT  2666.78 1383.36 2666.98 1400.18 ;
     RECT  2685.5 1389.26 2693.86 1400.18 ;
     RECT  2705.66 1395.96 2705.86 1400.18 ;
     RECT  3059.42 1385.9 3067.3 1400.38 ;
     RECT  3137.66 1380.02 3137.86 1400.38 ;
     RECT  2666.3 1400.18 2666.98 1400.6 ;
     RECT  3067.1 1400.38 3067.3 1400.8 ;
     RECT  2723.9 1393.04 2728.9 1403.54 ;
     RECT  1611.26 1396.82 1673.86 1403.96 ;
     RECT  1683.74 1398.5 1683.94 1403.96 ;
     RECT  2666.3 1400.6 2673.7 1403.96 ;
     RECT  2685.5 1400.18 2705.86 1403.96 ;
     RECT  3217.82 1382.54 3470 1404.16 ;
     RECT  1591.58 197.72 1591.78 1404.38 ;
     RECT  1611.26 1403.96 1683.94 1404.38 ;
     RECT  3083.42 1403.96 3083.62 1404.8 ;
     RECT  3102.4 1310.5 3107 1405.22 ;
     RECT  1702.94 803.78 1703.14 1406.06 ;
     RECT  3083.42 1404.8 3085.54 1406.48 ;
     RECT  3100.22 1405.22 3107 1408.16 ;
     RECT  3099.74 1408.16 3107 1408.58 ;
     RECT  1702.94 1406.06 1704.58 1409 ;
     RECT  1770.62 1396.18 1800.58 1409 ;
     RECT  3083.42 1406.48 3086.98 1409.42 ;
     RECT  3097.34 1408.58 3107 1409.42 ;
     RECT  2779.1 1409.82 2779.3 1410.24 ;
     RECT  2779.1 1410.24 2782.66 1410.66 ;
     RECT  1770.14 1409 1800.58 1411.1 ;
     RECT  1811.9 180 1812.1 1411.1 ;
     RECT  2755.58 1410.68 2764.9 1411.1 ;
     RECT  934.46 1393.04 1262.02 1411.52 ;
     RECT  1699.58 1409 1704.58 1411.94 ;
     RECT  1715.9 1390.94 1728.1 1411.94 ;
     RECT  1699.58 1411.94 1728.1 1412.14 ;
     RECT  1702.94 1412.14 1728.1 1412.56 ;
     RECT  2779.1 1410.66 2783.14 1412.76 ;
     RECT  1591.58 1404.38 1601.38 1412.78 ;
     RECT  1611.26 1404.38 1684.9 1412.78 ;
     RECT  2716.7 1403.54 2728.9 1412.78 ;
     RECT  1810.94 1411.1 1812.1 1412.98 ;
     RECT  2716.7 1412.78 2732.26 1413.6 ;
     RECT  2754.62 1411.1 2765.38 1413.6 ;
     RECT  2779.1 1412.76 2785.06 1413.6 ;
     RECT  2796.38 1412.78 2796.58 1413.6 ;
     RECT  1742.78 1380.86 1742.98 1413.62 ;
     RECT  -70 1379 178 1413.725 ;
     RECT  2716.7 1413.6 2765.38 1414.02 ;
     RECT  2779.1 1413.6 2796.58 1414.02 ;
     RECT  2631.74 1409 2631.94 1414.04 ;
     RECT  -70 1413.725 180 1414.225 ;
     RECT  2631.74 1414.04 2633.38 1414.46 ;
     RECT  3207.26 1410.26 3207.46 1414.88 ;
     RECT  934.46 1411.52 1262.98 1415.3 ;
     RECT  1559.9 1346.5 1581.7 1415.3 ;
     RECT  1591.58 1412.78 1684.9 1415.3 ;
     RECT  2549.66 1349.98 2549.86 1415.5 ;
     RECT  933.02 1415.3 1262.98 1415.72 ;
     RECT  1559.9 1415.3 1684.9 1416.56 ;
     RECT  2666.3 1403.96 2705.86 1417.5 ;
     RECT  3222 1404.16 3470 1419.08 ;
     RECT  2891.9 1382.32 2892.1 1419.92 ;
     RECT  2666.3 1417.5 2706.34 1421.16 ;
     RECT  2716.7 1414.02 2796.58 1421.16 ;
     RECT  2666.3 1421.16 2796.58 1422 ;
     RECT  2631.26 1414.46 2633.38 1422.02 ;
     RECT  2666.3 1422 2803.3 1422.42 ;
     RECT  3221.18 1419.08 3470 1423.7 ;
     RECT  3196.7 1412.78 3196.9 1423.9 ;
     RECT  3219.26 1423.7 3470 1423.9 ;
     RECT  932.54 1415.72 1263.46 1424.12 ;
     RECT  1559.9 1416.56 1690.18 1424.12 ;
     RECT  1702.94 1412.56 1704.58 1424.12 ;
     RECT  3220 1423.9 3470 1424.225 ;
     RECT  2666.3 1422.42 2805.7 1424.94 ;
     RECT  1715.9 1412.56 1728.1 1425.7 ;
     RECT  1739.9 1413.62 1742.98 1425.7 ;
     RECT  2666.3 1424.94 2809.06 1425.8 ;
     RECT  2588.06 180 2588.26 1426 ;
     RECT  2657.66 1425.8 2809.06 1426 ;
     RECT  2685.5 1426 2809.06 1426.2 ;
     RECT  932.54 1424.12 1269.7 1427.26 ;
     RECT  2685.5 1426.2 2810.02 1428.72 ;
     RECT  2631.26 1422.02 2642.5 1429.36 ;
     RECT  2841.5 1398.48 2841.7 1429.56 ;
     RECT  2161.82 183.64 2162.02 1429.78 ;
     RECT  2657.66 1426 2673.22 1430 ;
     RECT  2656.22 1430 2673.22 1430.2 ;
     RECT  932.54 1427.26 1264.9 1431.04 ;
     RECT  2441.66 1426.2 2441.86 1431.24 ;
     RECT  2656.22 1430.2 2672.74 1432.52 ;
     RECT  2685.5 1428.72 2816.74 1432.92 ;
     RECT  2426.78 1385.88 2426.98 1433.76 ;
     RECT  2441.66 1431.24 2444.26 1433.76 ;
     RECT  1559.9 1424.12 1704.58 1434.2 ;
     RECT  1715.9 1425.7 1727.62 1434.2 ;
     RECT  2685.5 1432.92 2824.42 1435.86 ;
     RECT  2836.22 1429.56 2841.7 1435.86 ;
     RECT  1769.18 1411.1 1800.58 1436.06 ;
     RECT  2685.5 1435.86 2841.7 1436.28 ;
     RECT  1559.9 1434.2 1727.62 1437.98 ;
     RECT  2006.3 181.96 2006.5 1438.18 ;
     RECT  2426.78 1433.76 2444.26 1438.8 ;
     RECT  3221.18 1424.225 3470 1439 ;
     RECT  2684.06 1436.28 2844.58 1439.1 ;
     RECT  2951.9 1419.5 2952.1 1439.44 ;
     RECT  1555.1 1437.98 1727.62 1439.66 ;
     RECT  1554.62 1439.66 1727.62 1440.5 ;
     RECT  1967.9 184.06 1968.1 1440.7 ;
     RECT  2200.22 180 2200.42 1441.12 ;
     RECT  2631.26 1429.36 2638.66 1441.32 ;
     RECT  1506.14 178 1506.34 1442.18 ;
     RECT  1554.14 1440.5 1727.62 1442.18 ;
     RECT  933.98 1431.04 1264.9 1443.02 ;
     RECT  2631.26 1441.32 2640.1 1443.02 ;
     RECT  2652.86 1432.52 2672.74 1443.02 ;
     RECT  2460.86 1403.52 2461.06 1443.86 ;
     RECT  2534.3 1429.16 2534.5 1444.06 ;
     RECT  2631.26 1443.02 2672.74 1444.26 ;
     RECT  2684.06 1439.1 2845.06 1444.26 ;
     RECT  1504.7 1442.18 1507.3 1444.7 ;
     RECT  1811.9 1412.98 1812.1 1444.9 ;
     RECT  915.26 1441.76 915.46 1445.12 ;
     RECT  928.22 1443.02 1264.9 1445.12 ;
     RECT  2394.14 180 2394.34 1445.32 ;
     RECT  915.26 1445.12 1264.9 1445.54 ;
     RECT  1491.26 769.34 1491.46 1445.54 ;
     RECT  1504.7 1444.7 1511.62 1445.54 ;
     RECT  1491.26 1445.54 1518.34 1445.96 ;
     RECT  1541.18 1445.12 1541.38 1445.96 ;
     RECT  1554.14 1442.18 1728.58 1445.96 ;
     RECT  1769.18 1436.06 1798.18 1445.96 ;
     RECT  1769.18 1445.96 1798.66 1446.36 ;
     RECT  1491.26 1445.96 1519.3 1446.8 ;
     RECT  1769.18 1446.36 1800.34 1446.8 ;
     RECT  915.26 1445.54 1267.3 1447.1 ;
     RECT  -70 1414.225 178 1449 ;
     RECT  1491.26 1446.8 1524.1 1449.1 ;
     RECT  1764.38 1446.8 1800.34 1449.74 ;
     RECT  2888.06 1419.92 2892.1 1451.42 ;
     RECT  2904.38 1451.4 2904.58 1451.42 ;
     RECT  2888.06 1451.42 2904.58 1451.62 ;
     RECT  1540.7 1445.96 1728.58 1453.52 ;
     RECT  1740.38 1425.7 1742.98 1453.52 ;
     RECT  914.3 1447.1 1267.3 1453.94 ;
     RECT  1537.34 1453.52 1728.58 1453.94 ;
     RECT  1739.42 1453.52 1742.98 1453.94 ;
     RECT  1763.42 1449.74 1800.34 1455.62 ;
     RECT  1537.34 1453.94 1742.98 1456.04 ;
     RECT  2460.86 1443.86 2464.42 1456.46 ;
     RECT  2457.02 1456.46 2464.42 1456.66 ;
     RECT  1535.42 1456.04 1742.98 1456.88 ;
     RECT  1756.7 1455.62 1800.34 1456.88 ;
     RECT  1535.42 1456.88 1800.34 1457.3 ;
     RECT  1534.46 1457.3 1800.34 1457.72 ;
     RECT  1533.5 1457.72 1800.34 1458.96 ;
     RECT  2631.26 1444.26 2845.06 1459.38 ;
     RECT  2856.86 1380.84 2857.06 1459.38 ;
     RECT  1491.26 1449.1 1520.26 1459.82 ;
     RECT  1533.5 1458.96 1800.58 1459.82 ;
     RECT  1287.74 925.16 1287.94 1461.08 ;
     RECT  914.3 1453.94 1267.78 1461.5 ;
     RECT  1279.1 1461.08 1287.94 1461.5 ;
     RECT  1491.26 1459.82 1800.58 1461.5 ;
     RECT  2631.26 1459.38 2857.06 1464 ;
     RECT  1487.42 1461.5 1800.58 1464.02 ;
     RECT  914.3 1461.5 1287.94 1464.44 ;
     RECT  2457.02 1456.66 2461.06 1465.06 ;
     RECT  2631.26 1464 2858.02 1466.1 ;
     RECT  2631.26 1466.1 2858.5 1467.8 ;
     RECT  2627.9 1467.8 2858.5 1467.9 ;
     RECT  2627.9 1467.9 2858.98 1468.22 ;
     RECT  1485.5 1464.02 1800.58 1468.64 ;
     RECT  2602.46 1456.44 2602.66 1469.06 ;
     RECT  2613.5 1454.36 2613.7 1469.06 ;
     RECT  2624.54 1468.22 2858.98 1471.14 ;
     RECT  1389.98 834.86 1472.26 1472 ;
     RECT  1484.06 1468.64 1800.58 1472 ;
     RECT  2889.5 1451.62 2904.58 1473.24 ;
     RECT  2602.46 1469.06 2613.7 1475.36 ;
     RECT  2624.54 1471.14 2868.1 1475.36 ;
     RECT  2368.7 1464.86 2368.9 1475.98 ;
     RECT  910.46 1464.44 1287.94 1479.56 ;
     RECT  2347.1 1475.78 2347.3 1483.12 ;
     RECT  2970.14 1439.24 2970.34 1483.54 ;
     RECT  2882.3 1473.24 2904.58 1486.06 ;
     RECT  2602.46 1475.36 2868.1 1486.26 ;
     RECT  2904.38 1486.06 2904.58 1486.68 ;
     RECT  2920.22 1445.1 2920.42 1486.68 ;
     RECT  909.5 1479.56 1288.9 1486.9 ;
     RECT  3055.58 1486.68 3055.78 1487.94 ;
     RECT  2602.46 1486.26 2868.58 1488.78 ;
     RECT  2882.3 1486.06 2892.1 1488.78 ;
     RECT  3055.58 1487.94 3060.1 1488.78 ;
     RECT  3055.58 1488.78 3063.46 1489.2 ;
     RECT  2314.94 1483.34 2315.14 1491.94 ;
     RECT  3053.18 1489.2 3063.46 1492.56 ;
     RECT  3053.18 1492.56 3073.06 1492.98 ;
     RECT  3047.9 1492.98 3073.06 1493.4 ;
     RECT  2602.46 1488.78 2892.1 1494.46 ;
     RECT  2554.46 1476.6 2554.66 1494.68 ;
     RECT  2602.46 1494.46 2612.74 1494.88 ;
     RECT  3018.14 1492.98 3028.9 1496.34 ;
     RECT  1389.98 1472 1800.58 1496.76 ;
     RECT  2997.02 1495.92 2997.22 1496.76 ;
     RECT  3018.14 1496.34 3030.34 1496.76 ;
     RECT  3044.06 1493.4 3073.06 1497.18 ;
     RECT  2997.02 1496.76 3030.34 1498.02 ;
     RECT  3040.7 1497.18 3073.06 1498.02 ;
     RECT  1389.98 1496.76 1807.3 1498.22 ;
     RECT  606.62 180 609.7 1499.5 ;
     RECT  1389.98 1498.22 1800.58 1499.92 ;
     RECT  2624.06 1494.46 2892.1 1500.96 ;
     RECT  606.62 1499.5 606.82 1501.6 ;
     RECT  2997.02 1498.02 3073.06 1501.8 ;
     RECT  3083.42 1409.42 3107 1501.8 ;
     RECT  2624.06 1500.96 2894.5 1503.48 ;
     RECT  2904.38 1486.68 2920.42 1503.48 ;
     RECT  2997.02 1501.8 3107 1504.94 ;
     RECT  3055.58 1504.94 3107 1505.36 ;
     RECT  2624.06 1503.48 2920.42 1508.94 ;
     RECT  2931.26 1508.52 2931.46 1508.94 ;
     RECT  2997.02 1504.94 3045.22 1508.94 ;
     RECT  2408.54 1428.72 2408.74 1509.36 ;
     RECT  2419.58 1438.8 2444.26 1509.36 ;
     RECT  1389.98 1499.92 1799.14 1511.88 ;
     RECT  2624.06 1508.94 2938.18 1513.14 ;
     RECT  1389.98 1511.88 1800.34 1513.78 ;
     RECT  909.5 1486.9 1287.94 1514.84 ;
     RECT  2552.06 1494.68 2554.66 1515.26 ;
     RECT  2552.06 1515.26 2556.1 1515.46 ;
     RECT  2588.06 1490.48 2588.26 1515.46 ;
     RECT  2460.86 1465.06 2461.06 1516.92 ;
     RECT  2995.58 1508.94 3045.22 1518.6 ;
     RECT  3055.58 1505.36 3072.1 1518.6 ;
     RECT  2480.54 1393.44 2495.14 1519.44 ;
     RECT  1422.62 1513.78 1800.34 1520.72 ;
     RECT  2552.06 1515.46 2555.62 1520.92 ;
     RECT  654.62 180 654.82 1521.34 ;
     RECT  909.5 1514.84 1288.9 1521.98 ;
     RECT  2984.06 1483.34 2984.26 1523.02 ;
     RECT  2995.58 1518.6 3072.1 1523.84 ;
     RECT  2477.66 1519.44 2495.14 1524.48 ;
     RECT  2508.38 1520.72 2508.58 1524.48 ;
     RECT  907.58 1521.98 1288.9 1524.5 ;
     RECT  1299.26 1343.48 1299.46 1524.5 ;
     RECT  1422.62 1520.72 1800.58 1524.5 ;
     RECT  1389.98 1513.78 1410.82 1526.5 ;
     RECT  2624.06 1513.14 2946.34 1526.58 ;
     RECT  2995.58 1523.84 3045.22 1527.42 ;
     RECT  907.58 1524.5 1299.46 1528.06 ;
     RECT  3084.86 1505.36 3107 1528.06 ;
     RECT  2624.06 1526.58 2955.94 1528.26 ;
     RECT  2554.46 1520.92 2555.62 1530.16 ;
     RECT  3097.34 1528.06 3107 1530.58 ;
     RECT  2624.06 1528.26 2959.3 1530.78 ;
     RECT  2969.66 1484.16 2969.86 1530.78 ;
     RECT  2584.7 1521.98 2584.9 1531.42 ;
     RECT  841.82 180 842.02 1531.84 ;
     RECT  2624.06 1530.78 2969.86 1532.04 ;
     RECT  907.58 1528.06 1288.9 1532.26 ;
     RECT  867.26 1414.04 867.46 1532.48 ;
     RECT  867.26 1532.48 876.58 1532.9 ;
     RECT  2460.86 1516.92 2461.54 1533.74 ;
     RECT  2568.38 1531.22 2568.58 1533.94 ;
     RECT  3084.86 1528.06 3087.46 1533.94 ;
     RECT  2454.62 1533.74 2461.54 1534.56 ;
     RECT  2984.06 1534.14 2984.26 1534.56 ;
     RECT  2995.1 1527.42 3045.22 1534.56 ;
     RECT  3056.06 1523.84 3072.1 1534.56 ;
     RECT  2541.5 1529.96 2541.7 1535.62 ;
     RECT  3084.86 1533.94 3086.98 1535.62 ;
     RECT  907.58 1532.26 1287.94 1536.68 ;
     RECT  3084.86 1535.62 3086.02 1538.14 ;
     RECT  2554.46 1530.16 2554.66 1539.9 ;
     RECT  2554.46 1539.9 2555.14 1540.1 ;
     RECT  3085.82 1538.14 3086.02 1541.08 ;
     RECT  2624.06 1532.04 2974.18 1541.7 ;
     RECT  2984.06 1534.56 3072.1 1541.7 ;
     RECT  2624.06 1541.7 3072.1 1542.32 ;
     RECT  3097.82 1530.58 3107 1543.18 ;
     RECT  2624.06 1542.32 3066.82 1544.44 ;
     RECT  2454.62 1534.56 2466.82 1544.64 ;
     RECT  2477.66 1524.48 2508.58 1544.64 ;
     RECT  2408.54 1509.36 2444.26 1544.66 ;
     RECT  2454.62 1544.64 2508.58 1544.66 ;
     RECT  2408.54 1544.66 2508.58 1544.86 ;
     RECT  2638.94 1544.44 3066.82 1546.94 ;
     RECT  867.26 1532.9 880.9 1547.18 ;
     RECT  907.1 1536.68 1287.94 1547.8 ;
     RECT  867.26 1547.18 889.54 1548.1 ;
     RECT  1422.62 1524.5 1801.06 1548.22 ;
     RECT  800.54 180 804.1 1549.48 ;
     RECT  2986.46 1546.94 3066.82 1550.3 ;
     RECT  803.9 1549.48 804.1 1550.32 ;
     RECT  3098.3 1543.18 3107 1558.3 ;
     RECT  2602.46 1494.88 2603.14 1558.72 ;
     RECT  3098.78 1558.3 3107 1558.94 ;
     RECT  907.58 1547.8 1287.94 1559.78 ;
     RECT  1373.18 1465.7 1373.38 1560.2 ;
     RECT  2638.94 1546.94 2975.14 1561.02 ;
     RECT  2638.94 1561.02 2979.46 1562.28 ;
     RECT  2991.74 1550.3 3066.82 1562.28 ;
     RECT  3098.78 1558.94 3110.98 1562.5 ;
     RECT  1339.1 1560.2 1373.38 1562.72 ;
     RECT  3221.18 1439 3400 1563 ;
     RECT  907.1 1559.78 1287.94 1563.14 ;
     RECT  1299.26 1528.06 1299.46 1563.14 ;
     RECT  2638.94 1562.28 3066.82 1564.38 ;
     RECT  2624.06 1544.44 2624.26 1565.86 ;
     RECT  2530.46 1535.42 2530.66 1566.28 ;
     RECT  907.1 1563.14 1299.46 1566.5 ;
     RECT  1336.7 1562.72 1373.38 1566.5 ;
     RECT  2408.54 1544.86 2500.9 1566.7 ;
     RECT  899.9 1566.5 1299.46 1567.12 ;
     RECT  2339.9 1558.94 2340.1 1567.54 ;
     RECT  1328.54 1566.5 1373.38 1567.76 ;
     RECT  1328.54 1567.76 1376.26 1568.18 ;
     RECT  1422.62 1548.22 1799.14 1569.42 ;
     RECT  1390.46 1526.5 1410.82 1569.44 ;
     RECT  1422.62 1569.42 1801.54 1569.84 ;
     RECT  1328.54 1568.18 1377.22 1569.86 ;
     RECT  1389.02 1569.44 1410.82 1569.86 ;
     RECT  867.74 1548.1 889.54 1570.48 ;
     RECT  889.34 1570.48 889.54 1570.7 ;
     RECT  899.9 1567.12 1287.94 1570.7 ;
     RECT  3099.5 1562.5 3110.98 1572.36 ;
     RECT  0 1449 178 1573 ;
     RECT  2638.94 1564.38 3071.14 1574.04 ;
     RECT  2638.94 1574.04 3072.58 1574.46 ;
     RECT  1328.54 1569.86 1410.82 1575.32 ;
     RECT  3221.18 1563 3470 1576.225 ;
     RECT  3220 1576.225 3470 1576.58 ;
     RECT  3207.26 1414.88 3207.94 1576.78 ;
     RECT  3219.26 1576.58 3470 1576.78 ;
     RECT  1326.14 1575.32 1410.82 1577 ;
     RECT  2638.94 1574.46 3073.54 1577.4 ;
     RECT  1317.02 1577 1410.82 1577.84 ;
     RECT  1422.62 1569.84 1805.38 1578.46 ;
     RECT  1425.98 1578.46 1805.38 1578.88 ;
     RECT  3207.26 1576.78 3207.46 1579.72 ;
     RECT  3220 1576.78 3470 1579.775 ;
     RECT  2638.46 1577.4 3073.54 1580.12 ;
     RECT  2638.46 1580.12 3071.62 1580.54 ;
     RECT  1316.06 1577.84 1410.82 1582.04 ;
     RECT  889.34 1570.7 1287.94 1582.24 ;
     RECT  2408.54 1566.7 2444.26 1582.44 ;
     RECT  1311.26 1582.04 1410.82 1584.76 ;
     RECT  2406.62 1582.44 2444.26 1590 ;
     RECT  2459.9 1566.7 2500.9 1590 ;
     RECT  2602.46 1558.72 2602.66 1592.1 ;
     RECT  925.82 1582.24 1287.94 1592.32 ;
     RECT  2602.46 1592.1 2609.38 1592.72 ;
     RECT  925.82 1592.32 1058.02 1593.16 ;
     RECT  1067.9 1592.32 1287.94 1596.1 ;
     RECT  925.82 1593.16 1051.78 1596.52 ;
     RECT  2638.46 1580.54 3067.3 1597.14 ;
     RECT  867.74 1570.48 876.58 1598 ;
     RECT  889.34 1582.24 909.22 1598 ;
     RECT  1425.98 1578.88 1453.54 1598 ;
     RECT  1463.42 1578.88 1805.38 1598 ;
     RECT  1425.98 1598 1805.38 1598.3 ;
     RECT  2635.1 1597.14 3067.3 1598.4 ;
     RECT  867.74 1598 914.5 1598.42 ;
     RECT  2635.1 1598.4 3069.22 1599.44 ;
     RECT  1067.9 1596.1 1268.74 1599.88 ;
     RECT  867.74 1598.42 914.98 1600.52 ;
     RECT  925.82 1596.52 1049.38 1600.52 ;
     RECT  1299.26 1567.12 1299.46 1600.52 ;
     RECT  1312.22 1584.76 1410.82 1600.52 ;
     RECT  1067.9 1599.88 1267.78 1600.72 ;
     RECT  867.74 1600.52 1049.38 1601.14 ;
     RECT  1067.9 1600.72 1266.34 1601.14 ;
     RECT  1067.9 1601.14 1262.5 1601.56 ;
     RECT  3081.5 1592.52 3081.7 1602.6 ;
     RECT  3095.9 1572.36 3110.98 1602.6 ;
     RECT  1080.38 1601.56 1262.5 1604.5 ;
     RECT  2554.94 1540.1 2555.14 1604.7 ;
     RECT  1425.02 1598.3 1805.38 1604.92 ;
     RECT  1299.26 1600.52 1410.82 1605.76 ;
     RECT  834.62 1605.56 834.82 1605.98 ;
     RECT  1041.98 1601.14 1049.38 1607.44 ;
     RECT  2609.18 1592.72 2609.38 1607.64 ;
     RECT  -70 1573 178 1607.725 ;
     RECT  1425.02 1604.92 1595.62 1607.86 ;
     RECT  834.62 1605.98 842.02 1608.08 ;
     RECT  852.38 1605.14 852.58 1608.08 ;
     RECT  -70 1607.725 180 1608.225 ;
     RECT  867.74 1601.14 1030.66 1608.28 ;
     RECT  1309.82 1605.76 1410.82 1608.28 ;
     RECT  829.82 1608.08 842.02 1608.5 ;
     RECT  1325.18 1608.28 1410.82 1609.12 ;
     RECT  2635.1 1599.44 3068.26 1610.16 ;
     RECT  822.14 1608.5 842.02 1611.02 ;
     RECT  852.38 1608.08 854.02 1611.02 ;
     RECT  867.74 1608.28 1029.7 1611.44 ;
     RECT  822.14 1611.02 854.02 1612.28 ;
     RECT  864.86 1611.44 1029.7 1612.28 ;
     RECT  1080.38 1604.5 1259.14 1612.48 ;
     RECT  822.14 1612.28 1029.7 1612.7 ;
     RECT  1080.38 1612.48 1255.78 1612.7 ;
     RECT  2633.66 1610.16 3068.26 1613.3 ;
     RECT  2633.66 1613.3 3064.9 1614.56 ;
     RECT  815.9 1612.7 1029.7 1615.64 ;
     RECT  1606.94 1604.92 1805.38 1615.64 ;
     RECT  1299.26 1605.76 1299.46 1616.26 ;
     RECT  1077.98 1612.7 1255.78 1616.68 ;
     RECT  1042.46 1607.44 1049.38 1616.9 ;
     RECT  2554.94 1604.7 2560.42 1617.72 ;
     RECT  3221.18 1579.775 3470 1617.725 ;
     RECT  2635.1 1614.56 3064.9 1617.92 ;
     RECT  3220 1617.725 3470 1618.225 ;
     RECT  3171.26 1587.5 3171.46 1618.36 ;
     RECT  808.7 1615.64 1029.7 1618.58 ;
     RECT  1042.46 1616.9 1053.7 1618.58 ;
     RECT  1067.9 1601.56 1068.1 1619 ;
     RECT  1309.82 1608.28 1314.82 1619.42 ;
     RECT  1325.66 1609.12 1410.82 1619.42 ;
     RECT  1603.1 1615.64 1805.38 1619.42 ;
     RECT  808.7 1618.58 1053.7 1619.84 ;
     RECT  1066.46 1619 1068.1 1619.84 ;
     RECT  1425.02 1607.86 1590.82 1619.84 ;
     RECT  1602.14 1619.42 1805.38 1619.84 ;
     RECT  1077.98 1616.68 1253.38 1620.04 ;
     RECT  1309.82 1619.42 1410.82 1620.26 ;
     RECT  2608.7 1607.64 2609.38 1620.66 ;
     RECT  1077.98 1620.04 1252.9 1622.56 ;
     RECT  1425.02 1619.84 1805.38 1622.78 ;
     RECT  3081.5 1602.6 3110.98 1622.96 ;
     RECT  808.7 1619.84 1068.1 1623.62 ;
     RECT  1077.98 1622.56 1242.82 1623.62 ;
     RECT  2541.02 1590.42 2541.22 1624.44 ;
     RECT  2553.5 1617.72 2560.42 1624.44 ;
     RECT  2541.02 1624.44 2560.42 1625.28 ;
     RECT  1279.1 1596.1 1287.94 1627.3 ;
     RECT  808.7 1623.62 1242.82 1627.6 ;
     RECT  2534.78 1625.28 2560.42 1627.8 ;
     RECT  2530.94 1627.8 2560.42 1629.06 ;
     RECT  2406.62 1590 2500.9 1629.48 ;
     RECT  2516.54 1629.06 2560.42 1629.48 ;
     RECT  3081.5 1622.96 3081.7 1630.1 ;
     RECT  1303.1 1620.26 1410.82 1631.6 ;
     RECT  1423.58 1622.78 1805.38 1631.6 ;
     RECT  808.7 1627.6 1235.14 1632.02 ;
     RECT  2406.62 1629.48 2560.42 1632.42 ;
     RECT  2636.54 1617.92 3064.9 1632.42 ;
     RECT  2598.62 1632.42 2598.82 1632.84 ;
     RECT  2608.7 1620.66 2612.26 1632.84 ;
     RECT  3221.18 1618.225 3470 1633 ;
     RECT  2598.62 1632.84 2612.26 1634.72 ;
     RECT  2406.62 1632.42 2562.34 1635.36 ;
     RECT  2636.54 1632.42 3066.82 1636.82 ;
     RECT  1279.58 1627.3 1287.94 1637.06 ;
     RECT  1303.1 1631.6 1805.38 1637.06 ;
     RECT  2406.14 1635.36 2562.34 1637.46 ;
     RECT  1279.58 1637.06 1805.38 1637.48 ;
     RECT  2637.98 1636.82 3066.82 1637.88 ;
     RECT  807.74 1632.02 1235.14 1638.1 ;
     RECT  1272.38 1637.48 1805.38 1638.3 ;
     RECT  1225.82 1638.1 1235.14 1638.32 ;
     RECT  1225.82 1638.32 1241.38 1638.52 ;
     RECT  2406.14 1637.46 2568.58 1640.4 ;
     RECT  1272.38 1638.3 1807.3 1640.6 ;
     RECT  2406.14 1640.4 2569.54 1640.82 ;
     RECT  2580.86 1621.92 2581.06 1640.82 ;
     RECT  807.74 1638.1 1215.94 1641.46 ;
     RECT  807.74 1641.46 1201.54 1642.52 ;
     RECT  3095.9 1622.96 3110.98 1642.92 ;
     RECT  -70 1608.225 178 1643 ;
     RECT  1272.38 1640.6 1805.38 1645.04 ;
     RECT  2406.14 1640.82 2581.06 1645.44 ;
     RECT  2637.98 1637.88 3070.66 1647.96 ;
     RECT  2606.78 1634.72 2612.26 1649.22 ;
     RECT  1265.18 1645.04 1805.38 1650.08 ;
     RECT  3090.62 1642.92 3110.98 1650.48 ;
     RECT  2637.98 1647.96 3072.1 1651.74 ;
     RECT  2629.82 1651.74 3072.1 1652.36 ;
     RECT  2406.14 1645.44 2587.78 1653 ;
     RECT  1230.14 1638.52 1241.38 1654.28 ;
     RECT  1252.7 1622.56 1252.9 1654.28 ;
     RECT  1215.74 1641.46 1215.94 1654.7 ;
     RECT  1230.14 1654.28 1252.9 1654.7 ;
     RECT  803.9 1642.52 1201.54 1656.8 ;
     RECT  3088.7 1650.48 3110.98 1658.24 ;
     RECT  1262.78 1650.08 1805.38 1659.32 ;
     RECT  3089.18 1658.24 3110.98 1659.5 ;
     RECT  803.9 1656.8 1202.5 1660.58 ;
     RECT  1262.78 1659.32 1805.86 1661.2 ;
     RECT  2406.14 1653 2590.18 1663.08 ;
     RECT  2601.5 1649.22 2612.26 1663.08 ;
     RECT  803.9 1660.58 1204.9 1663.1 ;
     RECT  1215.74 1654.7 1252.9 1663.1 ;
     RECT  803.9 1663.1 1252.9 1665.4 ;
     RECT  2282.3 1659.32 2282.5 1666.66 ;
     RECT  2629.82 1652.36 3070.66 1667.28 ;
     RECT  2406.14 1663.08 2612.26 1669.8 ;
     RECT  3089.66 1659.5 3110.98 1670.64 ;
     RECT  2406.14 1669.8 2613.22 1674.42 ;
     RECT  2629.82 1667.28 3071.14 1674.84 ;
     RECT  2406.14 1674.42 2614.66 1675.68 ;
     RECT  2627.42 1674.84 3071.62 1675.68 ;
     RECT  806.78 1665.4 1252.9 1675.9 ;
     RECT  807.74 1675.9 1252.9 1676.12 ;
     RECT  1262.78 1661.2 1805.38 1676.12 ;
     RECT  3081.5 1670.64 3110.98 1676.72 ;
     RECT  0 1643 178 1681.16 ;
     RECT  190.46 761.78 190.66 1681.16 ;
     RECT  807.74 1676.12 1805.38 1687.46 ;
     RECT  801.98 1687.46 1805.38 1687.88 ;
     RECT  2406.14 1675.68 3071.62 1693.32 ;
     RECT  3088.7 1676.72 3110.98 1698.56 ;
     RECT  2406.14 1693.32 3072.1 1700.88 ;
     RECT  799.1 1687.88 1805.38 1706.56 ;
     RECT  813.5 1706.56 1805.38 1715.58 ;
     RECT  2406.14 1700.88 3081.7 1717.04 ;
     RECT  2406.14 1717.04 3074.02 1720.4 ;
     RECT  799.1 1706.56 802.66 1721.48 ;
     RECT  813.5 1715.58 1807.3 1721.48 ;
     RECT  799.1 1721.48 1807.3 1721.68 ;
     RECT  3093.5 1698.56 3110.98 1723.56 ;
     RECT  803.9 1721.68 1807.3 1723.76 ;
     RECT  2406.14 1720.4 2943.94 1727.12 ;
     RECT  2651.9 1727.12 2943.94 1730.7 ;
     RECT  2953.82 1720.4 3074.02 1730.7 ;
     RECT  803.9 1723.76 1801.54 1733.44 ;
     RECT  247.58 1733.24 247.78 1734.08 ;
     RECT  813.02 1733.44 1801.54 1735.96 ;
     RECT  813.5 1735.96 1801.54 1736.16 ;
     RECT  247.58 1734.08 251.14 1736.6 ;
     RECT  233.18 1608.08 233.38 1736.8 ;
     RECT  813.5 1736.16 1804.42 1737.64 ;
     RECT  244.7 1736.6 251.14 1737.86 ;
     RECT  264.86 1736.6 265.06 1737.86 ;
     RECT  3088.7 1723.56 3110.98 1738.04 ;
     RECT  2051.42 1731.98 2051.62 1738.7 ;
     RECT  1994.3 1724.84 1994.5 1738.9 ;
     RECT  2076.86 1731.56 2077.06 1738.9 ;
     RECT  2406.14 1727.12 2640.58 1739.1 ;
     RECT  2406.14 1739.1 2642.02 1739.94 ;
     RECT  2651.9 1730.7 3074.02 1739.94 ;
     RECT  237.02 1737.86 265.06 1739.96 ;
     RECT  237.02 1739.96 265.54 1741.42 ;
     RECT  2048.06 1738.7 2051.62 1741.64 ;
     RECT  814.46 1737.64 1804.42 1741.84 ;
     RECT  2048.06 1741.64 2052.1 1741.84 ;
     RECT  250.94 1741.42 265.54 1743.94 ;
     RECT  250.94 1743.94 265.06 1744.36 ;
     RECT  712.7 1728.62 712.9 1744.36 ;
     RECT  237.02 1741.42 238.18 1744.78 ;
     RECT  250.94 1744.36 251.14 1745.2 ;
     RECT  2118.14 1738.7 2118.34 1746.04 ;
     RECT  814.46 1741.84 1372.42 1748.36 ;
     RECT  1384.7 1741.84 1804.42 1748.78 ;
     RECT  237.98 1744.78 238.18 1748.98 ;
     RECT  810.14 1748.36 1372.42 1749.7 ;
     RECT  810.62 1749.7 1372.42 1751.08 ;
     RECT  2406.14 1739.94 3074.02 1751.48 ;
     RECT  2406.14 1751.48 2602.18 1755.06 ;
     RECT  810.62 1751.08 1362.34 1756.12 ;
     RECT  2133.98 1745.84 2134.18 1756.54 ;
     RECT  3221.18 1633 3400 1757 ;
     RECT  810.62 1756.12 1233.22 1758.22 ;
     RECT  1245.02 1756.12 1362.34 1759.48 ;
     RECT  2405.66 1755.06 2602.18 1763.04 ;
     RECT  2405.66 1763.04 2603.14 1764.3 ;
     RECT  2613.5 1751.48 3074.02 1764.3 ;
     RECT  1246.46 1759.48 1362.34 1766.2 ;
     RECT  810.62 1758.22 1229.86 1766.84 ;
     RECT  0 1681.16 190.66 1767 ;
     RECT  3221.18 1757 3470 1770.2 ;
     RECT  3220.145 1770.2 3470 1770.225 ;
     RECT  1384.7 1748.78 1804.9 1771.24 ;
     RECT  1246.46 1766.2 1360.42 1772.5 ;
     RECT  3220 1770.225 3470 1773.775 ;
     RECT  2405.66 1764.3 3074.02 1776.26 ;
     RECT  2406.14 1776.26 3074.02 1777.52 ;
     RECT  2159.9 1756.34 2160.1 1778.8 ;
     RECT  2406.62 1777.52 3074.02 1779.62 ;
     RECT  2408.54 1779.62 3074.02 1780.88 ;
     RECT  2409.02 1780.88 3074.02 1781.3 ;
     RECT  2409.5 1781.3 3074.02 1781.72 ;
     RECT  2048.06 1741.84 2048.26 1782.16 ;
     RECT  805.34 1766.84 1229.86 1783 ;
     RECT  1387.1 1771.24 1804.9 1783.42 ;
     RECT  1388.06 1783.42 1804.9 1786.36 ;
     RECT  805.34 1783 1205.86 1789.52 ;
     RECT  1216.7 1783 1229.86 1789.52 ;
     RECT  1267.1 1772.5 1360.42 1791.4 ;
     RECT  1372.22 1751.08 1372.42 1791.4 ;
     RECT  2414.78 1781.72 3074.02 1791.8 ;
     RECT  2414.78 1791.8 2423.14 1792.02 ;
     RECT  2062.46 1741.64 2062.66 1793.08 ;
     RECT  802.46 1789.52 1205.86 1793.3 ;
     RECT  1216.7 1789.52 1231.3 1793.3 ;
     RECT  1246.46 1772.5 1252.9 1794.14 ;
     RECT  1388.06 1786.36 1390.66 1794.56 ;
     RECT  1267.1 1791.4 1297.06 1794.76 ;
     RECT  1307.42 1791.4 1360.42 1794.76 ;
     RECT  2181.5 1778.6 2181.7 1796.44 ;
     RECT  802.46 1793.3 1231.3 1797.08 ;
     RECT  2433.5 1791.8 2538.34 1798.52 ;
     RECT  2414.3 1792.02 2423.14 1799.36 ;
     RECT  801.5 1797.08 1234.66 1801.48 ;
     RECT  -70 1767 190.66 1801.9 ;
     RECT  2077.82 1792.88 2078.02 1801.9 ;
     RECT  2462.78 1798.52 2538.34 1802.94 ;
     RECT  2551.58 1791.8 3074.02 1803.56 ;
     RECT  2372.06 1803.36 2372.26 1803.78 ;
     RECT  2369.66 1803.78 2372.26 1804.2 ;
     RECT  801.5 1801.48 1233.7 1804.64 ;
     RECT  1311.74 1794.76 1360.42 1804.64 ;
     RECT  1311.74 1804.64 1360.9 1805.48 ;
     RECT  1267.1 1794.76 1296.58 1806.32 ;
     RECT  1307.9 1805.48 1360.9 1806.32 ;
     RECT  2414.3 1799.36 2414.5 1806.72 ;
     RECT  2433.5 1798.52 2452.42 1806.72 ;
     RECT  1382.3 1794.56 1390.66 1807.16 ;
     RECT  2109.5 1801.7 2109.7 1807.16 ;
     RECT  797.66 1804.64 1233.7 1807.36 ;
     RECT  2109.5 1807.16 2117.38 1807.36 ;
     RECT  801.5 1807.36 1233.7 1807.78 ;
     RECT  2369.66 1804.2 2381.38 1807.98 ;
     RECT  2395.58 1806.72 2397.22 1807.98 ;
     RECT  2410.94 1806.72 2414.5 1807.98 ;
     RECT  2462.78 1802.94 2540.74 1807.98 ;
     RECT  2551.58 1803.56 3073.54 1807.98 ;
     RECT  801.98 1807.78 1233.7 1809.04 ;
     RECT  1245.5 1794.14 1252.9 1809.04 ;
     RECT  1379.9 1807.16 1390.66 1809.26 ;
     RECT  1376.06 1809.26 1390.66 1809.68 ;
     RECT  2369.66 1807.98 2383.3 1810.5 ;
     RECT  2395.58 1807.98 2414.5 1810.5 ;
     RECT  2369.66 1810.5 2414.5 1810.92 ;
     RECT  2361.5 1810.92 2414.5 1811.34 ;
     RECT  2425.34 1806.72 2452.42 1811.34 ;
     RECT  2462.78 1807.98 3073.54 1811.34 ;
     RECT  1267.1 1806.32 1360.9 1811.36 ;
     RECT  3222 1773.775 3470 1811.725 ;
     RECT  768.86 1743.74 769.06 1811.98 ;
     RECT  3192.86 1760.12 3193.06 1811.98 ;
     RECT  1267.1 1811.36 1365.22 1812.2 ;
     RECT  1376.06 1809.68 1392.1 1812.2 ;
     RECT  3220 1811.725 3470 1812.225 ;
     RECT  1267.1 1812.2 1392.1 1813.46 ;
     RECT  1401.98 1786.36 1804.9 1813.46 ;
     RECT  2358.14 1811.34 2414.5 1813.86 ;
     RECT  2425.34 1811.34 3073.54 1814.06 ;
     RECT  2353.82 1813.86 2415.46 1814.28 ;
     RECT  2425.34 1814.06 2522.02 1814.28 ;
     RECT  701.66 1798.34 701.86 1817.66 ;
     RECT  2117.18 1807.36 2117.38 1817.86 ;
     RECT  801.98 1809.04 1231.3 1819.76 ;
     RECT  2533.34 1814.06 3073.54 1821.62 ;
     RECT  2353.82 1814.28 2522.02 1821.84 ;
     RECT  801.98 1819.76 1237.54 1822.9 ;
     RECT  801.98 1822.9 1231.3 1824.16 ;
     RECT  701.66 1817.66 703.3 1824.38 ;
     RECT  2348.06 1821.84 2522.02 1825.2 ;
     RECT  2533.34 1821.62 2577.22 1825.2 ;
     RECT  2098.46 1781.96 2098.66 1825.42 ;
     RECT  2209.82 1743.74 2210.02 1826.06 ;
     RECT  2181.5 1817.66 2181.7 1826.26 ;
     RECT  2203.1 1826.06 2210.02 1826.26 ;
     RECT  2588.06 1821.62 3073.54 1826.66 ;
     RECT  1888.22 1815.98 1888.42 1826.9 ;
     RECT  3222 1812.225 3470 1827 ;
     RECT  802.46 1824.16 1231.3 1827.52 ;
     RECT  803.42 1827.52 1227.94 1828.9 ;
     RECT  1267.1 1813.46 1804.9 1831.1 ;
     RECT  803.42 1828.9 1227.46 1831.3 ;
     RECT  699.74 1824.38 703.3 1832.36 ;
     RECT  806.78 1831.3 1227.46 1833.4 ;
     RECT  2348.06 1825.2 2577.22 1833.6 ;
     RECT  -70 1801.9 183.46 1837 ;
     RECT  2588.54 1826.66 3073.54 1837.38 ;
     RECT  806.78 1833.4 1224.58 1839.28 ;
     RECT  1266.62 1831.1 1804.9 1839.28 ;
     RECT  2347.1 1833.6 2577.22 1841.16 ;
     RECT  2588.54 1837.38 3074.02 1841.16 ;
     RECT  806.78 1839.28 1224.1 1841.8 ;
     RECT  806.78 1841.8 1223.62 1842.22 ;
     RECT  1182.62 1842.22 1223.62 1842.64 ;
     RECT  806.78 1842.22 1171.78 1843.06 ;
     RECT  2256.86 1796.24 2257.06 1843.28 ;
     RECT  1182.62 1842.64 1216.9 1843.48 ;
     RECT  2256.86 1843.28 2264.26 1843.48 ;
     RECT  2347.1 1841.16 3074.02 1844.72 ;
     RECT  1216.7 1843.48 1216.9 1845.58 ;
     RECT  1911.26 1775.66 1911.46 1845.8 ;
     RECT  1923.26 1838.66 1923.46 1845.8 ;
     RECT  1182.62 1843.48 1202.5 1846.42 ;
     RECT  1182.62 1846.42 1201.54 1846.84 ;
     RECT  1185.02 1846.84 1201.54 1849.36 ;
     RECT  806.78 1843.06 1142.02 1850.2 ;
     RECT  1185.02 1849.36 1194.34 1850.62 ;
     RECT  813.98 1850.2 1141.06 1851.04 ;
     RECT  1189.82 1850.62 1190.5 1853.14 ;
     RECT  1267.1 1839.28 1804.9 1853.36 ;
     RECT  1189.82 1853.14 1190.02 1854.4 ;
     RECT  699.74 1832.36 707.62 1854.62 ;
     RECT  723.74 1831.94 723.94 1855.46 ;
     RECT  694.94 1854.62 707.62 1855.88 ;
     RECT  717.98 1855.46 723.94 1855.88 ;
     RECT  1870.94 1838.24 1871.14 1857.56 ;
     RECT  814.46 1851.04 1141.06 1858.6 ;
     RECT  2347.1 1844.72 3067.78 1860.06 ;
     RECT  820.22 1858.6 1141.06 1860.28 ;
     RECT  2203.58 1826.26 2210.02 1860.5 ;
     RECT  2203.58 1860.5 2213.86 1860.7 ;
     RECT  1264.22 1853.36 1804.9 1861.76 ;
     RECT  2343.74 1860.06 3067.78 1863.62 ;
     RECT  1264.22 1861.76 1811.14 1865.54 ;
     RECT  1840.7 1860.92 1840.9 1868.9 ;
     RECT  820.22 1860.28 1135.78 1869.94 ;
     RECT  1262.78 1865.54 1811.14 1870.36 ;
     RECT  1263.74 1870.36 1811.14 1872.04 ;
     RECT  822.14 1869.94 1135.78 1872.88 ;
     RECT  3093.5 1738.04 3110.98 1874.34 ;
     RECT  822.62 1872.88 1135.78 1876.66 ;
     RECT  1263.74 1872.04 1774.66 1877.08 ;
     RECT  1122.62 1876.66 1135.78 1878.76 ;
     RECT  2343.74 1863.62 3065.86 1878.96 ;
     RECT  1785.02 1872.04 1811.14 1880.02 ;
     RECT  1252.7 1809.04 1252.9 1880.24 ;
     RECT  1263.74 1877.08 1327.78 1880.24 ;
     RECT  822.62 1876.66 1112.26 1880.44 ;
     RECT  2343.26 1878.96 3065.86 1882.32 ;
     RECT  3089.18 1874.34 3110.98 1882.74 ;
     RECT  1122.62 1878.76 1128.58 1883.38 ;
     RECT  827.42 1880.44 1112.26 1884.22 ;
     RECT  1339.1 1877.08 1774.66 1885.28 ;
     RECT  2339.9 1882.32 3067.3 1885.46 ;
     RECT  2264.06 1843.48 2264.26 1886.54 ;
     RECT  2339.9 1885.46 3065.38 1886.72 ;
     RECT  2264.06 1886.54 2271.46 1886.74 ;
     RECT  1252.7 1880.24 1327.78 1886.96 ;
     RECT  827.9 1884.22 1112.26 1887.16 ;
     RECT  1250.3 1886.96 1327.78 1887.8 ;
     RECT  1250.3 1887.8 1329.22 1888.22 ;
     RECT  1339.1 1885.28 1779.94 1888.22 ;
     RECT  827.9 1887.16 1094.5 1888.42 ;
     RECT  835.58 1888.42 1088.26 1888.84 ;
     RECT  835.58 1888.84 1073.86 1890.52 ;
     RECT  835.58 1890.52 866.02 1890.94 ;
     RECT  875.9 1890.52 1073.86 1890.94 ;
     RECT  835.58 1890.94 836.26 1891.78 ;
     RECT  1250.3 1888.22 1779.94 1891.78 ;
     RECT  835.58 1891.78 835.78 1892.2 ;
     RECT  847.1 1890.94 866.02 1892.2 ;
     RECT  847.1 1892.2 863.62 1893.46 ;
     RECT  847.1 1893.46 860.74 1894.72 ;
     RECT  694.94 1855.88 723.94 1894.94 ;
     RECT  852.38 1894.72 860.74 1895.14 ;
     RECT  1112.06 1887.16 1112.26 1895.36 ;
     RECT  1128.38 1883.38 1128.58 1895.36 ;
     RECT  852.38 1895.14 858.82 1895.56 ;
     RECT  875.9 1890.94 1072.42 1895.56 ;
     RECT  679.58 1894.1 679.78 1896.2 ;
     RECT  690.14 1894.94 723.94 1896.2 ;
     RECT  856.7 1895.56 856.9 1896.4 ;
     RECT  882.14 1895.56 1072.42 1896.4 ;
     RECT  3088.7 1882.74 3110.98 1897.64 ;
     RECT  1112.06 1895.36 1128.58 1898.3 ;
     RECT  1154.3 1843.06 1171.78 1898.3 ;
     RECT  1112.06 1898.3 1171.78 1898.72 ;
     RECT  884.54 1896.4 1072.42 1899.34 ;
     RECT  1111.58 1898.72 1171.78 1899.56 ;
     RECT  1252.7 1891.78 1779.94 1900.4 ;
     RECT  1790.3 1880.02 1811.14 1900.4 ;
     RECT  3098.3 1897.64 3110.98 1900.4 ;
     RECT  884.54 1899.34 1071.46 1902.28 ;
     RECT  2341.82 1886.72 3062.98 1902.48 ;
     RECT  1109.18 1899.56 1171.78 1902.5 ;
     RECT  899.9 1902.28 1071.46 1902.7 ;
     RECT  1101.98 1902.5 1171.78 1902.92 ;
     RECT  884.54 1902.28 889.06 1903.12 ;
     RECT  899.9 1902.7 926.98 1903.12 ;
     RECT  937.34 1902.7 1071.46 1903.12 ;
     RECT  888.38 1903.12 889.06 1903.54 ;
     RECT  899.9 1903.12 904.42 1903.54 ;
     RECT  920.54 1903.12 920.74 1903.54 ;
     RECT  941.18 1903.12 1071.46 1904.38 ;
     RECT  2341.82 1902.48 3072.1 1904.78 ;
     RECT  2341.82 1904.78 3067.3 1905 ;
     RECT  941.18 1904.38 1065.7 1905.64 ;
     RECT  679.58 1896.2 723.94 1905.86 ;
     RECT  941.18 1905.64 1058.98 1906.06 ;
     RECT  1101.98 1902.92 1172.26 1906.28 ;
     RECT  1252.7 1900.4 1811.14 1906.7 ;
     RECT  946.46 1906.06 1055.62 1906.9 ;
     RECT  1101.98 1906.28 1173.22 1907.12 ;
     RECT  948.38 1906.9 1055.62 1907.32 ;
     RECT  1101.5 1907.12 1173.22 1907.54 ;
     RECT  3098.3 1900.4 3113.38 1907.54 ;
     RECT  1084.7 1888.84 1088.26 1907.96 ;
     RECT  951.26 1907.32 1055.62 1909.84 ;
     RECT  1101.5 1907.54 1176.1 1910.48 ;
     RECT  952.22 1909.84 1055.62 1910.68 ;
     RECT  1084.22 1907.96 1088.26 1910.9 ;
     RECT  964.22 1910.68 1046.02 1911.1 ;
     RECT  1082.78 1910.9 1088.26 1911.74 ;
     RECT  2209.82 1860.7 2213.86 1912.78 ;
     RECT  1082.78 1911.74 1090.66 1914.26 ;
     RECT  1082.78 1914.26 1091.62 1914.68 ;
     RECT  1247.9 1906.7 1811.14 1914.68 ;
     RECT  1028.54 1911.1 1046.02 1914.88 ;
     RECT  1081.34 1914.68 1091.62 1915.52 ;
     RECT  1101.5 1910.48 1181.86 1915.52 ;
     RECT  1245.98 1914.68 1811.14 1916.78 ;
     RECT  1245.98 1916.78 1815.94 1917.4 ;
     RECT  1031.42 1914.88 1046.02 1918.24 ;
     RECT  1079.9 1915.52 1181.86 1918.46 ;
     RECT  2337.98 1905 3067.3 1919.48 ;
     RECT  899.9 1903.54 900.1 1920.34 ;
     RECT  1073.18 1918.46 1181.86 1921.4 ;
     RECT  3093.98 1907.54 3113.38 1921.4 ;
     RECT  1073.18 1921.4 1182.34 1922.24 ;
     RECT  741.5 1915.1 741.7 1922.44 ;
     RECT  1248.38 1917.4 1815.94 1923.28 ;
     RECT  3092.54 1921.4 3113.38 1923.92 ;
     RECT  1070.3 1922.24 1182.34 1924.76 ;
     RECT  1253.66 1923.28 1815.94 1924.96 ;
     RECT  675.26 1905.86 723.94 1925.6 ;
     RECT  2092.7 1846.22 2092.9 1926.02 ;
     RECT  2107.1 1879.4 2107.3 1926.02 ;
     RECT  2224.7 1912.58 2224.9 1926.02 ;
     RECT  964.7 1911.1 1018.66 1926.22 ;
     RECT  2224.7 1926.02 2232.1 1926.22 ;
     RECT  953.66 1910.68 953.86 1927.06 ;
     RECT  1070.3 1924.76 1184.74 1929.8 ;
     RECT  1065.5 1929.8 1184.74 1930 ;
     RECT  2271.26 1886.74 2271.46 1930 ;
     RECT  973.82 1926.22 1018.66 1933.36 ;
     RECT  1065.5 1930 1183.78 1933.36 ;
     RECT  624.86 1933.16 625.06 1934.42 ;
     RECT  1146.62 1933.36 1183.3 1936.3 ;
     RECT  675.26 1925.6 727.3 1936.72 ;
     RECT  1255.58 1924.96 1815.94 1937.36 ;
     RECT  1146.62 1936.3 1181.86 1937.56 ;
     RECT  1253.18 1937.36 1815.94 1937.78 ;
     RECT  973.82 1933.36 1010.02 1937.98 ;
     RECT  1250.78 1937.78 1815.94 1939.88 ;
     RECT  662.78 1938.2 662.98 1941.14 ;
     RECT  1249.82 1939.88 1815.94 1944.08 ;
     RECT  2231.9 1926.22 2232.1 1944.28 ;
     RECT  1065.5 1933.36 1135.78 1944.5 ;
     RECT  1146.62 1937.56 1180.9 1944.5 ;
     RECT  662.78 1941.14 663.46 1944.92 ;
     RECT  675.26 1936.72 723.94 1944.92 ;
     RECT  980.06 1937.98 1010.02 1945.12 ;
     RECT  981.98 1945.12 1010.02 1946.38 ;
     RECT  2341.82 1919.48 3067.3 1947.2 ;
     RECT  1244.06 1944.08 1815.94 1948.28 ;
     RECT  900.38 1920.56 900.58 1948.9 ;
     RECT  3222 1827 3400 1951 ;
     RECT  3091.58 1923.92 3113.38 1951.1 ;
     RECT  1065.5 1944.5 1180.9 1952.68 ;
     RECT  1065.5 1952.68 1176.1 1953.32 ;
     RECT  1238.3 1948.28 1815.94 1953.52 ;
     RECT  2120.06 1825.22 2120.26 1954.78 ;
     RECT  1245.02 1953.52 1247.14 1955.62 ;
     RECT  982.46 1946.38 1010.02 1956.46 ;
     RECT  0 1837 183.46 1961 ;
     RECT  1064.54 1953.32 1176.1 1961.08 ;
     RECT  3091.58 1951.1 3113.86 1961.28 ;
     RECT  2347.1 1947.2 3067.3 1962.32 ;
     RECT  1245.98 1955.62 1247.14 1963.4 ;
     RECT  1260.38 1953.52 1815.94 1963.4 ;
     RECT  1064.54 1961.08 1143.46 1963.6 ;
     RECT  3089.18 1961.28 3113.86 1963.8 ;
     RECT  1064.54 1963.6 1094.02 1964.02 ;
     RECT  2369.18 1962.32 3067.3 1964.22 ;
     RECT  3222 1951 3470 1964.225 ;
     RECT  2282.3 1929.8 2282.5 1965.7 ;
     RECT  3220 1964.225 3470 1967.6 ;
     RECT  1064.54 1964.02 1088.74 1967.8 ;
     RECT  1154.78 1961.08 1176.1 1967.8 ;
     RECT  3219.26 1967.6 3470 1967.8 ;
     RECT  982.94 1956.46 1010.02 1968.64 ;
     RECT  2348.54 1962.32 2359.3 1969.46 ;
     RECT  2349.02 1969.46 2359.3 1969.88 ;
     RECT  1104.38 1963.6 1143.46 1971.38 ;
     RECT  1154.78 1967.8 1167.94 1971.38 ;
     RECT  1064.54 1967.8 1073.86 1971.58 ;
     RECT  2369.18 1964.22 3069.22 1972.4 ;
     RECT  2355.74 1969.88 2359.3 1974.3 ;
     RECT  2369.18 1972.4 3068.26 1974.3 ;
     RECT  624.86 1934.42 626.5 1974.32 ;
     RECT  662.78 1944.92 723.94 1974.32 ;
     RECT  1104.38 1971.38 1167.94 1975.36 ;
     RECT  1245.98 1963.4 1815.94 1975.36 ;
     RECT  662.78 1974.32 724.42 1975.58 ;
     RECT  1246.46 1975.36 1815.94 1976.2 ;
     RECT  3088.7 1963.8 3113.86 1976.84 ;
     RECT  662.78 1975.58 725.86 1977.68 ;
     RECT  982.94 1968.64 1006.66 1977.88 ;
     RECT  1252.7 1976.2 1815.94 1977.88 ;
     RECT  1106.78 1975.36 1167.94 1978.52 ;
     RECT  1106.78 1978.52 1170.82 1978.72 ;
     RECT  1040.06 1918.24 1046.02 1979.56 ;
     RECT  1260.38 1977.88 1815.94 1981.66 ;
     RECT  1107.74 1978.72 1134.82 1982.5 ;
     RECT  662.78 1977.68 726.82 1982.92 ;
     RECT  982.94 1977.88 993.7 1982.92 ;
     RECT  1107.74 1982.5 1110.34 1982.92 ;
     RECT  1120.22 1982.5 1134.82 1982.92 ;
     RECT  1148.54 1978.72 1170.82 1982.92 ;
     RECT  1265.66 1981.66 1815.94 1982.92 ;
     RECT  624.86 1974.32 629.86 1983.14 ;
     RECT  1064.54 1971.58 1065.7 1983.76 ;
     RECT  1110.14 1982.92 1110.34 1983.76 ;
     RECT  2355.74 1974.3 3068.26 1984.8 ;
     RECT  3085.34 1976.84 3113.86 1984.82 ;
     RECT  1121.66 1982.92 1134.82 1985.44 ;
     RECT  1155.26 1982.92 1170.82 1985.44 ;
     RECT  1267.1 1982.92 1815.94 1985.44 ;
     RECT  982.94 1982.92 983.14 1985.86 ;
     RECT  662.78 1982.92 724.42 1986.28 ;
     RECT  1125.98 1985.44 1134.82 1986.28 ;
     RECT  1155.26 1985.44 1167.94 1986.28 ;
     RECT  1267.58 1985.44 1815.94 1986.28 ;
     RECT  1274.78 1986.28 1815.94 1986.7 ;
     RECT  2355.74 1984.8 3068.74 1986.92 ;
     RECT  3078.62 1984.82 3113.86 1986.92 ;
     RECT  1155.26 1986.28 1155.46 1987.12 ;
     RECT  1006.46 1977.88 1006.66 1988.8 ;
     RECT  759.74 1983.56 759.94 1989.64 ;
     RECT  1040.06 1979.56 1040.26 1990.06 ;
     RECT  888.86 1903.54 889.06 1990.48 ;
     RECT  993.5 1982.92 993.7 1990.48 ;
     RECT  1275.26 1986.7 1815.94 1991.32 ;
     RECT  -70 1961 183.46 1995.94 ;
     RECT  -70 1995.94 180 1996.225 ;
     RECT  2355.74 1986.92 3113.86 2000.12 ;
     RECT  662.78 1986.28 719.62 2001.2 ;
     RECT  762.62 1990.7 762.82 2001.4 ;
     RECT  657.5 2001.2 719.62 2001.5 ;
     RECT  1084.22 1967.8 1088.74 2001.5 ;
     RECT  1128.86 1986.28 1134.82 2001.5 ;
     RECT  2355.74 2000.12 3046.66 2001.7 ;
     RECT  3056.54 2000.12 3113.86 2003.06 ;
     RECT  2359.58 2001.7 3046.66 2003.48 ;
     RECT  3222 1967.8 3470 2005.725 ;
     RECT  3207.26 1967.6 3207.46 2005.82 ;
     RECT  3220 2005.725 3470 2006.225 ;
     RECT  1292.06 1991.32 1815.94 2009.8 ;
     RECT  1292.06 2009.8 1325.38 2010.64 ;
     RECT  1335.26 2009.8 1815.94 2011.9 ;
     RECT  432.86 831.92 433.06 2012.12 ;
     RECT  1083.74 2001.5 1088.74 2012.32 ;
     RECT  1128.38 2001.5 1134.82 2012.32 ;
     RECT  1335.26 2011.9 1362.34 2012.32 ;
     RECT  622.46 1983.14 629.86 2012.54 ;
     RECT  1088.54 2012.32 1088.74 2012.74 ;
     RECT  1335.26 2012.32 1360.9 2013.16 ;
     RECT  3057.5 2003.06 3113.86 2013.36 ;
     RECT  2359.58 2003.48 3046.18 2014.2 ;
     RECT  3056.06 2013.36 3113.86 2014.2 ;
     RECT  932.06 1980.62 932.26 2019.46 ;
     RECT  2292.86 1965.5 2293.06 2020.72 ;
     RECT  2303.9 2020.52 2304.58 2020.72 ;
     RECT  3222 2006.225 3470 2021 ;
     RECT  2249.66 1944.08 2249.86 2021.56 ;
     RECT  2359.58 2014.2 3113.86 2022.5 ;
     RECT  3044.06 2022.5 3113.86 2022.8 ;
     RECT  3047.9 2022.8 3113.86 2026.16 ;
     RECT  3057.02 2026.16 3113.86 2026.58 ;
     RECT  2192.06 1954.58 2192.26 2027.44 ;
     RECT  586.94 1983.98 587.14 2030.3 ;
     RECT  657.02 2001.5 719.62 2030.3 ;
     RECT  2359.58 2022.5 3034.18 2030.36 ;
     RECT  3062.3 2026.58 3113.86 2030.36 ;
     RECT  586.94 2030.3 587.62 2030.5 ;
     RECT  -70 1996.225 178 2031 ;
     RECT  3065.66 2030.36 3113.86 2033.72 ;
     RECT  2397.98 2030.36 3034.18 2037.92 ;
     RECT  2304.38 2020.72 2304.58 2037.94 ;
     RECT  1165.82 1986.28 1166.02 2039.2 ;
     RECT  2359.58 2030.36 2388.1 2041.08 ;
     RECT  2397.98 2037.92 3031.3 2041.08 ;
     RECT  920.22 2038.12 920.42 2043.58 ;
     RECT  1335.26 2013.16 1359.94 2044.04 ;
     RECT  3070.94 2033.72 3113.86 2044.46 ;
     RECT  2359.58 2041.08 3031.3 2045.06 ;
     RECT  3029.66 2045.06 3031.3 2045.48 ;
     RECT  3029.66 2045.48 3029.86 2046.32 ;
     RECT  920.22 2043.58 925.22 2046.52 ;
     RECT  1332.38 2044.04 1359.94 2046.56 ;
     RECT  1374.14 2011.9 1815.94 2046.56 ;
     RECT  953.82 2046.52 954.02 2046.94 ;
     RECT  562.46 1220 562.66 2046.98 ;
     RECT  575.9 2000.78 576.1 2046.98 ;
     RECT  1332.38 2046.56 1815.94 2046.98 ;
     RECT  2359.58 2045.06 3017.86 2049.26 ;
     RECT  562.46 2046.98 576.1 2049.5 ;
     RECT  587.42 2030.5 587.62 2049.5 ;
     RECT  3016.7 2049.26 3016.9 2049.68 ;
     RECT  1064.54 1983.76 1064.74 2049.7 ;
     RECT  920.22 2046.52 930.02 2050.3 ;
     RECT  562.46 2049.5 587.62 2050.54 ;
     RECT  806.94 2033.08 807.14 2050.72 ;
     RECT  920.22 2050.3 931.46 2050.72 ;
     RECT  1329.98 2046.98 1815.94 2050.76 ;
     RECT  886.62 2050.72 886.82 2051.14 ;
     RECT  857.82 2035.6 858.02 2051.56 ;
     RECT  868.86 2050.72 869.06 2051.56 ;
     RECT  953.82 2046.94 962.18 2051.56 ;
     RECT  915.9 2050.72 937.7 2053.24 ;
     RECT  949.5 2051.56 962.18 2053.24 ;
     RECT  882.3 2051.14 887.78 2054.08 ;
     RECT  899.58 2043.16 899.78 2054.08 ;
     RECT  833.34 2048.2 833.54 2054.5 ;
     RECT  857.82 2051.56 869.06 2054.5 ;
     RECT  882.3 2054.08 899.78 2054.5 ;
     RECT  803.1 2050.72 807.14 2054.92 ;
     RECT  819.9 2040.64 820.1 2054.92 ;
     RECT  833.34 2054.5 839.3 2054.92 ;
     RECT  857.82 2054.5 869.54 2054.92 ;
     RECT  881.34 2054.5 899.78 2054.92 ;
     RECT  915.9 2053.24 962.18 2054.92 ;
     RECT  833.34 2054.92 842.66 2055.76 ;
     RECT  2359.58 2049.26 3005.38 2055.98 ;
     RECT  2260.7 2021.36 2260.9 2058.1 ;
     RECT  803.1 2054.92 820.1 2058.28 ;
     RECT  833.34 2055.76 843.62 2058.28 ;
     RECT  2359.58 2055.98 3004.9 2058.5 ;
     RECT  792.54 2058.28 820.1 2058.7 ;
     RECT  829.98 2058.28 843.62 2058.7 ;
     RECT  857.82 2054.92 903.14 2058.7 ;
     RECT  915.9 2054.92 967.94 2059.12 ;
     RECT  856.38 2058.7 903.62 2059.54 ;
     RECT  914.94 2059.12 967.94 2059.54 ;
     RECT  2359.58 2058.5 3003.94 2059.98 ;
     RECT  2357.66 2059.98 3003.94 2060.4 ;
     RECT  2356.7 2060.4 3003.94 2060.6 ;
     RECT  1292.06 2010.64 1317.22 2061.68 ;
     RECT  1329.5 2050.76 1815.94 2061.68 ;
     RECT  792.54 2058.7 843.62 2062.06 ;
     RECT  2975.9 2060.6 3003.94 2062.28 ;
     RECT  765.18 2062.06 766.34 2062.48 ;
     RECT  791.1 2062.06 843.62 2062.48 ;
     RECT  761.82 2062.48 769.22 2063.32 ;
     RECT  791.1 2062.48 844.1 2063.32 ;
     RECT  2975.9 2062.28 3000.58 2063.54 ;
     RECT  2356.7 2060.6 2965.54 2063.76 ;
     RECT  761.82 2063.32 844.1 2063.94 ;
     RECT  2975.9 2063.54 2999.14 2063.96 ;
     RECT  856.38 2059.54 973.22 2065 ;
     RECT  2975.9 2063.96 2996.26 2065.64 ;
     RECT  744.06 2061.64 744.26 2065.84 ;
     RECT  761.82 2063.94 776.42 2065.84 ;
     RECT  789.18 2063.94 844.1 2065.84 ;
     RECT  856.38 2065 975.14 2065.84 ;
     RECT  657.02 2030.3 720.1 2066.5 ;
     RECT  789.18 2065.84 975.14 2066.68 ;
     RECT  789.18 2066.68 976.1 2067.1 ;
     RECT  987.9 2065.84 988.1 2067.1 ;
     RECT  2353.82 2063.76 2965.54 2067.54 ;
     RECT  789.18 2067.1 990.02 2068.36 ;
     RECT  587.42 2050.54 587.62 2068.4 ;
     RECT  587.42 2068.4 596.26 2068.82 ;
     RECT  587.42 2068.82 601.54 2069.24 ;
     RECT  587.42 2069.24 610.66 2070.5 ;
     RECT  622.46 2012.54 637.06 2070.5 ;
     RECT  2352.86 2067.54 2965.54 2071.32 ;
     RECT  2975.9 2065.64 2995.3 2071.32 ;
     RECT  569.18 2050.54 576.1 2073.44 ;
     RECT  587.42 2070.5 637.06 2073.44 ;
     RECT  744.06 2065.84 776.42 2073.82 ;
     RECT  744.06 2073.82 777.86 2074.66 ;
     RECT  744.06 2074.66 778.34 2075.92 ;
     RECT  789.18 2068.36 992.9 2075.92 ;
     RECT  554.3 2076.38 554.5 2076.8 ;
     RECT  569.18 2073.44 577.06 2076.8 ;
     RECT  744.06 2075.92 992.9 2077.18 ;
     RECT  2328.86 2037.74 2329.06 2077.22 ;
     RECT  2282.3 2057.9 2282.5 2077.42 ;
     RECT  744.06 2077.18 998.66 2078.44 ;
     RECT  2171.9 1877.3 2172.1 2078.48 ;
     RECT  3207.26 2005.82 3207.94 2079.1 ;
     RECT  2351.42 2071.32 2995.3 2079.72 ;
     RECT  554.3 2076.8 577.06 2080.79 ;
     RECT  586.94 2073.44 637.06 2080.79 ;
     RECT  741.18 2078.44 998.66 2080.96 ;
     RECT  2349.98 2079.72 2995.3 2083.5 ;
     RECT  741.18 2080.96 1001.54 2084.74 ;
     RECT  537.98 2084.36 538.18 2084.78 ;
     RECT  554.3 2080.79 637.06 2084.78 ;
     RECT  740.7 2084.74 1001.54 2086 ;
     RECT  738.3 2086 1001.54 2086.84 ;
     RECT  1011.26 1989.44 1011.46 2086.84 ;
     RECT  2349.02 2083.5 2995.3 2087.48 ;
     RECT  529.82 2084.78 538.18 2087.72 ;
     RECT  738.3 2086.84 1011.46 2088.1 ;
     RECT  525.02 2087.72 538.18 2088.14 ;
     RECT  525.02 2088.14 540.1 2088.56 ;
     RECT  552.38 2084.78 637.06 2088.56 ;
     RECT  646.94 2044.46 647.14 2088.98 ;
     RECT  657.02 2066.5 715.78 2088.98 ;
     RECT  729.66 2088.1 1011.46 2089.36 ;
     RECT  2349.98 2087.48 2995.3 2090.42 ;
     RECT  2351.42 2090.42 2995.3 2090.84 ;
     RECT  728.7 2089.36 1011.46 2091.7 ;
     RECT  2352.38 2090.84 2995.3 2093.58 ;
     RECT  523.58 2088.56 637.06 2095.28 ;
     RECT  523.1 2095.28 637.06 2096.12 ;
     RECT  522.14 2096.12 637.06 2096.32 ;
     RECT  728.7 2091.7 1002.98 2096.7 ;
     RECT  522.14 2096.32 589.06 2096.74 ;
     RECT  599.9 2096.32 637.06 2096.74 ;
     RECT  2352.38 2093.58 2996.74 2098.2 ;
     RECT  522.14 2096.74 588.58 2100.1 ;
     RECT  600.38 2096.74 637.06 2100.52 ;
     RECT  522.14 2100.1 587.62 2100.94 ;
     RECT  2352.38 2098.2 2997.7 2101.56 ;
     RECT  2352.38 2101.56 3000.58 2102.6 ;
     RECT  646.94 2088.98 715.78 2102.62 ;
     RECT  2352.38 2102.6 2992.42 2104.7 ;
     RECT  2352.38 2104.7 2990.5 2105.76 ;
     RECT  1134.62 2012.32 1134.82 2105.98 ;
     RECT  2350.46 2105.76 2990.5 2108.48 ;
     RECT  2325.02 2077.22 2329.06 2109.34 ;
     RECT  2350.46 2108.48 2988.1 2109.56 ;
     RECT  519.74 2108.3 519.94 2110.82 ;
     RECT  529.82 2100.94 587.62 2110.82 ;
     RECT  601.34 2100.52 637.06 2110.82 ;
     RECT  2343.26 2109.56 2988.1 2111 ;
     RECT  519.74 2110.82 587.62 2111.24 ;
     RECT  597.5 2110.82 637.06 2111.24 ;
     RECT  2343.26 2111 2986.66 2112.68 ;
     RECT  2343.26 2112.68 2984.74 2113.94 ;
     RECT  2343.26 2113.94 2984.26 2114.36 ;
     RECT  728.7 2096.7 1001.54 2114.56 ;
     RECT  2343.26 2114.36 2980.9 2114.78 ;
     RECT  519.74 2111.24 637.06 2114.8 ;
     RECT  574.94 2114.8 637.06 2115.44 ;
     RECT  646.94 2102.62 706.34 2115.44 ;
     RECT  2343.26 2114.78 2762.5 2116.88 ;
     RECT  1292.06 2061.68 1815.94 2116.9 ;
     RECT  3192.86 2078.9 3193.06 2116.9 ;
     RECT  519.74 2114.8 563.62 2118.8 ;
     RECT  511.1 2118.8 563.62 2119 ;
     RECT  725.34 2114.56 1001.54 2119.38 ;
     RECT  1296.86 2116.9 1815.94 2121.94 ;
     RECT  511.1 2119 562.66 2122.16 ;
     RECT  728.7 2119.38 1001.54 2122.32 ;
     RECT  574.94 2115.44 706.34 2122.36 ;
     RECT  728.7 2122.32 997.7 2122.74 ;
     RECT  616.22 2122.36 706.34 2122.78 ;
     RECT  2772.38 2114.78 2980.9 2124.44 ;
     RECT  730.62 2122.74 997.7 2124.84 ;
     RECT  2772.86 2124.44 2971.3 2125.28 ;
     RECT  618.62 2122.78 706.34 2126.74 ;
     RECT  1008.54 2122.54 1009.22 2127.16 ;
     RECT  1020.06 2125.06 1020.26 2127.16 ;
     RECT  3169.82 2116.7 3170.02 2127.82 ;
     RECT  574.94 2122.36 604.9 2129.5 ;
     RECT  507.26 2122.16 562.66 2129.72 ;
     RECT  574.94 2129.5 601.06 2129.72 ;
     RECT  1008.54 2127.16 1020.26 2130.1 ;
     RECT  1035.9 2127.58 1036.1 2130.1 ;
     RECT  1052.22 2126.74 1052.42 2130.1 ;
     RECT  1062.3 2129.68 1062.5 2130.1 ;
     RECT  1008.54 2130.1 1036.1 2130.52 ;
     RECT  1052.22 2130.1 1062.5 2130.52 ;
     RECT  1086.3 2130.1 1086.5 2130.52 ;
     RECT  1297.82 2121.94 1815.94 2131.18 ;
     RECT  1086.3 2130.52 1086.98 2131.36 ;
     RECT  507.26 2129.72 601.06 2133.28 ;
     RECT  1008.54 2130.52 1062.5 2133.88 ;
     RECT  1086.3 2131.36 1087.46 2133.88 ;
     RECT  618.62 2126.74 710.66 2134.12 ;
     RECT  1086.3 2133.88 1093.22 2134.3 ;
     RECT  3070.46 2044.46 3113.86 2134.54 ;
     RECT  621.02 2134.12 710.66 2134.96 ;
     RECT  2983.58 2132.66 2985.22 2134.96 ;
     RECT  1080.06 2134.3 1093.22 2135.14 ;
     RECT  1105.98 2134.3 1106.18 2135.14 ;
     RECT  730.62 2124.84 997.22 2135.56 ;
     RECT  1008.54 2133.88 1063.46 2135.56 ;
     RECT  1074.3 2135.14 1093.22 2135.56 ;
     RECT  2772.86 2125.28 2970.82 2136.42 ;
     RECT  730.62 2135.56 1063.46 2136.82 ;
     RECT  1073.82 2135.56 1093.22 2136.82 ;
     RECT  1105.5 2135.14 1106.18 2136.82 ;
     RECT  1117.02 2136.4 1117.22 2136.82 ;
     RECT  2983.58 2134.96 2984.74 2137.06 ;
     RECT  508.7 2133.28 601.06 2137.48 ;
     RECT  2984.06 2137.06 2984.74 2137.48 ;
     RECT  730.62 2136.82 1093.22 2137.66 ;
     RECT  1105.5 2136.82 1117.22 2137.66 ;
     RECT  1131.9 2137.24 1132.1 2137.66 ;
     RECT  2984.54 2137.48 2984.74 2137.9 ;
     RECT  725.82 2137.66 1093.22 2138.08 ;
     RECT  1105.5 2137.66 1132.58 2138.08 ;
     RECT  1142.46 2137.66 1142.66 2138.08 ;
     RECT  1153.02 2138.5 1153.22 2139.34 ;
     RECT  1174.62 2131.36 1174.82 2139.76 ;
     RECT  2770.94 2136.42 2970.82 2141.24 ;
     RECT  1152.54 2139.34 1153.22 2141.44 ;
     RECT  511.1 2137.48 601.06 2141.68 ;
     RECT  1152.54 2141.44 1154.18 2141.86 ;
     RECT  1166.46 2139.76 1174.82 2141.86 ;
     RECT  543.26 2141.68 601.06 2142.1 ;
     RECT  725.82 2138.08 1142.66 2142.7 ;
     RECT  1152.54 2141.86 1174.82 2142.7 ;
     RECT  2770.94 2141.24 2960.26 2143.34 ;
     RECT  547.1 2142.1 601.06 2143.58 ;
     RECT  2970.62 2141.24 2970.82 2144.6 ;
     RECT  2328.86 2109.34 2329.06 2144.62 ;
     RECT  621.02 2134.96 621.22 2144.84 ;
     RECT  632.54 2134.96 710.66 2144.84 ;
     RECT  3222 2021 3400 2145 ;
     RECT  511.1 2141.68 526.18 2145.04 ;
     RECT  513.02 2145.04 526.18 2145.88 ;
     RECT  2343.26 2116.88 2757.22 2146.92 ;
     RECT  547.1 2143.58 603.94 2147.98 ;
     RECT  725.82 2142.7 1174.82 2148.78 ;
     RECT  513.02 2145.88 520.9 2148.82 ;
     RECT  568.7 2147.98 603.94 2149.04 ;
     RECT  517.34 2148.82 520.9 2149.24 ;
     RECT  547.1 2147.98 555.94 2149.24 ;
     RECT  568.7 2149.04 605.38 2149.24 ;
     RECT  547.1 2149.24 547.3 2149.66 ;
     RECT  1298.3 2131.18 1815.94 2149.84 ;
     RECT  2343.26 2146.92 2758.18 2150.7 ;
     RECT  2770.94 2143.34 2959.78 2150.7 ;
     RECT  2343.26 2150.7 2959.78 2154.48 ;
     RECT  2343.26 2154.48 2960.74 2154.9 ;
     RECT  0 2031 178 2155 ;
     RECT  725.82 2148.78 1174.34 2156.56 ;
     RECT  621.02 2144.84 710.66 2156.6 ;
     RECT  459.74 635.78 459.94 2157.44 ;
     RECT  481.82 1033.1 482.02 2157.44 ;
     RECT  2343.26 2154.9 2963.14 2157.84 ;
     RECT  3222 2145 3470 2158.225 ;
     RECT  2343.26 2157.84 2963.62 2158.88 ;
     RECT  2914.46 2158.88 2963.62 2159.3 ;
     RECT  475.1 2157.44 482.02 2159.96 ;
     RECT  572.06 2149.24 605.38 2159.96 ;
     RECT  615.26 2156.6 710.66 2159.96 ;
     RECT  2822.78 2158.88 2902.18 2160.98 ;
     RECT  3207.26 2079.1 3207.46 2161.22 ;
     RECT  3220 2158.225 3470 2161.22 ;
     RECT  3219.26 2161.22 3470 2161.42 ;
     RECT  3220 2161.42 3470 2161.775 ;
     RECT  2789.18 2158.88 2810.98 2162.24 ;
     RECT  2914.46 2159.3 2963.14 2162.24 ;
     RECT  2914.94 2162.24 2963.14 2163.08 ;
     RECT  517.34 2149.24 518.98 2163.74 ;
     RECT  2919.26 2163.08 2963.14 2163.92 ;
     RECT  451.1 2157.44 459.94 2164.16 ;
     RECT  475.1 2159.96 491.62 2164.16 ;
     RECT  503.42 2163.74 503.62 2164.16 ;
     RECT  516.86 2163.74 518.98 2164.16 ;
     RECT  723.42 2156.56 1174.34 2164.96 ;
     RECT  2926.94 2163.92 2963.14 2166.02 ;
     RECT  2343.26 2158.88 2777.38 2166.04 ;
     RECT  2343.26 2166.04 2775.94 2166.44 ;
     RECT  2822.78 2160.98 2901.22 2166.44 ;
     RECT  2927.9 2166.02 2963.14 2166.44 ;
     RECT  2927.9 2166.44 2960.26 2166.86 ;
     RECT  428.06 2012.12 433.06 2167.1 ;
     RECT  2343.26 2166.44 2773.06 2167.28 ;
     RECT  2927.9 2166.86 2941.06 2167.28 ;
     RECT  723.42 2164.96 1174.82 2167.9 ;
     RECT  427.58 2167.1 433.06 2167.94 ;
     RECT  451.1 2164.16 518.98 2167.94 ;
     RECT  446.3 2167.94 518.98 2168.78 ;
     RECT  2927.9 2167.28 2939.62 2168.96 ;
     RECT  2791.1 2162.24 2810.98 2169.18 ;
     RECT  2822.78 2166.44 2898.82 2169.18 ;
     RECT  2950.94 2166.86 2960.26 2169.38 ;
     RECT  2930.3 2168.96 2939.62 2169.8 ;
     RECT  2950.94 2169.38 2956.9 2169.8 ;
     RECT  2930.3 2169.8 2938.18 2170.22 ;
     RECT  2930.3 2170.22 2933.38 2171.48 ;
     RECT  427.58 2167.94 436.42 2171.72 ;
     RECT  446.3 2168.78 525.7 2171.72 ;
     RECT  427.58 2171.72 525.7 2171.92 ;
     RECT  723.42 2167.9 1175.78 2172.1 ;
     RECT  2791.1 2169.18 2898.82 2172.14 ;
     RECT  572.06 2159.96 710.66 2172.56 ;
     RECT  723.42 2172.1 1177.22 2174.82 ;
     RECT  2343.26 2167.28 2767.3 2174.86 ;
     RECT  568.22 2172.56 710.66 2175.5 ;
     RECT  723.42 2174.82 1176.74 2175.66 ;
     RECT  2786.3 2172.14 2898.82 2176.74 ;
     RECT  562.46 2175.5 710.66 2176.92 ;
     RECT  2786.3 2176.74 2899.78 2176.94 ;
     RECT  2930.3 2171.48 2930.5 2176.94 ;
     RECT  2348.06 2174.86 2767.3 2177.16 ;
     RECT  2797.34 2176.94 2899.78 2177.16 ;
     RECT  2797.34 2177.16 2901.7 2177.78 ;
     RECT  428.06 2171.92 525.7 2178.86 ;
     RECT  537.5 2178.44 537.7 2178.86 ;
     RECT  723.42 2175.66 1175.3 2179.66 ;
     RECT  2797.34 2177.78 2896.42 2181.14 ;
     RECT  2348.06 2177.16 2769.22 2181.56 ;
     RECT  2867.42 2181.14 2895.94 2181.56 ;
     RECT  2868.38 2181.56 2874.34 2181.98 ;
     RECT  2874.14 2181.98 2874.34 2182.4 ;
     RECT  2887.1 2181.56 2894.5 2182.4 ;
     RECT  3207.26 2161.22 3207.94 2182.42 ;
     RECT  428.06 2178.86 537.7 2183.06 ;
     RECT  2797.34 2181.14 2856.58 2184.08 ;
     RECT  2800.22 2184.08 2856.58 2184.5 ;
     RECT  2851.1 2184.5 2856.58 2184.92 ;
     RECT  2348.06 2181.56 2541.7 2184.94 ;
     RECT  722.46 2179.66 1175.3 2186.38 ;
     RECT  428.06 2183.06 539.14 2186.84 ;
     RECT  562.46 2176.92 706.34 2187.04 ;
     RECT  562.46 2187.04 617.86 2187.68 ;
     RECT  -70 2155 178 2188.145 ;
     RECT  2786.3 2176.94 2786.5 2188.72 ;
     RECT  2805.98 2184.5 2840.26 2189.12 ;
     RECT  428.06 2186.84 546.34 2189.78 ;
     RECT  428.06 2189.78 550.66 2190.2 ;
     RECT  561.5 2187.68 617.86 2190.2 ;
     RECT  428.06 2190.2 617.86 2190.82 ;
     RECT  -70 2188.145 180 2191.46 ;
     RECT  1236.06 2166.64 1236.26 2191.84 ;
     RECT  2812.7 2189.12 2840.26 2192.48 ;
     RECT  2349.5 2184.94 2541.7 2192.9 ;
     RECT  2812.7 2192.48 2827.3 2192.9 ;
     RECT  2028.38 2062.94 2028.58 2193.14 ;
     RECT  2840.06 2192.48 2840.26 2193.32 ;
     RECT  440.06 2190.82 617.86 2194.6 ;
     RECT  722.46 2186.38 1176.26 2194.98 ;
     RECT  2815.1 2192.9 2821.06 2195 ;
     RECT  -70 2191.46 180.1 2195.86 ;
     RECT  2816.54 2195 2821.06 2196.26 ;
     RECT  2349.5 2192.9 2538.82 2196.28 ;
     RECT  2551.58 2181.56 2769.22 2196.48 ;
     RECT  2816.54 2196.26 2816.74 2196.68 ;
     RECT  442.46 2194.6 617.86 2197.76 ;
     RECT  627.74 2187.04 706.34 2197.76 ;
     RECT  2050.94 1912.58 2051.14 2198.6 ;
     RECT  2548.7 2196.48 2769.22 2199.2 ;
     RECT  1293.18 2149.84 1815.94 2199.44 ;
     RECT  1825.82 1846.64 1826.02 2199.44 ;
     RECT  3221.18 2161.775 3470 2199.725 ;
     RECT  3220 2199.725 3470 2200.07 ;
     RECT  442.46 2197.76 706.34 2202.16 ;
     RECT  3219.74 2200.07 3470 2203 ;
     RECT  2710.94 2199.2 2769.22 2204.24 ;
     RECT  723.9 2194.98 1176.26 2205.28 ;
     RECT  723.42 2205.28 1176.26 2205.9 ;
     RECT  2548.7 2199.2 2701.06 2206.76 ;
     RECT  2357.66 2196.28 2538.82 2207.82 ;
     RECT  2548.7 2206.76 2696.74 2207.82 ;
     RECT  723.42 2205.9 1173.86 2210.1 ;
     RECT  2710.94 2204.24 2760.1 2211.38 ;
     RECT  723.9 2210.1 1169.54 2212.2 ;
     RECT  3070.46 2134.54 3113.38 2212.24 ;
     RECT  2710.94 2211.38 2759.14 2214.32 ;
     RECT  446.3 2202.16 706.34 2214.52 ;
     RECT  2710.94 2214.32 2757.7 2214.96 ;
     RECT  3221.18 2203 3470 2215 ;
     RECT  446.3 2214.52 707.3 2216.86 ;
     RECT  1228.86 2191.84 1236.26 2217.04 ;
     RECT  2357.66 2207.82 2696.74 2217.9 ;
     RECT  454.46 2216.86 707.3 2219.98 ;
     RECT  2357.66 2217.9 2697.22 2220 ;
     RECT  2707.1 2214.96 2757.7 2220 ;
     RECT  1977.5 1872.26 1977.7 2221.28 ;
     RECT  2357.66 2220 2757.7 2221.88 ;
     RECT  723.9 2212.2 1167.62 2222.08 ;
     RECT  723.9 2222.08 1168.1 2222.28 ;
     RECT  2721.02 2221.88 2757.7 2223.56 ;
     RECT  2704.22 2221.88 2711.14 2223.98 ;
     RECT  454.46 2219.98 710.66 2224.84 ;
     RECT  3070.46 2212.24 3112.42 2224.84 ;
     RECT  -70 2195.86 178 2225 ;
     RECT  2721.02 2223.56 2750.98 2225.24 ;
     RECT  2357.66 2221.88 2693.38 2225.66 ;
     RECT  2704.22 2223.98 2709.22 2225.66 ;
     RECT  464.54 2224.84 710.66 2225.68 ;
     RECT  2357.66 2225.66 2623.78 2226.5 ;
     RECT  2635.1 2225.66 2693.38 2226.5 ;
     RECT  2636.06 2226.5 2693.38 2226.92 ;
     RECT  2705.18 2225.66 2708.26 2226.92 ;
     RECT  2750.78 2225.24 2750.98 2227.34 ;
     RECT  2636.54 2226.92 2691.94 2227.76 ;
     RECT  2708.06 2226.92 2708.26 2227.76 ;
     RECT  723.9 2222.28 1167.62 2228.16 ;
     RECT  2636.54 2227.76 2678.02 2228.18 ;
     RECT  2640.38 2228.18 2678.02 2229.86 ;
     RECT  2691.74 2227.76 2691.94 2229.86 ;
     RECT  2721.02 2225.24 2740.9 2229.86 ;
     RECT  2728.7 2229.86 2740.9 2230.7 ;
     RECT  2640.38 2229.86 2643.94 2231.12 ;
     RECT  2657.66 2229.86 2678.02 2231.12 ;
     RECT  472.22 2225.68 710.66 2232.4 ;
     RECT  2657.66 2231.12 2668.9 2233.22 ;
     RECT  2737.82 2230.7 2740.9 2233.22 ;
     RECT  2357.66 2226.5 2619.46 2234.06 ;
     RECT  2357.66 2234.06 2538.82 2234.48 ;
     RECT  2640.38 2231.12 2640.58 2234.48 ;
     RECT  2657.66 2233.22 2659.3 2234.48 ;
     RECT  2738.3 2233.22 2740.9 2234.48 ;
     RECT  723.9 2228.16 1051.94 2234.68 ;
     RECT  2740.7 2234.48 2740.9 2234.9 ;
     RECT  475.1 2232.4 710.66 2235.34 ;
     RECT  2519.42 2234.48 2538.82 2237 ;
     RECT  2519.42 2237 2537.86 2237.42 ;
     RECT  1062.3 2228.16 1167.62 2237.5 ;
     RECT  2532.86 2237.42 2537.86 2237.84 ;
     RECT  722.94 2234.68 1051.94 2238.04 ;
     RECT  1062.3 2237.5 1168.58 2238.04 ;
     RECT  2519.42 2237.42 2521.54 2238.26 ;
     RECT  2357.66 2234.48 2495.14 2238.68 ;
     RECT  486.62 2235.34 710.66 2238.7 ;
     RECT  2235.26 2027.24 2235.46 2239.12 ;
     RECT  486.62 2238.7 562.18 2239.54 ;
     RECT  475.1 2235.34 475.3 2239.96 ;
     RECT  487.1 2239.54 562.18 2240.38 ;
     RECT  2519.42 2238.26 2520.58 2240.78 ;
     RECT  2549.18 2234.06 2618.02 2240.78 ;
     RECT  722.94 2238.04 1168.58 2241.18 ;
     RECT  2357.66 2238.68 2485.54 2241.62 ;
     RECT  2357.66 2241.62 2480.74 2241.64 ;
     RECT  2358.62 2241.64 2480.74 2242.04 ;
     RECT  2549.18 2240.78 2617.54 2242.04 ;
     RECT  2358.62 2242.04 2476.42 2242.06 ;
     RECT  2520.38 2240.78 2520.58 2242.46 ;
     RECT  2362.46 2242.06 2476.42 2244.56 ;
     RECT  3221.18 2215 3400 2244.58 ;
     RECT  572.06 2238.7 710.66 2244.76 ;
     RECT  722.94 2241.18 1083.62 2244.76 ;
     RECT  2384.54 2244.56 2476.42 2244.98 ;
     RECT  2549.18 2242.04 2617.06 2244.98 ;
     RECT  2550.14 2244.98 2617.06 2245.4 ;
     RECT  2550.14 2245.4 2552.74 2245.82 ;
     RECT  1093.5 2241.18 1168.58 2247.28 ;
     RECT  2362.46 2244.56 2373.22 2248.34 ;
     RECT  496.7 2240.38 562.18 2248.36 ;
     RECT  1093.5 2247.28 1175.3 2248.54 ;
     RECT  2384.54 2244.98 2472.1 2249.18 ;
     RECT  2564.06 2245.4 2617.06 2249.18 ;
     RECT  2370.14 2248.34 2373.22 2249.6 ;
     RECT  2385.5 2249.18 2467.78 2249.6 ;
     RECT  2552.54 2245.82 2552.74 2249.6 ;
     RECT  2564.06 2249.18 2568.58 2249.6 ;
     RECT  2600.54 2249.18 2602.18 2249.6 ;
     RECT  2613.02 2249.18 2617.06 2249.6 ;
     RECT  501.02 2248.36 562.18 2249.62 ;
     RECT  2564.06 2249.6 2564.26 2250.02 ;
     RECT  2616.86 2249.6 2617.06 2250.02 ;
     RECT  501.02 2249.62 551.62 2250.04 ;
     RECT  3207.74 2182.42 3207.94 2250.04 ;
     RECT  2370.14 2249.6 2372.26 2250.46 ;
     RECT  561.98 2249.62 562.18 2250.88 ;
     RECT  572.06 2244.76 1083.62 2251.9 ;
     RECT  1093.5 2248.54 1182.98 2251.9 ;
     RECT  572.06 2251.9 1182.98 2252.32 ;
     RECT  3070.94 2224.84 3112.42 2252.56 ;
     RECT  2387.42 2249.6 2424.58 2252.96 ;
     RECT  2580.86 2249.18 2585.86 2252.96 ;
     RECT  3077.66 2252.56 3112.42 2252.98 ;
     RECT  2387.42 2252.96 2407.78 2253.8 ;
     RECT  2583.26 2252.96 2583.46 2253.8 ;
     RECT  3084.38 2252.98 3112.42 2253.82 ;
     RECT  2399.9 2253.8 2407.78 2254.22 ;
     RECT  2436.86 2249.6 2461.54 2254.22 ;
     RECT  501.02 2250.04 549.7 2255.5 ;
     RECT  2420.06 2252.96 2424.58 2255.9 ;
     RECT  2436.86 2254.22 2456.74 2255.9 ;
     RECT  2455.58 2255.9 2456.74 2256.32 ;
     RECT  2420.06 2255.9 2421.22 2256.74 ;
     RECT  2436.86 2255.9 2445.7 2256.74 ;
     RECT  2253.02 2238.92 2253.22 2256.98 ;
     RECT  2399.9 2254.22 2401.06 2257.16 ;
     RECT  2420.06 2256.74 2420.26 2257.16 ;
     RECT  2253.02 2256.98 2253.7 2257.18 ;
     RECT  2399.9 2257.16 2400.1 2257.58 ;
     RECT  2438.3 2256.74 2440.9 2257.58 ;
     RECT  2455.58 2256.32 2455.78 2257.58 ;
     RECT  572.06 2252.32 1186.34 2257.82 ;
     RECT  2372.06 2250.46 2372.26 2258.02 ;
     RECT  2387.42 2253.8 2387.62 2258.02 ;
     RECT  562.46 2257.82 1186.34 2258.62 ;
     RECT  3098.78 2253.82 3112.42 2259.7 ;
     RECT  3084.38 2253.82 3088.42 2262.64 ;
     RECT  562.46 2258.62 1189.22 2263.86 ;
     RECT  3084.86 2262.64 3088.42 2264.32 ;
     RECT  2440.7 2257.58 2440.9 2264.74 ;
     RECT  562.46 2263.86 1175.3 2266.22 ;
     RECT  505.34 2255.5 549.7 2267.06 ;
     RECT  3098.78 2259.7 3111.94 2267.26 ;
     RECT  503.9 2267.06 549.7 2267.9 ;
     RECT  561.5 2266.22 1175.3 2267.9 ;
     RECT  1958.78 1856.3 1958.98 2268.74 ;
     RECT  3098.78 2267.26 3111.46 2269.78 ;
     RECT  503.9 2267.9 1175.3 2270.16 ;
     RECT  503.9 2270.16 1174.34 2270.2 ;
     RECT  1293.18 2199.44 1826.02 2271.26 ;
     RECT  1185.66 2263.86 1189.22 2273.32 ;
     RECT  505.34 2270.2 1174.34 2273.52 ;
     RECT  1888.22 1826.9 1893.22 2276.3 ;
     RECT  505.34 2273.52 1173.86 2278.18 ;
     RECT  1185.66 2273.32 1192.1 2278.78 ;
     RECT  2868.86 2256.98 2869.06 2279.02 ;
     RECT  3098.78 2269.78 3110.98 2279.06 ;
     RECT  2411.9 2264.54 2412.1 2280.28 ;
     RECT  1184.7 2278.78 1192.1 2282.56 ;
     RECT  3110.78 2279.06 3110.98 2283.22 ;
     RECT  1911.26 1845.8 1923.46 2283.86 ;
     RECT  513.02 2278.18 1173.86 2284.66 ;
     RECT  1184.7 2282.56 1195.94 2284.66 ;
     RECT  1293.18 2271.26 1828.42 2284.9 ;
     RECT  2400.38 2280.92 2400.58 2284.9 ;
     RECT  1205.82 2262.4 1206.02 2285.08 ;
     RECT  513.02 2284.66 1195.94 2285.74 ;
     RECT  2901.5 2257.82 2901.7 2286.16 ;
     RECT  1205.82 2285.08 1211.3 2286.34 ;
     RECT  1228.86 2217.04 1243.46 2286.34 ;
     RECT  514.94 2285.74 1195.94 2286.76 ;
     RECT  1205.82 2286.34 1243.46 2286.76 ;
     RECT  2792.06 2285.96 2792.26 2289.74 ;
     RECT  2774.3 2264.54 2774.5 2289.94 ;
     RECT  3098.78 2279.06 3098.98 2292.46 ;
     RECT  1865.18 1857.56 1871.14 2296.46 ;
     RECT  514.94 2286.76 1243.46 2297.3 ;
     RECT  1976.06 2221.28 1977.7 2298.98 ;
     RECT  512.54 2297.3 1243.46 2300.02 ;
     RECT  2937.5 2285.96 2937.7 2300.44 ;
     RECT  3020.06 2300.24 3020.26 2300.66 ;
     RECT  2951.9 2278.82 2952.1 2300.86 ;
     RECT  2005.34 2005.4 2005.54 2301.5 ;
     RECT  1411.58 2284.9 1828.42 2302.96 ;
     RECT  1938.14 1871.84 1938.34 2303.18 ;
     RECT  1411.58 2302.96 1562.5 2303.38 ;
     RECT  518.78 2300.02 1243.46 2303.8 ;
     RECT  1575.74 2302.96 1596.1 2303.8 ;
     RECT  1605.98 2302.96 1615.3 2303.8 ;
     RECT  541.82 2303.8 1243.46 2304.22 ;
     RECT  1605.98 2303.8 1610.02 2305.9 ;
     RECT  518.78 2303.8 531.94 2306.74 ;
     RECT  1268.7 2300.2 1268.9 2307.12 ;
     RECT  1605.98 2305.9 1606.18 2307.16 ;
     RECT  1629.02 2302.96 1828.42 2307.58 ;
     RECT  527.9 2306.74 531.94 2308 ;
     RECT  1630.46 2307.58 1828.42 2310.52 ;
     RECT  550.46 2304.22 1243.46 2310.9 ;
     RECT  2792.06 2289.74 2793.7 2311.36 ;
     RECT  3084.86 2264.32 3085.06 2311.78 ;
     RECT  550.46 2310.9 1212.26 2312.16 ;
     RECT  1228.86 2310.9 1243.46 2313.84 ;
     RECT  1633.34 2310.52 1828.42 2315.14 ;
     RECT  1633.34 2315.14 1637.38 2315.98 ;
     RECT  1658.3 2315.14 1790.5 2315.98 ;
     RECT  1411.58 2303.38 1560.58 2317.24 ;
     RECT  1560.38 2317.24 1560.58 2318.3 ;
     RECT  1411.58 2317.24 1549.54 2318.5 ;
     RECT  1293.18 2284.9 1400.74 2319.52 ;
     RECT  1411.58 2318.5 1543.3 2322.7 ;
     RECT  550.46 2312.16 1209.86 2324.14 ;
     RECT  550.46 2324.14 1217.54 2327.08 ;
     RECT  3012.86 2300.66 3020.26 2328.58 ;
     RECT  1411.58 2322.7 1540.42 2329.42 ;
     RECT  550.46 2327.08 1218.02 2330.68 ;
     RECT  1290.78 2319.52 1400.74 2330.68 ;
     RECT  552.38 2330.68 1218.02 2331.06 ;
     RECT  1658.78 2315.98 1790.5 2331.52 ;
     RECT  1803.26 2315.14 1828.42 2332.7 ;
     RECT  1411.58 2329.42 1536.58 2332.9 ;
     RECT  1658.78 2331.52 1772.26 2332.9 ;
     RECT  1411.58 2332.9 1526.5 2333.2 ;
     RECT  1658.78 2332.9 1771.3 2333.62 ;
     RECT  818.94 2331.06 1218.02 2333.8 ;
     RECT  818.94 2333.8 1221.38 2334.42 ;
     RECT  552.38 2331.06 809.06 2334.46 ;
     RECT  820.38 2334.42 1221.38 2338.2 ;
     RECT  1236.06 2313.84 1243.46 2338.62 ;
     RECT  3222 2244.58 3400 2339 ;
     RECT  820.38 2338.2 1219.94 2339.04 ;
     RECT  3031.1 2328.38 3031.3 2339.92 ;
     RECT  1658.78 2333.62 1765.06 2340.76 ;
     RECT  552.38 2334.46 552.58 2342.02 ;
     RECT  563.42 2334.46 809.06 2342.02 ;
     RECT  570.62 2342.02 809.06 2342.86 ;
     RECT  2815.1 2311.16 2815.3 2343.7 ;
     RECT  3012.86 2328.58 3013.06 2343.7 ;
     RECT  571.1 2342.86 809.06 2345.56 ;
     RECT  820.38 2339.04 1211.3 2345.56 ;
     RECT  1290.78 2330.68 1360.9 2345.76 ;
     RECT  1658.78 2340.76 1735.3 2345.8 ;
     RECT  1292.22 2345.76 1360.9 2346.18 ;
     RECT  1658.78 2345.8 1730.5 2348.32 ;
     RECT  0 2225 178 2349 ;
     RECT  1669.82 2348.32 1730.5 2349.16 ;
     RECT  571.1 2345.56 1211.3 2350.6 ;
     RECT  3222 2339 3470 2352.225 ;
     RECT  571.1 2350.6 1218.02 2353.36 ;
     RECT  1370.78 2330.68 1400.74 2354.5 ;
     RECT  3052.7 2340.14 3052.9 2354.62 ;
     RECT  3220 2352.225 3470 2355.47 ;
     RECT  581.18 2353.36 1218.02 2357.1 ;
     RECT  581.18 2357.1 1208.42 2357.56 ;
     RECT  3160.22 2343.5 3160.42 2357.78 ;
     RECT  3160.22 2357.78 3160.9 2357.98 ;
     RECT  581.66 2357.56 1208.42 2360.04 ;
     RECT  581.66 2360.04 1088.9 2360.5 ;
     RECT  3218.3 2355.47 3470 2361.34 ;
     RECT  1411.58 2333.2 1522.66 2363.02 ;
     RECT  1099.74 2360.04 1208.42 2364.24 ;
     RECT  1292.7 2346.18 1360.9 2364.66 ;
     RECT  600.86 2360.5 1088.9 2365.92 ;
     RECT  1463.42 2363.02 1522.66 2365.96 ;
     RECT  600.86 2365.92 1087.94 2366.34 ;
     RECT  581.66 2360.5 588.1 2368.9 ;
     RECT  1153.5 2364.24 1208.42 2369.5 ;
     RECT  1099.74 2364.24 1139.78 2369.7 ;
     RECT  1102.62 2369.7 1139.78 2371.8 ;
     RECT  1293.18 2364.66 1360.9 2372.06 ;
     RECT  1371.26 2354.5 1400.74 2372.06 ;
     RECT  1104.06 2371.8 1139.78 2372.22 ;
     RECT  1153.5 2369.5 1209.38 2372.22 ;
     RECT  600.86 2366.34 1078.82 2373.9 ;
     RECT  600.86 2373.9 755.78 2375.58 ;
     RECT  600.86 2375.58 741.86 2375.62 ;
     RECT  1243.26 2338.62 1243.46 2376 ;
     RECT  755.58 2375.58 755.78 2376.42 ;
     RECT  766.62 2373.9 1078.82 2376.42 ;
     RECT  766.62 2376.42 766.82 2376.84 ;
     RECT  1154.94 2372.22 1209.38 2376.84 ;
     RECT  777.18 2376.42 777.38 2377.26 ;
     RECT  791.1 2376.42 1078.82 2377.26 ;
     RECT  633.98 2375.62 741.86 2378.1 ;
     RECT  1104.54 2372.22 1139.78 2378.1 ;
     RECT  791.1 2377.26 1066.82 2378.52 ;
     RECT  802.62 2378.52 1066.82 2379.36 ;
     RECT  2750.78 2364.92 2750.98 2379.62 ;
     RECT  1104.54 2378.1 1134.98 2379.78 ;
     RECT  817.98 2379.36 1066.82 2380.2 ;
     RECT  817.98 2380.2 1046.66 2380.62 ;
     RECT  1066.62 2380.2 1066.82 2381.04 ;
     RECT  585.5 2368.9 588.1 2383.1 ;
     RECT  824.7 2380.62 1046.66 2383.14 ;
     RECT  600.86 2375.62 621.22 2383.3 ;
     RECT  -70 2349 178 2383.725 ;
     RECT  824.7 2383.14 1031.78 2383.98 ;
     RECT  1041.66 2383.14 1046.66 2383.98 ;
     RECT  -70 2383.725 180 2384.225 ;
     RECT  824.7 2383.98 858.5 2384.4 ;
     RECT  871.26 2383.98 1020.74 2384.4 ;
     RECT  871.26 2384.4 876.26 2384.82 ;
     RECT  887.1 2384.4 1020.74 2384.82 ;
     RECT  1030.62 2383.98 1031.78 2384.82 ;
     RECT  891.9 2384.82 1020.74 2385.24 ;
     RECT  898.14 2385.24 1020.74 2386.5 ;
     RECT  1030.62 2384.82 1030.82 2386.5 ;
     RECT  898.14 2386.5 996.26 2386.92 ;
     RECT  1411.58 2363.02 1453.54 2386.96 ;
     RECT  905.34 2386.92 996.26 2387.76 ;
     RECT  1154.94 2376.84 1207.94 2387.76 ;
     RECT  1006.14 2386.5 1020.74 2390.28 ;
     RECT  943.74 2387.76 996.26 2391.33 ;
     RECT  905.34 2387.76 930.02 2391.54 ;
     RECT  944.7 2391.33 996.26 2391.54 ;
     RECT  1011.42 2390.28 1020.74 2391.54 ;
     RECT  1170.3 2387.76 1193.54 2391.54 ;
     RECT  1187.1 2391.54 1191.14 2391.96 ;
     RECT  600.86 2383.3 619.78 2392 ;
     RECT  944.7 2391.54 989.54 2392.38 ;
     RECT  1011.42 2391.54 1018.18 2392.38 ;
     RECT  905.34 2391.54 910.34 2393.22 ;
     RECT  3222 2361.34 3470 2393.725 ;
     RECT  3175.1 2357.78 3175.3 2394.1 ;
     RECT  3220 2393.725 3470 2394.225 ;
     RECT  946.62 2392.38 989.54 2394.48 ;
     RECT  973.98 2394.48 984.74 2394.9 ;
     RECT  973.98 2394.9 978.98 2395.74 ;
     RECT  1174.14 2391.54 1174.34 2396.16 ;
     RECT  633.98 2378.1 732.26 2396.2 ;
     RECT  585.02 2383.1 588.1 2396.62 ;
     RECT  571.1 2353.36 571.3 2397.04 ;
     RECT  600.86 2392 615.46 2397.88 ;
     RECT  633.98 2396.2 639.46 2398.3 ;
     RECT  973.98 2395.74 975.14 2398.68 ;
     RECT  639.26 2398.3 639.46 2398.72 ;
     RECT  974.46 2398.68 974.66 2399.1 ;
     RECT  585.02 2396.62 585.22 2399.14 ;
     RECT  1017.98 2392.38 1018.18 2400.82 ;
     RECT  1207.74 2387.76 1207.94 2401.2 ;
     RECT  2876.06 2343.5 2876.26 2401.24 ;
     RECT  649.34 2396.2 732.26 2402.5 ;
     RECT  1188.54 2391.96 1191.14 2403.72 ;
     RECT  1748.06 2340.76 1765.06 2404.7 ;
     RECT  609.02 2397.88 615.46 2404.9 ;
     RECT  1669.82 2349.16 1707.46 2404.9 ;
     RECT  656.06 2402.5 732.26 2405.86 ;
     RECT  1113.66 2379.78 1134.98 2408.18 ;
     RECT  609.02 2404.9 613.54 2408.8 ;
     RECT  3222 2394.225 3470 2409 ;
     RECT  1154.94 2387.76 1159.94 2409.02 ;
     RECT  662.78 2405.86 732.26 2412.58 ;
     RECT  3016.7 2401.04 3016.9 2413.42 ;
     RECT  675.26 2412.58 732.26 2415.32 ;
     RECT  1154.94 2409.02 1163.62 2415.74 ;
     RECT  1414.94 2386.96 1453.54 2415.94 ;
     RECT  1113.66 2408.18 1135.78 2416.16 ;
     RECT  871.26 2384.82 871.46 2417.5 ;
     RECT  920.7 2391.54 923.78 2417.5 ;
     RECT  1188.54 2403.72 1188.74 2417.5 ;
     RECT  828.06 2384.4 858.5 2417.7 ;
     RECT  870.78 2417.5 871.46 2417.7 ;
     RECT  1188.06 2417.5 1188.74 2417.7 ;
     RECT  1293.18 2372.06 1400.74 2418.88 ;
     RECT  -70 2384.225 178 2419 ;
     RECT  1113.66 2416.16 1141.06 2421.36 ;
     RECT  1293.18 2418.88 1349.86 2421.4 ;
     RECT  1293.18 2421.4 1333.54 2422.46 ;
     RECT  3063.26 2354.42 3063.46 2422.46 ;
     RECT  3045.5 2413.22 3045.7 2422.66 ;
     RECT  920.22 2417.5 923.78 2426.4 ;
     RECT  3063.26 2422.46 3065.86 2426.86 ;
     RECT  675.26 2415.32 733.06 2428.76 ;
     RECT  946.62 2394.48 962.66 2428.92 ;
     RECT  1288.7 2422.46 1333.54 2428.96 ;
     RECT  1330.94 2428.96 1333.54 2431.48 ;
     RECT  1333.34 2431.48 1333.54 2432.32 ;
     RECT  3081.5 2426.66 3081.7 2433.8 ;
     RECT  3063.26 2426.86 3063.46 2434 ;
     RECT  1288.7 2428.96 1321.06 2434.42 ;
     RECT  1293.18 2434.42 1321.06 2436.1 ;
     RECT  802.62 2379.36 805.7 2436.48 ;
     RECT  1464.86 2365.96 1522.66 2437.36 ;
     RECT  675.26 2428.76 737.86 2437.78 ;
     RECT  675.74 2437.78 737.86 2439 ;
     RECT  1154.94 2415.74 1168.42 2439.46 ;
     RECT  905.34 2393.22 905.54 2441.52 ;
     RECT  1113.66 2421.36 1122.98 2444.04 ;
     RECT  1188.06 2417.7 1188.26 2444.04 ;
     RECT  1414.94 2415.94 1453.06 2444.08 ;
     RECT  1046.46 2383.98 1046.66 2446.56 ;
     RECT  1364.06 2418.88 1400.74 2446.6 ;
     RECT  0 2419 178 2448.08 ;
     RECT  191.42 2387.6 191.62 2448.08 ;
     RECT  3074.3 2433.8 3081.7 2448.08 ;
     RECT  0 2448.08 191.62 2448.28 ;
     RECT  1293.18 2436.1 1320.58 2448.28 ;
     RECT  3074.3 2448.08 3085.06 2448.28 ;
     RECT  948.06 2428.92 962.66 2449.08 ;
     RECT  609.02 2408.8 609.22 2451.64 ;
     RECT  1414.94 2444.08 1442.02 2451.64 ;
     RECT  1118.46 2444.04 1122.98 2454.12 ;
     RECT  1419.26 2451.64 1442.02 2454.16 ;
     RECT  3081.5 2448.28 3085.06 2455.42 ;
     RECT  920.22 2426.4 920.42 2456.64 ;
     RECT  1134.78 2421.36 1141.06 2456.64 ;
     RECT  1154.94 2439.46 1163.62 2459.16 ;
     RECT  1389.02 2446.6 1400.74 2459.2 ;
     RECT  1293.18 2448.28 1313.38 2462.56 ;
     RECT  675.74 2439 726.02 2464.2 ;
     RECT  1162.46 2459.16 1163.62 2464.66 ;
     RECT  3114.62 2455.22 3114.82 2464.66 ;
     RECT  1400.54 2459.2 1400.74 2465.92 ;
     RECT  1118.46 2454.12 1118.66 2466.72 ;
     RECT  1140.86 2456.64 1141.06 2466.76 ;
     RECT  1419.26 2454.16 1430.5 2466.76 ;
     RECT  828.06 2417.7 858.02 2469.24 ;
     RECT  1293.18 2462.56 1307 2469.24 ;
     RECT  1162.46 2464.66 1162.66 2471.8 ;
     RECT  3146.3 2464.46 3146.5 2473.48 ;
     RECT  725.82 2464.2 726.02 2476.8 ;
     RECT  1298.94 2469.24 1307 2476.8 ;
     RECT  1419.26 2466.76 1429.54 2476.84 ;
     RECT  675.74 2464.2 710.66 2484.36 ;
     RECT  737.66 2439 737.86 2484.4 ;
     RECT  675.74 2484.36 705.86 2487.34 ;
     RECT  1299.74 2476.8 1307 2487.56 ;
     RECT  828.06 2469.24 845.54 2489.4 ;
     RECT  805.5 2436.48 805.7 2489.5 ;
     RECT  805.02 2489.5 805.7 2489.7 ;
     RECT  693 2487.34 705.86 2494.44 ;
     RECT  1441.82 2454.16 1442.02 2494.9 ;
     RECT  870.78 2417.7 870.98 2496.96 ;
     RECT  855.42 2469.24 858.02 2499.48 ;
     RECT  857.82 2499.48 858.02 2502 ;
     RECT  1349.66 2421.4 1349.86 2505.5 ;
     RECT  675.74 2487.34 676.9 2505.7 ;
     RECT  1349.18 2505.5 1349.86 2505.7 ;
     RECT  948.06 2449.08 950.66 2508.98 ;
     RECT  962.46 2449.08 962.66 2508.98 ;
     RECT  834.3 2489.4 845.54 2509.56 ;
     RECT  3084.86 2455.42 3085.06 2512.34 ;
     RECT  3084.86 2512.34 3092.26 2512.54 ;
     RECT  834.3 2509.56 834.5 2514.6 ;
     RECT  648.86 2512.76 649.06 2515.48 ;
     RECT  948.06 2508.98 962.66 2516.32 ;
     RECT  962.46 2516.32 962.66 2517.12 ;
     RECT  948.06 2516.32 948.26 2519.64 ;
     RECT  675.74 2505.7 676.42 2522.62 ;
     RECT  845.34 2509.56 845.54 2524.68 ;
     RECT  805.02 2489.7 805.22 2527.2 ;
     RECT  693 2494.44 699.94 2529.52 ;
     RECT  0 2448.28 190.66 2530.6 ;
     RECT  3222 2409 3400 2533 ;
     RECT  693 2529.52 700.66 2534.6 ;
     RECT  676.22 2522.62 676.42 2534.8 ;
     RECT  3171.26 2473.28 3171.46 2534.8 ;
     RECT  693 2534.6 701.38 2541.74 ;
     RECT  693 2541.74 702.34 2542.32 ;
     RECT  0 2530.6 178 2543 ;
     RECT  3222 2533 3470 2546.225 ;
     RECT  3220 2546.225 3470 2546.57 ;
     RECT  3218.3 2546.57 3470 2555.8 ;
     RECT  662.78 2412.58 662.98 2560.42 ;
     RECT  693 2542.32 701.38 2570.04 ;
     RECT  3192.86 2534.6 3193.06 2570.5 ;
     RECT  -70 2543 178 2576.145 ;
     RECT  3092.06 2512.54 3092.26 2577.02 ;
     RECT  3092.06 2577.02 3099.46 2577.22 ;
     RECT  -70 2576.145 180 2577.86 ;
     RECT  -70 2577.86 180.58 2578.06 ;
     RECT  428.06 2190.82 428.26 2578.06 ;
     RECT  693 2570.04 700.9 2578.06 ;
     RECT  -70 2578.06 180 2579.855 ;
     RECT  693 2578.06 697.6 2582.72 ;
     RECT  693 2582.72 695 2585.32 ;
     RECT  1293.98 2487.56 1307 2585.32 ;
     RECT  3222 2555.8 3470 2587.725 ;
     RECT  3203.9 2570.3 3204.1 2588.14 ;
     RECT  3220 2587.725 3470 2588.225 ;
     RECT  3222 2588.225 3470 2603 ;
     RECT  -70 2579.855 178 2613 ;
     RECT  3099.26 2577.22 3099.46 2666.48 ;
     RECT  3099.26 2666.48 3105.22 2666.68 ;
     RECT  3105.02 2666.68 3105.22 2691.88 ;
     RECT  1464.86 2437.36 1478.02 2692.94 ;
     RECT  1488.38 2437.36 1522.66 2692.94 ;
     RECT  1464.86 2692.94 1522.66 2693.14 ;
     RECT  3117.5 2691.68 3117.7 2718.34 ;
     RECT  2556.38 2372.06 2556.58 2724.86 ;
     RECT  3222 2603 3400 2727 ;
     RECT  1475.9 2693.14 1522.66 2727.16 ;
     RECT  3222 2727 3470 2736.2 ;
     RECT  0 2613 178 2737 ;
     RECT  2092.7 1926.02 2107.3 2739.56 ;
     RECT  3218.3 2736.2 3470 2740.39 ;
     RECT  1747.58 2404.7 1765.06 2742.5 ;
     RECT  3132.38 2718.14 3132.58 2743.54 ;
     RECT  3220 2740.39 3470 2743.775 ;
     RECT  3146.3 2743.34 3146.5 2757.82 ;
     RECT  -70 2737 178 2771.725 ;
     RECT  3165.5 2757.62 3165.7 2772.1 ;
     RECT  -70 2771.725 180 2772.225 ;
     RECT  190.46 2530.6 190.66 2772.52 ;
     RECT  209.18 2769.8 209.38 2772.52 ;
     RECT  3222 2743.775 3470 2781.725 ;
     RECT  3182.78 2771.9 3182.98 2782.18 ;
     RECT  3220 2781.725 3470 2782.225 ;
     RECT  3222 2782.225 3470 2797 ;
     RECT  -70 2772.225 178 2807 ;
     RECT  0 2807 178 2843.72 ;
     RECT  190.94 2773.16 191.14 2843.72 ;
     RECT  0 2843.72 191.14 2843.92 ;
     RECT  1782.14 2331.52 1790.5 2858.3 ;
     RECT  1719.74 2349.16 1730.5 2869.12 ;
     RECT  1803.26 2332.7 1828.9 2876.26 ;
     RECT  1428.86 2476.84 1429.54 2883.82 ;
     RECT  1719.74 2869.12 1723.78 2883.82 ;
     RECT  1364.06 2446.6 1375.3 2887.1 ;
     RECT  1815.74 2876.26 1828.9 2887.3 ;
     RECT  2028.38 2193.14 2030.5 2887.3 ;
     RECT  1815.74 2887.3 1828.42 2890.96 ;
     RECT  1560.38 2318.3 1565.86 2894.96 ;
     RECT  1669.82 2404.9 1706.5 2899.58 ;
     RECT  1865.18 2296.46 1872.1 2900.42 ;
     RECT  1888.22 2276.3 1897.06 2900.42 ;
     RECT  1452.86 2444.08 1453.06 2901.68 ;
     RECT  1669.82 2899.58 1708.42 2901.68 ;
     RECT  1719.74 2883.82 1719.94 2901.68 ;
     RECT  1464.86 2693.14 1465.54 2904.62 ;
     RECT  1477.82 2727.16 1522.66 2904.62 ;
     RECT  1745.66 2742.5 1765.06 2904.62 ;
     RECT  1782.14 2858.3 1790.98 2904.62 ;
     RECT  1865.18 2900.42 1897.06 2904.62 ;
     RECT  1907.42 2283.86 1923.46 2904.62 ;
     RECT  1428.86 2883.82 1429.06 2905.46 ;
     RECT  1658.78 2348.32 1658.98 2905.88 ;
     RECT  1669.82 2901.68 1719.94 2905.88 ;
     RECT  1464.86 2904.62 1522.66 2906.3 ;
     RECT  1364.06 2887.1 1375.78 2907.14 ;
     RECT  1389.02 2459.2 1389.22 2907.14 ;
     RECT  1637.18 2315.98 1637.38 2907.14 ;
     RECT  0 2843.92 183.46 2907.34 ;
     RECT  1536.38 2332.9 1536.58 2907.56 ;
     RECT  1607.42 2324.18 1607.62 2907.56 ;
     RECT  1618.46 2329.22 1618.66 2907.56 ;
     RECT  1629.02 2907.14 1638.82 2907.56 ;
     RECT  1658.78 2905.88 1719.94 2907.56 ;
     RECT  1745.66 2904.62 1790.98 2907.56 ;
     RECT  1825.82 2890.96 1828.42 2907.56 ;
     RECT  1970.78 2298.98 1977.7 2907.56 ;
     RECT  1988.06 2221.7 1988.26 2907.56 ;
     RECT  2028.38 2887.3 2030.02 2907.56 ;
     RECT  2050.94 2198.6 2051.62 2907.56 ;
     RECT  1555.1 2894.96 1565.86 2907.98 ;
     RECT  1583.42 2303.8 1596.1 2907.98 ;
     RECT  1607.42 2907.56 1719.94 2907.98 ;
     RECT  1733.18 2907.56 1790.98 2907.98 ;
     RECT  1803.26 2876.26 1803.94 2907.98 ;
     RECT  1815.74 2890.96 1815.94 2907.98 ;
     RECT  1825.82 2907.56 1830.82 2907.98 ;
     RECT  1840.7 1868.9 1849.06 2907.98 ;
     RECT  1865.18 2904.62 1923.46 2907.98 ;
     RECT  1954.94 2268.74 1958.98 2907.98 ;
     RECT  1450.46 2901.68 1453.06 2908.4 ;
     RECT  1464.86 2906.3 1526.5 2908.4 ;
     RECT  1536.38 2907.56 1539.94 2908.4 ;
     RECT  1555.1 2907.98 1566.34 2908.4 ;
     RECT  1583.42 2907.98 1719.94 2908.4 ;
     RECT  1803.26 2907.98 1815.94 2908.4 ;
     RECT  1825.82 2907.98 1923.46 2908.4 ;
     RECT  1335.74 2907.56 1335.94 2908.82 ;
     RECT  1349.18 2505.7 1349.38 2908.82 ;
     RECT  1424.06 2905.46 1429.06 2908.82 ;
     RECT  1449.5 2908.4 1453.06 2908.82 ;
     RECT  1464.86 2908.4 1566.34 2908.82 ;
     RECT  2040.86 1800.86 2041.06 2908.82 ;
     RECT  2050.94 2907.56 2052.1 2908.82 ;
     RECT  2066.78 1915.52 2066.98 2908.82 ;
     RECT  1364.06 2907.14 1389.22 2909.24 ;
     RECT  1412.06 2905.88 1412.26 2910.92 ;
     RECT  1938.14 2303.18 1940.26 2912.18 ;
     RECT  1970.78 2907.56 1990.66 2912.18 ;
     RECT  2005.34 2301.5 2008.9 2912.18 ;
     RECT  2066.78 2908.82 2067.46 2912.18 ;
     RECT  2079.74 2306.54 2079.94 2912.18 ;
     RECT  1360.22 2909.24 1389.22 2912.6 ;
     RECT  1400.54 2907.98 1400.74 2912.6 ;
     RECT  1938.14 2912.18 1943.62 2912.6 ;
     RECT  1954.94 2907.98 1960.42 2912.6 ;
     RECT  1970.78 2912.18 2012.74 2912.6 ;
     RECT  2028.38 2907.56 2030.5 2912.6 ;
     RECT  2040.86 2908.82 2056.9 2912.6 ;
     RECT  1411.58 2910.92 1412.26 2913.02 ;
     RECT  1424.06 2908.82 1435.78 2913.02 ;
     RECT  1577.18 2908.4 1719.94 2913.02 ;
     RECT  1801.82 2908.4 1923.46 2913.02 ;
     RECT  1322.78 2908.82 1322.98 2913.44 ;
     RECT  1411.1 2913.02 1435.78 2913.44 ;
     RECT  1449.5 2908.82 1566.34 2913.44 ;
     RECT  1576.7 2913.02 1719.94 2913.44 ;
     RECT  1732.7 2907.98 1790.98 2913.44 ;
     RECT  1801.82 2913.02 1923.94 2913.44 ;
     RECT  1935.74 2912.6 1944.58 2913.44 ;
     RECT  2066.78 2912.18 2080.42 2913.44 ;
     RECT  2092.7 2739.56 2109.22 2913.44 ;
     RECT  1320.38 2913.44 1322.98 2914.7 ;
     RECT  1319.9 2914.7 1322.98 2915.12 ;
     RECT  1335.74 2908.82 1349.38 2915.12 ;
     RECT  1360.22 2912.6 1400.74 2915.12 ;
     RECT  1411.1 2913.44 1719.94 2915.12 ;
     RECT  1732.7 2913.44 1944.58 2915.12 ;
     RECT  1954.94 2912.6 2012.74 2915.12 ;
     RECT  2028.38 2912.6 2056.9 2915.12 ;
     RECT  2066.78 2913.44 2109.22 2915.12 ;
     RECT  1316.54 2915.12 1719.94 2915.54 ;
     RECT  1293.98 2585.32 1300.42 2917.22 ;
     RECT  1310.3 2915.54 1720.9 2917.22 ;
     RECT  3222 2797 3400 2921 ;
     RECT  1293.98 2917.22 1720.9 2925.32 ;
     RECT  1732.7 2915.12 2109.22 2925.32 ;
     RECT  1293.98 2925.32 2109.22 2928.56 ;
     RECT  0 2907.34 178 2931 ;
     RECT  1292.54 2928.56 2109.22 2936.32 ;
     RECT  3222 2921 3470 2991 ;
     RECT  -70 2931 178 3001 ;
     RECT  1293.98 2936.32 2109.22 3022 ;
     RECT  1293.98 3022 2107.3 3044.1 ;
     RECT  2077.34 3044.1 2107.3 3045.32 ;
     RECT  1293.98 3044.1 1397.86 3045.74 ;
     RECT  2077.34 3045.32 2110.66 3048.26 ;
     RECT  1279.58 3048.26 1279.78 3048.68 ;
     RECT  1292.54 3045.74 1397.86 3048.68 ;
     RECT  2077.34 3048.26 2112.58 3049.1 ;
     RECT  2077.34 3049.1 2113.06 3050.78 ;
     RECT  1279.58 3048.68 1397.86 3052.46 ;
     RECT  2008.7 3044.1 2065.06 3055.82 ;
     RECT  2077.34 3050.78 2115.46 3055.82 ;
     RECT  1277.66 3052.46 1397.86 3056.66 ;
     RECT  2008.7 3055.82 2116.9 3057.08 ;
     RECT  1275.74 3056.66 1397.86 3059.1 ;
     RECT  1408.22 3044.1 1664.74 3059.1 ;
     RECT  1682.3 3044.1 1710.82 3059.1 ;
     RECT  1720.7 3044.1 1720.9 3059.1 ;
     RECT  1734.62 3044.1 1993.54 3059.1 ;
     RECT  2008.7 3057.08 2124.1 3059.1 ;
     RECT  1275.74 3059.1 2124.1 3063.58 ;
     RECT  1275.74 3063.58 2118.34 3064.84 ;
     RECT  1281.5 3064.84 2118.34 3066.1 ;
     RECT  1281.5 3066.1 2117.86 3066.52 ;
     RECT  1281.5 3066.52 2114.98 3067.78 ;
     RECT  1281.98 3067.78 2114.98 3074.5 ;
     RECT  2112.38 3074.5 2112.58 3074.92 ;
     RECT  1281.98 3074.5 2099.62 3078.7 ;
     RECT  1293.02 3078.7 2099.16 3079.12 ;
     RECT  1296.38 3079.12 2099.16 3079.54 ;
     RECT  1298.3 3079.54 2099.16 3110.3 ;
     RECT  3222 2991 3400 3115 ;
     RECT  0 3001 178 3125 ;
     RECT  1297.82 3110.3 2099.16 3177.88 ;
     RECT  1297.82 3177.88 1305.28 3180.48 ;
     RECT  2094.56 3177.88 2099.16 3180.48 ;
     RECT  1297.82 3180.48 1302.68 3183.08 ;
     RECT  2097.16 3180.48 2099.16 3183.08 ;
     RECT  3222 3115 3470 3185 ;
     RECT  1281.98 3078.7 1282.18 3187.06 ;
     RECT  1449.98 3177.88 1457.86 3187.48 ;
     RECT  1479.74 3177.88 1512.1 3187.48 ;
     RECT  1523.9 3177.88 1524.1 3187.48 ;
     RECT  1539.74 3177.88 1545.22 3187.48 ;
     RECT  1569.98 3177.88 1570.18 3187.48 ;
     RECT  1581.02 3177.88 1581.22 3187.48 ;
     RECT  1603.1 3177.88 1612.42 3187.48 ;
     RECT  1631.9 3177.88 1665.7 3187.48 ;
     RECT  1682.78 3177.88 1716.58 3187.48 ;
     RECT  1758.14 3177.88 1758.34 3187.48 ;
     RECT  1796.54 3177.88 1811.62 3187.48 ;
     RECT  1835.42 3177.88 1859.62 3187.48 ;
     RECT  1876.7 3177.88 1876.9 3187.48 ;
     RECT  1888.7 3177.88 1888.9 3187.48 ;
     RECT  1904.06 3177.88 1913.86 3187.48 ;
     RECT  1931.9 3177.88 1932.1 3187.48 ;
     RECT  1942.46 3177.88 1942.66 3187.48 ;
     RECT  1963.58 3177.88 1963.78 3187.48 ;
     RECT  1297.82 3183.08 1298.02 3188.32 ;
     RECT  1677.5 3188.54 1678.66 3189.8 ;
     RECT  1697.66 3187.48 1716.58 3191.48 ;
     RECT  1432.22 3177.88 1432.42 3192.1 ;
     RECT  1454.3 3187.48 1454.5 3192.1 ;
     RECT  1492.7 3187.48 1492.9 3192.1 ;
     RECT  1540.7 3187.48 1540.9 3192.1 ;
     RECT  1554.14 3187.7 1554.34 3192.1 ;
     RECT  1583.9 3187.7 1585.06 3192.1 ;
     RECT  1603.1 3187.48 1603.3 3192.1 ;
     RECT  1655.9 3187.48 1656.1 3192.1 ;
     RECT  1673.66 3189.8 1678.66 3192.1 ;
     RECT  1742.3 3177.88 1742.5 3192.1 ;
     RECT  1773.98 3177.88 1774.18 3192.1 ;
     RECT  1787.42 3187.7 1787.62 3192.1 ;
     RECT  1803.26 3187.48 1803.46 3192.1 ;
     RECT  1838.3 3187.48 1854.34 3192.1 ;
     RECT  1907.9 3187.48 1908.1 3192.1 ;
     RECT  1943.42 3188.54 1943.62 3192.1 ;
     RECT  1697.66 3191.48 1717.06 3193.36 ;
     RECT  -70 3125 178 3195 ;
     RECT  1673.66 3192.1 1674.34 3195.04 ;
     RECT  1699.58 3193.36 1717.06 3195.04 ;
     RECT  1964.54 3188.54 1964.74 3195.04 ;
     RECT  1674.14 3195.04 1674.34 3195.46 ;
     RECT  1701.02 3195.04 1701.22 3195.88 ;
     RECT  2168.54 2078.48 2172.1 3211.3 ;
     RECT  1583.9 3192.1 1584.1 3215.42 ;
     RECT  2750.78 2379.62 2753.86 3217.94 ;
     RECT  830.3 2515.28 830.5 3219.2 ;
     RECT  0 3195 178 3220 ;
     RECT  638.78 2516.12 638.98 3220 ;
     RECT  830.3 3219.2 833.86 3220 ;
     RECT  1024.22 3219.2 1024.42 3220 ;
     RECT  1218.14 3219.2 1218.34 3220 ;
     RECT  1397.18 3203.66 1397.38 3220 ;
     RECT  1436.06 3203.24 1436.26 3220 ;
     RECT  1583.9 3215.42 1587.46 3220 ;
     RECT  1778.3 3196.94 1778.5 3220 ;
     RECT  1972.7 3196.94 1972.9 3220 ;
     RECT  2168.54 3211.3 2171.775 3220 ;
     RECT  2209.82 1912.78 2210.02 3220 ;
     RECT  2362.46 2653.04 2362.66 3220 ;
     RECT  2404.22 2314.52 2404.42 3220 ;
     RECT  2556.38 2724.86 2559.94 3220 ;
     RECT  2598.14 2264.12 2598.34 3220 ;
     RECT  2750.54 3217.94 2753.86 3220 ;
     RECT  2792.06 2311.36 2792.26 3220 ;
     RECT  3222 3185 3400 3220 ;
     RECT  1627.725 3220 1628.225 3220.04 ;
     RECT  1821.725 3220 1822.225 3220.04 ;
     RECT  0 3220 180 3222 ;
     RECT  636.145 3220 639.855 3222 ;
     RECT  830.145 3220 833.86 3222 ;
     RECT  1024.145 3220 1027.855 3222 ;
     RECT  1218.14 3220 1221.855 3222 ;
     RECT  1392.225 3220 1397.38 3222 ;
     RECT  1433.725 3220 1436.26 3222 ;
     RECT  1583.9 3220 1589.775 3222 ;
     RECT  1627.725 3220.04 1630.18 3222 ;
     RECT  1778.3 3220 1783.775 3222 ;
     RECT  1821.725 3220.04 1824.58 3222 ;
     RECT  1972.7 3220 1977.775 3222 ;
     RECT  2015.725 3220 2016.225 3222 ;
     RECT  2168.225 3220 2171.775 3222 ;
     RECT  2209.725 3220 2210.225 3222 ;
     RECT  2362.225 3220 2365.775 3222 ;
     RECT  2403.725 3220 2404.42 3222 ;
     RECT  2556.225 3220 2559.94 3222 ;
     RECT  2597.725 3220 2598.34 3222 ;
     RECT  2750.225 3220 2753.86 3222 ;
     RECT  2791.725 3220 2792.26 3222 ;
     RECT  3220 3220 3400 3222 ;
     RECT  0 3222 3400 3400 ;
     RECT  215 3400 285 3470 ;
     RECT  409 3400 479 3470 ;
     RECT  603 3400 673 3470 ;
     RECT  797 3400 867 3470 ;
     RECT  991 3400 1061 3470 ;
     RECT  1185 3400 1255 3470 ;
     RECT  1379 3400 1449 3470 ;
     RECT  1573 3400 1643 3470 ;
     RECT  1767 3400 1837 3470 ;
     RECT  1961 3400 2031 3470 ;
     RECT  2155 3400 2225 3470 ;
     RECT  2349 3400 2419 3470 ;
     RECT  2543 3400 2613 3470 ;
     RECT  2737 3400 2807 3470 ;
     RECT  2931 3400 3001 3470 ;
     RECT  3125 3400 3195 3470 ;
    LAYER Metal4 ;
     RECT  -70 215 0 285 ;
     RECT  -70 409 0 479 ;
     RECT  -70 603 0 673 ;
     RECT  -70 797 0 867 ;
     RECT  -70 991 0 1061 ;
     RECT  -70 1185 0 1255 ;
     RECT  -70 1379 0 1449 ;
     RECT  -70 1573 0 1643 ;
     RECT  -70 1767 0 1837 ;
     RECT  -70 1961 0 2031 ;
     RECT  -70 2155 0 2225 ;
     RECT  -70 2349 0 2419 ;
     RECT  -70 2543 0 2613 ;
     RECT  -70 2737 0 2807 ;
     RECT  -70 2931 0 3001 ;
     RECT  -70 3125 0 3195 ;
     RECT  0 0 178 3400 ;
     RECT  178 0 180 180 ;
     RECT  178 3220 180 3400 ;
     RECT  178 2530.4 183.46 2530.6 ;
     RECT  178 2907.14 183.46 2907.34 ;
     RECT  178 2771.9 187.1 2772.1 ;
     RECT  187.1 2771.9 187.3 2772.52 ;
     RECT  178 1801.7 190.66 1801.9 ;
     RECT  187.3 2772.32 190.66 2772.52 ;
     RECT  178 1025.96 201.7 1026.16 ;
     RECT  180 0 205 178 ;
     RECT  180 3222 215 3400 ;
     RECT  178 1608.08 233.38 1608.28 ;
     RECT  205 -70 275 178 ;
     RECT  215 3222 285 3470 ;
     RECT  275 0 399 178 ;
     RECT  285 3222 409 3400 ;
     RECT  178 831.92 433.06 832.12 ;
     RECT  429.5 2179.28 441.02 2179.48 ;
     RECT  441.02 2175.08 441.7 2179.48 ;
     RECT  441.7 2175.08 452.26 2175.28 ;
     RECT  453.5 2181.38 463.3 2181.58 ;
     RECT  399 -70 469 178 ;
     RECT  409 3222 479 3470 ;
     RECT  467.9 2171.3 479.62 2171.5 ;
     RECT  485.18 2212.88 486.14 2213.08 ;
     RECT  178 2195.66 489.98 2195.86 ;
     RECT  486.14 2205.32 489.98 2213.08 ;
     RECT  489.98 2195.66 491.14 2213.08 ;
     RECT  491.14 2212.88 493.54 2213.08 ;
     RECT  491.14 2195.66 496.9 2201.32 ;
     RECT  503.9 2212.88 505.34 2213.08 ;
     RECT  496.7 2225.06 505.34 2225.26 ;
     RECT  496.9 2195.66 505.82 2195.86 ;
     RECT  505.34 2212.88 507.74 2225.26 ;
     RECT  507.74 2212.88 509.86 2228.2 ;
     RECT  505.82 2194.4 511.3 2195.86 ;
     RECT  509.86 2216.24 514.18 2228.2 ;
     RECT  514.18 2228 522.82 2228.2 ;
     RECT  520.22 2121.74 524.06 2121.94 ;
     RECT  524.06 2121.74 525.5 2122.36 ;
     RECT  514.18 2216.24 527.14 2216.86 ;
     RECT  526.94 2137.7 527.42 2137.9 ;
     RECT  525.5 2121.74 527.9 2122.78 ;
     RECT  527.42 2137.28 527.9 2137.9 ;
     RECT  511.3 2195.66 528.86 2195.86 ;
     RECT  525.02 2087.72 529.82 2087.92 ;
     RECT  527.9 2121.74 530.3 2138.32 ;
     RECT  528.86 2195.66 532.7 2197.96 ;
     RECT  530.3 2118.8 532.9 2138.32 ;
     RECT  527.14 2216.66 533.38 2216.86 ;
     RECT  532.9 2122.58 534.34 2138.32 ;
     RECT  529.82 2084.78 534.62 2087.92 ;
     RECT  534.34 2126.78 535.3 2138.32 ;
     RECT  535.3 2126.78 535.78 2137.48 ;
     RECT  534.62 2084.78 536.06 2088.34 ;
     RECT  535.78 2126.78 536.26 2134.54 ;
     RECT  532.7 2195.66 538.18 2203 ;
     RECT  536.26 2129.72 540.1 2134.54 ;
     RECT  536.06 2084.78 541.06 2088.76 ;
     RECT  542.3 2224.64 543.26 2224.84 ;
     RECT  541.06 2084.78 544.42 2084.98 ;
     RECT  540.1 2129.72 545.38 2129.92 ;
     RECT  543.26 2220.86 545.38 2224.84 ;
     RECT  545.38 2222.54 546.34 2224.84 ;
     RECT  534.62 2235.56 547.78 2235.76 ;
     RECT  545.18 2114.6 548.06 2114.8 ;
     RECT  546.34 2223.8 548.26 2224.84 ;
     RECT  548.06 2114.6 550.66 2118.58 ;
     RECT  548.26 2223.8 552.58 2224 ;
     RECT  550.66 2118.38 553.54 2118.58 ;
     RECT  543.74 2102.42 554.5 2102.62 ;
     RECT  551.42 2144.84 554.5 2145.04 ;
     RECT  552.86 2209.52 554.5 2209.72 ;
     RECT  551.9 2285.12 560.54 2285.32 ;
     RECT  178 1220 562.66 1220.2 ;
     RECT  550.46 2312 565.34 2312.2 ;
     RECT  563.9 2212.04 566.5 2212.24 ;
     RECT  557.66 2088.56 566.78 2088.76 ;
     RECT  565.34 2312 569.18 2318.92 ;
     RECT  538.18 2195.66 569.66 2195.86 ;
     RECT  567.74 2205.32 569.66 2205.52 ;
     RECT  569.66 2195.66 570.14 2205.52 ;
     RECT  566.78 2084.36 571.3 2088.76 ;
     RECT  560.54 2284.7 572.54 2285.32 ;
     RECT  551.9 2297.3 572.54 2297.5 ;
     RECT  572.54 2284.7 573.7 2297.5 ;
     RECT  561.5 2334.26 573.98 2334.46 ;
     RECT  569.18 2312 575.14 2323.54 ;
     RECT  570.14 2193.98 575.42 2205.52 ;
     RECT  575.14 2312 575.62 2318.92 ;
     RECT  575.42 2193.98 576.1 2209.3 ;
     RECT  571.3 2084.36 576.58 2085.4 ;
     RECT  561.98 2239.34 577.54 2239.54 ;
     RECT  575.62 2312 577.54 2313.88 ;
     RECT  573.98 2273.36 578.02 2273.56 ;
     RECT  576.1 2195.66 578.3 2209.3 ;
     RECT  578.3 2195.66 579.74 2209.72 ;
     RECT  573.98 2334.26 582.14 2337.4 ;
     RECT  573.7 2297.3 582.34 2297.5 ;
     RECT  579.74 2195.66 582.62 2211.4 ;
     RECT  568.7 2103.26 583.78 2103.46 ;
     RECT  571.1 2396.84 585.02 2397.04 ;
     RECT  585.02 2396.84 585.98 2399.14 ;
     RECT  582.62 2195.66 586.18 2216.86 ;
     RECT  579.74 2250.26 586.94 2250.46 ;
     RECT  581.66 2137.7 588.1 2137.9 ;
     RECT  576.58 2085.2 589.82 2085.4 ;
     RECT  585.98 2096.12 589.82 2096.74 ;
     RECT  588.86 2322.92 589.82 2323.12 ;
     RECT  573.7 2284.7 590.5 2284.9 ;
     RECT  589.82 2322.92 592.22 2325.64 ;
     RECT  582.14 2334.26 592.22 2337.82 ;
     RECT  577.54 2313.68 592.7 2313.88 ;
     RECT  592.22 2322.92 592.7 2337.82 ;
     RECT  586.18 2211.2 592.9 2216.86 ;
     RECT  469 0 593 178 ;
     RECT  586.94 2073.44 593.66 2073.64 ;
     RECT  589.82 2085.2 593.66 2096.74 ;
     RECT  592.7 2313.68 594.14 2337.82 ;
     RECT  591.26 2118.8 595.58 2119 ;
     RECT  593.66 2073.44 596.26 2096.74 ;
     RECT  591.26 2273.36 598.18 2273.56 ;
     RECT  586.18 2195.66 598.46 2201.32 ;
     RECT  595.58 2118.38 600.1 2119 ;
     RECT  584.54 2179.28 601.06 2179.48 ;
     RECT  479 3222 603 3400 ;
     RECT  600.1 2118.8 603.94 2119 ;
     RECT  586.46 2167.94 604.42 2168.14 ;
     RECT  598.46 2193.98 604.7 2201.32 ;
     RECT  592.9 2211.2 604.7 2211.4 ;
     RECT  604.7 2193.98 604.9 2211.4 ;
     RECT  594.14 2311.58 605.18 2337.82 ;
     RECT  596.26 2080.58 606.82 2096.74 ;
     RECT  604.9 2209.1 607.58 2211.4 ;
     RECT  586.94 2246.48 608.54 2250.46 ;
     RECT  606.82 2088.56 610.18 2096.74 ;
     RECT  605.18 2310.32 611.14 2337.82 ;
     RECT  610.18 2092.34 611.42 2096.74 ;
     RECT  607.58 2107.04 611.42 2107.24 ;
     RECT  611.9 2282.18 612.38 2282.38 ;
     RECT  610.46 2163.74 613.06 2163.94 ;
     RECT  604.9 2195.66 613.34 2198.38 ;
     RECT  611.42 2092.34 613.54 2107.24 ;
     RECT  601.82 2235.56 614.3 2235.76 ;
     RECT  613.54 2092.34 614.98 2100.94 ;
     RECT  607.58 2209.1 617.18 2216.44 ;
     RECT  613.34 2190.2 617.38 2198.38 ;
     RECT  615.74 2363.66 617.38 2363.86 ;
     RECT  612.38 2276.72 617.86 2282.38 ;
     RECT  610.46 2296.88 618.14 2297.08 ;
     RECT  617.38 2190.62 618.34 2198.38 ;
     RECT  611.9 2265.8 618.62 2266 ;
     RECT  618.14 2295.62 619.1 2297.08 ;
     RECT  611.14 2311.58 619.3 2337.82 ;
     RECT  178 2383.82 619.58 2384.02 ;
     RECT  585.98 2393.9 619.58 2399.14 ;
     RECT  614.98 2096.54 620.74 2096.74 ;
     RECT  614.3 2231.78 621.02 2235.76 ;
     RECT  608.54 2246.48 621.02 2254.66 ;
     RECT  617.86 2277.14 621.02 2282.38 ;
     RECT  621.02 2277.14 621.98 2282.8 ;
     RECT  621.98 2277.14 622.46 2283.22 ;
     RECT  619.1 2295.62 622.46 2300.02 ;
     RECT  617.18 2209.1 622.66 2221.06 ;
     RECT  621.02 2231.78 623.42 2254.66 ;
     RECT  618.62 2265.8 623.42 2266.42 ;
     RECT  623.42 2231.78 624.1 2266.42 ;
     RECT  619.3 2312 624.1 2337.82 ;
     RECT  624.1 2242.28 624.58 2266.42 ;
     RECT  622.66 2217.08 626.3 2221.06 ;
     RECT  624.1 2231.78 626.3 2231.98 ;
     RECT  618.34 2195.66 627.94 2198.38 ;
     RECT  626.3 2217.08 627.94 2231.98 ;
     RECT  627.94 2228.42 629.38 2231.98 ;
     RECT  624.58 2242.28 630.34 2263.06 ;
     RECT  622.46 2277.14 630.82 2300.02 ;
     RECT  629.38 2231.78 631.3 2231.98 ;
     RECT  624.1 2315.36 631.58 2337.82 ;
     RECT  631.58 2315.36 633.02 2338.24 ;
     RECT  630.82 2277.56 633.7 2300.02 ;
     RECT  633.02 2311.16 633.7 2338.24 ;
     RECT  633.7 2281.76 634.18 2300.02 ;
     RECT  630.34 2246.48 638.02 2263.06 ;
     RECT  627.94 2195.66 638.98 2195.86 ;
     RECT  619.58 2383.82 639.74 2399.14 ;
     RECT  613.34 2408.6 640.22 2408.8 ;
     RECT  634.18 2282.18 640.7 2300.02 ;
     RECT  633.7 2311.16 642.34 2337.82 ;
     RECT  642.34 2315.78 645.22 2337.82 ;
     RECT  640.7 2282.18 645.98 2302.54 ;
     RECT  627.94 2217.08 646.66 2217.28 ;
     RECT  645.98 2282.18 646.66 2303.8 ;
     RECT  577.82 2049.5 646.94 2049.7 ;
     RECT  638.02 2250.26 647.62 2263.06 ;
     RECT  639.74 2383.82 649.34 2399.56 ;
     RECT  640.22 2408.6 649.34 2412.16 ;
     RECT  604.7 2348.12 650.5 2348.32 ;
     RECT  647.62 2250.26 650.98 2258.86 ;
     RECT  650.3 2202.38 654.82 2202.58 ;
     RECT  646.66 2295.62 655.3 2303.8 ;
     RECT  655.3 2296.04 656.06 2303.8 ;
     RECT  645.22 2323.76 658.66 2337.82 ;
     RECT  650.98 2250.26 659.62 2250.46 ;
     RECT  656.06 2296.04 660.38 2310.94 ;
     RECT  649.34 2383.82 661.06 2412.16 ;
     RECT  660.38 2296.04 662.5 2319.34 ;
     RECT  593 -70 663 178 ;
     RECT  661.06 2391.8 665.66 2412.16 ;
     RECT  648.86 2515.28 668.54 2515.48 ;
     RECT  668.54 2515.28 669.02 2520.94 ;
     RECT  663.26 1941.14 670.94 1941.34 ;
     RECT  603 3222 673 3470 ;
     RECT  668.54 1955.42 676.22 1955.62 ;
     RECT  676.22 1955.42 681.02 1961.08 ;
     RECT  669.02 2507.3 681.02 2520.94 ;
     RECT  669.02 1910.06 681.5 1910.26 ;
     RECT  681.02 2507.3 681.5 2525.14 ;
     RECT  681.5 2128.88 681.7 2137.9 ;
     RECT  681.02 1955.42 681.98 1962.76 ;
     RECT  681.98 2553.5 682.46 2553.7 ;
     RECT  682.46 2170.88 682.94 2171.08 ;
     RECT  681.7 2128.88 683.14 2129.08 ;
     RECT  681.7 2137.7 683.14 2137.9 ;
     RECT  682.94 2170.88 683.14 2172.34 ;
     RECT  662.5 2296.04 686.5 2310.94 ;
     RECT  668.06 2375.84 686.98 2376.04 ;
     RECT  682.94 1899.14 687.26 1899.34 ;
     RECT  646.66 2282.18 687.46 2282.38 ;
     RECT  670.94 1941.14 687.74 1945.12 ;
     RECT  680.54 1930.22 688.22 1930.42 ;
     RECT  650.3 2422.46 688.22 2422.66 ;
     RECT  668.06 1982.3 688.7 1982.5 ;
     RECT  688.7 1982.3 689.18 1985.02 ;
     RECT  681.5 2506.46 689.18 2525.14 ;
     RECT  668.06 2537.54 689.18 2537.74 ;
     RECT  687.26 1896.2 689.66 1899.34 ;
     RECT  683.42 2565.68 690.14 2565.88 ;
     RECT  681.5 1910.06 690.62 1914.46 ;
     RECT  688.22 1930.22 690.62 1930.84 ;
     RECT  679.1 1971.38 690.62 1971.58 ;
     RECT  689.18 1982.3 690.62 1985.44 ;
     RECT  690.14 2565.26 690.62 2565.88 ;
     RECT  690.62 1971.38 691.1 1985.44 ;
     RECT  646.94 2044.46 691.1 2049.7 ;
     RECT  689.66 1896.2 691.58 1900.6 ;
     RECT  676.22 2361.56 691.58 2361.76 ;
     RECT  688.7 2484.2 691.58 2484.4 ;
     RECT  690.62 1910.06 692.06 1930.84 ;
     RECT  687.74 1941.14 692.06 1945.54 ;
     RECT  692.06 1910.06 692.54 1945.54 ;
     RECT  681.98 1954.16 692.54 1962.76 ;
     RECT  692.06 2226.32 692.54 2228.2 ;
     RECT  691.1 1971.38 693 1987.12 ;
     RECT  635.42 2012.12 693.135 2012.32 ;
     RECT  691.58 2022.62 693.135 2022.82 ;
     RECT  686.5 2296.04 693.135 2304.22 ;
     RECT  682.46 2553.5 693.135 2556.22 ;
     RECT  691.1 2152.4 693.22 2153.44 ;
     RECT  691.58 2357.78 693.22 2361.76 ;
     RECT  693.135 2012.12 694.865 2022.82 ;
     RECT  693.135 2283.28 694.865 2304.22 ;
     RECT  691.58 1892.84 695.42 1900.6 ;
     RECT  692.54 1910.06 695.42 1962.76 ;
     RECT  693 1971.38 695.6 1996.8 ;
     RECT  690.62 2565.26 695.6 2573.02 ;
     RECT  693 2583.32 695.6 2585.32 ;
     RECT  693.135 2547.76 695.735 2556.22 ;
     RECT  695.6 2565.26 695.735 2585.32 ;
     RECT  691.1 2044.46 697.34 2052.64 ;
     RECT  692.06 2065.04 697.34 2065.24 ;
     RECT  695.735 2027.92 697.465 2033.4 ;
     RECT  693.22 2361.56 698.5 2361.76 ;
     RECT  689.18 2506.46 698.5 2537.74 ;
     RECT  695.735 2547.76 698.5 2585.32 ;
     RECT  691.1 2376.68 698.78 2376.88 ;
     RECT  698.5 2507.3 698.98 2515.48 ;
     RECT  698.5 2527.04 698.98 2537.74 ;
     RECT  698.5 2547.76 698.98 2565.46 ;
     RECT  692.54 2105.78 699.26 2105.98 ;
     RECT  692.54 2226.32 699.26 2234.92 ;
     RECT  658.66 2330.06 699.26 2337.82 ;
     RECT  691.58 2484.2 699.46 2491.96 ;
     RECT  697.34 2044.46 699.74 2065.24 ;
     RECT  699.26 2102 699.74 2105.98 ;
     RECT  699.26 2226.32 699.74 2238.7 ;
     RECT  698.78 2376.26 699.74 2376.88 ;
     RECT  699.46 2484.2 699.94 2491.54 ;
     RECT  692.54 2084.36 700.22 2084.56 ;
     RECT  699.74 2094.44 700.22 2105.98 ;
     RECT  699.74 2217.08 700.22 2217.28 ;
     RECT  688.22 2422.46 700.22 2426.86 ;
     RECT  680.54 2448.08 700.22 2448.28 ;
     RECT  699.74 2472.86 700.22 2473.06 ;
     RECT  699.94 2484.2 700.22 2484.4 ;
     RECT  700.22 2217.08 700.38 2217.7 ;
     RECT  699.74 2226.32 700.38 2239.12 ;
     RECT  687.74 2256.14 700.38 2256.34 ;
     RECT  699.26 2330.06 700.38 2339.92 ;
     RECT  699.74 2044.46 700.46 2066.5 ;
     RECT  698.98 2529.56 700.46 2537.74 ;
     RECT  698.98 2547.76 700.46 2558.32 ;
     RECT  700.38 2255.68 701.34 2256.34 ;
     RECT  700.22 2267.9 701.34 2275.66 ;
     RECT  694.865 2284.66 701.34 2304.22 ;
     RECT  700.22 2421.62 701.34 2426.86 ;
     RECT  700.22 2439.26 701.34 2484.4 ;
     RECT  695.42 1892.84 701.38 1962.76 ;
     RECT  700.46 2036.48 701.86 2066.5 ;
     RECT  701.34 2421.62 702.02 2484.4 ;
     RECT  700.22 2174.66 702.14 2174.86 ;
     RECT  701.38 1892.84 702.34 1900.6 ;
     RECT  701.86 2039 702.34 2066.5 ;
     RECT  698.3 2124.26 702.78 2124.46 ;
     RECT  701.38 1910.06 702.82 1962.76 ;
     RECT  702.34 2041.52 702.82 2066.5 ;
     RECT  702.82 1930.64 703.1 1962.76 ;
     RECT  695.6 1971.38 703.1 1999.4 ;
     RECT  702.82 2044.04 703.26 2066.5 ;
     RECT  700.22 2083.94 703.26 2084.56 ;
     RECT  687.26 2201.54 703.26 2201.74 ;
     RECT  699.74 2376.26 703.26 2381.08 ;
     RECT  702.14 2174.66 703.74 2179.06 ;
     RECT  703.1 1930.64 703.78 1999.4 ;
     RECT  702.78 2124.26 703.78 2130.3 ;
     RECT  703.26 2044.04 704.74 2084.56 ;
     RECT  703.74 2172.52 705.02 2179.06 ;
     RECT  705.02 2172.52 705.5 2179.48 ;
     RECT  700.22 2188.94 705.5 2190.4 ;
     RECT  705.5 2172.52 705.66 2190.4 ;
     RECT  703.26 2201.54 705.66 2202.54 ;
     RECT  700.38 2322.88 705.66 2339.92 ;
     RECT  703.78 1930.64 705.7 1972.42 ;
     RECT  700.38 2217.08 706.46 2239.12 ;
     RECT  702.34 1892.84 706.66 1899.34 ;
     RECT  704.74 2044.46 707.1 2084.56 ;
     RECT  700.22 2094.44 707.1 2107.24 ;
     RECT  703.78 2130.1 707.1 2130.3 ;
     RECT  700.22 2141.48 707.1 2144.2 ;
     RECT  705.66 2172.52 707.1 2202.54 ;
     RECT  706.46 2217.08 707.1 2241.64 ;
     RECT  701.34 2255.68 707.1 2275.66 ;
     RECT  701.34 2284.66 707.1 2305.44 ;
     RECT  705.66 2316.16 707.1 2339.92 ;
     RECT  703.26 2373.28 707.1 2381.08 ;
     RECT  706.66 1899.14 707.62 1899.34 ;
     RECT  703.78 1982.3 708.38 1999.4 ;
     RECT  694.865 2012.12 708.38 2012.32 ;
     RECT  702.82 1910.06 708.58 1922.02 ;
     RECT  705.7 1930.64 708.58 1962.76 ;
     RECT  665.66 2391.8 708.86 2412.58 ;
     RECT  702.02 2421.62 708.86 2426.86 ;
     RECT  708.58 1935.68 709.06 1962.76 ;
     RECT  700.46 2529.56 709.06 2558.32 ;
     RECT  708.58 1914.26 712.9 1922.02 ;
     RECT  709.06 1941.14 712.9 1962.76 ;
     RECT  709.06 2558.12 712.9 2558.32 ;
     RECT  708.86 2391.8 713.38 2426.86 ;
     RECT  705.7 1971.38 714.14 1972.42 ;
     RECT  708.38 1982.3 714.14 2012.32 ;
     RECT  709.06 2529.56 714.34 2549.08 ;
     RECT  714.14 1971.38 714.82 2012.32 ;
     RECT  714.34 2541.74 714.82 2549.08 ;
     RECT  712.9 1960.88 716.06 1962.76 ;
     RECT  714.82 1971.38 716.06 1971.58 ;
     RECT  709.82 2025.98 717.02 2026.18 ;
     RECT  712.9 1914.26 717.7 1914.46 ;
     RECT  707.1 2044.46 717.7 2118.96 ;
     RECT  717.02 2022.62 719.9 2026.18 ;
     RECT  714.82 1982.3 720.1 1983.76 ;
     RECT  712.9 1941.14 721.82 1948.9 ;
     RECT  716.06 1960.88 721.82 1971.58 ;
     RECT  721.82 1941.14 722.3 1971.58 ;
     RECT  722.3 1936.52 722.78 1971.58 ;
     RECT  707.1 2350.6 722.94 2350.8 ;
     RECT  722.78 1935.68 724.7 1971.58 ;
     RECT  722.94 2350.6 724.86 2353.74 ;
     RECT  707.1 2365.72 724.86 2381.08 ;
     RECT  714.82 2543 724.9 2549.08 ;
     RECT  724.7 1935.68 729.98 1972 ;
     RECT  724.9 2543 730.18 2543.2 ;
     RECT  729.98 1935.68 731.62 1976.2 ;
     RECT  719.9 2022.62 731.9 2027.02 ;
     RECT  713.38 2391.8 732.86 2412.58 ;
     RECT  713.38 2421.62 732.86 2426.86 ;
     RECT  700.22 1832.36 736.7 1832.56 ;
     RECT  707.1 2130.1 736.86 2341.14 ;
     RECT  724.86 2350.6 736.86 2381.08 ;
     RECT  731.42 1985.24 737.66 1985.44 ;
     RECT  714.82 1994.8 737.66 2012.32 ;
     RECT  732.86 2391.8 737.66 2426.86 ;
     RECT  702.02 2439.26 737.86 2484.4 ;
     RECT  717.7 2044.46 741.7 2050.54 ;
     RECT  727.1 1925.6 744.86 1925.8 ;
     RECT  731.62 1935.68 744.86 1971.58 ;
     RECT  717.7 2060.8 756.06 2118.96 ;
     RECT  756.06 2060.8 761.82 2119.38 ;
     RECT  736.86 2130.1 761.82 2381.08 ;
     RECT  761.82 2060.8 786.82 2381.08 ;
     RECT  663 0 787 178 ;
     RECT  786.82 2060.8 796.38 2376.42 ;
     RECT  673 3222 797 3400 ;
     RECT  808.7 1657.64 819.94 1657.84 ;
     RECT  813.02 1703 827.14 1703.2 ;
     RECT  796.38 2060.8 829.5 2378.52 ;
     RECT  815.42 1733.24 830.02 1733.44 ;
     RECT  827.42 1771.04 834.34 1771.24 ;
     RECT  818.3 1676.12 837.22 1676.32 ;
     RECT  698.98 2511.88 842.3 2515.48 ;
     RECT  818.78 1713.92 844.42 1714.12 ;
     RECT  829.5 2060.8 848.22 2379.36 ;
     RECT  842.3 1741.22 856.42 1741.42 ;
     RECT  787 -70 857 178 ;
     RECT  741.7 2044.46 861.18 2050.12 ;
     RECT  848.22 2060.8 861.18 2380.2 ;
     RECT  797 3222 867 3470 ;
     RECT  178 1414.04 867.46 1414.24 ;
     RECT  871.1 1727.36 871.3 1727.98 ;
     RECT  869.18 1771.04 872.06 1771.24 ;
     RECT  871.3 1727.78 872.74 1727.98 ;
     RECT  872.06 1771.04 872.74 1774.18 ;
     RECT  857.18 1718.12 873.22 1718.32 ;
     RECT  872.74 1773.98 873.22 1774.18 ;
     RECT  870.62 1741.22 875.14 1741.42 ;
     RECT  875.42 1878.98 883.58 1879.18 ;
     RECT  883.58 1878.56 886.66 1879.18 ;
     RECT  855.74 1804.64 895.58 1804.84 ;
     RECT  878.78 1691.24 896.26 1691.44 ;
     RECT  861.18 2044.46 897.86 2380.2 ;
     RECT  900.38 1679.9 900.58 1680.94 ;
     RECT  856.7 1610.18 900.86 1610.38 ;
     RECT  900.86 1604.72 901.06 1610.38 ;
     RECT  895.58 1801.28 901.06 1804.84 ;
     RECT  900.58 1679.9 902.02 1680.1 ;
     RECT  891.74 1627.4 903.46 1627.6 ;
     RECT  901.06 1604.72 904.305 1604.92 ;
     RECT  890.3 1759.28 904.42 1759.48 ;
     RECT  886.66 1878.56 904.42 1878.76 ;
     RECT  897.86 2059.54 909.66 2380.2 ;
     RECT  737.66 2391.8 909.66 2428.96 ;
     RECT  901.06 1804.64 913.06 1804.84 ;
     RECT  883.1 1786.16 914.78 1786.36 ;
     RECT  892.22 1770.2 915.46 1770.4 ;
     RECT  897.86 2044.46 915.9 2050.12 ;
     RECT  909.66 2059.54 915.9 2428.96 ;
     RECT  914.78 1785.74 915.94 1786.36 ;
     RECT  915.9 2044.46 916.1 2428.96 ;
     RECT  889.34 1576.58 916.42 1576.78 ;
     RECT  910.94 1680.32 917.18 1680.52 ;
     RECT  883.58 1727.78 918.14 1727.98 ;
     RECT  917.18 1676.96 918.82 1680.52 ;
     RECT  918.14 1725.68 920.54 1728.82 ;
     RECT  920.54 1722.32 921.5 1728.82 ;
     RECT  744.86 1925.6 921.7 1971.58 ;
     RECT  921.5 1476.62 923.14 1476.82 ;
     RECT  916.1 2044.46 925.98 2050.12 ;
     RECT  916.1 2058.7 925.98 2428.96 ;
     RECT  841.82 1531.64 926.3 1531.84 ;
     RECT  919.1 1551.38 928.9 1551.58 ;
     RECT  918.82 1680.32 930.82 1680.52 ;
     RECT  925.98 2044.46 931.94 2428.96 ;
     RECT  910.94 1758.02 936.38 1758.22 ;
     RECT  936.38 1758.02 936.86 1764.52 ;
     RECT  920.54 1512.32 937.06 1512.52 ;
     RECT  931.94 2044.46 937.7 2111.82 ;
     RECT  936.86 1758.02 938.78 1767.04 ;
     RECT  937.7 2058.7 940.38 2111.82 ;
     RECT  931.94 2121.7 940.38 2428.96 ;
     RECT  940.38 2058.7 945.38 2428.96 ;
     RECT  945.38 2119.18 946.34 2428.96 ;
     RECT  606.62 1501.4 947.42 1501.6 ;
     RECT  938.78 1758.02 947.62 1771.66 ;
     RECT  941.18 1812.2 948.38 1812.4 ;
     RECT  945.38 2058.7 948.74 2105.1 ;
     RECT  946.34 2119.18 948.74 2380.2 ;
     RECT  950.78 1702.16 951.94 1702.78 ;
     RECT  947.62 1758.02 951.94 1767.04 ;
     RECT  949.34 1713.5 952.7 1713.7 ;
     RECT  921.5 1722.32 952.7 1729.24 ;
     RECT  948.38 1804.64 953.86 1812.4 ;
     RECT  948.74 2122.54 954.98 2380.2 ;
     RECT  953.66 1434.2 955.3 1434.4 ;
     RECT  926.3 1531.64 955.78 1536.88 ;
     RECT  951.94 1766.84 955.78 1767.04 ;
     RECT  915.94 1786.16 957.5 1786.36 ;
     RECT  842.3 2511.88 957.5 2516.32 ;
     RECT  953.86 1804.64 957.7 1804.84 ;
     RECT  957.5 2508.98 957.7 2516.32 ;
     RECT  948.74 2059.12 958.34 2105.1 ;
     RECT  937.7 2044.46 958.62 2050.12 ;
     RECT  947.42 1501.4 958.94 1509.16 ;
     RECT  654.62 1521.14 958.94 1521.34 ;
     RECT  958.34 2066.68 961.7 2105.1 ;
     RECT  954.98 2122.54 963.62 2129.04 ;
     RECT  961.7 2084.32 964.1 2105.1 ;
     RECT  957.5 1780.28 965.66 1786.36 ;
     RECT  965.18 1466.12 966.34 1466.32 ;
     RECT  958.62 2044.46 967.94 2055.12 ;
     RECT  954.98 2137.66 968.22 2380.2 ;
     RECT  946.34 2391.8 968.22 2428.96 ;
     RECT  968.22 2137.66 968.42 2428.96 ;
     RECT  964.7 1377.92 968.54 1378.12 ;
     RECT  961.7 2066.68 969.38 2070.24 ;
     RECT  957.5 1697.54 969.98 1697.74 ;
     RECT  958.94 1501.4 970.66 1521.34 ;
     RECT  961.34 1544.24 970.66 1544.44 ;
     RECT  969.38 2068.36 971.3 2070.24 ;
     RECT  969.98 1693.76 971.62 1697.74 ;
     RECT  959.9 1669.4 971.9 1669.6 ;
     RECT  965.66 1780.28 971.9 1793.92 ;
     RECT  736.7 1832.36 971.9 1838.02 ;
     RECT  971.9 1669.4 972.1 1678.42 ;
     RECT  968.42 2137.66 972.26 2223.96 ;
     RECT  972.38 1873.1 973.34 1873.3 ;
     RECT  971.9 1774.4 973.54 1793.92 ;
     RECT  964.1 2085.16 973.7 2105.1 ;
     RECT  973.34 1873.1 974.02 1879.6 ;
     RECT  951.94 1758.02 974.3 1758.22 ;
     RECT  972.1 1669.4 974.98 1678 ;
     RECT  971.9 1829 974.98 1838.02 ;
     RECT  974.02 1873.94 974.98 1879.6 ;
     RECT  974.98 1876.88 975.46 1879.6 ;
     RECT  974.3 1752.14 975.74 1758.22 ;
     RECT  973.54 1780.28 975.74 1793.92 ;
     RECT  974.78 1804.64 975.74 1804.84 ;
     RECT  739.1 1914.68 976.7 1914.88 ;
     RECT  952.7 1713.5 976.9 1729.24 ;
     RECT  974.98 1832.36 977.18 1838.02 ;
     RECT  968.54 1377.5 977.38 1378.12 ;
     RECT  977.18 790.76 977.66 790.96 ;
     RECT  970.66 1518.2 978.62 1521.34 ;
     RECT  955.78 1531.64 978.62 1531.84 ;
     RECT  973.7 2085.16 978.78 2099.22 ;
     RECT  968.42 2232.58 979.46 2428.96 ;
     RECT  975.74 1748.36 979.78 1758.22 ;
     RECT  972.26 2137.66 980.7 2223.12 ;
     RECT  979.46 2232.58 980.7 2380.2 ;
     RECT  857 0 981 178 ;
     RECT  978.62 1518.2 981.22 1531.84 ;
     RECT  979.78 1751.72 981.22 1758.22 ;
     RECT  959.9 1566.92 982.18 1567.12 ;
     RECT  974.98 1669.4 983.14 1669.6 ;
     RECT  978.14 776.06 983.42 776.26 ;
     RECT  977.66 790.76 983.42 791.38 ;
     RECT  983.42 776.06 984.38 791.38 ;
     RECT  975.74 1780.28 984.58 1804.84 ;
     RECT  984.38 769.76 984.86 791.38 ;
     RECT  977.18 1832.36 984.86 1846 ;
     RECT  983.42 1900.82 985.82 1901.02 ;
     RECT  978.78 2084.74 986.18 2099.22 ;
     RECT  976.7 1914.68 986.3 1917.4 ;
     RECT  921.7 1926.86 986.3 1971.58 ;
     RECT  977.38 1377.92 986.5 1378.12 ;
     RECT  970.46 1467.38 986.98 1467.58 ;
     RECT  981.22 1753.4 986.98 1758.22 ;
     RECT  984.06 2113.3 987.62 2114.34 ;
     RECT  976.9 1713.5 987.94 1718.32 ;
     RECT  980.7 2137.66 988.1 2380.2 ;
     RECT  976.22 1410.68 989.66 1410.88 ;
     RECT  970.66 1501.4 989.66 1509.16 ;
     RECT  985.82 1900.82 989.66 1901.44 ;
     RECT  986.3 1914.68 989.66 1971.58 ;
     RECT  989.66 1408.16 990.34 1410.88 ;
     RECT  981.22 1521.14 990.34 1531.84 ;
     RECT  990.14 841.58 990.62 841.78 ;
     RECT  968.54 1593.38 990.62 1593.58 ;
     RECT  990.62 1593.38 990.82 1596.94 ;
     RECT  963.62 2122.96 990.98 2129.04 ;
     RECT  867 3222 991 3400 ;
     RECT  956.54 1431.68 991.1 1431.88 ;
     RECT  984.86 1830.68 991.1 1846 ;
     RECT  989.66 1501.4 991.78 1512.1 ;
     RECT  986.18 2085.16 991.94 2099.22 ;
     RECT  979.46 2391.34 991.94 2428.96 ;
     RECT  991.1 758.42 992.06 758.62 ;
     RECT  971.62 1697.54 992.06 1697.74 ;
     RECT  957.5 1864.28 992.06 1864.48 ;
     RECT  990.98 2122.96 992.22 2126.52 ;
     RECT  992.22 2119.6 992.42 2126.52 ;
     RECT  992.06 1697.54 992.74 1699.42 ;
     RECT  971.3 2068.36 992.9 2068.56 ;
     RECT  983.9 960.02 993.135 960.22 ;
     RECT  992.74 1699.22 993.7 1699.42 ;
     RECT  993.135 947.2 993.98 960.22 ;
     RECT  992.42 2119.6 994.82 2119.8 ;
     RECT  993.135 616.6 994.865 622.08 ;
     RECT  993.98 947.2 994.865 964.84 ;
     RECT  991.58 804.62 994.94 804.82 ;
     RECT  993 984.24 994.94 986.24 ;
     RECT  991.94 2085.16 995.3 2092.5 ;
     RECT  994.865 952.04 995.42 964.84 ;
     RECT  993 594.8 995.6 596.8 ;
     RECT  994.94 984.24 995.6 987.1 ;
     RECT  984.86 769.76 995.735 793.9 ;
     RECT  994.94 804.62 995.735 806.08 ;
     RECT  995.3 2091.88 996.26 2092.5 ;
     RECT  995.42 952.04 996.38 966.52 ;
     RECT  994.94 1892 996.38 1892.2 ;
     RECT  989.66 1900.82 996.38 1971.58 ;
     RECT  988.1 2137.66 996.54 2223.96 ;
     RECT  988.1 2232.58 996.54 2380.2 ;
     RECT  984.58 1798.76 996.58 1804.84 ;
     RECT  991.1 1830.68 996.86 1849.36 ;
     RECT  996.38 1892 996.86 1971.58 ;
     RECT  995.735 769.76 997.34 806.08 ;
     RECT  986.98 1753.4 997.34 1757.8 ;
     RECT  984.38 1770.2 997.34 1770.4 ;
     RECT  995.735 628 997.465 633.48 ;
     RECT  996.58 1798.76 997.54 1798.96 ;
     RECT  994.94 1818.92 997.54 1819.12 ;
     RECT  996.86 928.52 998.02 928.72 ;
     RECT  997.34 1753.4 998.02 1770.4 ;
     RECT  996.86 1891.16 998.3 1971.58 ;
     RECT  997.34 769.76 998.5 806.5 ;
     RECT  995.6 981.64 998.98 987.1 ;
     RECT  998.5 771.68 999.26 806.5 ;
     RECT  998.78 870.14 999.26 870.34 ;
     RECT  976.7 741.2 999.46 741.4 ;
     RECT  984.58 1780.28 999.46 1786.36 ;
     RECT  998.3 1814.72 999.46 1814.92 ;
     RECT  999.26 771.68 999.74 812.8 ;
     RECT  999.74 771.68 1000.22 816.58 ;
     RECT  999.26 863.42 1000.22 870.34 ;
     RECT  996.38 952.04 1000.42 967.78 ;
     RECT  990.62 834.02 1000.46 841.78 ;
     RECT  1000.42 957.08 1000.46 967.78 ;
     RECT  1000.22 858.8 1000.7 870.34 ;
     RECT  996.86 1830.68 1000.7 1850.2 ;
     RECT  998.02 1753.4 1000.9 1757.8 ;
     RECT  999.46 1785.32 1000.9 1786.36 ;
     RECT  998.3 1886.54 1001.18 1971.58 ;
     RECT  1000.46 957.08 1001.86 971.98 ;
     RECT  975.46 1876.88 1001.86 1877.08 ;
     RECT  1000.46 826.88 1002.3 846.4 ;
     RECT  996.54 2137.66 1002.3 2380.2 ;
     RECT  991.94 2391.8 1002.3 2428.96 ;
     RECT  1001.86 964.64 1002.34 971.98 ;
     RECT  1001.18 1886.12 1002.62 1971.58 ;
     RECT  1000.22 771.68 1002.78 817.42 ;
     RECT  1002.3 826.88 1002.78 847.48 ;
     RECT  1000.46 921.38 1002.82 921.58 ;
     RECT  1000.9 1753.4 1002.82 1754.44 ;
     RECT  1000.46 745.4 1003.26 745.6 ;
     RECT  992.06 755.06 1003.26 758.62 ;
     RECT  1002.78 771.68 1003.26 847.48 ;
     RECT  1000.7 858.8 1003.26 871.18 ;
     RECT  998.02 1770.2 1003.3 1770.4 ;
     RECT  1000.7 1826.9 1003.3 1850.2 ;
     RECT  1002.62 1879.82 1003.3 1971.58 ;
     RECT  1000.46 931.88 1003.78 943 ;
     RECT  980.54 1388.84 1003.78 1389.04 ;
     RECT  990.34 1408.16 1003.78 1408.36 ;
     RECT  1002.34 970.1 1004.06 971.98 ;
     RECT  1004.06 970.1 1004.26 972.4 ;
     RECT  1002.82 1753.4 1004.26 1753.6 ;
     RECT  1003.78 931.88 1004.74 939.64 ;
     RECT  1003.3 1826.9 1004.74 1827.1 ;
     RECT  1003.3 1835.72 1005.22 1850.2 ;
     RECT  1005.22 1837.82 1005.98 1850.2 ;
     RECT  992.06 1860.92 1005.98 1864.48 ;
     RECT  1004.74 939.44 1006.66 939.64 ;
     RECT  990.82 1596.74 1006.66 1596.94 ;
     RECT  1003.26 745.4 1007.1 759.28 ;
     RECT  1003.26 771.68 1007.1 871.18 ;
     RECT  1006.46 1823.54 1007.62 1824.16 ;
     RECT  1005.98 1837.82 1007.9 1864.48 ;
     RECT  1007.9 1837.82 1008.1 1866.16 ;
     RECT  1003.3 1886.96 1008.58 1971.58 ;
     RECT  991.78 1501.4 1008.86 1509.16 ;
     RECT  1007.1 745.4 1009.06 871.18 ;
     RECT  1008.38 1571.54 1009.54 1571.74 ;
     RECT  1004.26 972.2 1010.02 972.4 ;
     RECT  1007.62 1823.96 1010.02 1824.16 ;
     RECT  1008.1 1861.76 1010.02 1866.16 ;
     RECT  1008.86 1500.98 1010.5 1509.16 ;
     RECT  1007.9 1808.42 1010.5 1809.88 ;
     RECT  1009.06 749 1010.98 871.18 ;
     RECT  1010.5 1501.4 1013.18 1509.16 ;
     RECT  1010.98 813.44 1013.38 871.18 ;
     RECT  1010.78 1362.8 1013.38 1363 ;
     RECT  1007.9 1461.08 1014.82 1461.28 ;
     RECT  1010.5 1809.68 1015.3 1809.88 ;
     RECT  1000.9 1786.16 1016.54 1786.36 ;
     RECT  987.94 1718.12 1016.74 1718.32 ;
     RECT  976.9 1729.04 1017.98 1729.24 ;
     RECT  1016.54 1779.86 1018.18 1786.36 ;
     RECT  1010.98 749 1018.66 802.12 ;
     RECT  1017.98 1729.04 1018.66 1734.7 ;
     RECT  1008.38 1763.9 1018.94 1764.1 ;
     RECT  1018.94 1457.3 1019.42 1457.5 ;
     RECT  1017.98 1686.2 1020.1 1686.4 ;
     RECT  1013.38 813.44 1020.58 863.62 ;
     RECT  1013.18 1501.4 1021.06 1510.84 ;
     RECT  1018.66 1732.82 1021.54 1734.7 ;
     RECT  990.34 1531.64 1021.82 1531.84 ;
     RECT  1008.58 1886.96 1022.02 1905.22 ;
     RECT  1000.46 911.72 1022.5 911.92 ;
     RECT  1002.3 2137.66 1022.66 2428.96 ;
     RECT  1021.34 1627.4 1022.98 1627.6 ;
     RECT  1018.94 1763.9 1022.98 1766.62 ;
     RECT  1021.82 1531.64 1023.46 1537.72 ;
     RECT  1022.78 1820.6 1023.74 1820.8 ;
     RECT  1018.18 1786.16 1023.94 1786.36 ;
     RECT  1023.74 1820.18 1023.94 1820.8 ;
     RECT  1022.98 1766.42 1025.66 1766.62 ;
     RECT  1025.18 1675.28 1025.86 1675.48 ;
     RECT  1025.66 1766.42 1026.34 1774.6 ;
     RECT  1007.9 1752.14 1028.06 1752.34 ;
     RECT  990.34 1521.14 1029.02 1521.34 ;
     RECT  1028.06 1469.06 1029.22 1469.26 ;
     RECT  1019.42 1456.88 1031.42 1457.5 ;
     RECT  1018.66 783.86 1031.58 802.12 ;
     RECT  1029.02 1521.14 1031.62 1521.76 ;
     RECT  1018.94 925.16 1032.86 925.36 ;
     RECT  1018.46 1810.1 1032.86 1810.3 ;
     RECT  1020.58 813.44 1033.06 855.04 ;
     RECT  1024.7 1794.14 1034.02 1794.34 ;
     RECT  1023.26 1562.72 1034.78 1562.92 ;
     RECT  1011.74 1479.98 1036.22 1480.18 ;
     RECT  1031.42 1456.88 1036.42 1460.86 ;
     RECT  1034.78 1562.72 1036.9 1570.48 ;
     RECT  1028.06 1750.46 1037.18 1752.34 ;
     RECT  1032.86 1810.1 1038.14 1817.86 ;
     RECT  1026.34 1766.42 1038.34 1766.62 ;
     RECT  1031.58 783.86 1038.78 802.54 ;
     RECT  1029.5 1582.04 1038.82 1582.24 ;
     RECT  1038.14 1804.64 1040.06 1817.86 ;
     RECT  1040.06 1804.64 1041.22 1826.26 ;
     RECT  1022.66 2137.66 1041.86 2380.62 ;
     RECT  1036.42 1457.3 1044.1 1460.86 ;
     RECT  1038.78 783.86 1045.22 806.32 ;
     RECT  1036.22 1479.56 1045.54 1480.18 ;
     RECT  1042.94 1829 1045.54 1829.2 ;
     RECT  1037.18 1744.58 1046.5 1752.34 ;
     RECT  1036.9 1570.28 1047.94 1570.48 ;
     RECT  1018.66 749 1050.3 771.88 ;
     RECT  1020.38 1328.78 1050.34 1328.98 ;
     RECT  991.1 1426.64 1050.34 1431.88 ;
     RECT  1041.86 2137.66 1050.98 2380.2 ;
     RECT  981 -70 1051 178 ;
     RECT  1050.98 2137.66 1051.46 2221.86 ;
     RECT  1045.54 1479.98 1052.26 1480.18 ;
     RECT  1043.42 1713.92 1052.26 1714.12 ;
     RECT  1051.46 2137.66 1052.9 2216.82 ;
     RECT  1050.98 2232.16 1052.9 2380.2 ;
     RECT  1046.5 1744.58 1053.98 1748.56 ;
     RECT  1052.9 2137.66 1054.14 2161.38 ;
     RECT  1041.22 1804.64 1055.14 1817.86 ;
     RECT  1050.34 1426.64 1055.62 1426.84 ;
     RECT  1053.98 1744.16 1056.1 1748.56 ;
     RECT  1033.06 817.88 1056.54 855.04 ;
     RECT  1056.1 1744.16 1057.54 1744.78 ;
     RECT  1044.1 1460.66 1058.3 1460.86 ;
     RECT  1058.3 1460.66 1058.5 1461.7 ;
     RECT  1057.54 1744.58 1058.5 1744.78 ;
     RECT  1055.14 1810.1 1058.5 1817.86 ;
     RECT  1022.02 1886.96 1058.5 1904.8 ;
     RECT  1023.46 1531.64 1060.22 1531.84 ;
     RECT  991 3222 1061 3470 ;
     RECT  1054.14 2133.88 1063.46 2161.38 ;
     RECT  1060.22 1531.64 1063.78 1532.26 ;
     RECT  1045.22 783.86 1064.7 804.64 ;
     RECT  1064.54 1430.42 1065.7 1430.62 ;
     RECT  1064.7 783.86 1066.14 805.48 ;
     RECT  1063.46 2137.66 1066.34 2161.38 ;
     RECT  1010.02 1861.76 1070.98 1861.96 ;
     RECT  1062.3 877.94 1073.34 878.14 ;
     RECT  1065.98 1641.68 1073.38 1641.88 ;
     RECT  1050.3 749 1073.82 774.4 ;
     RECT  1066.14 783.02 1073.82 805.48 ;
     RECT  1072.7 1309.88 1074.34 1310.08 ;
     RECT  1072.7 1780.28 1075.1 1780.48 ;
     RECT  1068.38 1562.72 1075.58 1562.92 ;
     RECT  1071.74 1445.54 1075.78 1445.74 ;
     RECT  1057.82 1734.92 1075.78 1735.12 ;
     RECT  1075.58 1562.72 1076.74 1563.34 ;
     RECT  1031.62 1521.14 1077.02 1521.34 ;
     RECT  1073.82 749 1078.62 805.48 ;
     RECT  1075.1 1780.28 1079.14 1785.94 ;
     RECT  1066.34 2154.46 1079.58 2161.38 ;
     RECT  1052.9 2170.42 1079.58 2216.82 ;
     RECT  1073.34 877.94 1080.06 885.28 ;
     RECT  1052.9 2232.16 1080.26 2379.78 ;
     RECT  1056.54 817.88 1080.54 858.82 ;
     RECT  1080.86 1489.22 1081.06 1491.94 ;
     RECT  1079.58 2154.46 1081.22 2221.44 ;
     RECT  1081.06 1491.74 1081.54 1491.94 ;
     RECT  1081.22 2170.42 1081.7 2221.44 ;
     RECT  1063.78 1531.64 1081.82 1531.84 ;
     RECT  1080.38 1634.96 1081.82 1635.16 ;
     RECT  1081.7 2187.22 1082.18 2221.44 ;
     RECT  1069.82 1743.74 1082.5 1743.94 ;
     RECT  1081.34 1771.04 1082.78 1771.24 ;
     RECT  1079.14 1780.28 1082.78 1780.48 ;
     RECT  1081.82 1531.22 1083.46 1531.84 ;
     RECT  737.66 1985.24 1083.94 2012.32 ;
     RECT  1066.34 2137.66 1084.1 2143.74 ;
     RECT  1026.14 1681.16 1084.22 1681.36 ;
     RECT  1062.62 1725.68 1084.42 1725.88 ;
     RECT  1080.54 817.88 1084.58 861.34 ;
     RECT  1021.06 1501.4 1086.14 1509.16 ;
     RECT  1077.02 1521.14 1086.14 1521.76 ;
     RECT  1081.82 1634.96 1086.14 1642.3 ;
     RECT  1086.14 1501.4 1086.34 1521.76 ;
     RECT  1080.06 877.94 1086.78 893.68 ;
     RECT  1074.14 1325 1087.3 1325.2 ;
     RECT  1081.22 2154.46 1088.9 2161.38 ;
     RECT  1081.7 2170.42 1088.9 2176.08 ;
     RECT  1084.22 1676.12 1089.02 1681.36 ;
     RECT  1086.14 1634.96 1089.22 1642.72 ;
     RECT  1070.78 1760.12 1089.5 1760.32 ;
     RECT  1082.78 1771.04 1089.5 1780.48 ;
     RECT  714.34 2529.56 1089.7 2529.76 ;
     RECT  1082.18 2187.22 1089.86 2197.08 ;
     RECT  1008.58 1914.26 1089.98 1971.58 ;
     RECT  1089.5 1661.42 1090.66 1661.62 ;
     RECT  1076.74 1563.14 1090.94 1563.34 ;
     RECT  1089.5 1760.12 1090.94 1780.48 ;
     RECT  1089.98 1913.84 1092.1 1971.58 ;
     RECT  1088.9 2175.88 1092.74 2176.08 ;
     RECT  1089.22 1642.52 1093.34 1642.72 ;
     RECT  1078.62 749 1093.5 805.9 ;
     RECT  1084.58 817.88 1093.5 855.88 ;
     RECT  1093.5 816.2 1094.66 855.88 ;
     RECT  1094.78 1456.88 1095.46 1457.08 ;
     RECT  1090.94 1563.14 1095.46 1570.48 ;
     RECT  1090.94 1760.12 1095.46 1786.36 ;
     RECT  1095.26 1695.86 1095.74 1696.06 ;
     RECT  1089.86 2192.26 1095.9 2197.08 ;
     RECT  1095.26 1446.8 1095.94 1447 ;
     RECT  1093.34 1642.52 1095.94 1650.28 ;
     RECT  1082.18 2206.96 1096.1 2221.44 ;
     RECT  1086.34 1501.4 1096.22 1521.34 ;
     RECT  1083.46 1531.64 1096.22 1531.84 ;
     RECT  1095.46 1771.04 1096.22 1786.36 ;
     RECT  1094.78 1580.78 1096.42 1580.98 ;
     RECT  1089.02 1671.5 1096.7 1681.36 ;
     RECT  1096.22 1443.44 1096.9 1446.16 ;
     RECT  1096.1 2221.24 1097.06 2221.44 ;
     RECT  1095.46 1570.28 1097.38 1570.48 ;
     RECT  1086.78 869.96 1098.02 893.68 ;
     RECT  1096.1 2206.96 1098.02 2212.2 ;
     RECT  1098.02 869.96 1098.5 881.92 ;
     RECT  1096.7 1671.5 1098.82 1683.46 ;
     RECT  1095.74 1695.44 1099.1 1696.06 ;
     RECT  1096.22 1501.4 1099.3 1531.84 ;
     RECT  1080.26 2236.36 1099.94 2379.78 ;
     RECT  1099.1 1691.24 1100.06 1696.06 ;
     RECT  1098.02 893.48 1100.9 893.68 ;
     RECT  1100.54 1555.58 1101.22 1555.78 ;
     RECT  1098.82 1671.5 1101.7 1681.36 ;
     RECT  1095.9 2192.26 1102.34 2198.34 ;
     RECT  1093.5 749 1102.62 806.74 ;
     RECT  1094.66 816.2 1102.62 855.46 ;
     RECT  1095.94 1650.08 1102.66 1650.28 ;
     RECT  1100.06 1691.24 1102.66 1699 ;
     RECT  1102.34 2192.26 1103.1 2194.56 ;
     RECT  1101.98 1425.8 1103.14 1426 ;
     RECT  1098.02 2209.06 1103.3 2212.2 ;
     RECT  1103.1 2186.8 1103.58 2194.56 ;
     RECT  1103.58 2183.44 1103.78 2194.56 ;
     RECT  1103.9 1710.98 1104.38 1711.18 ;
     RECT  1099.94 2238.88 1104.74 2379.78 ;
     RECT  1096.22 1771.04 1104.86 1789.72 ;
     RECT  1104.38 1558.1 1105.06 1558.3 ;
     RECT  1100.06 1823.96 1105.06 1824.16 ;
     RECT  1101.7 1672.34 1105.54 1681.36 ;
     RECT  1104.38 1710.56 1105.82 1711.18 ;
     RECT  1103.78 2183.44 1106.18 2187.42 ;
     RECT  1105.82 1703.42 1107.26 1711.18 ;
     RECT  1107.26 1703.42 1107.46 1713.28 ;
     RECT  1102.66 1691.24 1107.94 1691.44 ;
     RECT  1098.5 874.16 1108.38 881.92 ;
     RECT  1104.86 1770.62 1108.42 1789.72 ;
     RECT  1104.74 2238.88 1108.58 2377.26 ;
     RECT  1099.3 1501.4 1108.7 1521.34 ;
     RECT  1058.5 1810.1 1108.7 1810.3 ;
     RECT  1095.46 1760.12 1108.9 1760.32 ;
     RECT  1108.42 1770.62 1108.9 1782.58 ;
     RECT  1071.26 1877.72 1108.9 1877.92 ;
     RECT  1102.62 749 1109.06 855.46 ;
     RECT  1084.1 2140.18 1109.34 2143.74 ;
     RECT  1108.58 2239.3 1109.54 2377.26 ;
     RECT  1109.34 2140.18 1109.82 2145.84 ;
     RECT  1108.38 873.74 1110.3 881.92 ;
     RECT  1102.46 1583.3 1110.34 1583.5 ;
     RECT  1107.46 1709.72 1111.58 1713.28 ;
     RECT  1110.3 870.38 1112.22 881.92 ;
     RECT  1108.9 1770.62 1112.26 1770.82 ;
     RECT  1108.9 1782.38 1112.26 1782.58 ;
     RECT  1109.54 2239.3 1112.42 2376.84 ;
     RECT  1109.82 2140.18 1113.38 2147.1 ;
     RECT  1103.3 2209.48 1113.66 2212.2 ;
     RECT  1112.06 1797.08 1113.7 1797.28 ;
     RECT  1111.58 1709.72 1114.18 1714.54 ;
     RECT  1112.42 2244.34 1114.34 2376.84 ;
     RECT  1058.5 1886.96 1114.46 1904.38 ;
     RECT  1092.1 1914.26 1114.46 1971.58 ;
     RECT  1088.9 2161.18 1114.62 2161.38 ;
     RECT  1112.22 869.12 1115.1 881.92 ;
     RECT  1114.62 2157.4 1115.1 2161.38 ;
     RECT  1113.98 1747.94 1115.42 1748.14 ;
     RECT  1113.5 1557.26 1115.62 1557.46 ;
     RECT  1106.18 2183.44 1116.06 2183.64 ;
     RECT  1114.18 1714.34 1116.1 1714.54 ;
     RECT  1108.7 1810.1 1116.1 1816.6 ;
     RECT  1115.1 2157.4 1116.54 2167.68 ;
     RECT  1116.06 2183.44 1117.02 2191.62 ;
     RECT  1115.42 1742.9 1117.54 1748.14 ;
     RECT  1113.38 2140.18 1117.98 2145.84 ;
     RECT  1114.46 1886.96 1118.02 1971.58 ;
     RECT  1101.5 1351.04 1118.5 1351.24 ;
     RECT  1116.38 1394.72 1118.5 1394.92 ;
     RECT  1109.06 749 1118.94 805.48 ;
     RECT  1109.06 814.52 1118.94 855.46 ;
     RECT  1111.58 1863.02 1119.26 1863.22 ;
     RECT  1022.66 2391.8 1119.42 2428.96 ;
     RECT  737.86 2439.26 1119.42 2479.36 ;
     RECT  1119.26 1861.76 1120.22 1863.22 ;
     RECT  1116.54 2157.4 1120.86 2173.98 ;
     RECT  1117.02 2183.44 1120.86 2194.56 ;
     RECT  1120.86 2157.4 1121.34 2194.56 ;
     RECT  1120.22 1776.92 1121.38 1777.12 ;
     RECT  1113.98 1642.52 1121.66 1642.72 ;
     RECT  1121.34 2157.4 1121.82 2195.82 ;
     RECT  1113.66 2209.48 1121.82 2213.04 ;
     RECT  1121.66 1424.96 1122.82 1426 ;
     RECT  1114.34 2244.34 1123.26 2376.42 ;
     RECT  1117.98 2138.92 1123.74 2145.84 ;
     RECT  1121.82 2157.4 1123.74 2213.04 ;
     RECT  1120.22 1861.76 1124.26 1866.58 ;
     RECT  1124.06 1699.22 1124.54 1699.42 ;
     RECT  1105.54 1681.16 1125.02 1681.36 ;
     RECT  1124.26 1861.76 1125.22 1861.96 ;
     RECT  1117.02 896.42 1125.66 896.62 ;
     RECT  1124.06 1436.72 1125.7 1436.92 ;
     RECT  1124.54 1738.28 1126.94 1738.48 ;
     RECT  1117.54 1747.94 1126.94 1748.14 ;
     RECT  1121.66 1642.52 1127.42 1649.86 ;
     RECT  1123.26 2242.24 1128.06 2376.42 ;
     RECT  1123.74 2138.92 1129.02 2213.46 ;
     RECT  1126.94 1738.28 1130.78 1748.14 ;
     RECT  1115.1 869.12 1130.94 887.38 ;
     RECT  1125.66 896.42 1130.94 897.46 ;
     RECT  1127.42 1642.52 1130.98 1650.28 ;
     RECT  1124.54 1699.22 1130.98 1699.84 ;
     RECT  1128.06 2235.94 1131.14 2376.42 ;
     RECT  1008.1 1837.82 1131.26 1850.2 ;
     RECT  1128.86 1721.9 1132.9 1722.1 ;
     RECT  1130.78 1738.28 1133.18 1749.4 ;
     RECT  1133.18 1738.28 1133.66 1755.7 ;
     RECT  1130.98 1699.22 1134.34 1699.42 ;
     RECT  1131.14 2239.3 1134.5 2376.42 ;
     RECT  1125.02 1672.76 1134.62 1681.36 ;
     RECT  1127.42 1309.88 1134.82 1310.08 ;
     RECT  1130.98 1642.52 1134.82 1649.86 ;
     RECT  1116.1 1810.1 1135.58 1810.3 ;
     RECT  1134.62 1672.76 1135.78 1689.76 ;
     RECT  1134.5 2269.54 1135.94 2376.42 ;
     RECT  1118.94 749 1137.38 855.46 ;
     RECT  1137.02 1641.68 1137.7 1641.88 ;
     RECT  1135.78 1673.18 1137.7 1689.76 ;
     RECT  1125.02 1823.96 1138.18 1824.16 ;
     RECT  1137.7 1673.18 1138.66 1681.36 ;
     RECT  1130.78 1771.04 1138.66 1771.24 ;
     RECT  1134.5 2239.3 1138.82 2260.5 ;
     RECT  1129.34 1710.56 1139.42 1710.76 ;
     RECT  1133.66 1732.82 1140.1 1755.7 ;
     RECT  1126.46 1787.42 1140.1 1787.62 ;
     RECT  1131.26 1835.3 1140.58 1850.2 ;
     RECT  1140.58 1835.3 1144.42 1842.22 ;
     RECT  1130.94 869.12 1144.58 897.46 ;
     RECT  1139.42 1710.56 1144.9 1714.12 ;
     RECT  1108.7 1499.72 1145.38 1521.34 ;
     RECT  1142.78 1540.46 1145.38 1540.66 ;
     RECT  1137.38 749 1147.46 855.04 ;
     RECT  1147.46 814.52 1147.74 855.04 ;
     RECT  1135.58 1801.7 1148.26 1810.3 ;
     RECT  1144.22 1781.96 1148.54 1782.16 ;
     RECT  1130.78 1456.88 1148.74 1457.08 ;
     RECT  1147.74 814.52 1149.18 855.46 ;
     RECT  1145.38 1499.72 1149.22 1507.9 ;
     RECT  1140.1 1732.82 1149.22 1749.4 ;
     RECT  1146.62 1653.02 1149.5 1653.22 ;
     RECT  1148.54 1777.76 1149.98 1782.16 ;
     RECT  1129.02 2138.92 1150.14 2217.24 ;
     RECT  1144.58 869.12 1150.34 897.04 ;
     RECT  1149.22 1732.82 1150.66 1738.48 ;
     RECT  1148.26 1805.48 1150.94 1810.3 ;
     RECT  1139.9 1820.18 1150.94 1820.38 ;
     RECT  1149.5 1471.16 1151.14 1471.36 ;
     RECT  1144.7 1759.28 1151.14 1759.48 ;
     RECT  1149.18 814.52 1152.06 855.88 ;
     RECT  1150.94 1805.48 1152.1 1820.38 ;
     RECT  1152.06 814.52 1153.02 856.72 ;
     RECT  1150.34 869.12 1153.02 892.42 ;
     RECT  1150.66 1738.28 1153.06 1738.48 ;
     RECT  1149.98 1771.88 1153.54 1782.16 ;
     RECT  1138.82 2252.32 1153.7 2260.5 ;
     RECT  1118.02 1886.96 1154.78 1904.38 ;
     RECT  1118.02 1914.26 1154.78 1971.58 ;
     RECT  1149.5 1649.66 1154.98 1653.22 ;
     RECT  1153.02 814.52 1155.14 892.42 ;
     RECT  1135.94 2271.64 1155.42 2376.42 ;
     RECT  1144.9 1710.56 1155.46 1710.76 ;
     RECT  1153.54 1771.88 1155.46 1777.96 ;
     RECT  1154.98 1653.02 1155.94 1653.22 ;
     RECT  1149.22 1747.94 1155.94 1749.4 ;
     RECT  1152.1 1805.48 1155.94 1812.4 ;
     RECT  1152.38 1663.52 1156.42 1665.4 ;
     RECT  1155.94 1805.48 1156.42 1810.3 ;
     RECT  1155.42 2269.54 1156.58 2376.42 ;
     RECT  1155.46 1777.76 1156.9 1777.96 ;
     RECT  1155.14 869.12 1157.06 892.42 ;
     RECT  1150.14 2138.92 1157.54 2218.08 ;
     RECT  1156.42 1808.42 1158.34 1810.3 ;
     RECT  1157.06 887.18 1158.5 892.42 ;
     RECT  1149.22 1501.4 1159.1 1507.9 ;
     RECT  1145.38 1516.52 1159.1 1521.34 ;
     RECT  1099.3 1531.64 1159.1 1531.84 ;
     RECT  1159.1 1763.06 1159.3 1764.1 ;
     RECT  1147.46 749 1160.22 805.06 ;
     RECT  1156.7 1461.08 1160.26 1461.28 ;
     RECT  1083.94 1985.24 1160.74 2007.7 ;
     RECT  1096.9 1445.96 1161.98 1446.16 ;
     RECT  1159.1 1731.14 1162.46 1731.34 ;
     RECT  1119.42 2391.8 1162.66 2479.36 ;
     RECT  1151.42 1612.7 1162.94 1612.9 ;
     RECT  1162.66 2391.8 1163.62 2464.66 ;
     RECT  1157.06 869.12 1163.78 878.14 ;
     RECT  1159.1 1501.4 1163.9 1521.34 ;
     RECT  1162.46 1731.14 1163.9 1733.44 ;
     RECT  1155.14 814.52 1164.06 858.82 ;
     RECT  1163.78 869.12 1164.06 876.88 ;
     RECT  1164.06 814.52 1164.26 876.88 ;
     RECT  1163.42 1490.9 1164.38 1491.1 ;
     RECT  1163.9 1500.14 1164.38 1521.34 ;
     RECT  1161.98 1445.96 1164.58 1450.78 ;
     RECT  1154.78 1886.96 1164.58 1971.58 ;
     RECT  1162.94 1778.18 1164.86 1778.38 ;
     RECT  1161.02 1657.64 1165.06 1657.84 ;
     RECT  1162.94 1604.72 1165.34 1612.9 ;
     RECT  1160.22 749 1165.5 805.9 ;
     RECT  1164.26 814.52 1165.5 855.88 ;
     RECT  1138.66 1681.16 1166.3 1681.36 ;
     RECT  1155.94 1748.36 1166.3 1749.4 ;
     RECT  1157.54 2138.92 1166.46 2217.24 ;
     RECT  1158.5 888.44 1167.14 892.42 ;
     RECT  1166.3 1673.6 1167.46 1681.36 ;
     RECT  1159.1 1366.16 1168.22 1366.36 ;
     RECT  1166.3 1748.36 1168.22 1751.5 ;
     RECT  1153.7 2252.32 1168.38 2258.82 ;
     RECT  1156.58 2273.32 1168.38 2376.42 ;
     RECT  1163.62 2391.8 1168.42 2459.2 ;
     RECT  1164.86 1778.18 1169.38 1778.8 ;
     RECT  1168.22 1366.16 1170.14 1369.72 ;
     RECT  1164.86 1710.56 1170.14 1710.76 ;
     RECT  1170.14 1710.56 1170.62 1713.28 ;
     RECT  1158.34 1810.1 1170.62 1810.3 ;
     RECT  1170.14 1779.02 1170.82 1779.22 ;
     RECT  1168.38 2252.32 1170.98 2376.42 ;
     RECT  1159.3 1763.06 1171.1 1763.26 ;
     RECT  1170.98 2269.96 1171.46 2376.42 ;
     RECT  1165.5 749 1172.7 855.88 ;
     RECT  1164.26 864.92 1172.7 876.88 ;
     RECT  1168.22 1748.36 1173.22 1752.34 ;
     RECT  1163.9 1729.04 1173.5 1733.44 ;
     RECT  1173.22 1748.36 1173.5 1751.92 ;
     RECT  1170.62 1808.42 1173.7 1810.3 ;
     RECT  1165.5 902.72 1174.34 902.92 ;
     RECT  1166.46 2136.4 1174.34 2217.24 ;
     RECT  1164.38 1490.9 1174.94 1521.34 ;
     RECT  1159.1 1531.64 1174.94 1550.32 ;
     RECT  1051 0 1175 178 ;
     RECT  1172.7 749 1175.1 876.88 ;
     RECT  1167.14 888.44 1175.1 889.9 ;
     RECT  1170.14 1359.02 1175.14 1369.72 ;
     RECT  1174.94 1490.9 1175.14 1550.32 ;
     RECT  1171.46 2269.96 1175.3 2292.84 ;
     RECT  1171.1 1760.96 1175.42 1763.26 ;
     RECT  1160.54 1570.28 1175.9 1570.48 ;
     RECT  1174.34 2194.36 1176.26 2217.24 ;
     RECT  1176.26 2194.36 1176.74 2202.12 ;
     RECT  1175.9 1567.76 1176.86 1570.48 ;
     RECT  1170.62 1702.16 1177.06 1713.28 ;
     RECT  1175.14 1366.16 1177.54 1369.72 ;
     RECT  1176.86 1567.76 1177.54 1571.32 ;
     RECT  1177.06 1713.08 1177.82 1713.28 ;
     RECT  1175.14 1490.9 1178.5 1545.28 ;
     RECT  1178.5 1531.64 1178.98 1545.28 ;
     RECT  1165.34 1596.74 1179.94 1612.9 ;
     RECT  1177.54 1570.28 1180.22 1571.32 ;
     RECT  1162.94 1627.4 1180.42 1627.6 ;
     RECT  1177.82 1713.08 1181.18 1713.7 ;
     RECT  1178.5 1490.9 1181.86 1521.34 ;
     RECT  1179.94 1596.74 1182.34 1604.92 ;
     RECT  1180.22 1570.28 1183.3 1576.78 ;
     RECT  1164.38 1823.96 1183.58 1824.16 ;
     RECT  1173.5 1729.04 1184.74 1751.92 ;
     RECT  1175.1 749 1184.9 889.9 ;
     RECT  1061 3222 1185 3400 ;
     RECT  1184.9 749 1186.82 855.46 ;
     RECT  1183.58 1823.96 1186.94 1827.52 ;
     RECT  1171.1 1782.38 1187.14 1782.58 ;
     RECT  1184.9 864.92 1187.78 889.9 ;
     RECT  1167.46 1676.54 1187.9 1681.36 ;
     RECT  1175.42 1760.96 1188.1 1763.68 ;
     RECT  1181.86 1511.48 1188.58 1521.34 ;
     RECT  1170.98 2252.32 1189.22 2258.82 ;
     RECT  1175.3 2273.32 1189.22 2292.84 ;
     RECT  1187.9 1676.12 1189.82 1681.36 ;
     RECT  1186.94 1823.96 1190.5 1827.94 ;
     RECT  1184.74 1740.38 1190.78 1751.92 ;
     RECT  1189.82 1670.24 1190.98 1681.36 ;
     RECT  1181.18 1713.08 1191.26 1714.12 ;
     RECT  1184.74 1729.04 1191.26 1729.24 ;
     RECT  1190.98 1676.12 1191.46 1681.36 ;
     RECT  1188.86 1377.08 1191.94 1377.28 ;
     RECT  1187.78 864.92 1192.1 878.56 ;
     RECT  1189.22 2273.32 1192.1 2292.42 ;
     RECT  1188.06 896.42 1192.58 896.62 ;
     RECT  1186.82 749 1193.06 855.04 ;
     RECT  1193.06 749 1193.54 847.9 ;
     RECT  1193.66 1698.8 1194.34 1699 ;
     RECT  1191.26 1713.08 1194.82 1729.24 ;
     RECT  1194.82 1713.08 1195.3 1721.68 ;
     RECT  1164.58 1445.96 1196.06 1446.16 ;
     RECT  1195.1 1419.5 1196.26 1419.7 ;
     RECT  1190.78 1740.38 1196.26 1752.76 ;
     RECT  1188.58 1512.32 1196.74 1521.34 ;
     RECT  1192.1 2273.74 1197.66 2292.42 ;
     RECT  1171.46 2304.82 1197.66 2376.42 ;
     RECT  1196.06 1445.96 1197.7 1447 ;
     RECT  1196.54 1700.9 1197.7 1701.1 ;
     RECT  1194.14 1778.6 1198.18 1778.8 ;
     RECT  1196.26 1740.38 1199.42 1751.5 ;
     RECT  1197.7 1446.8 1200.58 1447 ;
     RECT  1195.58 1456.88 1200.58 1457.08 ;
     RECT  1197.66 2273.74 1201.22 2376.42 ;
     RECT  1193.54 814.52 1201.5 847.9 ;
     RECT  1195.3 1721.48 1201.54 1721.68 ;
     RECT  1192.1 864.92 1201.7 876.88 ;
     RECT  1193.54 749 1201.98 805.48 ;
     RECT  1181.86 1490.9 1202.5 1502.44 ;
     RECT  1199.42 1739.96 1202.98 1751.5 ;
     RECT  1178.98 1531.64 1203.94 1538.14 ;
     RECT  1182.34 1596.74 1203.94 1596.94 ;
     RECT  1177.54 1366.16 1205.38 1366.36 ;
     RECT  1202.5 1500.14 1205.38 1501.6 ;
     RECT  1193.66 1547.6 1205.38 1547.8 ;
     RECT  1202.98 1747.94 1205.38 1748.56 ;
     RECT  1189.22 2252.32 1205.82 2256.3 ;
     RECT  1201.22 2273.74 1206.5 2298.72 ;
     RECT  1206.5 2273.74 1206.98 2292.42 ;
     RECT  1187.42 1430.84 1208.26 1431.04 ;
     RECT  1202.5 1490.9 1209.22 1491.1 ;
     RECT  1188.1 1763.48 1209.5 1763.68 ;
     RECT  1209.5 1763.48 1209.7 1764.1 ;
     RECT  1201.7 869.12 1210.14 876.88 ;
     RECT  1183.3 1576.58 1210.66 1576.78 ;
     RECT  1210.14 866.6 1213.02 876.88 ;
     RECT  1201.98 741.44 1214.46 805.48 ;
     RECT  1201.5 814.52 1214.46 850.84 ;
     RECT  1213.02 866.18 1214.46 876.88 ;
     RECT  1211.9 1597.16 1214.78 1597.36 ;
     RECT  1196.74 1516.52 1214.98 1521.34 ;
     RECT  1214.78 1596.32 1215.94 1597.36 ;
     RECT  1214.46 741.44 1216.1 850.84 ;
     RECT  1214.46 865.76 1216.1 876.88 ;
     RECT  1209.5 1479.56 1216.42 1479.76 ;
     RECT  1216.1 866.18 1216.58 876.88 ;
     RECT  1144.42 1837.82 1217.18 1842.22 ;
     RECT  1210.62 895.58 1217.54 895.78 ;
     RECT  1176.74 2194.36 1218.3 2195.82 ;
     RECT  1218.14 1416.56 1219.58 1416.76 ;
     RECT  1219.58 1415.72 1219.78 1416.76 ;
     RECT  1201.22 2308.18 1220.06 2376.42 ;
     RECT  1220.54 1389.26 1221.02 1389.46 ;
     RECT  1220.06 1420.76 1221.7 1420.96 ;
     RECT  1221.02 1389.26 1222.18 1389.88 ;
     RECT  1215.94 1597.16 1222.18 1597.36 ;
     RECT  1222.18 1389.26 1223.14 1389.46 ;
     RECT  1209.5 1468.22 1223.62 1468.42 ;
     RECT  1220.54 1736.6 1223.62 1736.8 ;
     RECT  1191.46 1681.16 1224.86 1681.36 ;
     RECT  1224.86 1665.62 1225.34 1665.82 ;
     RECT  1222.94 1421.6 1225.54 1421.8 ;
     RECT  1216.58 869.12 1225.98 876.88 ;
     RECT  1217.18 1835.3 1226.02 1842.22 ;
     RECT  1220.06 2301.08 1227.26 2376.42 ;
     RECT  1223.9 1379.18 1227.94 1379.38 ;
     RECT  1216.1 749 1228.38 850.84 ;
     RECT  1224.86 1676.12 1228.42 1681.36 ;
     RECT  1227.26 2300.66 1229.06 2376.42 ;
     RECT  1214.98 1521.14 1231.1 1521.34 ;
     RECT  1225.34 1660.58 1236.1 1665.82 ;
     RECT  1229.06 2319.1 1236.26 2376.42 ;
     RECT  1205.38 1747.94 1237.34 1748.14 ;
     RECT  1228.38 749 1238.18 855.04 ;
     RECT  1220.06 1487.12 1240.42 1487.32 ;
     RECT  1231.1 1517.78 1240.42 1521.34 ;
     RECT  1237.34 1740.38 1240.9 1748.14 ;
     RECT  1222.46 1725.68 1241.18 1725.88 ;
     RECT  1240.9 1740.8 1241.18 1748.14 ;
     RECT  1241.18 1721.06 1242.62 1725.88 ;
     RECT  1228.42 1681.16 1243.1 1681.36 ;
     RECT  1176.26 2212 1243.46 2217.24 ;
     RECT  1175 -70 1245 178 ;
     RECT  1242.62 1720.64 1246.18 1725.88 ;
     RECT  1243.1 1681.16 1246.46 1683.88 ;
     RECT  1246.46 1680.32 1248.1 1683.88 ;
     RECT  1245.5 1706.78 1248.1 1706.98 ;
     RECT  1236.1 1665.62 1248.58 1665.82 ;
     RECT  1248.1 1680.32 1253.38 1681.36 ;
     RECT  1205.82 2252.32 1254.5 2262.6 ;
     RECT  1238.18 749 1254.78 852.1 ;
     RECT  1185 3222 1255 3470 ;
     RECT  1246.18 1721.06 1255.3 1725.88 ;
     RECT  1249.82 1561.46 1255.78 1561.66 ;
     RECT  1255.3 1725.68 1255.78 1725.88 ;
     RECT  1241.18 1740.8 1255.78 1756.12 ;
     RECT  1254.78 749 1256.9 855.46 ;
     RECT  1256.9 804.86 1257.66 855.46 ;
     RECT  1255.78 1747.94 1258.66 1756.12 ;
     RECT  1254.5 2252.32 1263.26 2256.3 ;
     RECT  1256.06 2264.96 1263.26 2265.16 ;
     RECT  1235.42 1425.8 1263.46 1426 ;
     RECT  1263.26 1864.7 1263.46 1865.32 ;
     RECT  1257.66 804.86 1263.62 856.3 ;
     RECT  1263.62 804.86 1264.1 848.74 ;
     RECT  1160.74 1990.7 1266.14 2007.7 ;
     RECT  1260.54 896.42 1267.26 896.62 ;
     RECT  1252.22 1476.2 1267.3 1476.4 ;
     RECT  1267.26 896.42 1267.46 897.04 ;
     RECT  1253.38 1681.16 1268.06 1681.36 ;
     RECT  1265.66 1721.48 1268.26 1721.68 ;
     RECT  1263.46 1865.12 1268.74 1865.32 ;
     RECT  1225.98 866.18 1270.62 876.88 ;
     RECT  1190.5 1823.96 1271.62 1824.16 ;
     RECT  1164.58 1886.96 1272.38 1904.38 ;
     RECT  1226.02 1837.82 1273.54 1842.22 ;
     RECT  1272.38 1886.54 1276.42 1904.38 ;
     RECT  1264.1 833.42 1278.98 848.74 ;
     RECT  1256.9 749 1279.94 793.72 ;
     RECT  1264.22 1698.8 1280.06 1699 ;
     RECT  1276.22 1771.46 1280.54 1771.66 ;
     RECT  1273.54 1837.82 1280.54 1839.28 ;
     RECT  1280.06 1698.8 1282.94 1706.14 ;
     RECT  1266.14 1986.08 1282.94 2007.7 ;
     RECT  1282.94 1698.8 1283.14 1710.76 ;
     RECT  1280.54 1770.62 1284.1 1771.66 ;
     RECT  1281.66 896 1284.26 896.2 ;
     RECT  957.7 2508.98 1284.58 2509.18 ;
     RECT  1280.54 1831.52 1285.82 1839.28 ;
     RECT  1268.06 1672.76 1286.5 1681.36 ;
     RECT  1284.1 1770.62 1286.5 1771.24 ;
     RECT  1283.14 1698.8 1286.98 1699 ;
     RECT  1286.5 1770.62 1286.98 1770.82 ;
     RECT  1285.82 1831.52 1287.26 1845.58 ;
     RECT  1032.86 918.02 1287.94 925.36 ;
     RECT  1270.62 866.18 1288.58 878.14 ;
     RECT  1168.42 2391.8 1288.7 2433.96 ;
     RECT  1288.7 2391.8 1288.9 2434.42 ;
     RECT  1288.58 869.12 1289.06 878.14 ;
     RECT  1283.14 1710.56 1290.34 1710.76 ;
     RECT  1174.34 2136.4 1290.5 2184.48 ;
     RECT  1218.3 2194.36 1290.5 2197.08 ;
     RECT  1243.46 2212 1290.5 2212.2 ;
     RECT  1138.82 2239.3 1290.5 2242.44 ;
     RECT  1263.26 2252.32 1290.5 2265.16 ;
     RECT  1206.98 2273.74 1290.5 2291.58 ;
     RECT  1236.26 2319.1 1290.5 2334.42 ;
     RECT  1290.5 2319.1 1290.98 2319.72 ;
     RECT  1236.26 2345.56 1292.7 2376.42 ;
     RECT  1292.7 2344.3 1292.9 2376.42 ;
     RECT  1284.86 1730.3 1293.98 1730.5 ;
     RECT  1162.66 2476.64 1293.98 2479.36 ;
     RECT  1288.7 3049.1 1293.98 3049.3 ;
     RECT  1287.74 3063.38 1293.98 3063.58 ;
     RECT  1287.26 1831.52 1294.46 1847.26 ;
     RECT  1290.5 2142.74 1294.82 2157.6 ;
     RECT  1279.94 751.94 1295.1 793.72 ;
     RECT  1264.1 804.86 1295.1 822.28 ;
     RECT  1290.5 2273.74 1295.3 2273.94 ;
     RECT  1292.9 2344.3 1295.3 2360.04 ;
     RECT  1293.98 3049.1 1295.42 3063.58 ;
     RECT  1293.98 1729.46 1295.62 1730.5 ;
     RECT  1229.06 2300.66 1295.78 2308.38 ;
     RECT  1295.42 3049.1 1295.9 3066.94 ;
     RECT  1290.5 2239.3 1296.26 2239.5 ;
     RECT  1290.5 2329.6 1296.26 2334.42 ;
     RECT  1295.3 2359.84 1296.26 2360.04 ;
     RECT  1290.98 2319.1 1296.74 2319.3 ;
     RECT  1293.98 1710.14 1297.06 1710.34 ;
     RECT  1294.46 1824.38 1297.06 1847.26 ;
     RECT  1296.26 2334.22 1297.22 2334.42 ;
     RECT  1295.62 1730.3 1298.02 1730.5 ;
     RECT  1290.5 2255.68 1298.18 2265.16 ;
     RECT  1294.82 2154.92 1298.66 2157.6 ;
     RECT  1276.42 1886.96 1298.78 1904.38 ;
     RECT  1297.82 2130.98 1298.78 2131.18 ;
     RECT  1296.38 2897.9 1298.78 2898.1 ;
     RECT  1295.3 2344.3 1298.94 2346.18 ;
     RECT  1282.94 1982.72 1298.98 2007.7 ;
     RECT  1298.18 2256.1 1299.14 2265.16 ;
     RECT  1298.94 2343.88 1299.14 2346.18 ;
     RECT  1134.62 2105.78 1299.26 2105.98 ;
     RECT  1168.42 2443.88 1299.26 2459.2 ;
     RECT  1295.9 3049.1 1299.26 3074.08 ;
     RECT  1292.06 2116.7 1299.46 2116.9 ;
     RECT  1298.3 1861.34 1300.22 1861.54 ;
     RECT  967.94 2044.46 1300.22 2050.12 ;
     RECT  1288.9 2428.76 1300.42 2434.42 ;
     RECT  1299.26 2443.88 1300.42 2459.62 ;
     RECT  1295.1 751.94 1300.58 822.28 ;
     RECT  1299.74 2919.32 1300.68 2919.52 ;
     RECT  1299.26 3040.7 1300.815 3074.08 ;
     RECT  1298.3 1705.52 1300.9 1707.4 ;
     RECT  1300.22 1861.34 1301.18 1861.96 ;
     RECT  1277.18 1872.26 1301.18 1872.46 ;
     RECT  1298.78 1881.5 1301.18 1904.38 ;
     RECT  1298.78 2130.14 1301.18 2131.18 ;
     RECT  1294.82 2142.74 1301.18 2142.94 ;
     RECT  1297.06 1824.38 1301.38 1839.28 ;
     RECT  1301.18 1861.34 1301.38 1862.8 ;
     RECT  1299.26 2105.78 1301.38 2106.4 ;
     RECT  1301.18 2130.14 1301.38 2142.94 ;
     RECT  1298.66 2154.92 1301.38 2155.12 ;
     RECT  1300.42 2428.76 1301.38 2434 ;
     RECT  1300.58 751.94 1301.54 793.72 ;
     RECT  1301.38 2130.14 1301.66 2136.22 ;
     RECT  1290.5 2167.48 1301.66 2167.68 ;
     RECT  1299.14 2261.6 1301.66 2265.16 ;
     RECT  1290.5 2285.5 1301.66 2291.58 ;
     RECT  1292.9 2370.38 1301.66 2376.42 ;
     RECT  1288.9 2391.8 1301.66 2416.36 ;
     RECT  1293.98 2476.64 1301.66 2487.76 ;
     RECT  1301.66 2124.26 1301.86 2136.22 ;
     RECT  1286.5 1675.28 1302.14 1681.36 ;
     RECT  731.9 2022.62 1302.535 2027.44 ;
     RECT  1300.22 2041.1 1302.535 2050.12 ;
     RECT  1301.66 2282.6 1302.535 2291.58 ;
     RECT  1295.78 2300.66 1302.535 2301.28 ;
     RECT  1302.14 1667.72 1302.62 1681.36 ;
     RECT  1300.68 2919.32 1303.28 2922.12 ;
     RECT  1300.68 3181.08 1303.28 3183.08 ;
     RECT  1300.815 2942.2 1303.415 2947.68 ;
     RECT  1300.815 3010.6 1303.415 3016.08 ;
     RECT  1300.815 3040.7 1303.415 3082.2 ;
     RECT  1300.815 3145.12 1303.415 3150.6 ;
     RECT  1301.18 1872.26 1303.58 1904.38 ;
     RECT  1299.26 1778.6 1304.26 1778.8 ;
     RECT  1301.38 1861.76 1304.26 1862.8 ;
     RECT  1302.535 2022.62 1304.265 2050.12 ;
     RECT  1302.535 2282.6 1304.265 2301.28 ;
     RECT  1302.535 2559.16 1304.265 2564.64 ;
     RECT  1298.98 1990.7 1304.4 2007.7 ;
     RECT  698.5 2580.72 1304.4 2585.32 ;
     RECT  1302.62 1665.2 1304.74 1681.36 ;
     RECT  1299.74 1736.6 1304.74 1736.8 ;
     RECT  1164.58 1914.26 1305.02 1971.58 ;
     RECT  1304.265 2022.62 1305.135 2027.44 ;
     RECT  1304.74 1665.2 1305.22 1665.4 ;
     RECT  1301.54 751.94 1306.14 774.82 ;
     RECT  1305.135 2016.52 1306.865 2027.44 ;
     RECT  1305.135 2547.76 1306.865 2553.24 ;
     RECT  1304.4 2583.32 1307 2585.32 ;
     RECT  1300.9 1707.2 1307.14 1707.4 ;
     RECT  1305.02 1914.26 1307.14 1972 ;
     RECT  1305.5 1722.32 1307.42 1722.52 ;
     RECT  1304.265 2041.1 1307.62 2050.12 ;
     RECT  1301.66 2261.6 1307.62 2271.88 ;
     RECT  1303.28 2919.32 1307.68 2924.72 ;
     RECT  1303.415 2942.2 1307.68 2959.08 ;
     RECT  1303.415 3010.6 1307.68 3027.48 ;
     RECT  1303.415 3040.7 1307.68 3093.6 ;
     RECT  1303.415 3145.12 1307.68 3162 ;
     RECT  1303.28 3178.48 1307.68 3183.08 ;
     RECT  1307.42 1721.06 1308.1 1722.52 ;
     RECT  1305.98 2217.5 1308.58 2217.7 ;
     RECT  1305.02 2338.88 1309.06 2339.08 ;
     RECT  1278.98 833.42 1309.7 847.48 ;
     RECT  1306.14 745.64 1310.18 774.82 ;
     RECT  1173.7 1810.1 1310.3 1810.3 ;
     RECT  1301.38 2105.78 1310.3 2105.98 ;
     RECT  1307.62 2261.6 1310.3 2265.16 ;
     RECT  1307.1 733.88 1310.46 734.08 ;
     RECT  1309.34 1662.68 1310.5 1662.88 ;
     RECT  1301.38 1824.38 1310.5 1826.68 ;
     RECT  1303.58 1871.42 1310.5 1904.38 ;
     RECT  1308.1 1721.06 1310.78 1721.26 ;
     RECT  1301.38 1837.82 1310.78 1839.28 ;
     RECT  1310.5 1871.42 1310.78 1877.08 ;
     RECT  1304.265 2282.6 1310.78 2289.94 ;
     RECT  1310.78 1864.28 1310.98 1877.08 ;
     RECT  1300.58 802.34 1311.62 822.28 ;
     RECT  1310.3 2255.72 1311.74 2265.16 ;
     RECT  1301.66 2321.24 1311.74 2325.22 ;
     RECT  1310.78 2280.92 1311.94 2289.94 ;
     RECT  1311.74 2250.68 1312.22 2265.16 ;
     RECT  1304.4 1990.7 1313.66 1996.8 ;
     RECT  1304.4 2005.4 1313.66 2007.7 ;
     RECT  1301.86 2124.26 1313.66 2135.38 ;
     RECT  1312.22 2248.58 1313.86 2265.16 ;
     RECT  1310.3 1805.9 1314.14 1810.3 ;
     RECT  1310.5 1826.48 1314.62 1826.68 ;
     RECT  1310.78 1837.82 1314.62 1846.84 ;
     RECT  1301.66 2164.16 1315.1 2179.48 ;
     RECT  1310.18 751.94 1315.26 774.82 ;
     RECT  1313.66 2124.26 1316.06 2141.68 ;
     RECT  1310.98 1864.28 1316.26 1876.66 ;
     RECT  1310.46 733.88 1316.42 737.86 ;
     RECT  1311.62 802.34 1317.38 819.76 ;
     RECT  1316.06 2124.26 1317.98 2142.1 ;
     RECT  1315.1 2156.6 1317.98 2179.48 ;
     RECT  1313.66 1990.7 1318.18 2007.7 ;
     RECT  1310.78 1720.64 1318.46 1721.26 ;
     RECT  1307.14 1914.26 1318.46 1971.58 ;
     RECT  1301.54 789.32 1319.58 793.72 ;
     RECT  1317.38 802.34 1319.58 817.24 ;
     RECT  1318.46 1720.64 1319.62 1728.4 ;
     RECT  1313.86 2250.68 1319.62 2265.16 ;
     RECT  1316.06 1600.52 1320.1 1600.72 ;
     RECT  1313.66 1767.68 1320.86 1767.88 ;
     RECT  1311.94 2282.6 1321.06 2289.94 ;
     RECT  1317.98 2124.26 1321.34 2179.48 ;
     RECT  1321.34 2124.26 1321.54 2179.9 ;
     RECT  1301.66 2367.86 1321.54 2416.36 ;
     RECT  1314.14 1805.9 1322.3 1810.72 ;
     RECT  1301.38 2429.18 1322.3 2434 ;
     RECT  1300.42 2443.88 1322.3 2459.2 ;
     RECT  1319.62 1728.2 1322.78 1728.4 ;
     RECT  1318.46 1914.26 1322.98 1972.84 ;
     RECT  1321.54 2124.26 1323.74 2124.46 ;
     RECT  1319.58 888.02 1323.9 888.22 ;
     RECT  1311.74 2321.24 1324.42 2326.48 ;
     RECT  1011.26 2091.5 1324.7 2091.7 ;
     RECT  1310.3 2101.16 1324.7 2105.98 ;
     RECT  1323.74 2118.8 1324.7 2124.46 ;
     RECT  1324.7 2118.38 1324.9 2124.46 ;
     RECT  1324.7 2091.5 1325.38 2105.98 ;
     RECT  1316.42 737.66 1325.54 737.86 ;
     RECT  1314.62 1826.48 1325.86 1846.84 ;
     RECT  1321.54 2392.22 1326.34 2416.36 ;
     RECT  1258.66 1747.94 1326.62 1748.14 ;
     RECT  1326.62 1747.94 1327.58 1756.12 ;
     RECT  1322.78 1728.2 1328.06 1730.5 ;
     RECT  1325.86 1826.48 1328.06 1839.28 ;
     RECT  1304.265 2300.66 1328.06 2301.28 ;
     RECT  1325.18 1650.08 1328.26 1650.28 ;
     RECT  1322.3 2429.18 1328.26 2459.2 ;
     RECT  1315.26 751.94 1328.42 779.86 ;
     RECT  1328.06 1728.2 1328.54 1735.12 ;
     RECT  1321.34 1793.3 1328.54 1793.5 ;
     RECT  1321.54 2367.86 1328.54 2383.6 ;
     RECT  1319.62 2255.72 1328.74 2265.16 ;
     RECT  1328.06 2300.66 1328.74 2307.58 ;
     RECT  1319.58 789.32 1328.9 817.24 ;
     RECT  1328.74 2255.72 1329.7 2262.64 ;
     RECT  1300.7 2077.22 1329.98 2077.42 ;
     RECT  1328.06 1825.22 1330.46 1839.28 ;
     RECT  1328.74 2303.18 1330.66 2307.58 ;
     RECT  1321.54 2133.5 1330.94 2142.1 ;
     RECT  1316.26 1865.12 1331.62 1876.66 ;
     RECT  1328.54 2361.98 1331.62 2383.6 ;
     RECT  1331.42 1698.8 1331.9 1699 ;
     RECT  1330.94 2133.08 1331.9 2142.1 ;
     RECT  1323.9 888.02 1332.06 894.1 ;
     RECT  1318.18 1990.7 1332.1 1993.42 ;
     RECT  1318.18 2005.4 1333.34 2007.7 ;
     RECT  1324.9 2122.16 1333.34 2124.46 ;
     RECT  1328.54 1721.48 1333.54 1735.12 ;
     RECT  1321.54 2153.66 1333.54 2179.9 ;
     RECT  1326.34 2392.64 1334.02 2416.36 ;
     RECT  1332.06 888.02 1334.18 900.82 ;
     RECT  1334.18 888.02 1334.66 888.22 ;
     RECT  1321.06 2282.6 1335.46 2288.68 ;
     RECT  1333.34 2119.22 1335.94 2124.46 ;
     RECT  1334.18 896.84 1336.1 900.82 ;
     RECT  1331.9 1698.8 1336.22 1703.2 ;
     RECT  1306.865 2022.62 1336.22 2027.44 ;
     RECT  1307.62 2041.1 1336.22 2041.3 ;
     RECT  1333.34 2005.4 1336.9 2008.96 ;
     RECT  1336.1 896.84 1338.02 897.04 ;
     RECT  1294.46 1566.92 1338.14 1567.12 ;
     RECT  1337.66 1665.62 1338.14 1665.82 ;
     RECT  1331.62 1865.12 1338.34 1872.46 ;
     RECT  1329.98 2077.22 1339.1 2080.78 ;
     RECT  1325.38 2091.5 1339.1 2091.7 ;
     RECT  1331.9 2133.08 1339.1 2144.2 ;
     RECT  1333.54 2153.66 1339.1 2179.48 ;
     RECT  1287.94 918.02 1339.78 918.22 ;
     RECT  1334.3 1634.54 1339.78 1634.74 ;
     RECT  1339.1 2133.08 1339.78 2179.48 ;
     RECT  1325.66 1592.96 1340.06 1593.16 ;
     RECT  1339.78 2133.5 1340.74 2179.48 ;
     RECT  1329.7 2262.44 1341.22 2262.64 ;
     RECT  1325.38 2101.16 1341.5 2105.98 ;
     RECT  1335.94 2119.22 1341.5 2122.36 ;
     RECT  1289.06 869.12 1341.86 876.88 ;
     RECT  1304.74 1681.16 1341.98 1681.36 ;
     RECT  1336.22 1695.44 1342.18 1703.2 ;
     RECT  1330.66 2303.18 1342.18 2303.38 ;
     RECT  1341.86 869.12 1342.34 869.32 ;
     RECT  1328.54 1785.74 1342.46 1793.5 ;
     RECT  1338.14 1664.78 1342.66 1665.82 ;
     RECT  1320.86 1767.68 1342.94 1773.76 ;
     RECT  1322.3 1805.9 1343.14 1812.4 ;
     RECT  1324.42 2321.24 1343.14 2325.22 ;
     RECT  1339.58 2065.46 1343.62 2065.66 ;
     RECT  1340.74 2133.92 1343.62 2179.48 ;
     RECT  1328.9 804.86 1343.78 817.24 ;
     RECT  1343.14 1808.42 1343.9 1812.4 ;
     RECT  1328.9 789.32 1344.26 793.72 ;
     RECT  1301.66 2189.36 1344.38 2189.56 ;
     RECT  1301.66 2202.38 1344.38 2202.58 ;
     RECT  1301.66 2468.66 1344.86 2487.76 ;
     RECT  1335.26 2214.56 1345.06 2214.76 ;
     RECT  1341.5 2101.16 1345.54 2122.36 ;
     RECT  1340.06 1592.54 1345.82 1593.16 ;
     RECT  1327.58 1744.16 1345.82 1756.12 ;
     RECT  1345.82 1739.96 1346.02 1756.12 ;
     RECT  1345.54 2120.9 1346.02 2122.36 ;
     RECT  1338.14 1566.92 1346.98 1574.68 ;
     RECT  1335.46 2288.48 1347.46 2288.68 ;
     RECT  1342.66 1665.62 1347.94 1665.82 ;
     RECT  1338.34 1865.54 1348.22 1872.46 ;
     RECT  1343.62 2133.92 1348.42 2142.1 ;
     RECT  1343.62 2152.4 1348.42 2179.48 ;
     RECT  1333.54 1721.48 1349.18 1730.5 ;
     RECT  1341.98 1674.86 1349.66 1681.36 ;
     RECT  1344.38 2189.36 1349.66 2202.58 ;
     RECT  1344.86 2468.66 1349.86 2494.9 ;
     RECT  1342.94 1767.26 1350.14 1773.76 ;
     RECT  1342.46 1783.22 1350.14 1793.5 ;
     RECT  1348.42 2156.18 1350.14 2179.48 ;
     RECT  1349.18 1718.12 1350.34 1730.5 ;
     RECT  1331.62 2367.86 1350.34 2383.6 ;
     RECT  1348.22 1865.12 1350.62 1872.46 ;
     RECT  1336.7 1645.88 1350.82 1646.08 ;
     RECT  1346.02 1739.96 1350.82 1748.14 ;
     RECT  1350.34 2370.38 1350.82 2383.6 ;
     RECT  1350.82 2375.42 1351.3 2383.6 ;
     RECT  1345.34 1604.72 1351.78 1604.92 ;
     RECT  1350.14 2156.18 1352.06 2180.74 ;
     RECT  1349.66 2189.36 1352.06 2208.46 ;
     RECT  1345.82 1589.6 1352.26 1593.16 ;
     RECT  1330.46 1823.96 1352.74 1839.28 ;
     RECT  1350.34 1718.12 1353.22 1728.4 ;
     RECT  1350.82 1744.16 1353.22 1748.14 ;
     RECT  1339.1 2077.22 1353.7 2091.7 ;
     RECT  1353.22 1718.12 1354.66 1718.32 ;
     RECT  1353.22 1728.2 1355.14 1728.4 ;
     RECT  1345.54 2101.16 1355.62 2112.28 ;
     RECT  1328.42 751.94 1355.78 774.82 ;
     RECT  1348.42 2133.92 1355.9 2138.32 ;
     RECT  1352.06 2156.18 1355.9 2208.46 ;
     RECT  1355.9 2156.18 1356.1 2210.14 ;
     RECT  1355.78 757.82 1356.74 774.82 ;
     RECT  1344.38 2303.6 1357.06 2303.8 ;
     RECT  1356.74 757.82 1357.22 766.84 ;
     RECT  1356.1 2164.16 1357.82 2210.14 ;
     RECT  1345.34 1627.4 1358.02 1627.6 ;
     RECT  1355.62 2101.16 1358.02 2105.98 ;
     RECT  1342.18 1695.44 1358.98 1695.64 ;
     RECT  1332.1 1990.7 1359.26 1990.9 ;
     RECT  1334.02 2395.58 1359.46 2416.36 ;
     RECT  1350.62 1865.12 1359.94 1877.92 ;
     RECT  1309.7 833.42 1360.1 847.06 ;
     RECT  1352.26 1592.96 1360.42 1593.16 ;
     RECT  1355.9 2130.98 1360.42 2138.32 ;
     RECT  1353.02 2060.84 1360.7 2061.04 ;
     RECT  1353.7 2077.22 1360.7 2083.72 ;
     RECT  1346.02 2120.9 1360.7 2121.1 ;
     RECT  1349.66 1668.56 1360.9 1681.36 ;
     RECT  1359.94 1865.96 1360.9 1877.92 ;
     RECT  1359.46 2395.58 1360.9 2398.72 ;
     RECT  1357.22 758.66 1361.06 766.84 ;
     RECT  1360.7 2060.84 1361.38 2083.72 ;
     RECT  1360.7 2115.02 1361.86 2121.1 ;
     RECT  1361.66 2149.88 1362.62 2150.08 ;
     RECT  1322.98 1914.26 1363.1 1971.58 ;
     RECT  1359.26 1986.08 1363.1 1990.9 ;
     RECT  1362.14 2232.2 1363.58 2232.4 ;
     RECT  1361.18 1714.34 1363.78 1714.96 ;
     RECT  1343.9 1808.42 1364.06 1812.82 ;
     RECT  1351.3 2375.42 1364.26 2378.14 ;
     RECT  1363.78 1714.76 1364.74 1714.96 ;
     RECT  1361.86 2120.9 1365.5 2121.1 ;
     RECT  1360.42 2130.98 1365.5 2136.22 ;
     RECT  1361.66 1667.72 1365.7 1667.92 ;
     RECT  1361.38 2069.24 1367.42 2083.72 ;
     RECT  1352.74 1825.22 1367.9 1839.28 ;
     RECT  1336.9 2005.4 1368.38 2007.7 ;
     RECT  1367.42 2069.24 1368.86 2084.98 ;
     RECT  1245 0 1369 178 ;
     RECT  1367.9 1825.22 1369.34 1841.8 ;
     RECT  1360.9 1681.16 1370.3 1681.36 ;
     RECT  1357.82 2164.16 1370.3 2213.5 ;
     RECT  1350.14 1767.26 1371.26 1793.5 ;
     RECT  1362.62 2148.62 1371.26 2150.08 ;
     RECT  1370.3 2159.12 1371.26 2213.5 ;
     RECT  1328.26 2433.8 1371.94 2459.2 ;
     RECT  1364.06 1808.42 1372.22 1816.6 ;
     RECT  1369.82 1604.3 1372.42 1604.5 ;
     RECT  1343.14 2325.02 1372.42 2325.22 ;
     RECT  1368.38 1585.82 1373.66 1586.02 ;
     RECT  1365.5 2120.9 1373.66 2136.22 ;
     RECT  1373.66 1585.82 1373.86 1589.38 ;
     RECT  1370.3 1680.32 1374.14 1681.36 ;
     RECT  1373.18 1718.12 1374.14 1718.32 ;
     RECT  1358.02 2105.78 1374.14 2105.98 ;
     RECT  1373.66 2118.38 1374.14 2136.22 ;
     RECT  1371.26 2148.62 1374.14 2213.5 ;
     RECT  1374.14 1717.28 1375.1 1718.32 ;
     RECT  1360.9 1869.32 1375.1 1877.08 ;
     RECT  1310.5 1886.96 1375.1 1904.38 ;
     RECT  1374.14 2102 1375.1 2105.98 ;
     RECT  1363.58 2224.64 1375.1 2232.4 ;
     RECT  1375.1 2224.64 1375.58 2233.24 ;
     RECT  1375.1 2102 1376.06 2109.76 ;
     RECT  1353.22 1747.94 1376.26 1748.14 ;
     RECT  1375.58 2224.64 1376.54 2236.18 ;
     RECT  1374.14 1680.32 1376.74 1683.88 ;
     RECT  1374.14 2118.38 1377.02 2213.5 ;
     RECT  1376.54 2224.22 1377.02 2236.18 ;
     RECT  1375.1 1861.34 1377.22 1904.38 ;
     RECT  1376.06 2099.48 1377.98 2109.76 ;
     RECT  1377.02 2118.38 1377.98 2236.18 ;
     RECT  1375.1 1717.28 1378.18 1719.16 ;
     RECT  1364.26 2377.94 1378.66 2378.14 ;
     RECT  1255 3222 1379 3400 ;
     RECT  1377.22 1861.34 1380.58 1877.08 ;
     RECT  1368.86 2069.24 1381.34 2088.76 ;
     RECT  1377.98 2099.48 1381.54 2236.18 ;
     RECT  1376.74 1680.32 1382.02 1683.04 ;
     RECT  1381.54 2130.14 1382.98 2236.18 ;
     RECT  1368.38 2005.4 1383.26 2013.16 ;
     RECT  1381.34 2069.24 1383.26 2089.6 ;
     RECT  1381.54 2099.48 1383.26 2121.1 ;
     RECT  1378.18 1717.28 1383.94 1717.48 ;
     RECT  1307.62 2049.92 1384.9 2050.12 ;
     RECT  1382.02 1680.32 1385.38 1681.36 ;
     RECT  1372.22 1805.06 1386.14 1816.6 ;
     RECT  1369.34 1825.22 1386.14 1850.2 ;
     RECT  1373.86 1589.18 1386.62 1589.38 ;
     RECT  1383.26 2004.98 1387.58 2013.16 ;
     RECT  1386.62 1612.28 1388.54 1612.48 ;
     RECT  1361.06 764.12 1388.9 766.84 ;
     RECT  1344.26 789.32 1388.9 789.52 ;
     RECT  1343.78 812 1388.9 817.24 ;
     RECT  1360.1 835.1 1388.9 847.06 ;
     RECT  1386.62 1585.4 1389.22 1589.38 ;
     RECT  1389.22 1585.4 1389.7 1585.6 ;
     RECT  1388.54 1610.6 1389.7 1612.48 ;
     RECT  1363.1 1914.26 1389.98 1990.9 ;
     RECT  1387.58 2004.98 1389.98 2013.58 ;
     RECT  1382.98 2152.82 1389.98 2236.18 ;
     RECT  1297.34 2876.06 1389.98 2876.26 ;
     RECT  1298.78 2890.76 1389.98 2898.1 ;
     RECT  1389.7 1610.6 1390.18 1610.8 ;
     RECT  1349.86 2476.64 1390.66 2494.9 ;
     RECT  1388.9 835.1 1391.78 835.3 ;
     RECT  1380.58 1868.48 1391.9 1877.08 ;
     RECT  1389.98 1914.26 1392.1 2013.58 ;
     RECT  1386.14 1805.06 1392.58 1850.2 ;
     RECT  1391.9 1865.12 1393.82 1877.08 ;
     RECT  1383.26 2069.24 1394.02 2121.1 ;
     RECT  1388.9 846.86 1394.18 847.06 ;
     RECT  1382.98 2130.14 1394.3 2144.2 ;
     RECT  1389.98 2152.82 1394.3 2243.32 ;
     RECT  1392.1 1914.26 1394.5 2013.16 ;
     RECT  1391.42 1665.2 1395.46 1665.4 ;
     RECT  1205.38 1501.4 1396.7 1501.6 ;
     RECT  1336.22 2022.62 1397.18 2041.3 ;
     RECT  1371.94 2437.16 1397.38 2459.2 ;
     RECT  1396.7 1498.46 1397.86 1501.6 ;
     RECT  1397.18 2022.62 1398.14 2044.66 ;
     RECT  1394.5 1984.82 1398.82 2013.16 ;
     RECT  1397.66 750.44 1399.54 750.64 ;
     RECT  1377.22 1886.96 1399.58 1904.38 ;
     RECT  1394.5 1914.26 1399.58 1975.36 ;
     RECT  1396.7 1661 1399.78 1661.2 ;
     RECT  1398.62 1712.66 1399.78 1717.48 ;
     RECT  1394.3 2130.14 1400.06 2243.32 ;
     RECT  1399.1 760.94 1400.26 761.14 ;
     RECT  1397.18 3203.66 1400.26 3203.86 ;
     RECT  1389.98 791.6 1401.02 791.8 ;
     RECT  1398.14 820.58 1401.02 820.78 ;
     RECT  1398.62 1702.58 1401.02 1702.78 ;
     RECT  1399.78 1712.66 1401.02 1713.28 ;
     RECT  1401.02 820.16 1401.22 822.04 ;
     RECT  1385.38 1681.16 1401.22 1681.36 ;
     RECT  1401.02 1702.58 1401.22 1713.28 ;
     RECT  1392.58 1805.06 1401.22 1847.68 ;
     RECT  1400.54 811.34 1401.7 811.54 ;
     RECT  1401.22 1702.58 1401.7 1705.72 ;
     RECT  1401.02 789.08 1401.98 791.8 ;
     RECT  1400.06 2129.72 1402.18 2243.32 ;
     RECT  1401.98 781.1 1402.535 791.8 ;
     RECT  1399.58 1886.96 1402.66 1975.36 ;
     RECT  1398.82 1985.24 1402.66 2013.16 ;
     RECT  1402.18 2129.72 1402.66 2239.96 ;
     RECT  1399.58 1622.36 1403.14 1622.56 ;
     RECT  1401.7 1702.58 1403.14 1702.78 ;
     RECT  1371.26 1758.86 1403.14 1793.5 ;
     RECT  1402.66 2151.56 1403.14 2239.96 ;
     RECT  1401.02 1728.62 1403.62 1728.82 ;
     RECT  1379.42 1631.18 1404.1 1631.38 ;
     RECT  1400.06 1642.52 1404.1 1642.72 ;
     RECT  1402.535 628 1404.265 633.48 ;
     RECT  1402.535 781.1 1404.265 799.92 ;
     RECT  1402.535 958.6 1404.265 964.08 ;
     RECT  1394.02 2116.28 1404.38 2121.1 ;
     RECT  1402.66 2129.72 1404.38 2136.64 ;
     RECT  995.6 594.8 1404.4 599.4 ;
     RECT  998.98 981.64 1404.4 986.24 ;
     RECT  1394.02 2069.24 1405.34 2103.46 ;
     RECT  1404.38 2116.28 1405.34 2136.64 ;
     RECT  1393.82 1861.76 1406.02 1877.08 ;
     RECT  1397.86 1501.4 1406.3 1501.6 ;
     RECT  1405.34 2069.24 1406.3 2136.64 ;
     RECT  1402.66 2004.98 1406.5 2013.16 ;
     RECT  1403.14 2151.56 1406.5 2232.82 ;
     RECT  1405.135 616.6 1406.865 622.08 ;
     RECT  1405.135 947.2 1406.865 952.68 ;
     RECT  1404.4 594.8 1407 596.8 ;
     RECT  1404.4 984.24 1407 986.24 ;
     RECT  1402.66 1901.66 1407.26 1975.36 ;
     RECT  1401.98 823.94 1407.46 824.14 ;
     RECT  1406.3 1501.4 1407.46 1510 ;
     RECT  1406.5 2232.2 1407.46 2232.82 ;
     RECT  1390.66 2476.64 1407.46 2479.36 ;
     RECT  1398.14 2022.62 1407.74 2051.8 ;
     RECT  1404.265 781.1 1407.94 789.28 ;
     RECT  1401.98 839.06 1408.42 839.26 ;
     RECT  1402.66 1985.24 1408.42 1994.26 ;
     RECT  1407.94 789.08 1408.9 789.28 ;
     RECT  1408.22 1652.6 1408.9 1652.8 ;
     RECT  1403.14 1781.96 1409.86 1793.5 ;
     RECT  1407.74 2022.62 1409.86 2054.32 ;
     RECT  1401.22 1808.42 1410.14 1842.64 ;
     RECT  1406.3 2066.3 1410.34 2136.64 ;
     RECT  1389.98 2876.06 1410.34 2898.1 ;
     RECT  1410.34 2066.3 1410.62 2124.46 ;
     RECT  1406.02 1861.76 1411.1 1872.46 ;
     RECT  1406.5 2151.56 1411.1 2222.74 ;
     RECT  1410.14 1733.24 1411.3 1733.44 ;
     RECT  1410.14 1801.7 1411.58 1842.64 ;
     RECT  1408.42 1990.28 1411.58 1994.26 ;
     RECT  1406.5 2004.98 1411.58 2007.7 ;
     RECT  1411.1 1855.88 1412.06 1872.46 ;
     RECT  1410.34 2136.02 1412.06 2136.64 ;
     RECT  1411.1 2145.26 1412.06 2222.74 ;
     RECT  1410.62 2061.26 1413.7 2124.46 ;
     RECT  1412.06 2136.02 1413.7 2222.74 ;
     RECT  1397.38 2437.16 1415.14 2451.64 ;
     RECT  1411.58 1801.7 1415.9 1843.06 ;
     RECT  1412.06 1852.94 1415.9 1872.46 ;
     RECT  1413.7 2136.02 1416.1 2221.06 ;
     RECT  1407.46 2232.2 1416.38 2232.4 ;
     RECT  1403.14 1758.86 1416.86 1767.88 ;
     RECT  1409.86 1781.96 1416.86 1790.56 ;
     RECT  1411.58 1990.28 1416.86 2007.7 ;
     RECT  1409.86 2022.62 1416.86 2051.8 ;
     RECT  1407.26 1901.66 1418.78 1976.62 ;
     RECT  1413.7 2118.8 1419.26 2124.46 ;
     RECT  1416.1 2136.02 1419.26 2136.22 ;
     RECT  1416.1 2145.26 1419.46 2221.06 ;
     RECT  1407.46 2476.64 1419.46 2476.84 ;
     RECT  1416.38 2232.2 1420.22 2236.6 ;
     RECT  1417.82 2246.48 1420.22 2246.68 ;
     RECT  1419.26 2118.8 1420.42 2136.22 ;
     RECT  1307.68 2919.32 1420.7 3183.08 ;
     RECT  1416.86 1990.28 1421.86 2051.8 ;
     RECT  1413.7 2061.26 1422.14 2104.3 ;
     RECT  1422.14 2059.16 1422.82 2104.3 ;
     RECT  1422.14 2275.46 1422.82 2280.7 ;
     RECT  1416.86 1758.86 1423.58 1790.56 ;
     RECT  1415.9 1801.7 1423.58 1872.46 ;
     RECT  1419.46 2152.4 1423.58 2221.06 ;
     RECT  1420.22 2232.2 1423.58 2246.68 ;
     RECT  1422.82 2061.26 1424.06 2104.3 ;
     RECT  1423.58 2152.4 1425.22 2246.68 ;
     RECT  1423.58 1758.86 1425.5 1872.46 ;
     RECT  1422.82 2280.5 1425.7 2280.7 ;
     RECT  1425.5 1688.3 1426.66 1688.5 ;
     RECT  1421.86 1990.28 1426.94 2045.5 ;
     RECT  1426.94 1989.86 1427.62 2045.5 ;
     RECT  1424.06 2061.26 1427.9 2106.82 ;
     RECT  1418.78 1734.5 1428.1 1734.7 ;
     RECT  1425.22 2152.4 1428.38 2221.06 ;
     RECT  1425.5 1757.18 1428.86 1872.46 ;
     RECT  1420.7 2911.34 1428.86 3183.08 ;
     RECT  1428.86 2911.34 1429.06 3187.06 ;
     RECT  1425.98 1645.88 1429.34 1646.08 ;
     RECT  1420.42 2118.8 1429.34 2123.62 ;
     RECT  1420.42 2132.24 1429.34 2136.22 ;
     RECT  1429.06 2920.12 1429.34 3187.06 ;
     RECT  1429.34 2118.8 1429.54 2136.22 ;
     RECT  1428.86 2295.2 1429.54 2295.4 ;
     RECT  1410.34 2876.06 1429.54 2890.96 ;
     RECT  1429.34 1645.88 1430.5 1652.8 ;
     RECT  1428.38 2147.36 1430.98 2221.06 ;
     RECT  1427.62 1990.28 1431.74 2045.5 ;
     RECT  1431.74 1990.28 1432.7 2050.96 ;
     RECT  1427.9 2061.26 1432.7 2107.24 ;
     RECT  1432.7 1737.44 1433.38 1742.26 ;
     RECT  1417.34 1672.34 1433.66 1672.54 ;
     RECT  1433.38 1740.38 1433.66 1742.26 ;
     RECT  1428.86 1751.3 1433.66 1872.46 ;
     RECT  1429.54 2135.18 1434.14 2136.22 ;
     RECT  1402.66 1886.96 1434.34 1893.04 ;
     RECT  1432.7 1990.28 1435.1 2107.24 ;
     RECT  1429.54 2118.8 1435.1 2124.46 ;
     RECT  1434.14 2135.18 1435.3 2138.32 ;
     RECT  1429.54 2890.76 1436.26 2890.96 ;
     RECT  1433.66 1669.4 1436.74 1672.54 ;
     RECT  1429.54 2876.06 1436.74 2876.26 ;
     RECT  1240.42 1521.14 1438.46 1521.34 ;
     RECT  1435.1 1990.28 1438.94 2124.46 ;
     RECT  1369 -70 1439 178 ;
     RECT  1407.46 1501.4 1439.42 1501.6 ;
     RECT  1430.3 2282.18 1439.42 2282.38 ;
     RECT  1434.34 1886.96 1439.62 1892.2 ;
     RECT  1430.98 2152.4 1439.9 2221.06 ;
     RECT  1439.42 1501.4 1440.1 1507.06 ;
     RECT  1438.46 1518.2 1440.1 1521.34 ;
     RECT  1434.62 1710.56 1440.1 1710.76 ;
     RECT  1438.94 1989.44 1440.1 2124.46 ;
     RECT  1418.78 1901.66 1440.38 1979.56 ;
     RECT  1440.1 1989.44 1440.38 2120.68 ;
     RECT  1440.38 1901.66 1440.58 2120.68 ;
     RECT  1433.66 1740.38 1441.06 1872.46 ;
     RECT  1441.06 1742.06 1441.34 1872.46 ;
     RECT  1435.3 2135.6 1442.02 2138.32 ;
     RECT  1390.66 2494.7 1442.02 2494.9 ;
     RECT  1439.9 2151.98 1442.3 2221.06 ;
     RECT  1440.1 1521.14 1442.5 1521.34 ;
     RECT  1442.02 2135.6 1443.74 2135.8 ;
     RECT  1440.58 1901.66 1443.94 2053.48 ;
     RECT  1415.14 2437.16 1444.42 2444.08 ;
     RECT  1441.34 1724.84 1444.9 1725.04 ;
     RECT  1425.22 2232.2 1445.18 2246.68 ;
     RECT  1439.42 2277.14 1446.62 2282.38 ;
     RECT  1439.62 1886.96 1447.3 1888.42 ;
     RECT  1440.58 2062.94 1448.74 2120.68 ;
     RECT  1379 3222 1449 3470 ;
     RECT  1443.94 1985.24 1449.02 2053.48 ;
     RECT  1448.74 2062.94 1449.02 2084.56 ;
     RECT  1441.34 1742.06 1449.98 1876.66 ;
     RECT  1447.3 1886.96 1449.98 1888 ;
     RECT  1436.06 3203.24 1450.66 3203.44 ;
     RECT  1443.74 2130.98 1451.42 2135.8 ;
     RECT  1430.5 1650.08 1451.62 1652.8 ;
     RECT  1451.42 2130.98 1451.9 2139.58 ;
     RECT  1442.3 2148.62 1451.9 2221.06 ;
     RECT  1436.74 1672.34 1452.1 1672.54 ;
     RECT  1451.9 2130.98 1452.1 2221.06 ;
     RECT  1449.98 1742.06 1452.38 1888 ;
     RECT  1426.94 1691.24 1452.58 1691.44 ;
     RECT  1429.34 2920.12 1452.58 3187.48 ;
     RECT  1448.74 2094.02 1452.86 2120.68 ;
     RECT  1452.1 2130.98 1452.86 2135.8 ;
     RECT  1443.94 1901.66 1453.34 1976.62 ;
     RECT  1449.02 1985.24 1453.34 2084.56 ;
     RECT  1451.62 1652.18 1454.02 1652.8 ;
     RECT  1447.58 1718.96 1454.78 1719.16 ;
     RECT  1450.46 1728.62 1454.78 1728.82 ;
     RECT  1443.26 1663.1 1454.98 1663.3 ;
     RECT  1454.3 1686.2 1455.46 1686.4 ;
     RECT  1454.02 1652.6 1456.42 1652.8 ;
     RECT  1452.1 2145.26 1456.7 2221.06 ;
     RECT  1445.18 2232.2 1456.7 2252.56 ;
     RECT  1452.38 1738.28 1457.66 1888 ;
     RECT  1456.7 2145.26 1457.66 2252.56 ;
     RECT  1454.78 1718.96 1458.34 1728.82 ;
     RECT  1457.66 1737.44 1458.82 1888 ;
     RECT  1455.74 1627.4 1460.06 1627.6 ;
     RECT  1453.34 1901.66 1460.06 2084.56 ;
     RECT  1452.86 2094.02 1460.06 2135.8 ;
     RECT  1457.66 2145.26 1460.26 2260.54 ;
     RECT  1446.62 2275.04 1460.74 2282.38 ;
     RECT  1460.06 1627.4 1461.7 1628.02 ;
     RECT  1460.74 2275.04 1462.66 2280.28 ;
     RECT  1452.58 2920.12 1462.94 3183.7 ;
     RECT  1458.82 1739.96 1464.1 1888 ;
     RECT  1464.1 1741.22 1464.38 1888 ;
     RECT  1460.26 2145.26 1464.38 2218.96 ;
     RECT  1458.34 1721.48 1465.06 1728.82 ;
     RECT  1449.02 2911.34 1465.34 2911.54 ;
     RECT  1462.94 2920.12 1465.34 3187.48 ;
     RECT  1464.38 1741.22 1465.54 1892.62 ;
     RECT  1465.34 2911.34 1466.02 3187.48 ;
     RECT  1461.7 1627.82 1467.26 1628.02 ;
     RECT  1467.26 1627.82 1467.46 1633.06 ;
     RECT  1464.38 1668.14 1467.46 1668.34 ;
     RECT  1467.46 1632.86 1467.94 1633.06 ;
     RECT  1466.02 2914.28 1468.7 3187.48 ;
     RECT  1468.7 2914.28 1468.9 3187.9 ;
     RECT  1464.38 2144.84 1469.18 2218.96 ;
     RECT  1468.9 2915.12 1470.62 3187.9 ;
     RECT  1468.7 1676.54 1470.82 1676.74 ;
     RECT  1460.06 1901.66 1471.1 2135.8 ;
     RECT  1465.06 1721.48 1472.26 1721.68 ;
     RECT  1440.1 1501.4 1472.54 1501.6 ;
     RECT  1470.62 2915.12 1472.74 3189.16 ;
     RECT  1460.26 2233.88 1473.02 2260.54 ;
     RECT  1468.7 2271.68 1473.02 2271.88 ;
     RECT  1472.54 1501.4 1473.5 1510 ;
     RECT  1465.54 1741.22 1473.5 1891.36 ;
     RECT  1473.5 1501.4 1475.14 1518.4 ;
     RECT  1474.46 2689.58 1475.62 2689.78 ;
     RECT  1473.5 1740.8 1475.9 1891.36 ;
     RECT  1469.18 2144.84 1475.9 2219.8 ;
     RECT  1461.5 1643.78 1476.38 1643.98 ;
     RECT  1475.9 1735.34 1476.86 1891.78 ;
     RECT  1475.9 2144.84 1477.06 2220.64 ;
     RECT  1475.9 2314.94 1477.54 2315.14 ;
     RECT  1461.5 1558.1 1477.82 1558.3 ;
     RECT  1346.98 1566.92 1477.82 1567.12 ;
     RECT  1463.9 2301.08 1477.82 2301.28 ;
     RECT  1471.1 1901.66 1478.78 2136.22 ;
     RECT  1477.06 2144.84 1478.78 2202.16 ;
     RECT  1469.18 1540.46 1479.26 1540.66 ;
     RECT  1472.74 2915.12 1479.26 3188.32 ;
     RECT  1478.78 2739.56 1479.46 2739.76 ;
     RECT  1444.42 2437.16 1479.94 2437.36 ;
     RECT  1480.22 1578.68 1481.86 1578.88 ;
     RECT  1478.78 1901.66 1482.34 2202.16 ;
     RECT  1481.66 1634.12 1482.82 1634.32 ;
     RECT  1477.82 2301.08 1483.78 2307.58 ;
     RECT  1475.14 1501.4 1484.06 1513.36 ;
     RECT  1476.38 1643.36 1484.06 1643.98 ;
     RECT  1484.06 1639.16 1484.54 1643.98 ;
     RECT  1481.66 1666.46 1484.54 1666.66 ;
     RECT  1476.86 1730.3 1484.54 1891.78 ;
     RECT  1463.9 1710.98 1485.5 1711.18 ;
     RECT  1484.54 1730.3 1485.5 1893.04 ;
     RECT  1482.34 1901.66 1485.5 2196.7 ;
     RECT  1485.02 1627.4 1486.18 1627.6 ;
     RECT  1485.5 1710.98 1486.18 1720.84 ;
     RECT  1465.82 1599.68 1487.42 1599.88 ;
     RECT  1486.94 1611.44 1487.42 1611.64 ;
     RECT  1484.06 1501.4 1488.1 1519.66 ;
     RECT  1477.06 2210.78 1489.34 2220.64 ;
     RECT  1487.42 1599.68 1490.02 1611.64 ;
     RECT  1485.5 1730.3 1490.02 2196.7 ;
     RECT  1486.18 1710.98 1490.3 1719.58 ;
     RECT  1484.54 1582.04 1490.78 1582.24 ;
     RECT  1490.3 1706.78 1490.78 1719.58 ;
     RECT  1489.34 2210.36 1490.78 2220.64 ;
     RECT  1473.02 2233.88 1490.78 2271.88 ;
     RECT  1483.78 2301.08 1490.98 2305.06 ;
     RECT  1484.54 1639.16 1491.26 1650.28 ;
     RECT  1490.02 1730.3 1491.26 1893.46 ;
     RECT  1479.26 1540.46 1491.46 1547.8 ;
     RECT  1490.78 1582.04 1492.42 1588.54 ;
     RECT  1490.78 2210.36 1492.42 2271.88 ;
     RECT  1484.54 1666.46 1492.7 1668.76 ;
     RECT  1491.26 1634.12 1492.9 1650.28 ;
     RECT  1492.42 2210.36 1493.38 2220.64 ;
     RECT  1490.02 1904.6 1493.66 2196.7 ;
     RECT  1493.38 2210.36 1493.66 2218.54 ;
     RECT  1491.26 1728.2 1493.86 1893.46 ;
     RECT  1492.9 1639.16 1494.34 1650.28 ;
     RECT  1490.98 2301.08 1494.34 2301.28 ;
     RECT  1479.26 2908.82 1495.3 3188.32 ;
     RECT  1491.46 1547.6 1495.78 1547.8 ;
     RECT  1493.18 1625.3 1495.78 1625.5 ;
     RECT  1479.74 1491.32 1496.06 1491.52 ;
     RECT  1496.06 1491.32 1496.54 1494.04 ;
     RECT  1495.3 2908.82 1496.74 3187.9 ;
     RECT  1496.54 1487.12 1497.02 1494.04 ;
     RECT  1492.7 1666.46 1497.02 1675.06 ;
     RECT  1488.1 1506.02 1497.22 1519.66 ;
     RECT  1490.78 1699.22 1497.5 1719.58 ;
     RECT  1493.66 1904.6 1498.46 2218.54 ;
     RECT  1497.5 1695.44 1498.66 1719.58 ;
     RECT  1493.86 1729.88 1498.94 1893.46 ;
     RECT  1497.22 1506.86 1499.14 1519.66 ;
     RECT  1492.42 1582.04 1499.42 1584.76 ;
     RECT  1490.02 1599.68 1499.42 1600.72 ;
     RECT  1492.42 2233.04 1499.9 2271.88 ;
     RECT  1498.46 1902.92 1500.1 2218.54 ;
     RECT  1496.74 2917.22 1500.58 3187.9 ;
     RECT  1499.14 1507.7 1500.86 1519.66 ;
     RECT  1203.94 1531.64 1500.86 1531.84 ;
     RECT  1497.02 1475.78 1501.06 1494.04 ;
     RECT  1499.42 1599.68 1501.06 1601.56 ;
     RECT  1497.02 1658.48 1501.06 1675.06 ;
     RECT  1500.58 2917.22 1501.06 3184.12 ;
     RECT  1498.66 1695.44 1501.54 1695.64 ;
     RECT  1500.86 1507.7 1501.82 1531.84 ;
     RECT  1494.34 1639.16 1502.78 1643.98 ;
     RECT  1498.66 1706.78 1502.98 1719.58 ;
     RECT  1477.82 1558.1 1503.46 1567.12 ;
     RECT  1499.9 2233.04 1503.46 2278.6 ;
     RECT  1499.42 1576.58 1503.94 1584.76 ;
     RECT  1501.82 1507.7 1504.42 1533.52 ;
     RECT  1359.46 2408.18 1504.42 2416.36 ;
     RECT  1502.98 1717.7 1504.7 1719.58 ;
     RECT  1502.98 1706.78 1504.9 1707.82 ;
     RECT  1502.78 1639.16 1505.18 1646.92 ;
     RECT  1501.06 1475.78 1505.38 1491.52 ;
     RECT  1504.7 2295.2 1505.86 2299.18 ;
     RECT  1505.86 2298.98 1506.34 2299.18 ;
     RECT  1504.7 1717.7 1506.62 1721.26 ;
     RECT  1498.94 1729.88 1506.62 1894.3 ;
     RECT  1500.1 1902.92 1506.62 2013.16 ;
     RECT  1505.38 1475.78 1506.82 1487.32 ;
     RECT  1504.42 1529.12 1506.82 1533.52 ;
     RECT  1501.06 1599.68 1506.82 1600.72 ;
     RECT  1503.46 1563.56 1507.78 1567.12 ;
     RECT  1500.1 2021.78 1508.06 2218.54 ;
     RECT  1506.82 1475.78 1508.26 1483.96 ;
     RECT  1505.18 1630.76 1508.26 1646.92 ;
     RECT  1506.82 1529.12 1508.74 1531.84 ;
     RECT  1508.26 1631.18 1509.5 1646.92 ;
     RECT  1508.06 2021.78 1510.18 2219.8 ;
     RECT  1508.74 1529.54 1510.66 1531.84 ;
     RECT  1509.5 1631.18 1511.9 1649.86 ;
     RECT  1501.06 1666.46 1511.9 1675.06 ;
     RECT  1504.42 1509.8 1512.1 1519.66 ;
     RECT  1507.78 1563.98 1512.1 1567.12 ;
     RECT  1511.9 1631.18 1512.1 1650.28 ;
     RECT  1511.9 1666.46 1512.1 1683.46 ;
     RECT  1512.1 1566.92 1512.38 1567.12 ;
     RECT  1503.94 1576.58 1512.38 1576.78 ;
     RECT  1512.1 1666.46 1512.38 1670.86 ;
     RECT  1506.62 1717.7 1512.38 2013.16 ;
     RECT  1510.18 2021.78 1512.38 2202.16 ;
     RECT  1512.38 1717.7 1513.06 2202.16 ;
     RECT  1512.1 1509.8 1513.54 1511.68 ;
     RECT  1512.1 1680.32 1514.78 1683.46 ;
     RECT  1501.06 2920.12 1514.78 3184.12 ;
     RECT  1514.78 1680.32 1515.46 1691.44 ;
     RECT  1512.38 1661 1515.94 1670.86 ;
     RECT  1504.9 1707.62 1516.22 1707.82 ;
     RECT  1513.06 1717.7 1516.22 2085.4 ;
     RECT  1503.46 2233.04 1516.7 2271.88 ;
     RECT  1513.34 1548.02 1517.66 1548.22 ;
     RECT  1513.54 1509.8 1517.86 1510 ;
     RECT  1512.1 1631.18 1517.86 1639.36 ;
     RECT  1514.78 2912.6 1518.14 3184.12 ;
     RECT  1512.1 1650.08 1518.62 1650.28 ;
     RECT  1513.06 2095.7 1518.62 2202.16 ;
     RECT  1510.18 2210.78 1518.62 2219.8 ;
     RECT  1512.38 1566.92 1519.1 1576.78 ;
     RECT  1517.18 1585.82 1519.1 1586.02 ;
     RECT  1515.46 1683.26 1519.3 1683.46 ;
     RECT  1510.66 1529.54 1519.58 1529.74 ;
     RECT  1519.1 1566.92 1520.06 1586.02 ;
     RECT  1506.82 1599.68 1520.06 1599.88 ;
     RECT  1518.62 2095.7 1520.54 2219.8 ;
     RECT  1515.94 1665.2 1521.7 1670.86 ;
     RECT  1516.22 1707.62 1521.7 2085.4 ;
     RECT  1519.58 1529.54 1522.66 1536.46 ;
     RECT  1521.7 1670.66 1522.66 1670.86 ;
     RECT  1521.7 1713.5 1523.42 2085.4 ;
     RECT  1520.54 2095.7 1523.42 2221.06 ;
     RECT  1516.7 2232.2 1523.42 2271.88 ;
     RECT  1522.66 1529.54 1524.1 1531.42 ;
     RECT  1523.42 1713.5 1524.1 2271.88 ;
     RECT  1518.14 2912.6 1524.1 3187.48 ;
     RECT  1508.26 1475.78 1525.06 1475.98 ;
     RECT  1524.1 2912.6 1525.06 3184.12 ;
     RECT  1520.06 1566.92 1526.02 1599.88 ;
     RECT  1517.66 1548.02 1526.5 1555.36 ;
     RECT  1518.62 1650.08 1526.5 1653.64 ;
     RECT  1524.1 1713.92 1526.5 2271.88 ;
     RECT  1526.02 1566.92 1526.78 1585.18 ;
     RECT  1526.5 1713.92 1527.94 2013.16 ;
     RECT  1527.74 1698.38 1528.42 1699.42 ;
     RECT  1526.5 2021.78 1528.42 2271.88 ;
     RECT  1528.42 2201.96 1528.9 2271.88 ;
     RECT  1526.78 1559.36 1529.38 1585.18 ;
     RECT  1528.42 2021.78 1529.86 2192.08 ;
     RECT  1529.86 2094.44 1533.7 2192.08 ;
     RECT  1524.1 1531.22 1534.46 1531.42 ;
     RECT  1524.38 1679.9 1534.46 1680.1 ;
     RECT  1525.06 2915.12 1534.94 3184.12 ;
     RECT  1526.5 1548.02 1535.14 1548.22 ;
     RECT  1527.94 1715.6 1536.86 2013.16 ;
     RECT  1529.86 2021.78 1536.86 2085.4 ;
     RECT  1513.34 1498.46 1537.06 1499.08 ;
     RECT  1537.06 1498.46 1537.34 1498.66 ;
     RECT  1534.46 1528.7 1537.82 1531.42 ;
     RECT  1534.46 1679.9 1538.78 1684.72 ;
     RECT  1529.38 1559.36 1540.22 1567.12 ;
     RECT  1529.38 1576.58 1540.22 1585.18 ;
     RECT  1540.22 1559.36 1540.7 1585.18 ;
     RECT  1511.42 1444.7 1541.18 1444.9 ;
     RECT  1533.7 2169.62 1541.18 2192.08 ;
     RECT  1528.9 2202.8 1541.18 2271.88 ;
     RECT  1536.86 1715.6 1541.66 2085.4 ;
     RECT  1541.18 2169.62 1541.86 2274.82 ;
     RECT  1534.94 2915.12 1541.86 3187.48 ;
     RECT  1541.66 1711.82 1542.14 2085.4 ;
     RECT  1533.7 2094.44 1542.14 2159.74 ;
     RECT  1540.7 1559.36 1542.82 1586.02 ;
     RECT  1529.66 1695.44 1543.1 1695.64 ;
     RECT  1537.34 1494.68 1543.3 1498.66 ;
     RECT  1537.82 1528.28 1544.06 1531.42 ;
     RECT  1542.82 1566.92 1544.54 1586.02 ;
     RECT  1542.14 1711.82 1544.54 2159.74 ;
     RECT  1542.14 1510.22 1545.22 1510.42 ;
     RECT  1538.78 1675.7 1545.5 1684.72 ;
     RECT  1541.86 2915.12 1545.7 3184.12 ;
     RECT  1526.5 1650.08 1545.98 1650.28 ;
     RECT  1545.5 1671.92 1546.94 1684.72 ;
     RECT  1543.1 1695.44 1546.94 1696.9 ;
     RECT  1544.54 1566.92 1547.9 1589.38 ;
     RECT  1526.02 1599.68 1547.9 1599.88 ;
     RECT  1546.94 1671.92 1547.9 1696.9 ;
     RECT  1541.86 2204.48 1548.1 2274.82 ;
     RECT  1541.18 1444.7 1549.34 1445.32 ;
     RECT  1490.02 1611.44 1549.34 1611.64 ;
     RECT  1544.54 1709.72 1549.34 2159.74 ;
     RECT  1547.9 1566.92 1549.82 1599.88 ;
     RECT  1547.9 1668.56 1549.82 1696.9 ;
     RECT  1549.34 1709.72 1549.82 2163.94 ;
     RECT  1548.1 2212.46 1549.82 2274.82 ;
     RECT  1545.7 2920.12 1550.78 3184.12 ;
     RECT  1549.34 1611.44 1550.98 1613.74 ;
     RECT  1549.82 1566.92 1551.46 1601.98 ;
     RECT  1545.98 1650.08 1552.22 1654.06 ;
     RECT  1549.82 1668.56 1552.42 2163.94 ;
     RECT  1549.82 2212.46 1552.42 2277.76 ;
     RECT  1552.22 1650.08 1552.7 1656.58 ;
     RECT  1552.42 2069.66 1553.38 2163.94 ;
     RECT  1544.06 1528.28 1553.66 1531.84 ;
     RECT  1528.7 1459.82 1554.14 1460.02 ;
     RECT  1553.38 2094.44 1554.14 2163.94 ;
     RECT  1541.86 2172.98 1554.14 2192.08 ;
     RECT  1517.86 1639.16 1554.62 1639.36 ;
     RECT  1550.78 2920.12 1554.62 3187.48 ;
     RECT  1554.62 1637.9 1555.1 1639.36 ;
     RECT  1555.1 1637.9 1555.3 1640.2 ;
     RECT  1544.06 2894.96 1555.3 2895.16 ;
     RECT  1552.7 1649.66 1555.58 1656.58 ;
     RECT  1552.42 1668.56 1555.58 2012.32 ;
     RECT  1551.46 1576.58 1556.26 1599.88 ;
     RECT  1551.46 1566.92 1556.54 1567.12 ;
     RECT  1552.42 2212.46 1556.54 2271.88 ;
     RECT  1554.14 2094.44 1557.5 2192.08 ;
     RECT  1556.54 2212.04 1557.5 2271.88 ;
     RECT  1556.26 1576.58 1557.7 1589.38 ;
     RECT  1557.5 2211.62 1558.94 2271.88 ;
     RECT  1558.94 2207.42 1559.14 2271.88 ;
     RECT  1552.42 2021.78 1560.1 2058.1 ;
     RECT  1553.66 1525.34 1560.38 1531.84 ;
     RECT  1559.14 2207.42 1560.58 2261.38 ;
     RECT  1554.14 1459.82 1561.06 1465.06 ;
     RECT  1556.26 1599.68 1561.34 1599.88 ;
     RECT  1561.34 1599.68 1562.3 1600.72 ;
     RECT  1555.58 1649.66 1562.3 2012.32 ;
     RECT  1560.1 2021.78 1562.3 2051.8 ;
     RECT  1553.38 2069.66 1562.3 2084.14 ;
     RECT  1557.5 2094.44 1562.3 2196.28 ;
     RECT  1557.7 1577.84 1562.5 1589.38 ;
     RECT  1562.3 1649.66 1562.5 2051.8 ;
     RECT  1543.3 1498.46 1562.78 1498.66 ;
     RECT  1560.38 1521.98 1562.78 1531.84 ;
     RECT  1439 0 1563 178 ;
     RECT  1555.3 1639.16 1563.74 1640.2 ;
     RECT  1562.5 1649.66 1563.74 1873.72 ;
     RECT  1563.74 1639.16 1564.22 1873.72 ;
     RECT  1564.22 1638.32 1564.7 1873.72 ;
     RECT  1564.7 1637.48 1564.9 1873.72 ;
     RECT  1562.78 1498.46 1565.18 1499.08 ;
     RECT  1561.34 1476.62 1565.38 1476.82 ;
     RECT  1562.78 1521.98 1565.38 1532.68 ;
     RECT  1562.3 2069.66 1565.66 2196.28 ;
     RECT  1556.54 1562.72 1566.62 1567.12 ;
     RECT  1562.3 1599.68 1566.82 1601.56 ;
     RECT  1564.9 1637.48 1566.82 1695.64 ;
     RECT  1565.66 2069.66 1566.82 2198.38 ;
     RECT  1566.62 1551.8 1567.1 1567.12 ;
     RECT  1562.5 1577.84 1567.1 1585.6 ;
     RECT  1566.82 2094.86 1567.78 2198.38 ;
     RECT  1565.18 1628.24 1568.06 1628.44 ;
     RECT  1567.78 2098.22 1569.02 2198.38 ;
     RECT  1567.1 1551.8 1569.7 1585.6 ;
     RECT  1560.58 2210.78 1570.94 2261.38 ;
     RECT  1559.14 2271.26 1570.94 2271.88 ;
     RECT  1568.06 1624.46 1572.1 1628.44 ;
     RECT  1449 3222 1573 3400 ;
     RECT  1566.82 2069.66 1573.34 2085.4 ;
     RECT  1566.82 1648.4 1574.78 1695.64 ;
     RECT  1564.9 1705.1 1574.78 1873.72 ;
     RECT  1569.7 1562.72 1575.74 1585.6 ;
     RECT  1569.02 2098.22 1575.94 2202.16 ;
     RECT  1570.94 2210.78 1576.22 2271.88 ;
     RECT  1565.38 1524.92 1576.42 1532.68 ;
     RECT  1572.38 1486.28 1577.38 1486.48 ;
     RECT  1554.62 2915.54 1577.66 3187.48 ;
     RECT  1573.34 2067.98 1578.14 2085.4 ;
     RECT  1562.5 1883.18 1578.34 2051.8 ;
     RECT  1574.78 1648.4 1578.62 1873.72 ;
     RECT  1573 3222 1579.1 3470 ;
     RECT  1578.14 2062.1 1579.3 2085.4 ;
     RECT  1576.22 2208.68 1579.3 2271.88 ;
     RECT  1579.1 1548.44 1580.54 1548.64 ;
     RECT  1504.42 2408.18 1580.74 2415.94 ;
     RECT  1577.66 1487.54 1581.98 1487.74 ;
     RECT  1565.18 1498.46 1581.98 1503.7 ;
     RECT  1566.82 1637.48 1581.98 1639.36 ;
     RECT  1578.62 1648.4 1581.98 1874.14 ;
     RECT  1575.74 1562.72 1582.46 1586.44 ;
     RECT  1571.42 1425.8 1583.42 1426 ;
     RECT  1549.34 1437.98 1583.42 1445.32 ;
     RECT  1580.06 3196.94 1584.1 3197.14 ;
     RECT  1572.1 1626.14 1584.38 1628.44 ;
     RECT  1581.98 1637.48 1584.38 1874.14 ;
     RECT  1578.34 1883.18 1585.06 2050.54 ;
     RECT  1584.38 1626.14 1585.82 1874.14 ;
     RECT  1585.06 1883.18 1585.82 2041.72 ;
     RECT  1580.54 1544.24 1586.02 1548.64 ;
     RECT  1577.66 2915.12 1586.3 3187.48 ;
     RECT  1581.98 1487.54 1586.5 1503.7 ;
     RECT  1585.82 1626.14 1586.5 2041.72 ;
     RECT  1580.74 2408.18 1586.5 2409.64 ;
     RECT  1575.94 2098.22 1586.78 2198.38 ;
     RECT  1579.3 2208.68 1586.78 2271.46 ;
     RECT  1586.3 1514 1587.46 1514.2 ;
     RECT  1586.78 2098.22 1587.46 2271.46 ;
     RECT  1579.1 3215.42 1587.46 3470 ;
     RECT  1586.5 1487.54 1587.94 1499.08 ;
     RECT  1566.82 1599.68 1588.22 1600.3 ;
     RECT  1550.98 1611.44 1588.22 1611.64 ;
     RECT  1587.46 2098.22 1588.22 2198.38 ;
     RECT  1587.94 1492.58 1588.42 1499.08 ;
     RECT  1579.3 2067.98 1588.7 2085.4 ;
     RECT  1588.42 1495.1 1588.9 1499.08 ;
     RECT  1576.42 1528.28 1589.18 1532.68 ;
     RECT  1586.5 1626.14 1589.38 2041.3 ;
     RECT  1582.46 1562.72 1590.14 1589.38 ;
     RECT  1588.9 1498.46 1590.34 1499.08 ;
     RECT  1589.38 1993.64 1590.34 2041.3 ;
     RECT  1588.7 2066.72 1590.34 2085.4 ;
     RECT  1578.14 1476.2 1590.82 1476.4 ;
     RECT  1588.22 1599.68 1591.3 1611.64 ;
     RECT  1588.22 2096.96 1591.58 2198.38 ;
     RECT  1590.34 1498.88 1591.78 1499.08 ;
     RECT  1590.14 1555.16 1591.78 1589.38 ;
     RECT  1589.18 1528.28 1593.7 1541.08 ;
     RECT  1591.58 2092.34 1593.7 2198.38 ;
     RECT  1590.34 2066.72 1594.18 2082.46 ;
     RECT  1589.38 1626.14 1595.14 1985.02 ;
     RECT  1590.34 1993.64 1596.1 2027.86 ;
     RECT  1590.34 2037.32 1597.82 2041.3 ;
     RECT  1585.06 2050.34 1597.82 2050.54 ;
     RECT  1595.14 1883.18 1598.02 1985.02 ;
     RECT  1561.06 1459.82 1599.26 1460.02 ;
     RECT  1595.14 1626.14 1599.46 1874.14 ;
     RECT  1360.9 2395.58 1599.94 2395.78 ;
     RECT  1591.3 1611.44 1600.22 1611.64 ;
     RECT  1599.46 1626.14 1600.22 1696.9 ;
     RECT  1596.1 2009.18 1600.7 2027.86 ;
     RECT  1597.82 2037.32 1600.7 2050.54 ;
     RECT  1594.18 2066.72 1601.18 2081.62 ;
     RECT  1600.7 2009.18 1601.38 2050.54 ;
     RECT  1593.7 2096.96 1601.38 2198.38 ;
     RECT  1586.5 2409.02 1601.86 2409.64 ;
     RECT  1601.38 2111.66 1602.14 2198.38 ;
     RECT  1587.46 2208.68 1602.14 2271.46 ;
     RECT  1591.78 1555.16 1602.34 1567.12 ;
     RECT  1601.18 2062.1 1602.34 2081.62 ;
     RECT  1602.34 1555.16 1603.3 1555.36 ;
     RECT  1596.1 1993.64 1603.3 1999.72 ;
     RECT  1603.3 1998.26 1603.78 1999.72 ;
     RECT  1589.18 2339.72 1603.78 2339.92 ;
     RECT  1602.34 2069.66 1604.06 2081.62 ;
     RECT  1599.26 1456.88 1605.02 1460.02 ;
     RECT  1604.06 2069.66 1605.02 2087.5 ;
     RECT  1601.38 2096.96 1605.02 2098.84 ;
     RECT  1602.14 2111.66 1605.7 2271.46 ;
     RECT  1598.02 1883.18 1606.46 1890.1 ;
     RECT  1598.02 1899.14 1606.46 1985.02 ;
     RECT  1601.38 2050.34 1606.46 2050.54 ;
     RECT  1606.46 1883.18 1606.94 1985.02 ;
     RECT  1595.42 2324.18 1607.62 2324.38 ;
     RECT  1605.7 2201.96 1608.58 2271.46 ;
     RECT  1601.86 2409.02 1608.58 2409.22 ;
     RECT  1593.02 1517.36 1609.06 1517.56 ;
     RECT  1599.46 1706.36 1609.34 1874.14 ;
     RECT  1606.94 1883.18 1609.34 1985.44 ;
     RECT  1606.46 2050.34 1609.54 2058.94 ;
     RECT  1586.3 2912.6 1609.54 3187.48 ;
     RECT  1600.22 1611.44 1609.82 1696.9 ;
     RECT  1609.34 1706.36 1609.82 1985.44 ;
     RECT  1609.82 1611.44 1610.02 1985.44 ;
     RECT  1609.54 2050.34 1610.98 2054.32 ;
     RECT  1610.02 1611.44 1611.94 1948.06 ;
     RECT  1611.94 1935.68 1612.42 1948.06 ;
     RECT  1591.78 1577.84 1612.9 1589.38 ;
     RECT  1611.94 1611.44 1612.9 1926.64 ;
     RECT  1601.38 2009.18 1612.9 2041.3 ;
     RECT  1605.7 2111.66 1612.9 2190.4 ;
     RECT  1605.02 2069.66 1613.18 2098.84 ;
     RECT  1612.9 2111.66 1613.18 2113.12 ;
     RECT  1612.42 1936.1 1614.82 1948.06 ;
     RECT  1613.18 2069.66 1616.54 2113.12 ;
     RECT  1612.9 2127.2 1617.98 2190.4 ;
     RECT  1609.54 2912.6 1617.98 3183.7 ;
     RECT  1617.98 2127.2 1618.46 2190.82 ;
     RECT  1608.58 2202.38 1618.46 2271.46 ;
     RECT  1612.9 1619.84 1620.1 1926.64 ;
     RECT  1620.1 1899.14 1621.06 1926.64 ;
     RECT  1612.9 2012.12 1622.5 2041.3 ;
     RECT  1558.94 2284.7 1622.78 2284.9 ;
     RECT  1616.54 2063.78 1622.98 2113.12 ;
     RECT  1612.9 1577.84 1623.26 1584.76 ;
     RECT  1610.02 1958.78 1623.26 1985.44 ;
     RECT  1603.78 1998.26 1623.26 1998.46 ;
     RECT  1622.98 2096.96 1623.46 2113.12 ;
     RECT  1605.02 1454.78 1623.74 1460.02 ;
     RECT  1621.06 1899.98 1623.74 1926.64 ;
     RECT  1614.82 1937.78 1623.74 1948.06 ;
     RECT  1623.26 1958.78 1623.94 1998.46 ;
     RECT  1622.3 1479.98 1624.7 1480.18 ;
     RECT  1624.7 1478.72 1625.18 1480.18 ;
     RECT  1623.74 1454.36 1625.38 1460.02 ;
     RECT  1623.46 2096.96 1625.38 2098.84 ;
     RECT  1617.98 2912.6 1625.86 3187.48 ;
     RECT  1602.34 1566.92 1626.14 1567.12 ;
     RECT  1625.18 1477.04 1626.62 1480.18 ;
     RECT  1622.5 2012.12 1626.62 2027.44 ;
     RECT  1623.46 2111.66 1626.62 2113.12 ;
     RECT  1618.46 2127.2 1626.62 2271.46 ;
     RECT  1623.94 1958.78 1626.82 1985.44 ;
     RECT  1591.3 1599.68 1627.1 1599.88 ;
     RECT  1622.78 2284.7 1627.1 2286.16 ;
     RECT  1593.7 1540.88 1627.3 1541.08 ;
     RECT  1627.1 1599.26 1627.3 1599.88 ;
     RECT  1626.82 1958.78 1627.3 1985.02 ;
     RECT  1625.38 1454.78 1628.54 1460.02 ;
     RECT  1626.62 1477.04 1628.54 1484.8 ;
     RECT  1623.26 1577.84 1628.54 1589.38 ;
     RECT  1627.3 1599.26 1628.54 1599.46 ;
     RECT  1628.54 1477.04 1629.02 1491.94 ;
     RECT  1626.62 2111.66 1629.02 2271.46 ;
     RECT  1627.1 2280.08 1629.02 2286.16 ;
     RECT  1629.02 2111.66 1629.22 2286.16 ;
     RECT  1593.7 1528.28 1629.7 1531.84 ;
     RECT  1629.02 1476.2 1629.98 1491.94 ;
     RECT  1629.22 2122.58 1630.66 2286.16 ;
     RECT  1623.94 1998.26 1631.14 1998.46 ;
     RECT  1610.98 2050.34 1631.14 2050.54 ;
     RECT  1629.98 1476.2 1631.62 1492.36 ;
     RECT  1628.54 1577.84 1631.62 1599.46 ;
     RECT  1623.74 1899.98 1632.1 1948.06 ;
     RECT  1622.5 2041.1 1632.1 2041.3 ;
     RECT  1631.62 1584.56 1632.58 1599.46 ;
     RECT  1629.22 2111.66 1632.58 2113.12 ;
     RECT  1563 -70 1633 178 ;
     RECT  1631.62 1476.2 1633.06 1491.94 ;
     RECT  1628.54 1454.78 1633.34 1464.22 ;
     RECT  1622.98 2063.78 1633.34 2088.34 ;
     RECT  1625.38 2096.96 1633.34 2098.42 ;
     RECT  1625.86 2916.8 1633.54 3187.48 ;
     RECT  1633.34 2063.78 1634.02 2098.42 ;
     RECT  1634.02 2063.78 1634.3 2088.34 ;
     RECT  1620.1 1619.84 1634.5 1890.1 ;
     RECT  1634.5 1668.14 1634.98 1890.1 ;
     RECT  1634.02 2098.22 1635.74 2098.42 ;
     RECT  1633.54 2920.12 1635.94 3187.48 ;
     RECT  1635.26 1506.44 1636.7 1506.64 ;
     RECT  1633.06 1477.04 1637.86 1491.94 ;
     RECT  1634.3 2058.32 1637.86 2088.34 ;
     RECT  1634.5 1619.84 1638.82 1657.42 ;
     RECT  1637.86 1484.6 1639.3 1491.94 ;
     RECT  1583.42 1425.8 1640.06 1445.32 ;
     RECT  1633.34 1454.78 1640.06 1465.06 ;
     RECT  1632.1 1900.82 1640.06 1948.06 ;
     RECT  1627.3 1960.46 1640.06 1985.02 ;
     RECT  1638.82 1638.74 1640.26 1657.42 ;
     RECT  1634.98 1668.14 1640.26 1696.48 ;
     RECT  1637.86 2058.32 1642.46 2058.52 ;
     RECT  1636.7 1506.44 1642.66 1513.78 ;
     RECT  1629.7 1528.7 1642.94 1531.84 ;
     RECT  1635.74 2098.22 1642.94 2098.84 ;
     RECT  1632.58 2111.66 1642.94 2111.86 ;
     RECT  1587.46 3222 1643 3470 ;
     RECT  1632.58 1584.56 1643.9 1589.38 ;
     RECT  1632.58 1599.26 1643.9 1599.46 ;
     RECT  1642.46 2054.96 1644.58 2058.52 ;
     RECT  1640.06 1900.82 1644.86 1985.02 ;
     RECT  1644.86 1900.4 1645.34 1985.02 ;
     RECT  1630.66 2127.62 1645.54 2286.16 ;
     RECT  1643.9 1584.56 1646.5 1599.46 ;
     RECT  1638.82 1619.84 1646.98 1627.18 ;
     RECT  1642.94 2098.22 1647.46 2115.22 ;
     RECT  1647.26 1474.94 1647.74 1475.14 ;
     RECT  1642.66 1506.44 1647.74 1506.64 ;
     RECT  1640.06 1425.8 1648.22 1465.06 ;
     RECT  1647.74 1474.94 1648.22 1475.98 ;
     RECT  1640.26 1668.14 1648.7 1672.96 ;
     RECT  1640.26 1683.26 1648.7 1696.48 ;
     RECT  1648.22 1425.8 1649.38 1475.98 ;
     RECT  1645.54 2127.62 1649.86 2271.46 ;
     RECT  1645.34 1900.4 1650.14 1990.48 ;
     RECT  1647.74 1501.4 1651.3 1506.64 ;
     RECT  1649.86 2235.14 1651.78 2271.46 ;
     RECT  1585.82 1406.06 1652.06 1406.26 ;
     RECT  1601.66 1415.3 1652.06 1415.5 ;
     RECT  1634.98 1705.1 1652.06 1890.1 ;
     RECT  1650.14 1899.14 1652.06 1990.48 ;
     RECT  1638.62 2364.92 1652.06 2365.12 ;
     RECT  1637.18 2379.62 1652.06 2379.82 ;
     RECT  1637.86 2069.66 1652.74 2088.34 ;
     RECT  1649.38 1425.8 1653.22 1465.06 ;
     RECT  1648.7 1668.14 1653.22 1696.48 ;
     RECT  1644.58 2054.96 1653.5 2055.16 ;
     RECT  1635.94 2920.12 1653.5 3184.12 ;
     RECT  1647.26 1396.4 1653.98 1396.6 ;
     RECT  1652.06 1406.06 1653.98 1415.5 ;
     RECT  1640.26 1639.16 1653.98 1657.42 ;
     RECT  1642.94 1528.7 1654.18 1536.88 ;
     RECT  1652.06 1705.1 1654.18 1990.48 ;
     RECT  1653.5 2915.54 1654.18 3191.68 ;
     RECT  1653.5 2051.18 1654.46 2055.16 ;
     RECT  1647.46 2098.64 1654.66 2115.22 ;
     RECT  1645.54 2285.96 1655.9 2286.16 ;
     RECT  1646.98 1626.14 1656.1 1627.18 ;
     RECT  1654.18 1733.24 1656.1 1990.48 ;
     RECT  1653.98 1639.16 1656.58 1657.84 ;
     RECT  1653.22 1683.26 1658.5 1696.48 ;
     RECT  1656.1 1626.98 1659.26 1627.18 ;
     RECT  1656.58 1639.16 1659.26 1651.12 ;
     RECT  1626.62 2010.44 1659.46 2027.44 ;
     RECT  1654.66 2104.1 1659.46 2115.22 ;
     RECT  1659.26 1626.98 1659.94 1651.12 ;
     RECT  1654.46 2050.34 1659.94 2055.16 ;
     RECT  1659.46 2110.82 1659.94 2115.22 ;
     RECT  1646.5 1599.26 1660.22 1599.46 ;
     RECT  1659.94 2051.18 1660.42 2055.16 ;
     RECT  1656.1 1733.24 1661.38 1985.02 ;
     RECT  1659.94 1626.98 1661.86 1627.18 ;
     RECT  1655.9 2280.08 1662.34 2286.16 ;
     RECT  1662.34 2284.7 1662.62 2286.16 ;
     RECT  1639.3 1491.74 1663.1 1491.94 ;
     RECT  1654.18 1705.1 1663.1 1717.06 ;
     RECT  1661.38 1756.76 1663.3 1985.02 ;
     RECT  1654.18 1528.7 1664.06 1531.84 ;
     RECT  1649.86 2127.62 1664.06 2226.52 ;
     RECT  1651.78 2235.56 1664.06 2271.46 ;
     RECT  1660.22 1599.26 1664.26 1604.92 ;
     RECT  1663.1 1705.1 1664.26 1724.62 ;
     RECT  1664.06 2127.62 1664.54 2271.46 ;
     RECT  1652.74 2070.08 1666.18 2088.34 ;
     RECT  1665.5 2040.26 1666.66 2040.46 ;
     RECT  1649.38 1474.94 1667.42 1475.98 ;
     RECT  1653.22 1668.14 1667.42 1672.12 ;
     RECT  1661.38 1733.24 1667.62 1747.3 ;
     RECT  1659.94 2110.82 1668.38 2113.96 ;
     RECT  1664.54 2127.62 1668.38 2273.98 ;
     RECT  1664.06 1527.44 1668.86 1531.84 ;
     RECT  1663.3 1756.76 1669.06 1773.34 ;
     RECT  1667.42 1474.94 1669.34 1478.92 ;
     RECT  1626.14 1566.5 1669.34 1567.12 ;
     RECT  1646.5 1584.56 1669.34 1589.38 ;
     RECT  1664.26 1599.26 1669.34 1599.46 ;
     RECT  1667.62 1743.32 1669.82 1747.3 ;
     RECT  1669.06 1756.76 1669.82 1771.66 ;
     RECT  1659.46 2012.12 1669.82 2027.44 ;
     RECT  1669.34 1474.94 1670.02 1483.12 ;
     RECT  1668.38 2110.82 1670.02 2273.98 ;
     RECT  1669.34 1562.72 1670.3 1567.12 ;
     RECT  1667.42 1668.14 1670.3 1673.38 ;
     RECT  1659.94 1639.16 1670.78 1651.12 ;
     RECT  1670.3 1562.3 1670.98 1567.12 ;
     RECT  1669.82 2005.82 1671.26 2027.44 ;
     RECT  1670.3 2098.64 1671.26 2098.84 ;
     RECT  1670.02 2111.66 1671.26 2273.98 ;
     RECT  1654.94 1543.4 1671.46 1543.6 ;
     RECT  1653.22 1425.8 1671.74 1460.02 ;
     RECT  1654.18 2920.12 1672.7 3191.68 ;
     RECT  1671.26 2111.66 1672.9 2274.82 ;
     RECT  1670.98 1562.72 1673.66 1567.12 ;
     RECT  1662.62 2284.7 1674.62 2289.94 ;
     RECT  1672.22 2299.82 1674.62 2300.02 ;
     RECT  1669.82 1743.32 1674.82 1771.66 ;
     RECT  1670.02 1474.94 1675.58 1482.7 ;
     RECT  1670.78 1638.32 1675.58 1651.12 ;
     RECT  1666.18 2078.06 1675.58 2088.34 ;
     RECT  1671.26 2097.38 1675.58 2098.84 ;
     RECT  1674.62 2284.7 1675.78 2300.02 ;
     RECT  1663.1 1491.74 1676.06 1496.14 ;
     RECT  1651.3 1506.44 1676.06 1506.64 ;
     RECT  1676.06 1491.74 1676.54 1512.52 ;
     RECT  1675.58 2078.06 1677.02 2098.84 ;
     RECT  1676.54 1491.74 1677.22 1515.04 ;
     RECT  1673.66 1562.72 1677.22 1574.68 ;
     RECT  1668.86 1608.5 1677.5 1609.54 ;
     RECT  1670.3 1668.14 1677.5 1675.48 ;
     RECT  1658.5 1690.4 1677.5 1696.48 ;
     RECT  1663.3 1783.22 1677.5 1945.12 ;
     RECT  1664.26 1705.1 1677.7 1720.42 ;
     RECT  1668.86 1524.92 1677.98 1531.84 ;
     RECT  1674.82 1743.32 1678.46 1767.46 ;
     RECT  1677.5 1777.76 1678.46 1945.12 ;
     RECT  1677.5 1688.72 1678.66 1696.48 ;
     RECT  1672.9 2111.66 1678.66 2273.98 ;
     RECT  1672.7 2915.54 1678.66 3191.68 ;
     RECT  1677.98 1524.92 1678.94 1539.82 ;
     RECT  1663.3 1955 1678.94 1985.02 ;
     RECT  1678.94 1521.98 1679.14 1539.82 ;
     RECT  1677.5 1668.14 1679.14 1678.42 ;
     RECT  1678.66 2111.66 1679.14 2206.78 ;
     RECT  1671.26 2005.4 1679.42 2027.44 ;
     RECT  1677.5 1608.5 1679.62 1612.9 ;
     RECT  1667.62 1733.24 1679.9 1733.44 ;
     RECT  1678.46 1777.76 1680.1 1945.54 ;
     RECT  1678.46 1742.48 1680.58 1767.46 ;
     RECT  1678.94 1954.58 1680.58 1985.02 ;
     RECT  1677.02 2073.02 1680.86 2098.84 ;
     RECT  1680.1 1783.22 1682.02 1945.54 ;
     RECT  1679.62 1608.5 1682.5 1609.12 ;
     RECT  1675.58 1473.26 1682.78 1482.7 ;
     RECT  1677.22 1491.74 1682.78 1512.52 ;
     RECT  1680.86 2072.18 1683.26 2098.84 ;
     RECT  1679.14 2111.66 1683.26 2197.12 ;
     RECT  1680.58 1742.48 1683.46 1747.3 ;
     RECT  1680.58 1955 1683.46 1985.02 ;
     RECT  1678.66 2217.08 1683.94 2273.98 ;
     RECT  1671.74 1425.8 1684.42 1462.96 ;
     RECT  1669.34 1584.56 1684.42 1599.46 ;
     RECT  1679.14 1521.98 1684.9 1531.84 ;
     RECT  1675.78 2285.96 1684.9 2300.02 ;
     RECT  1679.9 1732.82 1685.66 1733.44 ;
     RECT  1683.26 2072.18 1685.86 2197.12 ;
     RECT  1684.42 1599.26 1686.82 1599.46 ;
     RECT  1682.78 1473.26 1687.3 1512.52 ;
     RECT  1685.66 1728.2 1687.3 1733.44 ;
     RECT  1683.46 1743.74 1687.78 1747.3 ;
     RECT  1679.42 1998.68 1687.78 2027.44 ;
     RECT  1675.58 1634.12 1688.26 1651.12 ;
     RECT  1678.66 1690.4 1688.26 1696.48 ;
     RECT  1682.02 1783.22 1688.54 1922.44 ;
     RECT  1687.3 1506.02 1689.02 1512.52 ;
     RECT  1684.9 1521.98 1689.02 1528.9 ;
     RECT  1688.54 1780.7 1689.02 1922.44 ;
     RECT  1689.02 1506.02 1689.22 1528.9 ;
     RECT  1685.86 2072.18 1689.22 2196.7 ;
     RECT  1687.3 1728.2 1689.7 1733.02 ;
     RECT  1684.42 1584.56 1689.98 1588.12 ;
     RECT  1678.66 2915.54 1689.98 3184.12 ;
     RECT  1688.26 1690.4 1690.66 1690.6 ;
     RECT  1689.98 2884.88 1690.66 2885.08 ;
     RECT  1689.02 1779.86 1691.14 1922.44 ;
     RECT  1679.14 2206.58 1691.42 2206.78 ;
     RECT  1683.94 2217.08 1691.42 2271.88 ;
     RECT  1679.14 1668.14 1691.9 1675.48 ;
     RECT  1689.22 2076.38 1692.1 2196.7 ;
     RECT  1691.9 1668.14 1692.58 1680.52 ;
     RECT  1682.02 1933.16 1692.58 1945.54 ;
     RECT  1687.3 1473.26 1692.86 1494.88 ;
     RECT  1688.26 1634.12 1693.06 1650.7 ;
     RECT  1691.42 2206.58 1693.54 2271.88 ;
     RECT  1692.1 2078.48 1694.3 2196.7 ;
     RECT  1693.54 2206.58 1694.3 2266.42 ;
     RECT  1680.58 1758.02 1694.5 1767.46 ;
     RECT  1681.82 2314.94 1694.78 2315.14 ;
     RECT  1694.3 2078.48 1694.98 2266.42 ;
     RECT  1694.5 1763.9 1695.46 1767.46 ;
     RECT  1684.9 2285.96 1695.46 2293.3 ;
     RECT  1683.46 1958.78 1695.74 1985.02 ;
     RECT  1692.86 1469.48 1695.94 1494.88 ;
     RECT  1689.22 1506.44 1695.94 1528.9 ;
     RECT  1677.22 1562.72 1695.94 1567.54 ;
     RECT  1691.14 1779.86 1695.94 1918.66 ;
     RECT  1694.98 2078.48 1695.94 2265.58 ;
     RECT  1689.7 1728.62 1696.22 1733.02 ;
     RECT  1687.78 1743.74 1696.22 1745.2 ;
     RECT  1696.22 1728.62 1696.7 1745.2 ;
     RECT  1682.5 1608.92 1697.18 1609.12 ;
     RECT  1695.94 1521.98 1697.66 1528.9 ;
     RECT  1660.42 2054.96 1697.86 2055.16 ;
     RECT  1697.66 2301.08 1698.14 2301.28 ;
     RECT  1694.78 2314.94 1698.14 2318.08 ;
     RECT  1689.98 2915.54 1699.1 3191.26 ;
     RECT  1689.98 1577.42 1699.3 1588.12 ;
     RECT  1695.94 2095.7 1699.78 2265.58 ;
     RECT  1684.42 1425.8 1700.06 1460.02 ;
     RECT  1699.3 1577.42 1700.26 1587.28 ;
     RECT  1695.74 1955.42 1700.26 1985.02 ;
     RECT  1699.1 2908.82 1700.26 3192.52 ;
     RECT  1695.46 2285.96 1700.54 2286.16 ;
     RECT  1692.58 1933.16 1701.02 1933.36 ;
     RECT  1700.54 2285.54 1701.02 2286.16 ;
     RECT  1699.78 2095.7 1701.7 2135.38 ;
     RECT  1700.06 1425.8 1702.18 1460.86 ;
     RECT  1693.34 1684.52 1702.18 1685.14 ;
     RECT  1695.94 1779.86 1702.18 1885.9 ;
     RECT  1692.58 1668.14 1702.46 1675.48 ;
     RECT  1695.94 1470.32 1702.66 1494.88 ;
     RECT  1701.02 1932.32 1702.66 1933.36 ;
     RECT  1701.7 2097.38 1702.66 2135.38 ;
     RECT  1701.02 2056.22 1703.14 2056.42 ;
     RECT  1696.7 1728.62 1703.42 1753.18 ;
     RECT  1702.18 1779.86 1703.42 1885.06 ;
     RECT  1700.26 2916.8 1704.38 3192.52 ;
     RECT  1699.78 2144 1704.58 2265.58 ;
     RECT  1677.7 1705.1 1704.86 1717.06 ;
     RECT  1703.42 1726.1 1704.86 1753.18 ;
     RECT  1697.66 1521.98 1705.06 1533.52 ;
     RECT  1704.38 2916.8 1705.06 3195.04 ;
     RECT  1704.58 2188.1 1705.54 2265.58 ;
     RECT  1704.38 2332.16 1705.54 2332.36 ;
     RECT  1701.5 2754.68 1705.54 2754.88 ;
     RECT  1705.06 2920.12 1705.54 3195.04 ;
     RECT  1703.42 1779.02 1705.82 1885.06 ;
     RECT  1701.02 2282.6 1705.82 2286.16 ;
     RECT  1704.86 1691.24 1706.02 1691.44 ;
     RECT  1702.66 1482.5 1706.5 1494.88 ;
     RECT  1697.18 1608.08 1706.78 1609.12 ;
     RECT  1695.46 1763.9 1706.78 1765.78 ;
     RECT  1705.82 1775.24 1706.78 1885.06 ;
     RECT  1702.66 1933.16 1706.78 1933.36 ;
     RECT  1700.26 1955.84 1706.98 1985.02 ;
     RECT  1702.46 1668.14 1707.26 1680.1 ;
     RECT  1695.94 2078.48 1707.26 2081.2 ;
     RECT  1705.54 2231.78 1707.26 2265.58 ;
     RECT  1705.82 2275.46 1707.26 2286.16 ;
     RECT  1687.78 2005.4 1708.22 2027.44 ;
     RECT  1706.5 1487.96 1708.9 1494.88 ;
     RECT  1708.22 2001.62 1708.9 2027.44 ;
     RECT  1704.58 2160.8 1708.9 2178.22 ;
     RECT  1695.94 1506.44 1709.66 1512.52 ;
     RECT  1705.06 1521.98 1709.66 1525.54 ;
     RECT  1704.86 1705.1 1709.66 1753.18 ;
     RECT  1706.78 1763.9 1709.66 1885.06 ;
     RECT  1708.22 2747.12 1709.86 2747.32 ;
     RECT  1704.58 2144 1710.34 2150.08 ;
     RECT  1706.78 1933.16 1710.82 1940.08 ;
     RECT  1698.14 2301.08 1710.82 2318.08 ;
     RECT  1700.26 1577.42 1711.58 1586.02 ;
     RECT  1705.54 2188.1 1711.78 2220.22 ;
     RECT  1706.78 1603.88 1712.06 1609.12 ;
     RECT  1702.66 2097.38 1712.26 2098.84 ;
     RECT  1710.82 2306.12 1712.26 2318.08 ;
     RECT  1709.66 1762.22 1712.54 1885.06 ;
     RECT  1695.94 1894.94 1712.54 1918.66 ;
     RECT  1707.26 2071.34 1712.74 2081.2 ;
     RECT  1707.26 2231.78 1712.74 2286.16 ;
     RECT  1712.26 2306.12 1712.74 2308.84 ;
     RECT  1709.66 1703 1713.5 1753.18 ;
     RECT  1711.58 1576.16 1713.7 1586.02 ;
     RECT  1710.14 1952.48 1713.7 1952.68 ;
     RECT  1712.26 2317.88 1713.7 2318.08 ;
     RECT  1708.9 2001.62 1713.98 2016.1 ;
     RECT  1712.74 2280.08 1713.98 2286.16 ;
     RECT  1709.66 1521.56 1714.46 1525.54 ;
     RECT  1713.5 1697.12 1714.46 1753.18 ;
     RECT  1712.54 1762.22 1714.46 1918.66 ;
     RECT  1706.98 1963.4 1714.94 1985.02 ;
     RECT  1709.66 1505.18 1715.42 1512.52 ;
     RECT  1714.46 1521.56 1715.42 1526.8 ;
     RECT  1714.46 1697.12 1715.62 1918.66 ;
     RECT  1713.98 2280.08 1715.62 2293.72 ;
     RECT  1712.06 1600.52 1715.9 1609.12 ;
     RECT  1713.98 2001.2 1715.9 2016.1 ;
     RECT  1714.46 1943.66 1716.1 1944.28 ;
     RECT  1715.62 1697.12 1716.38 1848.1 ;
     RECT  1714.46 1471.58 1716.58 1471.78 ;
     RECT  1705.54 2920.12 1716.86 3192.1 ;
     RECT  1715.42 1505.18 1717.06 1526.8 ;
     RECT  1715.9 2000.36 1717.06 2016.1 ;
     RECT  1714.94 2036.06 1717.06 2036.26 ;
     RECT  1713.98 2901.68 1717.06 2901.88 ;
     RECT  1695.94 1566.5 1717.34 1567.54 ;
     RECT  1713.7 1576.16 1717.34 1580.98 ;
     RECT  1713.5 2066.72 1717.34 2069.44 ;
     RECT  1717.34 1566.5 1717.54 1580.98 ;
     RECT  1717.06 1506.44 1718.02 1526.8 ;
     RECT  1681.82 1551.38 1719.26 1551.58 ;
     RECT  1716.86 2920.12 1719.74 3195.04 ;
     RECT  1717.34 2065.04 1719.94 2069.44 ;
     RECT  1719.26 1543.82 1720.22 1551.58 ;
     RECT  1716.38 1695.02 1720.42 1848.1 ;
     RECT  1708.9 1487.96 1720.7 1494.04 ;
     RECT  1708.9 2167.94 1720.7 2178.22 ;
     RECT  1714.94 1963.4 1720.9 1988.8 ;
     RECT  1717.06 2001.2 1720.9 2016.1 ;
     RECT  1715.9 1597.58 1721.18 1609.12 ;
     RECT  1715.62 1862.6 1721.18 1918.66 ;
     RECT  1712.26 2098.64 1721.18 2098.84 ;
     RECT  1702.66 2111.66 1721.18 2135.38 ;
     RECT  1720.7 2164.58 1721.18 2178.22 ;
     RECT  1711.78 2194.4 1721.18 2220.22 ;
     RECT  1712.74 2231.78 1721.18 2268.94 ;
     RECT  1720.9 2005.4 1721.38 2016.1 ;
     RECT  1720.9 1963.4 1721.66 1986.28 ;
     RECT  1717.54 1566.5 1722.14 1577.62 ;
     RECT  1719.94 2066.72 1722.34 2069.44 ;
     RECT  1721.18 1862.6 1722.82 1924.12 ;
     RECT  1721.18 2098.64 1723.1 2135.38 ;
     RECT  1721.18 2157.86 1723.1 2178.22 ;
     RECT  1721.18 2194.4 1723.1 2268.94 ;
     RECT  1723.1 2096.54 1723.58 2135.38 ;
     RECT  1721.66 1962.98 1723.78 1986.28 ;
     RECT  1722.82 1877.3 1724.06 1924.12 ;
     RECT  1710.82 1933.16 1724.06 1933.36 ;
     RECT  1723.58 2095.7 1724.54 2135.38 ;
     RECT  1724.06 1877.3 1725.7 1933.36 ;
     RECT  1725.02 1943.24 1725.98 1943.44 ;
     RECT  1720.22 1540.04 1726.46 1551.58 ;
     RECT  1722.14 1562.72 1726.46 1577.62 ;
     RECT  1693.06 1634.12 1728.1 1646.5 ;
     RECT  1728.1 1634.12 1729.06 1634.32 ;
     RECT  1715.62 2280.08 1729.34 2286.16 ;
     RECT  1719.26 2296.46 1729.34 2296.66 ;
     RECT  1719.74 2912.18 1729.34 3195.04 ;
     RECT  1720.42 1733.66 1729.54 1848.1 ;
     RECT  1721.18 1597.16 1729.82 1609.12 ;
     RECT  1726.46 1540.04 1730.02 1577.62 ;
     RECT  1729.82 1594.64 1730.02 1609.12 ;
     RECT  1723.1 2157.86 1730.02 2268.94 ;
     RECT  1721.66 1478.72 1730.3 1478.92 ;
     RECT  1730.02 2157.86 1730.98 2232.82 ;
     RECT  1724.54 2091.08 1731.94 2135.38 ;
     RECT  1708.9 2027.24 1732.22 2027.44 ;
     RECT  1730.02 1594.64 1732.42 1600.3 ;
     RECT  1722.34 2069.24 1732.42 2069.44 ;
     RECT  1712.74 2308.64 1733.66 2308.84 ;
     RECT  1730.3 1472 1734.62 1478.92 ;
     RECT  1723.78 1962.98 1734.82 1985.02 ;
     RECT  1729.34 2280.08 1735.1 2296.66 ;
     RECT  1733.66 2307.38 1735.1 2308.84 ;
     RECT  1731.94 2091.08 1735.3 2120.26 ;
     RECT  1734.82 1962.98 1735.58 1964.86 ;
     RECT  1712.74 2078.48 1735.58 2081.2 ;
     RECT  1725.7 1887.38 1735.78 1933.36 ;
     RECT  1729.54 1733.66 1736.06 1847.26 ;
     RECT  1730.02 1543.82 1736.26 1577.62 ;
     RECT  1730.98 2194.4 1736.26 2232.82 ;
     RECT  1725.98 1942.82 1736.54 1948.06 ;
     RECT  1735.58 1957.1 1736.54 1964.86 ;
     RECT  1732.22 2023.46 1737.98 2027.44 ;
     RECT  1733.66 2036.06 1737.98 2036.26 ;
     RECT  1736.06 1732.82 1738.18 1847.26 ;
     RECT  1736.26 2194.4 1738.66 2228.62 ;
     RECT  1737.98 2023.46 1739.14 2036.26 ;
     RECT  1710.34 2144 1739.62 2144.2 ;
     RECT  1730.98 2157.86 1740.1 2178.22 ;
     RECT  1721.38 2005.4 1740.58 2014 ;
     RECT  1734.62 1471.16 1741.06 1478.92 ;
     RECT  1735.78 1891.58 1741.06 1933.36 ;
     RECT  1736.54 1942.82 1741.06 1964.86 ;
     RECT  1738.66 2203.64 1741.06 2226.52 ;
     RECT  1735.58 2073.86 1741.34 2081.2 ;
     RECT  1722.82 1862.6 1741.82 1862.8 ;
     RECT  1736.26 1543.82 1742.02 1551.58 ;
     RECT  1739.14 2023.46 1742.02 2028.28 ;
     RECT  1735.1 2280.08 1742.02 2308.84 ;
     RECT  1740.1 2164.58 1742.5 2178.22 ;
     RECT  1741.82 1862.6 1742.78 1864.48 ;
     RECT  1725.7 1877.3 1742.78 1877.5 ;
     RECT  1729.34 2908.82 1742.98 3195.04 ;
     RECT  1718.02 1512.32 1743.26 1526.8 ;
     RECT  1730.02 2241.44 1743.26 2268.94 ;
     RECT  1742.02 2280.08 1743.26 2307.58 ;
     RECT  1738.18 1732.82 1743.46 1827.1 ;
     RECT  1738.18 1835.72 1743.46 1847.26 ;
     RECT  1741.06 1959.62 1743.46 1964.86 ;
     RECT  1743.46 1732.82 1744.42 1820.38 ;
     RECT  1744.42 1732.82 1744.7 1817.02 ;
     RECT  1720.42 1695.02 1745.18 1723.36 ;
     RECT  1744.7 1732.4 1745.18 1817.02 ;
     RECT  1738.46 2050.34 1745.38 2050.54 ;
     RECT  1744.7 2148.62 1745.38 2148.82 ;
     RECT  1735.3 2111.66 1745.86 2120.26 ;
     RECT  1743.46 1838.24 1746.14 1847.26 ;
     RECT  1741.34 2073.44 1746.14 2081.2 ;
     RECT  1741.06 2203.64 1746.82 2204.68 ;
     RECT  1742.98 2912.18 1746.82 3195.04 ;
     RECT  1742.02 2027.24 1747.58 2028.28 ;
     RECT  1736.26 1566.5 1747.78 1577.62 ;
     RECT  1743.26 2241.44 1747.78 2307.58 ;
     RECT  1745.86 2111.66 1748.54 2111.86 ;
     RECT  1731.94 2133.5 1748.54 2135.38 ;
     RECT  1738.66 2194.4 1748.74 2194.6 ;
     RECT  1741.06 1478.72 1749.5 1478.92 ;
     RECT  1720.7 1487.96 1749.5 1494.46 ;
     RECT  1729.82 2317.88 1749.5 2318.08 ;
     RECT  1747.58 2027.24 1749.7 2035.84 ;
     RECT  1748.54 2130.98 1749.7 2135.38 ;
     RECT  1747.78 2241.44 1749.7 2280.28 ;
     RECT  1749.5 2317.88 1749.7 2318.5 ;
     RECT  1743.46 1962.98 1750.46 1964.86 ;
     RECT  1734.82 1976.42 1750.46 1985.02 ;
     RECT  1746.14 2070.5 1750.46 2081.2 ;
     RECT  1746.14 1838.24 1750.66 1850.62 ;
     RECT  1750.66 1838.24 1752.1 1842.22 ;
     RECT  1746.82 2912.18 1752.58 3187.48 ;
     RECT  1745.18 1695.02 1753.34 1817.02 ;
     RECT  1741.06 1892 1753.54 1933.36 ;
     RECT  1652.06 2364.92 1753.82 2379.82 ;
     RECT  1748.54 2109.56 1754.02 2111.86 ;
     RECT  1754.02 2110.4 1754.5 2111.86 ;
     RECT  1735.3 2091.92 1754.98 2098.84 ;
     RECT  1749.02 1469.06 1755.46 1469.26 ;
     RECT  1742.02 1543.82 1755.46 1544.86 ;
     RECT  1732.42 1597.58 1756.22 1600.3 ;
     RECT  1740.58 2005.4 1756.42 2012.74 ;
     RECT  1742.5 2167.52 1756.9 2178.22 ;
     RECT  1633 0 1757 178 ;
     RECT  1747.78 1577.42 1757.18 1577.62 ;
     RECT  1749.02 1829.42 1757.38 1829.62 ;
     RECT  1741.06 2220.02 1757.38 2226.52 ;
     RECT  1743.26 1511.48 1757.66 1526.8 ;
     RECT  1756.22 1591.28 1757.66 1600.3 ;
     RECT  1730.02 1608.92 1757.66 1609.12 ;
     RECT  1753.34 1695.02 1758.34 1819.12 ;
     RECT  1754.98 2091.92 1758.34 2097.16 ;
     RECT  1752.1 1838.24 1758.82 1838.44 ;
     RECT  1750.46 1962.98 1758.82 1985.02 ;
     RECT  1758.34 1725.68 1759.3 1819.12 ;
     RECT  1753.54 1892 1759.78 1927.48 ;
     RECT  1750.46 2068.4 1759.78 2081.2 ;
     RECT  1757.66 1508.96 1760.06 1526.8 ;
     RECT  1757.66 1591.28 1760.26 1609.12 ;
     RECT  1760.06 1508.96 1760.74 1529.32 ;
     RECT  1759.3 1765.58 1761.22 1819.12 ;
     RECT  1761.22 1765.58 1761.7 1807.78 ;
     RECT  1757.18 1577.42 1761.98 1582.24 ;
     RECT  1760.26 1591.28 1761.98 1600.3 ;
     RECT  1761.7 1765.58 1762.18 1786.78 ;
     RECT  1761.98 1577.42 1762.66 1600.3 ;
     RECT  1759.78 1892 1762.66 1895.14 ;
     RECT  1758.34 2096.12 1762.66 2097.16 ;
     RECT  1760.74 1508.96 1763.14 1526.8 ;
     RECT  1762.18 1767.26 1763.14 1786.78 ;
     RECT  1742.78 1862.6 1763.14 1877.5 ;
     RECT  1761.22 1818.92 1763.62 1819.12 ;
     RECT  1758.82 1974.74 1763.62 1985.02 ;
     RECT  1759.78 2073.44 1763.9 2081.2 ;
     RECT  1749.7 2241.44 1763.9 2278.6 ;
     RECT  1757.38 2224.22 1764.1 2226.52 ;
     RECT  1752.58 2912.18 1764.38 3183.7 ;
     RECT  1702.18 1425.8 1764.58 1460.02 ;
     RECT  1763.14 1511.48 1764.58 1526.8 ;
     RECT  1653.98 1396.4 1764.86 1415.5 ;
     RECT  1762.66 1589.6 1765.06 1600.3 ;
     RECT  1764.38 2904.62 1765.06 3183.7 ;
     RECT  1763.9 2241.44 1765.54 2283.22 ;
     RECT  1763.9 2073.44 1766.02 2084.14 ;
     RECT  1763.14 1770.62 1766.5 1786.78 ;
     RECT  1763.62 1976.42 1766.5 1985.02 ;
     RECT  1766.5 1770.62 1766.98 1782.16 ;
     RECT  1761.7 1796.24 1766.98 1807.78 ;
     RECT  1765.82 2055.38 1766.98 2055.58 ;
     RECT  1643 3222 1767 3400 ;
     RECT  1765.06 2912.18 1767.74 3183.7 ;
     RECT  1758.82 1962.98 1768.7 1963.6 ;
     RECT  1766.5 1976.42 1768.9 1982.92 ;
     RECT  1766.02 2073.44 1769.38 2078.68 ;
     RECT  1763.14 1872.68 1769.86 1877.5 ;
     RECT  1765.82 1847.06 1770.14 1847.26 ;
     RECT  1768.7 1962.98 1770.14 1964.86 ;
     RECT  1768.7 2097.8 1770.62 2098 ;
     RECT  1759.78 1904.18 1770.82 1927.48 ;
     RECT  1765.06 1591.28 1771.1 1600.3 ;
     RECT  1760.26 1608.92 1771.1 1609.12 ;
     RECT  1759.3 1725.68 1771.1 1753.18 ;
     RECT  1770.62 2097.8 1771.1 2099.26 ;
     RECT  1765.54 2241.44 1771.1 2276.5 ;
     RECT  1768.7 1626.98 1771.3 1627.18 ;
     RECT  1766.98 1796.24 1771.3 1801.06 ;
     RECT  1771.1 1591.28 1772.06 1609.12 ;
     RECT  1741.06 1942.82 1772.06 1948.06 ;
     RECT  1764.58 1512.32 1772.54 1526.8 ;
     RECT  1749.7 2027.24 1773.5 2027.44 ;
     RECT  1758.34 1695.02 1773.7 1714.96 ;
     RECT  1686.62 2736.2 1774.46 2736.4 ;
     RECT  1773.7 1695.02 1774.66 1714.12 ;
     RECT  1749.5 1478.72 1774.94 1494.46 ;
     RECT  1771.1 1724.84 1774.94 1756.54 ;
     RECT  1771.1 2241.02 1775.14 2276.5 ;
     RECT  1772.06 1591.28 1775.62 1612.06 ;
     RECT  1770.14 1847.06 1775.62 1850.2 ;
     RECT  1769.18 1992.8 1775.9 1993 ;
     RECT  1756.9 2167.52 1775.9 2173.18 ;
     RECT  1767 3222 1775.9 3470 ;
     RECT  1775.62 1600.1 1776.1 1612.06 ;
     RECT  1771.3 1798.34 1776.1 1801.06 ;
     RECT  1776.1 1600.1 1776.58 1609.12 ;
     RECT  1773.5 2039 1776.86 2039.2 ;
     RECT  1772.06 1942.82 1777.06 1953.94 ;
     RECT  1764.1 2224.22 1777.34 2224.42 ;
     RECT  1774.66 1709.72 1777.54 1714.12 ;
     RECT  1763.9 1835.3 1777.54 1835.5 ;
     RECT  1763.14 1862.6 1777.54 1862.8 ;
     RECT  1775.9 1992.8 1777.82 1993.84 ;
     RECT  1756.42 2005.4 1777.82 2008.54 ;
     RECT  1777.34 1789.1 1778.5 1789.3 ;
     RECT  1771.1 2097.8 1778.5 2102.62 ;
     RECT  1773.5 3196.94 1778.5 3197.14 ;
     RECT  1747.78 1566.5 1778.78 1567.54 ;
     RECT  1762.66 1577.42 1778.78 1577.62 ;
     RECT  1775.62 1591.28 1778.78 1591.48 ;
     RECT  1774.94 1724.84 1778.78 1759.48 ;
     RECT  1766.98 1770.62 1778.78 1779.64 ;
     RECT  1762.66 1894.94 1779.26 1895.14 ;
     RECT  1770.82 1906.28 1779.26 1927.48 ;
     RECT  1774.94 1470.74 1779.46 1494.46 ;
     RECT  1779.26 1894.94 1779.46 1927.48 ;
     RECT  1770.14 1962.98 1779.46 1967.8 ;
     RECT  1776.86 2039 1779.46 2042.56 ;
     RECT  1778.78 1577.42 1780.42 1591.48 ;
     RECT  1773.5 2023.04 1780.7 2027.44 ;
     RECT  1777.54 1709.72 1781.86 1713.7 ;
     RECT  1775.9 3220.04 1781.86 3470 ;
     RECT  1774.66 1695.02 1782.34 1695.22 ;
     RECT  1775.62 1850 1782.34 1850.2 ;
     RECT  1772.54 1512.32 1782.62 1532.68 ;
     RECT  1777.82 1992.8 1782.82 2008.54 ;
     RECT  1778.5 2097.8 1783.3 2099.68 ;
     RECT  1782.82 1992.8 1783.58 1993 ;
     RECT  1770.14 2088.56 1783.78 2088.76 ;
     RECT  1782.62 1512.32 1784.26 1533.1 ;
     RECT  1768.9 1976.42 1784.74 1976.62 ;
     RECT  1755.46 1543.82 1785.02 1544.02 ;
     RECT  1779.46 2039 1785.7 2039.2 ;
     RECT  1783.3 2099.06 1786.18 2099.68 ;
     RECT  1777.34 2224.22 1786.46 2228.62 ;
     RECT  1776.1 1798.34 1787.9 1800.64 ;
     RECT  1777.06 1942.82 1787.9 1948.48 ;
     RECT  1778.78 1724.84 1788.1 1779.64 ;
     RECT  1787.9 1798.34 1789.06 1804 ;
     RECT  1786.18 2099.48 1789.06 2099.68 ;
     RECT  1786.46 2224.22 1789.06 2231.98 ;
     RECT  1788.1 1724.84 1789.54 1772.08 ;
     RECT  1786.46 2050.34 1789.54 2050.54 ;
     RECT  1789.06 1798.34 1789.82 1800.64 ;
     RECT  1789.54 1763.9 1790.5 1772.08 ;
     RECT  1789.82 1793.3 1790.5 1800.64 ;
     RECT  1780.7 2020.52 1790.78 2027.44 ;
     RECT  1775.9 2164.16 1791.74 2173.18 ;
     RECT  1790.5 1771.88 1792.42 1772.08 ;
     RECT  1790.5 1793.3 1792.42 1798.54 ;
     RECT  1775.14 2241.02 1793 2268.94 ;
     RECT  1781.66 2285.96 1793 2286.16 ;
     RECT  1793.135 1017.88 1794.865 1023.36 ;
     RECT  1793.135 1628.92 1794.865 1634.4 ;
     RECT  1793 994.8 1795.6 996.8 ;
     RECT  1728.1 1646.3 1795.735 1646.5 ;
     RECT  1747.78 2296.46 1796.26 2307.58 ;
     RECT  1795.735 1029.28 1797.465 1034.76 ;
     RECT  1795.735 1640.32 1797.465 1646.5 ;
     RECT  1787.9 1942.4 1797.98 1948.48 ;
     RECT  1779.46 1962.98 1797.98 1963.18 ;
     RECT  1791.26 2069.24 1797.98 2069.44 ;
     RECT  1677.5 2548.46 1797.98 2548.66 ;
     RECT  1707.26 1667.72 1798.18 1680.1 ;
     RECT  1789.06 2227.16 1798.46 2231.98 ;
     RECT  1776.58 1608.92 1799.14 1609.12 ;
     RECT  1764.86 1396.4 1799.9 1416.76 ;
     RECT  1767.74 2912.18 1800.1 3187.48 ;
     RECT  1784.26 1512.32 1800.34 1532.68 ;
     RECT  1780.42 1577.42 1800.34 1583.92 ;
     RECT  1789.54 1724.84 1800.34 1753.18 ;
     RECT  1799.42 1658.48 1800.38 1658.68 ;
     RECT  1798.18 1667.72 1800.38 1675.48 ;
     RECT  1779.46 1470.74 1800.58 1478.92 ;
     RECT  1799.9 1395.98 1801.06 1416.76 ;
     RECT  1778.78 1558.52 1801.34 1567.54 ;
     RECT  1800.34 1577.42 1801.34 1583.9 ;
     RECT  1764.58 1425.8 1803.26 1451.62 ;
     RECT  1800.58 1471.56 1803.26 1478.92 ;
     RECT  1779.46 1487.54 1803.26 1494.46 ;
     RECT  1800.34 1512.32 1803.26 1515.04 ;
     RECT  1800.34 1524.08 1803.26 1532.68 ;
     RECT  1785.02 1543.82 1803.26 1544.44 ;
     RECT  1801.34 1558.52 1803.26 1583.9 ;
     RECT  1776.58 1600.1 1803.26 1600.3 ;
     RECT  1800.86 1626.12 1803.26 1626.32 ;
     RECT  1797.465 1642.92 1803.26 1646.5 ;
     RECT  1800.38 1658.48 1803.26 1675.48 ;
     RECT  1781.86 1713.5 1803.26 1713.7 ;
     RECT  1800.34 1724.84 1803.26 1743.94 ;
     RECT  1800.1 2912.18 1805.86 3184.12 ;
     RECT  1803.26 1622.76 1807.1 1626.32 ;
     RECT  1803.26 1642.92 1807.1 1675.48 ;
     RECT  1730.3 2868.92 1810.46 2869.12 ;
     RECT  1723.58 2883.62 1810.46 2883.82 ;
     RECT  1805.86 2912.18 1814.78 3183.7 ;
     RECT  1779.46 1894.94 1824.58 1911.94 ;
     RECT  1810.46 2868.92 1824.86 2883.82 ;
     RECT  1757 -70 1827 178 ;
     RECT  1793 2241.02 1828.9 2286.16 ;
     RECT  1781.86 3222 1837 3470 ;
     RECT  1824.86 2868.92 1875.46 2890.96 ;
     RECT  1814.78 2912.18 1882.66 3187.48 ;
     RECT  1882.66 2912.18 1893.5 3183.7 ;
     RECT  1755.74 2343.5 1898.02 2343.7 ;
     RECT  1875.46 2890.76 1920.58 2890.96 ;
     RECT  1796.26 2298.98 1925.86 2307.58 ;
     RECT  1925.86 2303.6 1947.94 2307.58 ;
     RECT  1827 0 1951 178 ;
     RECT  1792.42 1798.34 1954.66 1798.54 ;
     RECT  1828.9 2243.96 1955.14 2286.16 ;
     RECT  1837 3222 1961 3400 ;
     RECT  1893.5 2912.18 1970.98 3187.48 ;
     RECT  1954.46 3196.94 1972.9 3197.14 ;
     RECT  1970.98 2912.18 1976.26 3183.7 ;
     RECT  1790.78 2020.52 1977.7 2034.16 ;
     RECT  1782.82 2005.4 2005.54 2008.54 ;
     RECT  1961 3222 2015.9 3470 ;
     RECT  1800.34 1752.98 2016.58 1753.18 ;
     RECT  2015.9 3220.04 2016.58 3470 ;
     RECT  1951 -70 2021 178 ;
     RECT  1976.26 2912.18 2021.38 3183.08 ;
     RECT  2016.58 3222 2031 3470 ;
     RECT  1749.5 2193.14 2049.22 2193.34 ;
     RECT  1875.46 2868.92 2055.46 2876.26 ;
     RECT  1803.26 1685.76 2077.06 1743.94 ;
     RECT  1947.94 2307.38 2077.54 2307.58 ;
     RECT  1792.22 1849.16 2091.46 1849.36 ;
     RECT  1769.86 1876.46 2091.94 1877.5 ;
     RECT  2021.38 2915.54 2092.16 3183.08 ;
     RECT  2092.16 2942.2 2096.425 2959.08 ;
     RECT  2092.16 3010.6 2096.425 3068.2 ;
     RECT  2092.16 3076.72 2096.425 3093.6 ;
     RECT  2092.16 3145.12 2096.425 3162 ;
     RECT  2092.16 2915.54 2096.56 2924.72 ;
     RECT  2092.16 3178.48 2096.56 3183.08 ;
     RECT  2096.425 2942.2 2099.025 2947.68 ;
     RECT  2096.425 3010.6 2099.025 3016.08 ;
     RECT  2096.425 3076.72 2099.025 3082.2 ;
     RECT  2096.425 3145.12 2099.025 3150.6 ;
     RECT  2096.56 2915.54 2099.16 2922.12 ;
     RECT  2096.56 3181.08 2099.16 3183.08 ;
     RECT  2099.16 2915.54 2101.06 2915.74 ;
     RECT  2096.425 3032.3 2101.06 3068.2 ;
     RECT  2055.46 2876.06 2101.54 2876.26 ;
     RECT  2101.06 3032.3 2102.02 3032.5 ;
     RECT  2101.06 3045.32 2102.02 3061.06 ;
     RECT  2102.02 3052.88 2104.42 3061.06 ;
     RECT  2104.42 3052.88 2106.34 3059.38 ;
     RECT  2106.34 3053.3 2109.7 3059.38 ;
     RECT  2109.7 3053.3 2110.18 3053.5 ;
     RECT  2021 0 2145 178 ;
     RECT  2031 3222 2155 3400 ;
     RECT  1769.38 2078.48 2168.74 2078.68 ;
     RECT  2091.94 1877.3 2172.1 1877.5 ;
     RECT  1803.26 1425.8 2200.42 1454.12 ;
     RECT  2077.06 1736.16 2210.02 1743.94 ;
     RECT  2145 -70 2215 178 ;
     RECT  2155 3222 2225 3470 ;
     RECT  1977.7 2020.52 2315.42 2023.24 ;
     RECT  1977.7 2033.96 2315.42 2034.16 ;
     RECT  2215 0 2339 178 ;
     RECT  1824.58 1894.94 2341.82 1911.52 ;
     RECT  2225 3222 2349 3400 ;
     RECT  1779.46 1923.92 2354.3 1927.48 ;
     RECT  1797.98 1942.4 2354.3 1963.18 ;
     RECT  1797.98 2064.62 2354.3 2069.44 ;
     RECT  1754.5 2111.66 2354.3 2111.86 ;
     RECT  2354.3 1923.92 2355.94 1963.18 ;
     RECT  2354.3 2111.66 2356.7 2116.88 ;
     RECT  1955.14 2243.96 2357.66 2264.32 ;
     RECT  2354.3 2064.62 2358.14 2071.96 ;
     RECT  1807.1 1638.3 2358.34 1675.48 ;
     RECT  2315.42 2020.52 2358.62 2034.16 ;
     RECT  2358.14 2060.4 2359.1 2071.96 ;
     RECT  2341.82 1894.08 2361.02 1911.52 ;
     RECT  1666.46 2653.04 2362.66 2653.24 ;
     RECT  2361.5 2044.86 2362.94 2045.06 ;
     RECT  2355.94 1923.92 2363.14 1955.2 ;
     RECT  2358.62 2020.1 2364.86 2034.16 ;
     RECT  2356.7 2111.66 2365.54 2120.66 ;
     RECT  1749.7 2133.5 2365.54 2135.38 ;
     RECT  2365.54 2120.46 2366.78 2120.66 ;
     RECT  1783.58 1985.66 2367.26 1993 ;
     RECT  1746.82 2204.48 2367.74 2204.68 ;
     RECT  2364.86 1869.72 2367.94 1869.92 ;
     RECT  2362.94 2044.86 2367.94 2049.26 ;
     RECT  1803.26 1471.56 2368.7 1515.04 ;
     RECT  2361.02 1890.72 2368.7 1911.52 ;
     RECT  2359.1 2060.4 2368.7 2072.38 ;
     RECT  2368.22 2082.66 2368.7 2082.86 ;
     RECT  2368.7 1886.52 2369.18 1911.52 ;
     RECT  2366.78 2120.46 2369.18 2124.44 ;
     RECT  2365.54 2133.5 2369.18 2133.7 ;
     RECT  1791.74 2163.74 2370.14 2173.18 ;
     RECT  2361.98 1841.16 2371.1 1841.36 ;
     RECT  2364.38 1855.86 2371.58 1860.26 ;
     RECT  2363.14 1923.92 2371.58 1932.5 ;
     RECT  2369.18 2120.46 2371.78 2133.7 ;
     RECT  2357.66 2241.44 2372.26 2264.32 ;
     RECT  2371.58 1922.22 2373.02 1932.5 ;
     RECT  2368.7 2060.4 2373.7 2086.22 ;
     RECT  2373.7 2086.02 2373.98 2086.22 ;
     RECT  2369.66 1965.48 2374.46 1965.68 ;
     RECT  2367.26 1981.02 2374.46 1993 ;
     RECT  1798.46 2220.86 2374.94 2231.98 ;
     RECT  2373.98 2086.02 2375.42 2088.32 ;
     RECT  2375.42 2086.02 2375.9 2091.68 ;
     RECT  2354.3 2101.98 2375.9 2102.18 ;
     RECT  2365.54 2111.66 2375.9 2111.86 ;
     RECT  2369.18 1885.68 2376.38 1911.52 ;
     RECT  2364.38 1818.9 2376.86 1819.1 ;
     RECT  2362.94 1829.4 2376.86 1829.6 ;
     RECT  2371.1 1841.16 2376.86 1841.78 ;
     RECT  2373.02 1921.8 2376.86 1932.5 ;
     RECT  2363.14 1941.96 2376.86 1955.2 ;
     RECT  2374.46 1965.48 2377.06 1993 ;
     RECT  2376.86 1818.48 2377.34 1819.1 ;
     RECT  2005.54 2008.34 2378.3 2008.54 ;
     RECT  2376.38 1881.9 2378.78 1911.52 ;
     RECT  2376.86 1921.8 2378.78 1955.2 ;
     RECT  2375.9 2086.02 2378.78 2092.52 ;
     RECT  2367.94 2044.86 2378.98 2045.48 ;
     RECT  2371.78 2123.82 2380.22 2133.7 ;
     RECT  2380.22 2123.4 2382.14 2133.7 ;
     RECT  2370.14 2188.5 2382.34 2188.7 ;
     RECT  2373.7 2060.4 2382.62 2072.38 ;
     RECT  2377.34 1814.28 2384.06 1819.1 ;
     RECT  2376.86 1829.4 2384.06 1841.78 ;
     RECT  2370.14 2163.74 2384.06 2177.36 ;
     RECT  2384.06 1814.28 2384.26 1841.78 ;
     RECT  2374.94 2220.86 2384.74 2234.06 ;
     RECT  2378.3 2150.7 2385.02 2150.9 ;
     RECT  2384.06 2163.74 2385.02 2181.98 ;
     RECT  2371.58 1852.5 2385.22 1860.26 ;
     RECT  2374.94 1870.98 2385.5 1871.18 ;
     RECT  2382.62 2056.62 2386.46 2072.38 ;
     RECT  2385.5 1870.98 2387.42 1871.6 ;
     RECT  2378.78 1881.9 2387.42 1955.2 ;
     RECT  2386.46 2056.2 2389.34 2072.38 ;
     RECT  2375.9 2101.98 2389.54 2111.86 ;
     RECT  2378.98 2045.28 2390.02 2045.48 ;
     RECT  2367.74 2201.94 2390.5 2204.68 ;
     RECT  2385.22 1852.5 2390.98 1856.48 ;
     RECT  2387.42 1870.98 2391.94 1955.2 ;
     RECT  2382.14 2120.88 2391.94 2133.7 ;
     RECT  2389.34 2056.2 2392.42 2075.3 ;
     RECT  2392.42 2056.2 2392.7 2072.38 ;
     RECT  2391.94 1871.4 2393.38 1955.2 ;
     RECT  2393.38 1873.92 2393.86 1955.2 ;
     RECT  2200.42 1445.12 2394.34 1454.12 ;
     RECT  2391.94 2122.98 2396.26 2133.7 ;
     RECT  2390.98 1855.86 2397.5 1856.48 ;
     RECT  2384.26 1837.8 2399.9 1841.78 ;
     RECT  2377.06 1973.04 2399.9 1973.24 ;
     RECT  2377.06 1984.38 2399.9 1993 ;
     RECT  2378.3 2007.48 2400.1 2008.54 ;
     RECT  2384.26 1814.28 2400.86 1822.04 ;
     RECT  2389.54 2103.68 2400.86 2111.86 ;
     RECT  2399.9 1973.04 2402.02 1993 ;
     RECT  2384.74 2220.86 2402.3 2231.98 ;
     RECT  2393.86 1873.92 2404.7 1951.4 ;
     RECT  2402.02 1973.04 2404.7 1976.18 ;
     RECT  2390.78 2192.28 2404.7 2192.48 ;
     RECT  2390.5 2201.94 2404.7 2202.14 ;
     RECT  2402.3 2214.54 2404.7 2231.98 ;
     RECT  2404.7 1873.92 2404.9 1976.18 ;
     RECT  2392.7 2052.84 2404.9 2072.38 ;
     RECT  2385.02 2150.7 2404.9 2181.98 ;
     RECT  2404.9 2052.84 2405.18 2070.28 ;
     RECT  2404.9 1905.86 2405.38 1976.18 ;
     RECT  2404.7 2192.28 2406.14 2193.32 ;
     RECT  2404.7 2201.94 2406.14 2231.98 ;
     RECT  2405.38 1965.48 2406.34 1976.18 ;
     RECT  2406.14 2192.28 2407.1 2231.98 ;
     RECT  2399.9 1835.28 2407.78 1841.78 ;
     RECT  2378.78 2086.02 2408.06 2093.36 ;
     RECT  2400.86 2103.26 2408.06 2111.86 ;
     RECT  2077.06 1685.76 2408.54 1723.34 ;
     RECT  2210.02 1736.16 2408.54 1736.36 ;
     RECT  2405.18 2050.32 2408.54 2070.28 ;
     RECT  2339 -70 2409 178 ;
     RECT  2402.02 1984.8 2409.02 1993 ;
     RECT  2400.1 2007.92 2409.02 2008.54 ;
     RECT  2408.06 2086.02 2409.5 2111.86 ;
     RECT  2404.9 2162.04 2409.5 2181.98 ;
     RECT  2407.1 2192.28 2409.5 2234.48 ;
     RECT  2408.54 1685.76 2409.7 1736.36 ;
     RECT  2372.26 2243.96 2411.9 2264.32 ;
     RECT  2400.86 1814.28 2413.34 1826.24 ;
     RECT  2407.78 1835.28 2413.34 1840.1 ;
     RECT  2409.02 1984.8 2413.34 2008.54 ;
     RECT  2413.34 1981.86 2415.26 2008.54 ;
     RECT  2364.86 2017.16 2415.26 2034.16 ;
     RECT  2404.9 2150.7 2415.26 2150.9 ;
     RECT  2409.5 2162.04 2415.26 2234.48 ;
     RECT  2396.26 2122.98 2415.46 2124.44 ;
     RECT  2411.9 2243.96 2415.74 2264.74 ;
     RECT  2397.5 1855.86 2416.22 1859 ;
     RECT  2416.22 1855.02 2417.18 1859 ;
     RECT  2415.26 2150.7 2417.18 2234.48 ;
     RECT  2413.34 1814.28 2418.62 1840.1 ;
     RECT  2349 3222 2419 3470 ;
     RECT  2418.62 1814.28 2419.1 1840.94 ;
     RECT  2404.9 1873.92 2419.1 1894.28 ;
     RECT  2405.38 1905.86 2419.1 1954.76 ;
     RECT  2417.18 2143.56 2420.54 2234.48 ;
     RECT  2415.74 2243.12 2420.54 2264.74 ;
     RECT  2200.42 1425.8 2423.42 1436.06 ;
     RECT  2394.34 1445.54 2423.42 1454.12 ;
     RECT  2420.54 2143.56 2423.9 2264.74 ;
     RECT  2419.1 1873.92 2424.1 1954.76 ;
     RECT  2417.18 1854.6 2424.38 1859 ;
     RECT  2424.38 1854.6 2424.58 1863.62 ;
     RECT  2409.7 1685.76 2424.86 1723.34 ;
     RECT  2396.26 2133.5 2424.86 2133.7 ;
     RECT  2423.9 2142.3 2424.86 2264.74 ;
     RECT  2406.34 1965.48 2425.34 1973.24 ;
     RECT  2415.26 1981.86 2425.34 2034.16 ;
     RECT  2419.1 1814.28 2425.82 1841.36 ;
     RECT  2409.5 2084.76 2425.82 2111.86 ;
     RECT  2415.46 2124.24 2425.82 2124.44 ;
     RECT  2406.62 1750.44 2426.3 1750.64 ;
     RECT  2424.1 1905.86 2426.98 1954.76 ;
     RECT  2419.58 1784.04 2427.74 1784.24 ;
     RECT  2424.86 1685.76 2429.38 1727.54 ;
     RECT  2407.58 1765.98 2429.66 1766.18 ;
     RECT  2358.34 1638.3 2430.14 1672.12 ;
     RECT  2429.38 1685.76 2430.14 1723.34 ;
     RECT  2426.3 1746.24 2431.1 1750.64 ;
     RECT  2408.54 2044.02 2431.1 2070.28 ;
     RECT  2425.82 2084.76 2431.1 2124.44 ;
     RECT  2427.74 1784.04 2431.58 1791.8 ;
     RECT  2426.98 1905.86 2432.26 1939.64 ;
     RECT  2431.1 1746.24 2432.54 1752.32 ;
     RECT  2429.66 1765.14 2432.54 1766.18 ;
     RECT  2425.34 1965.48 2432.54 2034.16 ;
     RECT  2431.1 2044.02 2432.54 2072.78 ;
     RECT  2431.1 2082.66 2432.54 2124.44 ;
     RECT  2424.1 1873.92 2432.74 1894.28 ;
     RECT  2432.54 1746.24 2433.02 1766.18 ;
     RECT  2433.02 1746.24 2433.5 1769.12 ;
     RECT  2431.58 1783.62 2433.5 1791.8 ;
     RECT  2433.5 1746.24 2433.98 1791.8 ;
     RECT  2426.98 1950.78 2434.18 1954.76 ;
     RECT  2424.58 1855.44 2434.46 1863.62 ;
     RECT  2432.74 1873.92 2434.46 1890.08 ;
     RECT  2425.82 1813.86 2434.94 1841.36 ;
     RECT  2434.46 1855.44 2434.94 1890.08 ;
     RECT  2433.98 1746.24 2436.86 1796 ;
     RECT  2424.86 2133.5 2437.54 2264.74 ;
     RECT  2430.14 1638.3 2439.94 1723.34 ;
     RECT  2434.94 1813.86 2440.42 1890.08 ;
     RECT  2436.86 1746.24 2440.7 1796.42 ;
     RECT  2439.94 1638.3 2440.9 1675.06 ;
     RECT  2432.26 1905.86 2441.66 1934.6 ;
     RECT  2440.7 1746.24 2446.46 1798.1 ;
     RECT  2446.46 1746.24 2446.66 1803.56 ;
     RECT  2441.66 1905.86 2447.42 1935.86 ;
     RECT  2434.18 1950.78 2447.42 1951.4 ;
     RECT  2437.54 2138.52 2447.62 2264.74 ;
     RECT  2447.42 1905.86 2448.86 1951.4 ;
     RECT  2432.54 1965.06 2448.86 2034.16 ;
     RECT  2448.86 1905.86 2449.06 2034.16 ;
     RECT  2446.66 1759.68 2450.02 1803.56 ;
     RECT  2432.54 2044.02 2450.3 2124.44 ;
     RECT  2439.94 1685.76 2451.26 1723.34 ;
     RECT  2409.7 1736.16 2451.26 1736.36 ;
     RECT  2449.06 1905.86 2453.38 1985 ;
     RECT  2450.3 2044.02 2453.86 2128.22 ;
     RECT  2440.9 1638.3 2455.1 1660.76 ;
     RECT  2440.9 1670.64 2455.1 1675.06 ;
     RECT  2453.86 2044.02 2455.1 2093.78 ;
     RECT  2451.26 1685.76 2455.3 1736.36 ;
     RECT  2447.62 2138.52 2455.3 2211.8 ;
     RECT  2447.62 2222.52 2455.3 2264.74 ;
     RECT  2450.02 1759.68 2455.58 1793.48 ;
     RECT  2423.42 1425.8 2457.02 1454.12 ;
     RECT  2368.7 1464.86 2457.02 1515.04 ;
     RECT  2455.58 1758 2457.02 1793.48 ;
     RECT  2457.02 1425.8 2457.22 1515.04 ;
     RECT  2453.86 2103.26 2457.22 2128.22 ;
     RECT  2455.3 2201.94 2457.5 2211.8 ;
     RECT  2455.3 2222.52 2457.5 2224.84 ;
     RECT  2457.02 1757.58 2458.94 1793.48 ;
     RECT  2450.02 1803.36 2458.94 1803.56 ;
     RECT  2457.22 2115.84 2461.34 2128.22 ;
     RECT  2455.3 2138.52 2461.34 2192.48 ;
     RECT  2453.38 1965.06 2461.82 1985 ;
     RECT  2449.06 1994.88 2461.82 2034.16 ;
     RECT  2453.38 1905.86 2463.46 1951.4 ;
     RECT  2458.94 1757.58 2463.74 1803.56 ;
     RECT  2463.46 1916.76 2463.74 1951.4 ;
     RECT  2455.3 2234.28 2463.94 2264.74 ;
     RECT  2457.22 1425.8 2464.42 1456.66 ;
     RECT  2440.42 1814.28 2465.86 1890.08 ;
     RECT  2461.82 1965.06 2466.14 2034.16 ;
     RECT  2455.3 1736.16 2467.1 1736.36 ;
     RECT  2457.22 2103.26 2467.1 2105.96 ;
     RECT  2461.34 2115.84 2467.1 2192.48 ;
     RECT  2455.1 2043.6 2467.58 2093.78 ;
     RECT  2467.1 2103.26 2467.58 2192.48 ;
     RECT  2463.74 1757.58 2468.26 1803.98 ;
     RECT  2455.3 1685.76 2468.54 1723.76 ;
     RECT  2467.1 1736.16 2468.54 1743.08 ;
     RECT  2467.58 2043.6 2469.7 2192.48 ;
     RECT  2463.94 2237.64 2469.7 2264.74 ;
     RECT  2468.54 1685.76 2470.18 1743.08 ;
     RECT  2466.14 1962.54 2470.46 2034.16 ;
     RECT  2465.86 1818.48 2471.14 1890.08 ;
     RECT  2463.46 1905.86 2472.86 1906.48 ;
     RECT  2470.46 1962.12 2473.06 2034.16 ;
     RECT  2473.06 1962.12 2474.5 2034.14 ;
     RECT  2472.86 1905.86 2474.78 1907.3 ;
     RECT  2463.74 1916.76 2474.78 1951.82 ;
     RECT  2470.18 1685.76 2474.98 1736.36 ;
     RECT  2471.14 1818.48 2476.42 1864.46 ;
     RECT  2474.98 1685.76 2477.38 1723.76 ;
     RECT  2474.78 1905.86 2479.1 1951.82 ;
     RECT  2474.5 1994.88 2479.3 2034.14 ;
     RECT  2479.3 2019.26 2481.98 2034.14 ;
     RECT  2469.7 2043.6 2481.98 2104.72 ;
     RECT  2468.26 1760.52 2484.58 1803.98 ;
     RECT  2481.98 2019.26 2484.58 2104.72 ;
     RECT  2476.42 1825.62 2485.06 1864.46 ;
     RECT  2469.7 2241.42 2485.54 2264.74 ;
     RECT  2479.1 1899.12 2486.78 1951.82 ;
     RECT  2474.5 1962.12 2486.78 1983.74 ;
     RECT  2484.58 1760.52 2487.74 1803.56 ;
     RECT  2479.3 1994.88 2487.74 2010.2 ;
     RECT  2455.1 1638.3 2489.18 1675.06 ;
     RECT  2477.38 1685.76 2489.18 1723.34 ;
     RECT  2469.7 2113.32 2489.86 2192.48 ;
     RECT  2487.74 1758 2491.3 1803.56 ;
     RECT  2486.78 1899.12 2491.78 1983.74 ;
     RECT  2489.86 2138.52 2492.06 2192.48 ;
     RECT  2457.5 2201.94 2492.06 2224.84 ;
     RECT  2491.78 1899.12 2492.26 1951.4 ;
     RECT  2489.18 1638.3 2493.22 1723.34 ;
     RECT  2487.74 1994.04 2493.5 2010.2 ;
     RECT  2484.58 2019.26 2495.14 2058.08 ;
     RECT  2493.22 1638.3 2496.1 1675.06 ;
     RECT  2485.06 1825.62 2498.3 1829.6 ;
     RECT  2485.06 1844.52 2498.3 1864.46 ;
     RECT  2489.86 2113.32 2498.3 2124.44 ;
     RECT  2496.1 1660.56 2499.46 1675.06 ;
     RECT  2471.14 1873.92 2500.22 1890.08 ;
     RECT  2491.3 1760.52 2501.66 1803.56 ;
     RECT  2493.98 1813.44 2501.66 1813.64 ;
     RECT  2500.22 1873.92 2501.86 1896.38 ;
     RECT  2492.26 1905.86 2501.86 1951.4 ;
     RECT  2501.86 1906.28 2502.34 1951.4 ;
     RECT  2502.34 1924.32 2502.62 1951.4 ;
     RECT  2491.78 1961.28 2502.62 1983.74 ;
     RECT  2502.62 1924.32 2502.82 1983.74 ;
     RECT  2492.06 2138.52 2504.54 2224.84 ;
     RECT  2493.22 1685.76 2505.5 1723.34 ;
     RECT  2495.14 2019.26 2505.5 2031.62 ;
     RECT  2495.14 2041.08 2505.5 2058.08 ;
     RECT  2484.58 2069.24 2505.5 2104.72 ;
     RECT  2498.3 2113.32 2505.5 2126.96 ;
     RECT  2504.54 2136 2505.5 2224.84 ;
     RECT  2505.5 2018.84 2505.7 2031.62 ;
     RECT  2498.3 1825.62 2505.98 1864.46 ;
     RECT  2501.86 1873.92 2505.98 1890.08 ;
     RECT  2505.5 2041.08 2506.46 2058.92 ;
     RECT  2505.5 2069.24 2506.46 2224.84 ;
     RECT  2506.46 2041.08 2507.14 2224.84 ;
     RECT  2501.66 1760.52 2508.38 1813.64 ;
     RECT  2508.38 1755.06 2509.06 1813.64 ;
     RECT  2502.34 1906.28 2509.06 1915.7 ;
     RECT  2509.06 1764.72 2510.3 1813.64 ;
     RECT  2505.98 1825.62 2510.3 1890.08 ;
     RECT  2502.82 1934.4 2512.7 1983.74 ;
     RECT  2493.5 1992.36 2512.7 2010.2 ;
     RECT  2509.06 1908.36 2515.1 1915.7 ;
     RECT  2502.82 1924.32 2515.1 1924.52 ;
     RECT  2496.1 1638.3 2516.06 1650.68 ;
     RECT  2499.46 1660.56 2516.06 1660.76 ;
     RECT  2510.3 1764.72 2516.06 1890.08 ;
     RECT  2515.1 1908.36 2516.06 1924.52 ;
     RECT  2512.7 1934.4 2516.06 2010.2 ;
     RECT  2516.06 1764.72 2516.54 1897.22 ;
     RECT  2516.06 1908.36 2518.18 2010.2 ;
     RECT  2505.7 2018.84 2518.66 2030.36 ;
     RECT  2507.14 2041.08 2518.66 2126.96 ;
     RECT  2509.06 1755.06 2518.94 1755.26 ;
     RECT  2516.54 1764.72 2518.94 1897.64 ;
     RECT  2505.5 1685.76 2519.9 1727.54 ;
     RECT  2474.98 1736.16 2519.9 1736.36 ;
     RECT  2518.94 1755.06 2521.82 1897.64 ;
     RECT  2519.9 1685.76 2522.3 1743.08 ;
     RECT  2521.82 1753.8 2522.3 1897.64 ;
     RECT  2518.18 1908.36 2522.3 1924.52 ;
     RECT  2522.3 1685.76 2522.5 1924.52 ;
     RECT  2518.66 2070.48 2524.9 2126.96 ;
     RECT  2522.5 1873.92 2527.1 1924.52 ;
     RECT  2518.18 1934.4 2527.1 2010.2 ;
     RECT  2524.9 2115.84 2528.06 2126.96 ;
     RECT  2507.14 2136 2528.06 2224.84 ;
     RECT  1807.1 1622.76 2531.14 1628 ;
     RECT  2409 0 2533 178 ;
     RECT  2518.66 2018.84 2533.82 2029.94 ;
     RECT  2518.66 2041.08 2533.82 2058.92 ;
     RECT  2524.9 2070.48 2534.3 2105.96 ;
     RECT  2528.06 2115.84 2534.3 2224.84 ;
     RECT  2534.3 2070.48 2537.18 2224.84 ;
     RECT  2533.82 2018.84 2537.38 2058.92 ;
     RECT  2527.1 1873.92 2539.3 2010.2 ;
     RECT  2537.18 2068.8 2539.58 2224.84 ;
     RECT  2539.58 2068.8 2541.7 2230.7 ;
     RECT  2539.3 1873.92 2542.18 2008.54 ;
     RECT  2537.38 2031.84 2542.66 2058.92 ;
     RECT  2419 3222 2543 3400 ;
     RECT  2522.5 1685.76 2544.86 1864.46 ;
     RECT  2537.38 2018.84 2545.54 2022.8 ;
     RECT  2516.06 1638.3 2546.02 1660.76 ;
     RECT  2541.7 2071.32 2546.78 2230.7 ;
     RECT  2546.02 1660.56 2547.26 1660.76 ;
     RECT  2499.46 1670.64 2547.26 1675.06 ;
     RECT  2542.66 2031.84 2547.26 2058.08 ;
     RECT  2542.18 1873.92 2547.46 1903.1 ;
     RECT  2531.14 1622.76 2547.74 1626.32 ;
     RECT  2546.02 1638.3 2547.74 1650.68 ;
     RECT  2544.86 1685.34 2548.22 1864.46 ;
     RECT  2547.46 1873.92 2548.22 1889.66 ;
     RECT  2547.26 1660.56 2549.38 1675.06 ;
     RECT  2547.26 2031 2549.38 2058.08 ;
     RECT  2546.78 2071.32 2550.34 2234.48 ;
     RECT  2542.18 1912.98 2553.22 2008.54 ;
     RECT  2550.34 2234.28 2553.5 2234.48 ;
     RECT  2485.54 2243.12 2553.5 2264.74 ;
     RECT  2547.74 1622.76 2554.18 1650.68 ;
     RECT  2553.22 2007.92 2554.46 2008.54 ;
     RECT  2545.54 2018.84 2554.46 2021.98 ;
     RECT  2548.22 1685.34 2555.14 1889.66 ;
     RECT  2549.38 1670.64 2555.9 1675.06 ;
     RECT  2547.46 1902.9 2555.9 1903.1 ;
     RECT  2553.22 1912.98 2555.9 1998.44 ;
     RECT  2550.34 2071.32 2556.1 2224.84 ;
     RECT  1753.82 2361.14 2556.58 2379.82 ;
     RECT  2555.9 1670.64 2557.34 1675.48 ;
     RECT  2555.14 1685.34 2557.34 1864.46 ;
     RECT  2555.14 1873.92 2559.26 1889.66 ;
     RECT  1629.02 2724.86 2559.94 2725.06 ;
     RECT  2557.34 1670.64 2560.9 1864.46 ;
     RECT  2559.26 1873.92 2561.18 1890.92 ;
     RECT  2555.9 1902.9 2561.18 1998.44 ;
     RECT  2554.46 2007.92 2563.1 2021.98 ;
     RECT  2549.38 2031.84 2563.1 2058.08 ;
     RECT  2561.18 1873.92 2563.58 1998.44 ;
     RECT  2563.1 2007.92 2563.58 2058.08 ;
     RECT  2556.1 2071.32 2565.02 2158.46 ;
     RECT  2556.1 2167.52 2565.02 2224.84 ;
     RECT  2560.9 1685.76 2568.38 1864.46 ;
     RECT  2563.58 1873.92 2568.38 2058.08 ;
     RECT  2568.38 1685.76 2571.94 2058.08 ;
     RECT  2571.94 1907.94 2577.02 2058.08 ;
     RECT  2565.02 2071.32 2577.02 2224.84 ;
     RECT  2577.02 1907.94 2579.9 2224.84 ;
     RECT  2553.5 2234.28 2579.9 2264.74 ;
     RECT  2560.9 1670.64 2587.1 1675.48 ;
     RECT  2571.94 1685.76 2587.1 1897.64 ;
     RECT  2464.42 1425.8 2588.26 1454.12 ;
     RECT  2587.1 1670.64 2596.9 1897.64 ;
     RECT  2579.9 1907.94 2597.86 2264.74 ;
     RECT  2596.9 1670.64 2598.34 1864.46 ;
     RECT  2598.34 1670.64 2599.3 1751.48 ;
     RECT  2597.86 1907.94 2600.26 2058.92 ;
     RECT  2599.3 1670.64 2600.54 1749.4 ;
     RECT  2598.34 1760.94 2601.7 1864.46 ;
     RECT  2533 -70 2603 178 ;
     RECT  1803.26 1524.08 2603.14 1583.9 ;
     RECT  2596.9 1873.92 2604.38 1897.64 ;
     RECT  2600.26 1907.94 2604.38 1998.44 ;
     RECT  2597.86 2071.32 2606.5 2264.74 ;
     RECT  2606.5 2071.32 2608.22 2224.84 ;
     RECT  2604.38 1873.92 2608.42 1998.44 ;
     RECT  2608.42 1873.92 2609.38 1951.82 ;
     RECT  2600.54 1669.8 2609.86 1749.4 ;
     RECT  2609.38 1950.78 2610.82 1951.82 ;
     RECT  2606.5 2234.28 2611.78 2264.74 ;
     RECT  2554.18 1622.76 2612.06 1626.32 ;
     RECT  2601.7 1761.78 2612.06 1864.46 ;
     RECT  2609.38 1873.92 2612.06 1942.16 ;
     RECT  2608.22 2070.9 2612.26 2224.84 ;
     RECT  2543 3222 2613 3470 ;
     RECT  2609.86 1669.8 2613.22 1670.84 ;
     RECT  2612.26 2108.7 2613.22 2224.84 ;
     RECT  2609.86 1685.76 2613.5 1749.4 ;
     RECT  2612.06 1761.78 2613.5 1942.16 ;
     RECT  2611.78 2235.54 2614.18 2264.74 ;
     RECT  2600.26 2010 2615.42 2058.92 ;
     RECT  2614.18 2236.8 2615.62 2264.74 ;
     RECT  2613.5 1685.76 2617.54 1942.16 ;
     RECT  2613.22 1670.64 2618.3 1670.84 ;
     RECT  2617.54 1685.76 2618.3 1864.46 ;
     RECT  2610.82 1950.78 2620.22 1950.98 ;
     RECT  2608.42 1961.28 2620.22 1998.44 ;
     RECT  2612.26 2070.9 2620.7 2098.84 ;
     RECT  2613.22 2108.7 2620.7 2181.14 ;
     RECT  2615.42 2010 2623.58 2060.6 ;
     RECT  2620.7 2070.9 2623.58 2181.14 ;
     RECT  2603.14 1565.66 2624.26 1583.9 ;
     RECT  2617.54 1873.92 2624.74 1942.16 ;
     RECT  2623.58 2008.74 2628.1 2060.6 ;
     RECT  2549.38 1660.56 2630.78 1660.76 ;
     RECT  2618.3 1670.64 2630.78 1864.46 ;
     RECT  2624.74 1873.92 2630.78 1938.8 ;
     RECT  2624.26 1566.92 2631.46 1583.9 ;
     RECT  2603.14 1524.08 2631.94 1554.92 ;
     RECT  2623.58 2070.9 2633.38 2181.56 ;
     RECT  2628.1 2008.74 2634.14 2058.08 ;
     RECT  2630.78 1660.56 2634.62 1938.8 ;
     RECT  2634.14 2008.32 2634.82 2058.08 ;
     RECT  2634.82 2033.1 2637.98 2058.08 ;
     RECT  2634.82 2008.32 2638.66 2023.24 ;
     RECT  2634.62 1660.56 2638.94 1939.22 ;
     RECT  2638.94 1660.56 2640.1 1940.48 ;
     RECT  2633.38 2109.12 2641.34 2181.56 ;
     RECT  2613.22 2191.44 2641.34 2224.84 ;
     RECT  2620.22 1950.78 2642.02 1998.44 ;
     RECT  1801.06 1396.4 2642.3 1416.76 ;
     RECT  2588.26 1429.16 2642.3 1454.12 ;
     RECT  2637.98 2033.1 2642.98 2060.6 ;
     RECT  2612.06 1620.66 2643.74 1626.32 ;
     RECT  2554.18 1638.3 2643.74 1650.68 ;
     RECT  2643.74 1620.66 2644.22 1650.68 ;
     RECT  2640.1 1660.56 2644.22 1938.82 ;
     RECT  2644.22 1620.66 2644.42 1938.82 ;
     RECT  2631.94 1524.5 2645.86 1554.92 ;
     RECT  2644.42 1901.64 2645.86 1938.82 ;
     RECT  2633.38 2070.9 2645.86 2098.84 ;
     RECT  2642.98 2036.46 2646.14 2060.6 ;
     RECT  2645.86 2071.32 2646.62 2098.84 ;
     RECT  2641.34 2109.12 2646.62 2224.84 ;
     RECT  2644.42 1620.66 2649.5 1889.66 ;
     RECT  2649.5 1618.56 2649.7 1889.66 ;
     RECT  2646.14 2036.46 2649.7 2061.02 ;
     RECT  2649.7 2040.24 2650.66 2061.02 ;
     RECT  2645.86 1524.92 2656.7 1554.92 ;
     RECT  1803.26 1597.56 2656.7 1607.84 ;
     RECT  2649.7 1618.56 2656.7 1889.24 ;
     RECT  2645.86 1901.64 2656.7 1938.38 ;
     RECT  2638.66 2008.32 2656.7 2022.8 ;
     RECT  2631.46 1569.42 2657.18 1583.9 ;
     RECT  2656.7 1597.56 2657.18 1889.24 ;
     RECT  2457.22 1471.56 2657.66 1515.04 ;
     RECT  2642.02 1953.74 2657.86 1998.44 ;
     RECT  2656.7 1524.92 2659.1 1557.02 ;
     RECT  2656.7 2007.9 2659.3 2022.8 ;
     RECT  2659.1 1524.92 2660.06 1557.44 ;
     RECT  2657.18 1569 2660.06 1583.9 ;
     RECT  2657.18 1593.78 2660.26 1889.24 ;
     RECT  2650.66 2040.24 2660.54 2060.6 ;
     RECT  2646.62 2071.32 2660.54 2224.84 ;
     RECT  2657.66 1471.56 2661.02 1515.86 ;
     RECT  2660.06 1524.92 2661.02 1583.9 ;
     RECT  2660.26 1593.78 2661.02 1691 ;
     RECT  2660.26 1701.3 2661.7 1889.24 ;
     RECT  2661.7 1851.24 2661.98 1889.24 ;
     RECT  2656.7 1901.64 2661.98 1945.1 ;
     RECT  2660.54 2040.24 2663.9 2224.84 ;
     RECT  2661.02 1471.56 2664.1 1691 ;
     RECT  2663.9 2033.52 2664.1 2224.84 ;
     RECT  2659.3 2007.9 2666.98 2015.66 ;
     RECT  2661.98 1851.24 2669.18 1945.1 ;
     RECT  2657.86 1954.14 2669.18 1998.44 ;
     RECT  2669.18 1851.24 2670.14 1998.44 ;
     RECT  2666.98 2007.9 2670.14 2014.82 ;
     RECT  2670.14 1851.24 2671.58 2014.82 ;
     RECT  2664.1 2033.52 2672.54 2116.04 ;
     RECT  2664.1 2125.08 2672.54 2224.84 ;
     RECT  2661.7 1701.3 2673.02 1841.78 ;
     RECT  2671.58 1850.82 2673.02 2014.82 ;
     RECT  2642.3 1396.4 2678.02 1454.12 ;
     RECT  2664.1 1593.78 2678.3 1691 ;
     RECT  2673.02 1701.3 2678.3 2014.82 ;
     RECT  2664.1 1471.56 2678.78 1583.9 ;
     RECT  2678.3 1593.78 2678.78 2014.82 ;
     RECT  2678.78 1471.56 2678.98 2014.82 ;
     RECT  2678.98 1471.56 2679.74 1527.2 ;
     RECT  2678.98 1539.6 2679.74 2014.82 ;
     RECT  2679.74 1539.6 2681.18 2021.54 ;
     RECT  2672.54 2033.52 2681.18 2224.84 ;
     RECT  2679.74 1466.52 2681.66 1527.2 ;
     RECT  2681.18 1539.6 2683.3 2224.84 ;
     RECT  2683.3 1951.2 2684.74 2224.84 ;
     RECT  2678.02 1396.4 2685.5 1420.54 ;
     RECT  2678.02 1429.16 2685.7 1454.12 ;
     RECT  2684.74 1954.14 2685.7 2224.84 ;
     RECT  2685.7 1435.86 2687.42 1454.12 ;
     RECT  2681.66 1464 2687.42 1527.2 ;
     RECT  2685.7 1954.14 2690.98 2184.92 ;
     RECT  2685.7 2196.9 2690.98 2224.84 ;
     RECT  2687.42 1435.86 2691.26 1527.2 ;
     RECT  2683.3 1539.6 2692.22 1938.38 ;
     RECT  2690.98 1954.14 2693.38 1981.64 ;
     RECT  2691.26 1435.86 2696.26 1528.88 ;
     RECT  2696.26 1471.56 2699.62 1528.88 ;
     RECT  2690.98 1991.94 2701.06 2184.92 ;
     RECT  2696.26 1435.86 2702.02 1462.94 ;
     RECT  2692.22 1537.92 2702.02 1938.38 ;
     RECT  2702.02 1537.92 2703.94 1890.08 ;
     RECT  2702.02 1901.64 2704.7 1938.38 ;
     RECT  2693.38 1954.14 2706.62 1980.8 ;
     RECT  2701.06 2115.84 2707.1 2184.92 ;
     RECT  2690.98 2196.9 2707.1 2203 ;
     RECT  2707.1 2115.84 2707.3 2203 ;
     RECT  2704.7 1901.64 2708.54 1939.64 ;
     RECT  2702.02 1462.74 2709.02 1462.94 ;
     RECT  2699.62 1471.56 2709.02 1527.2 ;
     RECT  2707.3 2127.18 2711.62 2203 ;
     RECT  2702.02 1435.86 2715.26 1454.12 ;
     RECT  2709.02 1462.74 2715.26 1527.2 ;
     RECT  2706.62 1949.94 2715.46 1980.8 ;
     RECT  2711.62 2127.18 2715.74 2181.56 ;
     RECT  2685.5 1389.26 2716.22 1420.54 ;
     RECT  2715.26 1435.86 2716.22 1527.2 ;
     RECT  2716.22 1389.26 2716.9 1527.2 ;
     RECT  2708.54 1901.64 2718.62 1941.32 ;
     RECT  2718.62 1901.64 2719.3 1948.46 ;
     RECT  2711.62 2192.28 2720.54 2203 ;
     RECT  2690.98 2211.62 2720.54 2224.84 ;
     RECT  2715.74 2126.76 2720.74 2181.56 ;
     RECT  2715.46 1957.08 2721.5 1980.8 ;
     RECT  2720.54 2192.28 2721.7 2224.84 ;
     RECT  2701.06 1991.94 2723.42 2105.96 ;
     RECT  2721.5 1957.08 2723.62 1981.64 ;
     RECT  2719.3 1902.06 2723.9 1948.46 ;
     RECT  2720.74 2127.18 2723.9 2181.56 ;
     RECT  2723.9 1902.06 2725.54 1950.14 ;
     RECT  2723.42 1991.52 2725.82 2105.96 ;
     RECT  2707.3 2115.84 2725.82 2118.14 ;
     RECT  2603 0 2727 178 ;
     RECT  2725.82 1991.52 2727.46 2118.14 ;
     RECT  2725.54 1902.06 2729.38 1948.46 ;
     RECT  2729.38 1902.06 2729.86 1941.32 ;
     RECT  2727.46 1991.94 2730.34 2118.14 ;
     RECT  2730.34 2115.84 2730.62 2118.14 ;
     RECT  2723.9 2127.18 2730.62 2182.42 ;
     RECT  2716.9 1428.72 2731.58 1527.2 ;
     RECT  2729.86 1902.06 2731.78 1939.64 ;
     RECT  2730.62 2115.84 2732.06 2182.42 ;
     RECT  2721.7 2192.28 2732.06 2203 ;
     RECT  2730.34 1991.94 2733.22 2105.96 ;
     RECT  2731.58 1428.72 2733.5 1527.62 ;
     RECT  2731.78 1902.06 2733.7 1938.38 ;
     RECT  2733.22 2061.24 2735.62 2105.96 ;
     RECT  2703.94 1537.92 2735.9 1889.66 ;
     RECT  2732.06 2115.84 2736.1 2203 ;
     RECT  2613 3222 2737 3400 ;
     RECT  2736.1 2122.56 2737.06 2203 ;
     RECT  2716.9 1389.26 2738.3 1416.76 ;
     RECT  2733.5 1425.36 2738.3 1527.62 ;
     RECT  2737.06 2199.84 2738.5 2203 ;
     RECT  2738.3 1389.26 2738.78 1527.62 ;
     RECT  2735.9 1537.5 2738.78 1889.66 ;
     RECT  2738.78 1389.26 2739.46 1889.66 ;
     RECT  2737.06 2122.56 2739.94 2189.98 ;
     RECT  2735.62 2081.82 2740.7 2105.96 ;
     RECT  2739.94 2143.56 2742.34 2189.98 ;
     RECT  2733.7 1903.32 2742.82 1938.38 ;
     RECT  2739.94 2122.56 2744.26 2134.94 ;
     RECT  2739.46 1467.36 2744.74 1889.66 ;
     RECT  2742.34 2158.26 2748.86 2189.98 ;
     RECT  2738.5 2202.8 2748.86 2203 ;
     RECT  2744.26 2127.18 2750.3 2134.94 ;
     RECT  2742.34 2143.56 2750.3 2149.64 ;
     RECT  2739.46 1389.26 2750.5 1458.34 ;
     RECT  2556.58 2361.14 2750.98 2365.12 ;
     RECT  2723.62 1960.86 2752.22 1981.64 ;
     RECT  2733.22 1991.94 2752.22 2051.78 ;
     RECT  2750.5 1389.26 2752.9 1456.22 ;
     RECT  2750.3 2127.18 2753.38 2149.64 ;
     RECT  2748.86 2158.26 2753.86 2203 ;
     RECT  2556.58 2379.62 2753.86 2379.82 ;
     RECT  2752.22 1960.86 2754.14 2051.78 ;
     RECT  2753.86 2182.22 2755.3 2203 ;
     RECT  2744.74 1467.78 2756.06 1889.66 ;
     RECT  2754.14 1954.56 2756.06 2051.78 ;
     RECT  2753.86 2158.26 2756.26 2173.18 ;
     RECT  2756.06 1467.78 2757.98 1893.02 ;
     RECT  2742.82 1903.32 2757.98 1928.72 ;
     RECT  2742.82 1938.18 2757.98 1938.38 ;
     RECT  2756.06 1950.36 2758.46 2051.78 ;
     RECT  2752.9 1432.5 2758.94 1456.22 ;
     RECT  2757.98 1467.78 2758.94 1938.38 ;
     RECT  2758.46 1950.36 2758.94 2052.62 ;
     RECT  2758.94 1432.5 2760.1 2052.62 ;
     RECT  2760.1 1497.6 2763.26 2052.62 ;
     RECT  2735.62 2063.34 2763.26 2070.68 ;
     RECT  2740.7 2081.82 2764.7 2112.26 ;
     RECT  2753.38 2127.18 2764.7 2134.94 ;
     RECT  2753.38 2143.56 2764.7 2149.64 ;
     RECT  2763.26 1497.6 2766.82 2070.68 ;
     RECT  2764.7 2081.82 2768.74 2113.1 ;
     RECT  2766.82 1497.6 2769.7 1981.64 ;
     RECT  2760.1 1432.5 2771.42 1488.98 ;
     RECT  2769.7 1497.6 2771.42 1944.68 ;
     RECT  2764.7 2127.18 2772.38 2149.64 ;
     RECT  2752.9 1389.26 2773.34 1421.36 ;
     RECT  2766.82 1992.36 2774.78 2070.68 ;
     RECT  2771.42 1432.5 2774.98 1944.68 ;
     RECT  2774.78 1992.36 2775.74 2071.52 ;
     RECT  2768.74 2111.64 2775.74 2113.1 ;
     RECT  2772.38 2123.4 2775.74 2149.64 ;
     RECT  2769.7 1955.4 2778.62 1981.64 ;
     RECT  2775.74 2111.64 2778.82 2149.64 ;
     RECT  2778.82 2123.4 2780.74 2149.64 ;
     RECT  2773.34 1389.26 2781.02 1422.2 ;
     RECT  2774.98 1432.5 2781.02 1930.82 ;
     RECT  2778.62 1953.3 2781.02 1981.64 ;
     RECT  2775.74 1992.36 2781.02 2072.36 ;
     RECT  2781.02 1953.3 2781.22 2072.36 ;
     RECT  2781.22 2070.48 2781.5 2072.36 ;
     RECT  2768.74 2081.82 2781.5 2101.76 ;
     RECT  2755.3 2182.22 2782.66 2189.98 ;
     RECT  2774.98 1941.54 2782.94 1944.68 ;
     RECT  2781.22 1953.3 2782.94 2058.08 ;
     RECT  2778.82 2111.64 2783.62 2113.52 ;
     RECT  2780.74 2127.18 2787.26 2149.64 ;
     RECT  2781.5 2070.48 2788.9 2101.76 ;
     RECT  2781.02 1389.26 2791.58 1930.82 ;
     RECT  2782.94 1941.54 2791.58 2058.08 ;
     RECT  1955.14 2274.46 2792.26 2286.16 ;
     RECT  2787.26 2127.18 2793.7 2153.84 ;
     RECT  2791.58 1389.26 2794.18 2058.08 ;
     RECT  2794.18 1389.26 2795.14 1985 ;
     RECT  2756.26 2162.9 2796.38 2173.18 ;
     RECT  2727 -70 2797 178 ;
     RECT  2782.66 2184.32 2797.34 2189.98 ;
     RECT  2794.18 1995.3 2797.82 2058.08 ;
     RECT  2788.9 2070.48 2797.82 2073.2 ;
     RECT  2795.14 1389.26 2802.34 1436.9 ;
     RECT  2802.34 1389.26 2803.3 1436.48 ;
     RECT  2795.14 1451.4 2803.58 1981.64 ;
     RECT  2796.38 2162.9 2803.58 2174.42 ;
     RECT  2797.34 2183.88 2803.58 2189.98 ;
     RECT  2803.58 2162.9 2806.66 2189.98 ;
     RECT  2737 3222 2807 3470 ;
     RECT  2803.3 1429.14 2807.14 1436.48 ;
     RECT  2806.66 2162.9 2807.14 2174 ;
     RECT  2783.62 2111.64 2807.9 2111.84 ;
     RECT  2803.58 1451.4 2808.38 1986.68 ;
     RECT  2797.82 1995.3 2808.38 2073.2 ;
     RECT  2808.38 1451.4 2809.34 2073.2 ;
     RECT  2788.9 2081.82 2809.34 2101.76 ;
     RECT  2807.14 1429.98 2809.54 1436.48 ;
     RECT  2809.34 1451.4 2811.74 2101.76 ;
     RECT  2807.9 2111.64 2811.74 2116.88 ;
     RECT  2811.74 1451.4 2813.38 2116.88 ;
     RECT  2813.38 1466.1 2814.14 2116.88 ;
     RECT  2793.7 2127.18 2814.62 2149.64 ;
     RECT  2807.14 2162.9 2815.58 2173.18 ;
     RECT  2806.66 2183.9 2815.58 2189.98 ;
     RECT  2814.14 1466.1 2815.78 2118.14 ;
     RECT  2815.78 1466.94 2816.26 2118.14 ;
     RECT  2809.54 1433.34 2818.66 1436.48 ;
     RECT  2816.26 1467.78 2819.9 2118.14 ;
     RECT  2814.62 2126.76 2819.9 2149.64 ;
     RECT  2819.9 1467.78 2820.86 2149.64 ;
     RECT  2815.58 2162.9 2820.86 2189.98 ;
     RECT  2820.86 1467.78 2821.54 2189.98 ;
     RECT  2821.54 1467.78 2823.46 2173.18 ;
     RECT  2823.46 1467.78 2823.94 2150.06 ;
     RECT  2823.94 1467.78 2828.06 1472.18 ;
     RECT  2813.38 1451.4 2831.9 1454.12 ;
     RECT  2831.9 1451.4 2834.02 1455.8 ;
     RECT  2823.94 1481.22 2836.9 2150.06 ;
     RECT  2823.46 2162.9 2839.1 2173.18 ;
     RECT  2821.54 2181.8 2839.1 2189.98 ;
     RECT  2839.1 2162.9 2839.58 2189.98 ;
     RECT  2818.66 1435.44 2839.78 1436.48 ;
     RECT  2828.06 1465.68 2841.22 1472.18 ;
     RECT  2836.9 1481.64 2843.14 2150.06 ;
     RECT  2843.14 1481.64 2844.1 2129.48 ;
     RECT  2843.14 2142.3 2844.38 2150.06 ;
     RECT  2839.58 2158.68 2844.38 2189.98 ;
     RECT  2839.78 1436.28 2844.58 1436.48 ;
     RECT  2844.1 1484.16 2855.62 2129.48 ;
     RECT  2841.22 1468.2 2857.54 1472.18 ;
     RECT  2855.62 1484.16 2857.54 1492.34 ;
     RECT  2855.62 1505.16 2857.54 2129.48 ;
     RECT  2844.38 2142.3 2858.5 2189.98 ;
     RECT  2857.54 1507.68 2858.78 2129.48 ;
     RECT  2858.5 2142.3 2858.78 2150.06 ;
     RECT  2858.78 1507.68 2860.42 2150.06 ;
     RECT  2857.54 1484.16 2864.74 1489.4 ;
     RECT  2860.42 1507.68 2865.98 2129.48 ;
     RECT  2865.98 1500.96 2870.78 2129.48 ;
     RECT  2870.78 1493.4 2870.98 2129.48 ;
     RECT  2858.5 2159.12 2871.26 2189.98 ;
     RECT  2870.98 1511.46 2872.22 2129.48 ;
     RECT  2871.26 2158.68 2873.38 2189.98 ;
     RECT  2870.98 1493.4 2873.86 1501.16 ;
     RECT  2872.22 1511.46 2875.3 2131.58 ;
     RECT  2875.3 1511.88 2877.5 2131.58 ;
     RECT  2860.42 2141.48 2877.5 2150.06 ;
     RECT  2877.5 1511.88 2877.7 2150.06 ;
     RECT  2877.7 1511.88 2879.62 2053.88 ;
     RECT  2877.7 2063.76 2883.74 2150.06 ;
     RECT  2873.38 2159.12 2883.74 2189.98 ;
     RECT  2879.62 1511.88 2885.38 2053.04 ;
     RECT  2873.86 1500.96 2886.82 1501.16 ;
     RECT  2803.3 1389.26 2888.26 1420.12 ;
     RECT  2834.02 1451.4 2889.7 1454.12 ;
     RECT  2885.38 1511.88 2891.14 2048.84 ;
     RECT  2883.74 2063.76 2901.22 2189.98 ;
     RECT  2864.74 1484.16 2901.5 1484.36 ;
     RECT  2901.22 2063.76 2901.7 2162.24 ;
     RECT  2891.14 1516.08 2903.14 2048.84 ;
     RECT  2903.14 1516.08 2903.62 2045.9 ;
     RECT  2901.22 2174.64 2904.1 2189.98 ;
     RECT  2889.7 1451.4 2904.58 1451.6 ;
     RECT  2903.62 1516.08 2905.06 2045.48 ;
     RECT  2901.7 2063.76 2905.54 2153.84 ;
     RECT  2905.06 1516.08 2913.7 2041.7 ;
     RECT  2913.7 1533.72 2914.46 2041.7 ;
     RECT  2905.54 2083.5 2914.46 2153.84 ;
     RECT  2914.46 1533.72 2915.9 2048 ;
     RECT  2905.54 2063.76 2915.9 2074.46 ;
     RECT  2914.46 2083.5 2916.58 2159.72 ;
     RECT  2915.9 1533.72 2916.86 2074.46 ;
     RECT  2916.58 2083.5 2916.86 2101.76 ;
     RECT  2916.86 1533.72 2919.46 2101.76 ;
     RECT  2797 0 2921 178 ;
     RECT  2919.46 1533.72 2925.7 2098.4 ;
     RECT  2916.58 2111.66 2927.9 2159.72 ;
     RECT  2925.7 2065.86 2928.1 2098.4 ;
     RECT  2807 3222 2931 3400 ;
     RECT  2925.7 1533.72 2931.46 2056.82 ;
     RECT  2928.1 2070.48 2932.22 2098.4 ;
     RECT  2913.7 1516.08 2933.66 1524.68 ;
     RECT  2901.5 1484.16 2933.86 1486.06 ;
     RECT  2931.46 1536.66 2934.34 2056.82 ;
     RECT  2927.9 2111.66 2934.82 2166.44 ;
     RECT  2933.66 1515.26 2935.3 1524.68 ;
     RECT  2934.34 1563.96 2936.54 2056.82 ;
     RECT  2936.54 1563.96 2937.02 2060.18 ;
     RECT  2932.22 2070.48 2937.02 2098.84 ;
     RECT  2937.02 1563.96 2937.7 2098.84 ;
     RECT  2934.82 2111.66 2938.66 2162.24 ;
     RECT  2935.3 1524.48 2944.42 1524.68 ;
     RECT  2937.7 1563.96 2944.42 2098.4 ;
     RECT  2938.66 2124.24 2944.7 2162.24 ;
     RECT  2944.7 2124.24 2947.58 2165.18 ;
     RECT  2947.58 2124.24 2947.78 2166.44 ;
     RECT  2944.42 2070.48 2949.7 2098.4 ;
     RECT  2934.34 1536.66 2951.14 1554.08 ;
     RECT  2949.7 2070.48 2951.62 2091.26 ;
     RECT  2888.26 1389.26 2952.1 1419.7 ;
     RECT  2951.62 2071.32 2952.1 2091.26 ;
     RECT  2947.78 2124.24 2952.86 2136.64 ;
     RECT  2944.42 1563.96 2954.98 2060.6 ;
     RECT  2947.78 2149.86 2955.46 2166.44 ;
     RECT  2952.86 2122.56 2955.94 2136.64 ;
     RECT  2954.98 1583.7 2956.42 2060.6 ;
     RECT  2956.42 2052.42 2956.9 2060.6 ;
     RECT  2956.9 2052.84 2957.38 2060.6 ;
     RECT  2957.38 2053.68 2958.34 2060.6 ;
     RECT  2955.46 2154.48 2958.82 2166.44 ;
     RECT  2951.14 1541.7 2959.1 1554.08 ;
     RECT  2938.66 2111.66 2959.1 2111.86 ;
     RECT  2959.1 1541.7 2959.3 1554.5 ;
     RECT  2959.1 2111.66 2959.3 2113.54 ;
     RECT  2958.82 2155.74 2959.78 2166.44 ;
     RECT  2954.98 1563.96 2960.26 1567.52 ;
     RECT  2959.78 2155.74 2961.22 2165.18 ;
     RECT  2952.1 2071.32 2962.66 2071.52 ;
     RECT  2961.22 2155.74 2962.66 2162.66 ;
     RECT  2962.66 2158.68 2963.14 2161.82 ;
     RECT  2963.14 2158.68 2964.58 2159.72 ;
     RECT  2952.1 2082.26 2965.06 2090.84 ;
     RECT  2964.58 2159.52 2965.06 2159.72 ;
     RECT  2958.34 2053.68 2966.02 2056.82 ;
     RECT  2959.3 2113.34 2966.78 2113.54 ;
     RECT  2955.94 2127.62 2966.78 2136.64 ;
     RECT  2966.02 2053.68 2966.98 2053.88 ;
     RECT  2933.86 1484.16 2969.86 1484.36 ;
     RECT  2956.42 1583.7 2970.34 2041.28 ;
     RECT  2970.34 1983.54 2971.78 2041.28 ;
     RECT  2965.06 2082.26 2972.54 2084.98 ;
     RECT  2970.34 1583.7 2973.7 1973.24 ;
     RECT  2971.78 1983.96 2974.46 2041.28 ;
     RECT  2959.3 1541.7 2974.66 1549.04 ;
     RECT  2972.54 2078.88 2975.9 2084.98 ;
     RECT  2975.9 2078.88 2977.34 2090.42 ;
     RECT  2977.34 2070.48 2977.54 2090.42 ;
     RECT  2977.54 2070.48 2978.3 2072.36 ;
     RECT  2974.46 1983.96 2979.94 2042.12 ;
     RECT  2966.78 2113.34 2979.94 2136.64 ;
     RECT  2974.66 1541.7 2980.42 1541.9 ;
     RECT  2979.94 2113.34 2980.7 2113.54 ;
     RECT  2977.54 2082.26 2981.38 2090.42 ;
     RECT  2979.94 2127.62 2983.58 2136.64 ;
     RECT  2935.3 1515.26 2984.06 1515.46 ;
     RECT  2980.7 2105.76 2984.06 2113.54 ;
     RECT  2983.58 2127.62 2984.06 2137.06 ;
     RECT  2984.06 2127.62 2984.54 2137.48 ;
     RECT  2978.3 2063.76 2986.94 2072.36 ;
     RECT  2984.06 2102.4 2986.94 2113.54 ;
     RECT  2986.94 2056.2 2987.14 2072.36 ;
     RECT  2987.14 2056.2 2987.9 2057.24 ;
     RECT  2921 -70 2991 178 ;
     RECT  2986.94 2094 2992.42 2113.54 ;
     RECT  2973.7 1583.7 2992.7 1641.44 ;
     RECT  2979.94 1983.96 2992.9 2041.28 ;
     RECT  2987.14 2071.32 2993.38 2071.52 ;
     RECT  2992.7 1579.92 2993.66 1641.44 ;
     RECT  2987.9 2052.84 2993.86 2057.24 ;
     RECT  2992.9 2037.3 2994.82 2041.28 ;
     RECT  2960.26 1565.64 2995.1 1567.52 ;
     RECT  2993.66 1576.56 2995.1 1641.44 ;
     RECT  2984.06 1515.26 2995.58 1523.02 ;
     RECT  2994.82 2038.56 2996.26 2041.28 ;
     RECT  2995.1 1557.66 2996.74 1641.44 ;
     RECT  2993.86 2053.26 2997.98 2057.24 ;
     RECT  2992.42 2094 2998.66 2102.6 ;
     RECT  2996.74 1564.8 2998.94 1641.44 ;
     RECT  2973.7 1650.48 2998.94 1973.24 ;
     RECT  2998.94 1564.8 3000.1 1973.24 ;
     RECT  2996.26 2041.08 3000.58 2041.28 ;
     RECT  2998.66 2102.4 3000.58 2102.6 ;
     RECT  2931 3222 3001 3470 ;
     RECT  3000.1 1564.8 3001.54 1748.96 ;
     RECT  3000.1 1758.42 3001.54 1973.24 ;
     RECT  3001.54 1761.36 3002.5 1973.24 ;
     RECT  2997.98 2053.26 3002.98 2060.6 ;
     RECT  3002.98 2053.26 3003.74 2055.98 ;
     RECT  3001.54 1579.92 3004.42 1748.96 ;
     RECT  3003.74 2045.28 3004.42 2055.98 ;
     RECT  3004.42 2055.78 3005.38 2055.98 ;
     RECT  3002.5 1765.56 3005.66 1973.24 ;
     RECT  2992.9 1983.96 3005.66 2026.58 ;
     RECT  2995.58 1508.94 3006.34 1523.02 ;
     RECT  3004.42 2045.28 3006.34 2045.48 ;
     RECT  3005.66 1765.56 3007.3 2026.58 ;
     RECT  3001.54 1564.8 3007.78 1567.52 ;
     RECT  3007.3 1765.56 3008.74 2022.8 ;
     RECT  2992.42 2113.34 3009.5 2113.54 ;
     RECT  3004.42 1579.92 3009.7 1635.98 ;
     RECT  3008.74 1765.56 3009.7 1964 ;
     RECT  3008.74 1973.04 3009.7 2022.8 ;
     RECT  3009.5 2111.66 3009.7 2113.54 ;
     RECT  3007.58 1504.32 3013.82 1504.52 ;
     RECT  3004.42 1647.54 3014.78 1706.12 ;
     RECT  3013.34 1538.34 3015.74 1538.54 ;
     RECT  3009.7 1983.96 3016.42 2022.8 ;
     RECT  3015.74 1538.34 3017.38 1539.8 ;
     RECT  3014.78 1647.12 3017.66 1706.12 ;
     RECT  3004.42 1716.42 3017.66 1748.96 ;
     RECT  3009.7 1765.56 3022.66 1887.14 ;
     RECT  3009.7 1579.92 3023.9 1633.88 ;
     RECT  3022.66 1765.56 3024.1 1886.3 ;
     RECT  3017.66 1647.12 3025.54 1748.96 ;
     RECT  3013.82 1496.76 3026.98 1504.52 ;
     RECT  3007.78 1565.64 3029.66 1567.52 ;
     RECT  3025.54 1647.12 3030.14 1727.12 ;
     RECT  3029.66 1565.64 3031.58 1568.78 ;
     RECT  3009.7 1896.18 3032.06 1964 ;
     RECT  3009.7 1973.04 3032.06 1973.24 ;
     RECT  3016.42 1983.96 3032.54 2018.6 ;
     RECT  3023.9 1578.66 3033.5 1633.88 ;
     RECT  3030.14 1646.28 3033.5 1727.12 ;
     RECT  3031.58 1565.64 3033.98 1569.2 ;
     RECT  3033.5 1578.66 3033.98 1727.12 ;
     RECT  3032.06 1896.18 3034.66 1973.24 ;
     RECT  3025.54 1739.1 3037.06 1748.96 ;
     RECT  3024.1 1765.56 3038.98 1885.88 ;
     RECT  3017.38 1538.34 3039.46 1538.54 ;
     RECT  3033.98 1565.64 3040.42 1727.12 ;
     RECT  3038.98 1822.68 3040.9 1885.88 ;
     RECT  3032.54 1983.54 3040.9 2018.6 ;
     RECT  3038.98 1765.56 3041.38 1812.38 ;
     RECT  3040.9 1836.96 3041.38 1885.88 ;
     RECT  3041.38 1840.74 3042.34 1885.88 ;
     RECT  3042.34 1854.6 3045.02 1885.88 ;
     RECT  3045.02 1854.6 3045.22 1886.72 ;
     RECT  3006.34 1515.26 3045.5 1523.02 ;
     RECT  3045.5 1515.26 3045.7 1530.16 ;
     RECT  3041.38 1765.56 3045.7 1802.72 ;
     RECT  3040.9 1983.96 3046.18 2018.6 ;
     RECT  3046.18 1983.96 3046.66 2015.66 ;
     RECT  3045.22 1870.98 3048.58 1886.72 ;
     RECT  3040.9 1822.68 3049.06 1825.82 ;
     RECT  3040.42 1565.64 3049.82 1580.12 ;
     RECT  3040.42 1592.94 3050.02 1727.12 ;
     RECT  3050.02 1592.94 3050.3 1633.88 ;
     RECT  3037.06 1742.88 3050.3 1748.96 ;
     RECT  3042.34 1840.74 3050.98 1845.98 ;
     RECT  3048.58 1870.98 3050.98 1885.88 ;
     RECT  3049.82 1565.64 3051.26 1581.38 ;
     RECT  3050.3 1591.68 3051.26 1633.88 ;
     RECT  3034.66 1896.18 3051.46 1964 ;
     RECT  3050.3 1736.58 3052.9 1748.96 ;
     RECT  3051.26 1565.64 3053.38 1633.88 ;
     RECT  3052.9 1736.58 3053.38 1746.02 ;
     RECT  3050.98 1870.98 3053.86 1882.94 ;
     RECT  3053.38 1565.64 3054.82 1633.04 ;
     RECT  3050.02 1647.54 3055.3 1727.12 ;
     RECT  3045.7 1765.98 3056.26 1802.72 ;
     RECT  3051.46 1897.86 3056.54 1964 ;
     RECT  3034.66 1973.04 3056.54 1973.24 ;
     RECT  3055.3 1647.96 3056.74 1727.12 ;
     RECT  3056.54 1897.86 3056.74 1973.24 ;
     RECT  3053.38 1736.58 3057.22 1743.08 ;
     RECT  3054.82 1565.64 3057.7 1577.18 ;
     RECT  3054.82 1585.8 3057.7 1633.04 ;
     RECT  3057.7 1586.64 3058.18 1633.04 ;
     RECT  3057.22 1736.58 3058.18 1742.24 ;
     RECT  3057.7 1565.64 3058.66 1574.24 ;
     RECT  3056.74 1897.86 3058.66 1923.68 ;
     RECT  3056.74 1935.26 3058.66 1973.24 ;
     RECT  3058.66 1565.64 3059.14 1573.82 ;
     RECT  3041.38 1812.18 3059.14 1812.38 ;
     RECT  3059.14 1565.64 3059.62 1570.46 ;
     RECT  3058.18 1613.52 3059.62 1633.04 ;
     RECT  3058.66 1903.32 3059.62 1923.68 ;
     RECT  3059.62 1615.62 3060.1 1633.04 ;
     RECT  3056.74 1647.96 3060.1 1705.7 ;
     RECT  3045.22 1854.6 3060.1 1862.36 ;
     RECT  3059.62 1903.32 3060.1 1911.5 ;
     RECT  3045.7 1522.82 3060.86 1530.16 ;
     RECT  3059.62 1920.12 3061.06 1923.68 ;
     RECT  3050.98 1845.78 3061.54 1845.98 ;
     RECT  3060.86 1522.82 3063.46 1535.18 ;
     RECT  3058.18 1586.64 3063.46 1597.76 ;
     RECT  3063.46 1587.48 3063.94 1597.76 ;
     RECT  3056.26 1765.98 3065.86 1797.26 ;
     RECT  3063.94 1587.5 3066.34 1588.1 ;
     RECT  3061.06 1923.48 3066.34 1923.68 ;
     RECT  3046.66 1983.96 3066.34 2014.82 ;
     RECT  3058.18 1742.04 3066.82 1742.24 ;
     RECT  3060.1 1903.32 3067.3 1907.72 ;
     RECT  3049.06 1822.68 3067.78 1822.88 ;
     RECT  3066.34 1983.96 3067.78 1999.28 ;
     RECT  3067.78 1983.96 3068.26 1985 ;
     RECT  3068.26 1984.8 3068.74 1985 ;
     RECT  2721.7 2211.62 3070.66 2224.84 ;
     RECT  3026.98 1504.32 3070.94 1504.52 ;
     RECT  3058.66 1973.04 3070.94 1973.24 ;
     RECT  3070.46 2044.46 3070.94 2044.66 ;
     RECT  3063.46 1522.82 3071.14 1530.16 ;
     RECT  3058.66 1950.36 3071.42 1964 ;
     RECT  3070.66 2211.62 3071.62 2216.44 ;
     RECT  3070.94 1504.32 3071.9 1512.52 ;
     RECT  3058.66 1935.26 3071.9 1935.46 ;
     RECT  3060.1 1647.96 3072.1 1703.6 ;
     RECT  3067.78 1993.62 3072.1 1999.28 ;
     RECT  3072.1 1999.08 3072.58 1999.28 ;
     RECT  3070.94 2042.36 3072.86 2044.66 ;
     RECT  3066.34 2008.34 3073.06 2014.82 ;
     RECT  3059.62 1565.64 3073.34 1567.52 ;
     RECT  3072.86 2039.84 3073.34 2047.6 ;
     RECT  3071.62 2211.62 3073.54 2216.02 ;
     RECT  3067.3 1907.52 3077.66 1907.72 ;
     RECT  3077.66 1986.92 3078.62 1987.12 ;
     RECT  3060.1 1615.62 3081.7 1631.36 ;
     RECT  3072.1 1652.58 3081.7 1703.6 ;
     RECT  3069.98 1492.58 3083.42 1492.78 ;
     RECT  3071.9 1504.32 3083.42 1515.46 ;
     RECT  3073.06 2008.34 3083.9 2012.32 ;
     RECT  2904.1 2178.44 3084.1 2189.98 ;
     RECT  3083.42 1492.58 3084.38 1515.46 ;
     RECT  3071.14 1529.96 3084.86 1530.16 ;
     RECT  3077.66 1907.52 3084.86 1911.94 ;
     RECT  3083.9 2008.34 3084.86 2019.88 ;
     RECT  2857.54 1469.04 3085.34 1472.18 ;
     RECT  3084.38 1487.54 3085.34 1515.46 ;
     RECT  3070.46 1898.72 3085.34 1898.92 ;
     RECT  3084.86 1907.52 3085.34 1916.56 ;
     RECT  3070.94 1973.04 3085.34 1974.52 ;
     RECT  3078.62 1984.82 3085.34 1987.12 ;
     RECT  2981.38 2082.26 3085.54 2084.98 ;
     RECT  3084.86 1529.96 3085.82 1538.14 ;
     RECT  3084.86 1548.44 3085.82 1548.64 ;
     RECT  3071.9 1934 3085.82 1935.46 ;
     RECT  3071.42 1949.12 3085.82 1964 ;
     RECT  3084.86 2004.56 3085.82 2019.88 ;
     RECT  3085.34 1468.22 3086.3 1515.46 ;
     RECT  3085.82 1529.96 3086.3 1548.64 ;
     RECT  3085.34 1973.04 3086.3 1987.12 ;
     RECT  3085.82 1999.52 3086.3 2019.88 ;
     RECT  3073.34 2032.7 3086.3 2047.6 ;
     RECT  3086.3 1973.04 3086.78 1990.9 ;
     RECT  3086.3 1999.52 3086.78 2047.6 ;
     RECT  3086.3 1468.22 3088.9 1548.64 ;
     RECT  3073.34 1563.14 3088.9 1567.52 ;
     RECT  3063.94 1597.56 3088.9 1597.76 ;
     RECT  3081.7 1615.62 3088.9 1621.7 ;
     RECT  3081.7 1652.58 3088.9 1673.36 ;
     RECT  3081.7 1683.24 3088.9 1703.6 ;
     RECT  3060.1 1862.16 3088.9 1862.36 ;
     RECT  3053.86 1874.34 3088.9 1882.94 ;
     RECT  3085.82 1934 3088.9 1964 ;
     RECT  3086.78 1973.04 3088.9 2047.6 ;
     RECT  3088.9 1468.22 3089.38 1502.86 ;
     RECT  3088.9 1656.78 3089.38 1671.26 ;
     RECT  3088.9 1874.34 3089.38 1874.54 ;
     RECT  3088.9 1934 3089.38 1961.48 ;
     RECT  3089.38 1666.44 3089.86 1671.26 ;
     RECT  3089.38 1656.78 3090.34 1656.98 ;
     RECT  3085.34 1898.72 3091.58 1916.56 ;
     RECT  3085.54 2082.68 3091.78 2084.98 ;
     RECT  3088.9 1512.32 3092.06 1548.64 ;
     RECT  3088.9 1563.14 3092.06 1563.34 ;
     RECT  3091.58 1898.72 3092.54 1924.12 ;
     RECT  3092.54 1893.26 3093.02 1924.12 ;
     RECT  3089.38 1934 3093.02 1958.14 ;
     RECT  3084.1 2178.86 3093.22 2189.98 ;
     RECT  3093.02 1893.26 3093.5 1958.14 ;
     RECT  3093.22 2181.8 3093.7 2189.98 ;
     RECT  3056.74 1716.42 3094.18 1727.12 ;
     RECT  3065.86 1789.08 3094.18 1797.26 ;
     RECT  3065.86 1765.98 3094.66 1777.1 ;
     RECT  3009.7 2111.66 3094.66 2111.86 ;
     RECT  3094.66 1773.12 3095.14 1777.1 ;
     RECT  3091.78 2082.68 3095.14 2084.56 ;
     RECT  3094.18 1789.08 3095.62 1789.28 ;
     RECT  3094.18 1723.14 3097.06 1727.12 ;
     RECT  2984.54 2127.62 3097.06 2137.9 ;
     RECT  3095.14 2082.68 3097.54 2082.88 ;
     RECT  3088.9 1685.76 3098.02 1702.34 ;
     RECT  3097.06 2127.62 3098.02 2137.48 ;
     RECT  3089.38 1469.06 3098.3 1502.86 ;
     RECT  3092.06 1512.32 3098.3 1563.34 ;
     RECT  3098.02 1685.76 3098.5 1694.36 ;
     RECT  3095.14 1776.9 3098.5 1777.1 ;
     RECT  3093.7 2182.22 3098.5 2189.98 ;
     RECT  3093.5 1891.16 3098.78 1958.14 ;
     RECT  2952.1 1389.26 3098.98 1419.28 ;
     RECT  3089.86 1671.06 3098.98 1671.26 ;
     RECT  3097.06 1726.92 3098.98 1727.12 ;
     RECT  3098.02 2127.62 3098.98 2136.64 ;
     RECT  3098.98 1389.26 3099.46 1396.6 ;
     RECT  3098.3 1469.06 3099.46 1563.34 ;
     RECT  2615.62 2243.12 3099.46 2264.74 ;
     RECT  3099.46 1477.46 3099.7 1563.34 ;
     RECT  3098.78 1889.06 3099.7 1958.14 ;
     RECT  3088.9 1974.32 3099.7 2047.6 ;
     RECT  3099.7 1512.32 3099.94 1512.52 ;
     RECT  3099.7 1916.36 3099.94 1916.56 ;
     RECT  3099.7 2017.16 3099.94 2017.36 ;
     RECT  3098.98 1405.22 3100.42 1419.28 ;
     RECT  3099.7 1529.96 3100.42 1530.16 ;
     RECT  3073.54 2211.62 3100.42 2213.92 ;
     RECT  3100.42 1406.9 3101.38 1419.28 ;
     RECT  3101.38 1407.74 3101.86 1419.28 ;
     RECT  3099.46 2243.12 3102.14 2259.7 ;
     RECT  3102.535 1029.28 3104.265 1034.76 ;
     RECT  3102.535 1640.32 3104.265 1645.8 ;
     RECT  3102.14 2241.44 3104.265 2259.7 ;
     RECT  1795.6 994.8 3104.4 999.4 ;
     RECT  2792.26 2274.46 3104.4 2279.06 ;
     RECT  3081.7 1631.16 3105.135 1631.36 ;
     RECT  3105.135 1017.88 3106.865 1023.36 ;
     RECT  3105.135 1628.92 3106.865 1634.4 ;
     RECT  3104.4 994.8 3107 996.8 ;
     RECT  3104.4 2277.06 3107 2279.06 ;
     RECT  3098.98 2127.62 3107.62 2134.96 ;
     RECT  2755.3 2202.8 3110.3 2203 ;
     RECT  3100.42 2211.62 3110.3 2212.24 ;
     RECT  3104.265 2241.44 3110.5 2250.04 ;
     RECT  3110.3 1999.94 3111.94 2003.08 ;
     RECT  3104.265 2259.5 3112.42 2259.7 ;
     RECT  3111.94 2000.78 3112.9 2003.08 ;
     RECT  3110.3 2050.76 3112.9 2052.64 ;
     RECT  3110.3 2101.58 3112.9 2103.04 ;
     RECT  3110.3 2202.38 3112.9 2212.24 ;
     RECT  3112.9 2000.78 3113.38 2000.98 ;
     RECT  3112.9 2051.18 3113.38 2051.8 ;
     RECT  3112.9 2102.84 3113.38 2103.04 ;
     RECT  3110.3 2152.4 3113.38 2153.44 ;
     RECT  3112.9 2202.38 3113.38 2203 ;
     RECT  3112.9 2212.04 3113.38 2212.24 ;
     RECT  3107.62 2127.62 3113.86 2134.54 ;
     RECT  2991 0 3115 178 ;
     RECT  3001 3222 3125 3400 ;
     RECT  3113.86 2127.62 3170.02 2127.82 ;
     RECT  3066.34 1587.5 3171.46 1587.7 ;
     RECT  3115 -70 3185 178 ;
     RECT  3125 3222 3195 3470 ;
     RECT  3101.86 1410.26 3207.46 1419.28 ;
     RECT  3098.5 2182.22 3207.46 2182.42 ;
     RECT  3207.46 1414.88 3207.94 1419.28 ;
     RECT  3110.5 2244.38 3207.94 2250.04 ;
     RECT  3185 0 3220 178 ;
     RECT  3195 3222 3220 3400 ;
     RECT  3220 0 3222 180 ;
     RECT  3099.46 1389.26 3222 1389.46 ;
     RECT  3207.94 1419.08 3222 1419.28 ;
     RECT  3207.26 1771.88 3222 1772.08 ;
     RECT  3207.26 1965.08 3222 1965.28 ;
     RECT  3113.38 2202.8 3222 2203 ;
     RECT  3207.94 2244.38 3222 2244.58 ;
     RECT  2750.98 2361.14 3222 2361.34 ;
     RECT  1797.98 2548.46 3222 2555.8 ;
     RECT  1774.46 2736.2 3222 2743.54 ;
     RECT  3220 3220 3222 3400 ;
     RECT  3222 0 3400 3400 ;
     RECT  3400 205 3470 275 ;
     RECT  3400 399 3470 469 ;
     RECT  3400 593 3470 663 ;
     RECT  3400 787 3470 857 ;
     RECT  3400 981 3470 1051 ;
     RECT  3400 1175 3470 1245 ;
     RECT  3400 1369 3470 1439 ;
     RECT  3400 1563 3470 1633 ;
     RECT  3400 1757 3470 1827 ;
     RECT  3400 1951 3470 2021 ;
     RECT  3400 2145 3470 2215 ;
     RECT  3400 2339 3470 2409 ;
     RECT  3400 2533 3470 2603 ;
     RECT  3400 2727 3470 2797 ;
     RECT  3400 2921 3470 2991 ;
     RECT  3400 3115 3470 3185 ;
    LAYER Metal5 ;
     RECT  205 -70 275 0 ;
     RECT  399 -70 469 0 ;
     RECT  593 -70 663 0 ;
     RECT  787 -70 857 0 ;
     RECT  981 -70 1051 0 ;
     RECT  1175 -70 1245 0 ;
     RECT  1369 -70 1439 0 ;
     RECT  1563 -70 1633 0 ;
     RECT  1757 -70 1827 0 ;
     RECT  1951 -70 2021 0 ;
     RECT  2145 -70 2215 0 ;
     RECT  2339 -70 2409 0 ;
     RECT  2533 -70 2603 0 ;
     RECT  2727 -70 2797 0 ;
     RECT  2921 -70 2991 0 ;
     RECT  3115 -70 3185 0 ;
     RECT  0 0 3400 178 ;
     RECT  0 178 180 180 ;
     RECT  3220 178 3400 180 ;
     RECT  3222 180 3400 205 ;
     RECT  0 180 178 215 ;
     RECT  3222 205 3470 275 ;
     RECT  -70 215 178 285 ;
     RECT  3222 275 3400 399 ;
     RECT  0 285 178 409 ;
     RECT  3222 399 3470 469 ;
     RECT  -70 409 178 479 ;
     RECT  3222 469 3400 593 ;
     RECT  0 479 178 603 ;
     RECT  993.18 616.555 994.82 622.125 ;
     RECT  1405.18 616.555 1406.82 622.125 ;
     RECT  995.78 627.955 997.42 633.525 ;
     RECT  1402.58 627.955 1404.22 633.525 ;
     RECT  3222 593 3470 663 ;
     RECT  -70 603 178 673 ;
     RECT  992.06 755.06 992.26 758.42 ;
     RECT  1397.66 750.44 1397.86 760.94 ;
     RECT  1397.66 760.94 1399.3 763.04 ;
     RECT  976.7 741.2 976.9 769.76 ;
     RECT  991.1 758.42 992.26 769.76 ;
     RECT  1008.86 745.4 1009.06 777.32 ;
     RECT  1008.38 777.32 1009.06 778.16 ;
     RECT  1188.54 764.54 1188.74 779.44 ;
     RECT  1250.46 760.34 1250.66 779.86 ;
     RECT  1397.66 763.04 1399.78 781.1 ;
     RECT  976.7 769.76 992.26 782.995 ;
     RECT  976.7 782.995 994.82 783.62 ;
     RECT  1008.38 778.16 1018.66 783.62 ;
     RECT  3222 663 3400 787 ;
     RECT  1397.66 781.1 1407.94 789.08 ;
     RECT  0 673 178 797 ;
     RECT  1252.86 802.34 1253.06 802.76 ;
     RECT  1252.86 802.76 1253.54 809.9 ;
     RECT  976.7 783.62 1018.66 816.38 ;
     RECT  1032.86 813.44 1033.06 816.38 ;
     RECT  1252.38 809.9 1253.54 818.08 ;
     RECT  1252.86 818.08 1253.54 833.2 ;
     RECT  1252.86 833.2 1253.06 851.68 ;
     RECT  1153.98 843.92 1154.18 856.72 ;
     RECT  3222 787 3470 857 ;
     RECT  -70 797 178 867 ;
     RECT  976.7 816.38 1033.06 918.22 ;
     RECT  3222 857 3400 981 ;
     RECT  0 867 178 991 ;
     RECT  1793.18 1017.835 1794.82 1023.405 ;
     RECT  3105.18 1017.835 3106.82 1023.405 ;
     RECT  1795.78 1029.235 1797.42 1034.805 ;
     RECT  3102.58 1029.235 3104.22 1034.805 ;
     RECT  3222 981 3470 1051 ;
     RECT  -70 991 178 1061 ;
     RECT  3222 1051 3400 1175 ;
     RECT  0 1061 178 1185 ;
     RECT  3222 1175 3470 1245 ;
     RECT  -70 1185 178 1255 ;
     RECT  3222 1245 3400 1369 ;
     RECT  0 1255 178 1379 ;
     RECT  3099.26 1396.4 3099.46 1404.38 ;
     RECT  2681.66 1403.96 2681.86 1404.8 ;
     RECT  2660.54 1403.96 2660.74 1405.64 ;
     RECT  3098.78 1404.38 3099.46 1406.06 ;
     RECT  2675.42 1404.8 2681.86 1406.48 ;
     RECT  2660.54 1405.64 2661.22 1406.9 ;
     RECT  2674.46 1406.48 2681.86 1406.9 ;
     RECT  2660.54 1406.9 2681.86 1407.32 ;
     RECT  3084.86 1405.64 3085.06 1407.32 ;
     RECT  3097.82 1406.06 3099.46 1407.32 ;
     RECT  1767.74 1409.42 1767.94 1409.84 ;
     RECT  3070.94 1403.54 3071.14 1410.4 ;
     RECT  1760.06 1409.84 1767.94 1411.52 ;
     RECT  1760.06 1411.52 1776.1 1411.94 ;
     RECT  2757.02 1412.68 2763.94 1413.2 ;
     RECT  2652.86 1407.32 2681.86 1413.62 ;
     RECT  2757.02 1413.2 2765.38 1415.92 ;
     RECT  2757.98 1415.92 2765.38 1416.98 ;
     RECT  2757.98 1416.98 2774.5 1417.44 ;
     RECT  2763.26 1417.44 2774.5 1418.24 ;
     RECT  2763.26 1418.24 2782.66 1419.08 ;
     RECT  1585.82 1406.06 1586.02 1429.16 ;
     RECT  3222 1369 3470 1439 ;
     RECT  1692.86 1423.28 1693.06 1439.24 ;
     RECT  1653.98 1403.54 1654.18 1439.66 ;
     RECT  2729.18 1437.76 2735.14 1440.04 ;
     RECT  2763.26 1419.08 2786.5 1441.12 ;
     RECT  2729.18 1440.04 2735.62 1442.18 ;
     RECT  2729.18 1442.18 2736.58 1442.32 ;
     RECT  2764.7 1441.12 2786.5 1442.38 ;
     RECT  2728.22 1442.32 2736.58 1442.52 ;
     RECT  1104.86 1418.66 1105.06 1443.44 ;
     RECT  2422.46 1414.88 2422.66 1443.44 ;
     RECT  2728.22 1442.52 2735.62 1444.48 ;
     RECT  2696.06 1404.38 2696.26 1444.7 ;
     RECT  2774.3 1442.38 2786.5 1444.9 ;
     RECT  2782.46 1444.9 2786.5 1445.74 ;
     RECT  1653.98 1439.66 1663.78 1446.38 ;
     RECT  1086.14 1445.96 1086.34 1446.8 ;
     RECT  1096.22 1443.44 1105.06 1446.8 ;
     RECT  1689.98 1439.24 1693.06 1446.88 ;
     RECT  3070.94 1410.4 3073.54 1446.88 ;
     RECT  2696.06 1444.7 2696.74 1447.84 ;
     RECT  2696.06 1447.84 2696.26 1448.26 ;
     RECT  -70 1379 178 1449 ;
     RECT  2729.66 1444.48 2735.62 1449.36 ;
     RECT  1653.98 1446.38 1670.98 1449.52 ;
     RECT  1653.98 1449.52 1654.18 1450.58 ;
     RECT  1649.18 1450.58 1654.18 1454.36 ;
     RECT  1625.18 1393.04 1625.38 1454.56 ;
     RECT  1670.78 1449.52 1670.98 1456.88 ;
     RECT  1684.7 1446.88 1693.06 1456.88 ;
     RECT  3084.86 1407.32 3099.46 1458.28 ;
     RECT  2750.3 1453.72 2750.5 1458.34 ;
     RECT  2783.42 1445.74 2786.5 1458.48 ;
     RECT  2733.5 1449.36 2735.62 1462.74 ;
     RECT  2783.42 1458.48 2783.62 1463.16 ;
     RECT  2774.78 1463.16 2783.62 1465.32 ;
     RECT  1670.78 1456.88 1693.06 1469.68 ;
     RECT  2645.66 1413.62 2681.86 1472.4 ;
     RECT  1670.78 1469.68 1690.18 1473.46 ;
     RECT  1670.78 1473.46 1684.9 1482.92 ;
     RECT  1759.58 1411.94 1776.1 1483.76 ;
     RECT  3084.86 1458.28 3100.42 1484.8 ;
     RECT  1584.86 1429.16 1586.02 1487.12 ;
     RECT  2645.66 1472.4 2688.1 1488.16 ;
     RECT  2733.5 1462.74 2739.46 1491.92 ;
     RECT  1641.98 1454.36 1654.18 1492.16 ;
     RECT  3069.98 1446.88 3073.54 1492.78 ;
     RECT  2681.66 1488.16 2688.1 1494.04 ;
     RECT  2774.78 1465.32 2774.98 1495.5 ;
     RECT  1629.98 1492.16 1630.18 1495.52 ;
     RECT  1397.66 789.08 1408.9 1498.66 ;
     RECT  2774.78 1495.5 2777.86 1502.84 ;
     RECT  2687.9 1494.04 2688.1 1504.1 ;
     RECT  2777.18 1502.84 2777.86 1504.74 ;
     RECT  3084.86 1484.8 3099.46 1507.9 ;
     RECT  2735.9 1491.92 2739.46 1508.1 ;
     RECT  1669.82 1482.92 1684.9 1509.16 ;
     RECT  1513.34 1498.88 1513.54 1511.68 ;
     RECT  3070.94 1492.78 3073.54 1512.52 ;
     RECT  1584.86 1487.12 1586.5 1514.2 ;
     RECT  2645.66 1488.16 2667.46 1515.04 ;
     RECT  2933.66 1485.86 2933.86 1515.46 ;
     RECT  1439.42 1506.86 1439.62 1518.2 ;
     RECT  2751.26 1511.46 2751.46 1518.6 ;
     RECT  3084.86 1507.9 3096.1 1519.66 ;
     RECT  2731.58 1508.1 2739.46 1520.28 ;
     RECT  2777.18 1504.74 2778.82 1520.9 ;
     RECT  1641.98 1492.16 1658.02 1521.34 ;
     RECT  1086.14 1446.8 1105.06 1521.76 ;
     RECT  2777.18 1520.9 2778.34 1522.16 ;
     RECT  3071.9 1512.52 3073.54 1522.82 ;
     RECT  2645.66 1515.04 2645.86 1524.7 ;
     RECT  2751.26 1518.6 2759.62 1524.9 ;
     RECT  2660.06 1515.04 2667.46 1525.12 ;
     RECT  1657.82 1521.34 1658.02 1527.44 ;
     RECT  1669.82 1509.16 1681.06 1527.44 ;
     RECT  1537.34 1494.68 1537.54 1528.28 ;
     RECT  2731.1 1520.28 2739.46 1528.46 ;
     RECT  1621.82 1495.52 1630.18 1528.7 ;
     RECT  1547.9 1495.94 1548.1 1528.9 ;
     RECT  3045.5 1515.26 3045.7 1530.16 ;
     RECT  2660.06 1525.12 2661.22 1531.42 ;
     RECT  1537.34 1528.28 1538.02 1531.64 ;
     RECT  1572.38 1479.56 1572.58 1532.48 ;
     RECT  2660.06 1531.42 2660.26 1532.68 ;
     RECT  1697.18 1507.28 1697.38 1533.32 ;
     RECT  2789.66 1521.54 2789.86 1535.6 ;
     RECT  1177.34 1521.56 1177.54 1535.84 ;
     RECT  1749.98 1483.76 1776.1 1536.88 ;
     RECT  2777.18 1522.16 2777.38 1537.28 ;
     RECT  2735.9 1528.46 2739.46 1538.96 ;
     RECT  1584.86 1514.2 1586.02 1540.88 ;
     RECT  1697.18 1533.32 1697.86 1541.3 ;
     RECT  2735.9 1538.96 2737.06 1541.48 ;
     RECT  1584.86 1540.88 1589.38 1544.44 ;
     RECT  1657.82 1527.44 1681.06 1547.6 ;
     RECT  1697.18 1541.3 1706.5 1547.6 ;
     RECT  3084.86 1519.66 3088.42 1548.64 ;
     RECT  1738.46 1536.68 1738.66 1551.58 ;
     RECT  1749.98 1536.88 1775.14 1552 ;
     RECT  2751.26 1524.9 2760.58 1558.08 ;
     RECT  1094.78 1521.76 1105.06 1558.3 ;
     RECT  2736.38 1541.48 2737.06 1561.64 ;
     RECT  1565.18 1532.48 1572.58 1562.5 ;
     RECT  3222 1439 3400 1563 ;
     RECT  3070.94 1522.82 3073.54 1563.34 ;
     RECT  2829.98 1540.02 2830.18 1565 ;
     RECT  2718.62 1549.68 2718.82 1567.1 ;
     RECT  2631.26 1410.4 2631.46 1567.12 ;
     RECT  1173.98 1535.84 1177.54 1567.96 ;
     RECT  2751.26 1558.08 2768.26 1569.2 ;
     RECT  1173.98 1567.96 1174.18 1569.64 ;
     RECT  2736.86 1561.64 2737.06 1572.78 ;
     RECT  0 1449 178 1573 ;
     RECT  1521.98 1555.16 1522.18 1574.06 ;
     RECT  1537.34 1531.64 1544.26 1574.06 ;
     RECT  2794.46 1563.12 2794.66 1577.82 ;
     RECT  2767.58 1569.2 2768.26 1578.24 ;
     RECT  1473.5 1518.2 1473.7 1578.68 ;
     RECT  2659.1 1554.3 2659.3 1579.7 ;
     RECT  2736.86 1572.78 2739.94 1579.92 ;
     RECT  2734.94 1579.92 2739.94 1580.34 ;
     RECT  2751.26 1569.2 2756.74 1580.34 ;
     RECT  2767.58 1578.24 2769.22 1580.34 ;
     RECT  2779.1 1562.28 2779.3 1580.34 ;
     RECT  2907.74 1576.98 2907.94 1580.54 ;
     RECT  1094.78 1558.3 1094.98 1580.98 ;
     RECT  2734.94 1580.34 2756.74 1581.18 ;
     RECT  2767.58 1580.34 2779.3 1581.18 ;
     RECT  1657.82 1547.6 1706.5 1582.24 ;
     RECT  2734.94 1581.18 2779.3 1583.28 ;
     RECT  1104.86 1558.3 1105.06 1583.5 ;
     RECT  2794.46 1577.82 2798.5 1583.7 ;
     RECT  1753.34 1552 1775.14 1583.72 ;
     RECT  2706.62 1583.28 2706.82 1584.12 ;
     RECT  2706.62 1584.12 2716.42 1584.54 ;
     RECT  2733.02 1583.28 2779.3 1584.54 ;
     RECT  1566.62 1562.5 1572.58 1584.56 ;
     RECT  1589.18 1544.44 1589.38 1584.56 ;
     RECT  1521.98 1574.06 1551.46 1585.4 ;
     RECT  1566.62 1584.56 1589.38 1585.4 ;
     RECT  1753.34 1583.72 1778.98 1586.66 ;
     RECT  1788.86 1465.12 1789.06 1586.66 ;
     RECT  3070.94 1563.34 3071.14 1587.7 ;
     RECT  2706.62 1584.54 2779.3 1588.1 ;
     RECT  2794.46 1583.7 2798.98 1591.68 ;
     RECT  1521.98 1585.4 1589.38 1596.1 ;
     RECT  2998.94 1553.88 2999.14 1597.56 ;
     RECT  2706.62 1588.1 2753.38 1597.98 ;
     RECT  2706.62 1597.98 2753.86 1599.02 ;
     RECT  2789.66 1591.68 2798.98 1599.02 ;
     RECT  1473.5 1578.68 1480.42 1599.68 ;
     RECT  2764.7 1588.1 2779.3 1600.08 ;
     RECT  2789.66 1599.02 2798.5 1600.08 ;
     RECT  3050.78 1582.02 3050.98 1600.28 ;
     RECT  2898.14 1600.08 2898.34 1600.5 ;
     RECT  2716.22 1599.02 2753.86 1600.7 ;
     RECT  2764.7 1600.08 2798.5 1601.12 ;
     RECT  2898.14 1600.5 2899.3 1601.2 ;
     RECT  1503.74 1574.9 1503.94 1601.36 ;
     RECT  2909.18 1602.18 2909.38 1604.28 ;
     RECT  1657.82 1582.24 1697.86 1604.5 ;
     RECT  2716.22 1600.7 2740.42 1604.9 ;
     RECT  2951.9 1602.18 2952.1 1604.9 ;
     RECT  1524.38 1596.1 1589.38 1607.86 ;
     RECT  2764.7 1601.12 2785.54 1608.26 ;
     RECT  1621.82 1528.7 1631.14 1608.92 ;
     RECT  1524.38 1607.86 1524.58 1609.54 ;
     RECT  2753.18 1600.7 2753.86 1611 ;
     RECT  1465.82 1599.68 1480.42 1611.44 ;
     RECT  2909.18 1604.28 2917.54 1611.62 ;
     RECT  2909.18 1611.62 2914.18 1612.04 ;
     RECT  2937.5 1600.92 2937.7 1612.26 ;
     RECT  1151.42 1508.96 1151.62 1612.9 ;
     RECT  2764.7 1608.26 2780.74 1614.56 ;
     RECT  2929.82 1612.26 2937.7 1614.56 ;
     RECT  2724.86 1604.9 2740.42 1615.62 ;
     RECT  2752.22 1611 2753.86 1615.62 ;
     RECT  2881.34 1602.18 2881.54 1620.02 ;
     RECT  2910.14 1612.04 2914.18 1620.02 ;
     RECT  2724.86 1615.62 2754.82 1621.28 ;
     RECT  2839.1 1614.36 2839.3 1621.5 ;
     RECT  2726.3 1621.28 2754.82 1623.6 ;
     RECT  2798.3 1601.12 2798.5 1623.6 ;
     RECT  2726.3 1623.6 2755.3 1624.44 ;
     RECT  2767.58 1614.56 2780.74 1624.44 ;
     RECT  1499.42 1601.36 1503.94 1624.46 ;
     RECT  2910.14 1620.02 2912.74 1625.48 ;
     RECT  2726.3 1624.44 2780.74 1626.12 ;
     RECT  2792.06 1623.6 2798.5 1626.12 ;
     RECT  2726.3 1626.12 2798.5 1627.58 ;
     RECT  2767.1 1627.58 2798.5 1628.42 ;
     RECT  1753.34 1586.66 1789.06 1628.875 ;
     RECT  1737.5 1600.1 1737.7 1630.12 ;
     RECT  1499.42 1624.46 1513.54 1631.18 ;
     RECT  2958.62 1625.7 2958.82 1632.62 ;
     RECT  2834.78 1621.5 2839.3 1632.84 ;
     RECT  3222 1563 3470 1633 ;
     RECT  1465.82 1611.44 1487.14 1634.12 ;
     RECT  1499.42 1631.18 1516.42 1634.12 ;
     RECT  1657.82 1604.5 1658.02 1634.12 ;
     RECT  3105.18 1628.875 3106.82 1634.445 ;
     RECT  2767.1 1628.42 2767.78 1637.66 ;
     RECT  1614.62 1608.92 1631.14 1637.68 ;
     RECT  2726.3 1627.58 2753.86 1638.08 ;
     RECT  1621.82 1637.68 1631.14 1638.74 ;
     RECT  1641.98 1521.34 1647.94 1638.74 ;
     RECT  1753.34 1628.875 1794.82 1640.275 ;
     RECT  3045.98 1631.16 3046.18 1640.4 ;
     RECT  2910.14 1625.48 2910.34 1640.6 ;
     RECT  1600.22 1619.84 1600.42 1641.68 ;
     RECT  -70 1573 178 1643 ;
     RECT  2833.82 1632.84 2839.3 1643.54 ;
     RECT  2998.94 1597.56 3002.02 1643.54 ;
     RECT  2834.3 1643.54 2839.3 1644.38 ;
     RECT  1753.34 1640.275 1797.42 1645.845 ;
     RECT  3102.58 1640.275 3104.22 1645.845 ;
     RECT  2779.1 1628.42 2798.5 1646.06 ;
     RECT  2834.3 1644.38 2838.34 1646.06 ;
     RECT  2834.78 1646.06 2838.34 1648.16 ;
     RECT  1455.74 1627.4 1455.94 1650.08 ;
     RECT  2726.3 1638.08 2734.18 1650.68 ;
     RECT  2726.3 1650.68 2729.86 1651.94 ;
     RECT  3001.82 1643.54 3002.02 1652.36 ;
     RECT  1621.82 1638.74 1647.94 1653.02 ;
     RECT  2726.3 1651.94 2726.5 1654.04 ;
     RECT  2745.02 1638.08 2753.86 1655.3 ;
     RECT  3044.06 1640.4 3046.18 1655.3 ;
     RECT  2929.82 1614.56 2930.02 1655.94 ;
     RECT  2834.78 1648.16 2834.98 1656.56 ;
     RECT  2912.06 1657.2 2912.26 1657.62 ;
     RECT  1537.34 1607.86 1589.38 1658.48 ;
     RECT  1600.22 1641.68 1603.78 1658.48 ;
     RECT  1620.86 1653.02 1647.94 1658.48 ;
     RECT  2929.82 1655.94 2934.34 1659.72 ;
     RECT  2884.22 1654.68 2884.42 1660.76 ;
     RECT  1619.42 1658.48 1647.94 1661.42 ;
     RECT  1657.82 1634.12 1659.46 1661.42 ;
     RECT  1438.46 1518.2 1439.62 1663.1 ;
     RECT  1450.94 1650.08 1455.94 1663.1 ;
     RECT  2779.1 1646.06 2793.22 1666.44 ;
     RECT  2440.22 1666.46 2440.42 1667.72 ;
     RECT  1438.46 1663.1 1455.94 1668.14 ;
     RECT  1465.82 1634.12 1516.42 1668.14 ;
     RECT  2314.46 1668.14 2314.66 1668.56 ;
     RECT  2929.82 1659.72 2936.74 1669.16 ;
     RECT  2779.1 1666.44 2799.94 1670 ;
     RECT  2929.82 1669.16 2934.34 1670 ;
     RECT  3050.78 1656.36 3050.98 1670 ;
     RECT  2749.82 1655.3 2753.86 1670.42 ;
     RECT  1438.46 1668.14 1516.42 1670.66 ;
     RECT  2422.46 1443.44 2423.62 1671.7 ;
     RECT  2422.46 1671.7 2422.66 1672.12 ;
     RECT  1619.42 1661.42 1659.46 1672.54 ;
     RECT  1753.34 1645.845 1789.06 1672.54 ;
     RECT  3012.38 1669.38 3016.42 1672.74 ;
     RECT  1537.34 1658.48 1603.78 1672.76 ;
     RECT  1619.42 1672.54 1631.14 1672.76 ;
     RECT  2831.42 1660.98 2831.62 1673.16 ;
     RECT  2440.22 1667.72 2440.9 1674.64 ;
     RECT  2586.14 1674.44 2586.34 1674.86 ;
     RECT  2440.22 1674.64 2440.42 1675.06 ;
     RECT  2357.66 1408.16 2357.86 1675.28 ;
     RECT  2912.06 1657.62 2915.14 1676.52 ;
     RECT  2586.14 1674.86 2590.66 1677.36 ;
     RECT  2602.46 1674.86 2602.66 1677.38 ;
     RECT  1101.02 1672.76 1101.22 1677.58 ;
     RECT  2590.46 1677.36 2590.66 1677.58 ;
     RECT  1537.34 1672.76 1631.14 1679.26 ;
     RECT  2912.06 1676.52 2922.82 1679.88 ;
     RECT  976.7 918.22 1026.34 1681.36 ;
     RECT  2831.42 1673.16 2835.94 1682.18 ;
     RECT  1669.82 1604.5 1697.86 1684.52 ;
     RECT  3011.9 1672.74 3016.42 1685.96 ;
     RECT  2779.1 1670 2793.22 1687.02 ;
     RECT  2835.74 1682.18 2835.94 1688.48 ;
     RECT  1537.34 1679.26 1606.66 1689.56 ;
     RECT  1617.98 1679.26 1631.14 1689.56 ;
     RECT  1137.02 1641.68 1137.22 1689.76 ;
     RECT  2779.1 1687.02 2799.46 1690.16 ;
     RECT  1669.82 1684.52 1702.18 1691.24 ;
     RECT  2779.1 1690.16 2793.22 1692.68 ;
     RECT  2910.62 1679.88 2922.82 1693.32 ;
     RECT  2934.14 1670 2934.34 1694.36 ;
     RECT  1753.34 1672.54 1779.46 1695.02 ;
     RECT  1438.46 1670.66 1522.66 1695.44 ;
     RECT  1537.34 1689.56 1631.14 1695.44 ;
     RECT  2909.18 1693.32 2922.82 1696.04 ;
     RECT  2767.58 1637.66 2767.78 1696.68 ;
     RECT  2779.1 1692.68 2790.34 1696.68 ;
     RECT  2753.18 1670.42 2753.86 1698.14 ;
     RECT  2767.58 1696.68 2790.34 1698.14 ;
     RECT  1201.34 1695.86 1201.54 1698.8 ;
     RECT  1438.46 1695.44 1631.14 1698.8 ;
     RECT  1669.82 1691.24 1705.06 1698.8 ;
     RECT  1728.86 1698.38 1729.06 1698.8 ;
     RECT  1438.46 1698.8 1631.62 1705.52 ;
     RECT  1641.98 1672.54 1659.46 1705.52 ;
     RECT  1669.82 1698.8 1729.06 1705.52 ;
     RECT  2779.1 1698.14 2790.34 1705.7 ;
     RECT  2808.38 1702.14 2808.58 1705.7 ;
     RECT  2874.62 1679.88 2874.82 1705.7 ;
     RECT  2910.62 1696.04 2922.82 1705.7 ;
     RECT  3011.9 1685.96 3012.1 1705.7 ;
     RECT  1398.14 1498.66 1408.9 1705.72 ;
     RECT  1669.82 1705.52 1734.34 1706.36 ;
     RECT  2721.02 1692.9 2721.22 1708.64 ;
     RECT  2914.46 1705.7 2922.82 1710.54 ;
     RECT  1438.46 1705.52 1659.46 1710.56 ;
     RECT  1669.82 1706.36 1742.02 1710.56 ;
     RECT  1753.34 1695.02 1782.34 1710.56 ;
     RECT  1134.14 1695.44 1134.34 1710.76 ;
     RECT  2914.46 1710.54 2927.62 1711.8 ;
     RECT  2707.58 1683.66 2707.78 1712.22 ;
     RECT  2767.58 1698.14 2767.78 1713.26 ;
     RECT  1399.1 1705.72 1408.9 1713.28 ;
     RECT  2779.1 1705.7 2784.1 1715.78 ;
     RECT  1399.58 1713.28 1408.9 1717.48 ;
     RECT  2707.58 1712.22 2708.26 1719.14 ;
     RECT  2783.9 1715.78 2784.1 1719.36 ;
     RECT  2783.9 1719.36 2784.58 1719.98 ;
     RECT  2656.22 1717.26 2656.42 1720.82 ;
     RECT  2784.38 1719.98 2784.58 1720.82 ;
     RECT  3045.02 1719.78 3045.22 1720.82 ;
     RECT  2914.46 1711.8 2929.06 1722.5 ;
     RECT  2584.22 1728.18 2584.42 1729.02 ;
     RECT  2670.62 1722.3 2670.82 1730.9 ;
     RECT  2530.94 1733.64 2531.14 1734.06 ;
     RECT  1434.62 1710.56 1659.46 1734.08 ;
     RECT  1669.82 1710.56 1782.34 1734.08 ;
     RECT  2914.46 1722.5 2928.1 1734.26 ;
     RECT  2528.54 1734.06 2531.14 1734.48 ;
     RECT  2528.54 1734.48 2531.62 1734.9 ;
     RECT  1400.06 1717.48 1408.9 1734.92 ;
     RECT  1434.62 1734.08 1782.34 1737.44 ;
     RECT  2581.34 1729.02 2584.42 1738.68 ;
     RECT  2528.54 1734.9 2532.58 1739.52 ;
     RECT  2775.26 1739.1 2775.46 1741.62 ;
     RECT  2942.78 1728.18 2942.98 1741.62 ;
     RECT  2942.78 1741.62 2943.46 1745.4 ;
     RECT  2528.54 1739.52 2537.38 1745.82 ;
     RECT  1193.66 1698.8 1201.54 1746.04 ;
     RECT  2773.34 1741.62 2775.46 1748.54 ;
     RECT  1193.66 1746.04 1193.86 1748.56 ;
     RECT  1432.7 1737.44 1782.34 1749.4 ;
     RECT  2602.46 1677.38 2609.86 1749.4 ;
     RECT  2635.58 1749.2 2635.78 1749.5 ;
     RECT  2635.58 1749.5 2640.58 1749.7 ;
     RECT  2790.62 1746.24 2790.82 1750.44 ;
     RECT  2922.62 1734.26 2928.1 1750.44 ;
     RECT  2528.54 1745.82 2543.14 1750.64 ;
     RECT  2707.58 1719.14 2707.78 1751.28 ;
     RECT  2942.78 1745.4 2947.3 1755.26 ;
     RECT  2581.34 1738.68 2589.22 1755.9 ;
     RECT  2790.62 1750.44 2791.3 1755.9 ;
     RECT  2901.98 1753.38 2902.18 1755.9 ;
     RECT  2922.62 1750.44 2932.42 1756.1 ;
     RECT  2572.7 1755.9 2589.22 1756.32 ;
     RECT  3222 1633 3400 1757 ;
     RECT  1797.98 1679.9 1798.18 1757.18 ;
     RECT  2753.18 1698.14 2753.38 1757.36 ;
     RECT  2528.54 1750.64 2541.22 1758 ;
     RECT  2927.9 1756.1 2932.42 1758 ;
     RECT  2947.1 1755.26 2947.3 1758 ;
     RECT  1400.06 1734.92 1416.58 1758.64 ;
     RECT  2705.18 1751.28 2707.78 1760.94 ;
     RECT  2705.18 1760.94 2712.1 1761.36 ;
     RECT  2947.1 1758 2949.22 1761.36 ;
     RECT  2947.1 1761.36 2954.98 1761.56 ;
     RECT  2705.18 1761.36 2713.06 1761.78 ;
     RECT  2527.58 1758 2541.22 1761.98 ;
     RECT  2927.9 1758 2935.78 1764.08 ;
     RECT  2790.62 1755.9 2809.06 1765.34 ;
     RECT  2774.3 1748.54 2775.46 1765.56 ;
     RECT  2790.62 1765.34 2805.22 1765.56 ;
     RECT  2572.7 1756.32 2590.66 1765.76 ;
     RECT  2901.98 1755.9 2905.06 1766.4 ;
     RECT  2561.66 1753.8 2561.86 1766.6 ;
     RECT  942.62 1763.9 942.82 1766.62 ;
     RECT  0 1643 178 1767 ;
     RECT  2572.7 1765.76 2572.9 1767.02 ;
     RECT  1432.7 1749.4 1659.46 1767.26 ;
     RECT  1669.82 1749.4 1782.34 1767.26 ;
     RECT  1408.7 1758.64 1416.58 1767.88 ;
     RECT  2737.34 1765.98 2737.54 1768.08 ;
     RECT  2949.02 1761.56 2954.98 1769.34 ;
     RECT  2585.66 1765.76 2590.66 1769.76 ;
     RECT  2529.98 1761.98 2541.22 1770.18 ;
     RECT  2585.66 1769.76 2592.1 1770.18 ;
     RECT  2935.58 1764.08 2935.78 1770.38 ;
     RECT  2529.98 1770.18 2544.1 1770.8 ;
     RECT  1342.94 1767.26 1343.14 1771.04 ;
     RECT  2537.66 1770.8 2544.1 1771.22 ;
     RECT  2585.66 1770.18 2593.06 1771.22 ;
     RECT  2737.34 1768.08 2739.94 1771.22 ;
     RECT  1432.7 1767.26 1782.34 1771.88 ;
     RECT  1792.22 1757.18 1798.18 1771.88 ;
     RECT  3207.26 1453.72 3207.46 1772.08 ;
     RECT  2760.86 1769.76 2761.06 1772.7 ;
     RECT  2996.06 1768.5 2996.26 1773.54 ;
     RECT  1313.66 1767.68 1313.86 1773.56 ;
     RECT  2537.66 1771.22 2541.22 1774.16 ;
     RECT  976.7 1681.36 1025.86 1774.6 ;
     RECT  2589.02 1771.22 2593.06 1775.84 ;
     RECT  2737.34 1771.22 2737.54 1775.84 ;
     RECT  2436.86 1765.98 2437.06 1776.26 ;
     RECT  2589.02 1775.84 2592.1 1778.78 ;
     RECT  1170.14 1733.24 1170.34 1779.22 ;
     RECT  2757.98 1772.7 2761.06 1780.68 ;
     RECT  2774.3 1765.56 2805.22 1780.68 ;
     RECT  2874.14 1755.9 2874.34 1780.68 ;
     RECT  2591.9 1778.78 2592.1 1780.88 ;
     RECT  1342.94 1771.04 1349.86 1781.96 ;
     RECT  1342.94 1781.96 1350.34 1783.22 ;
     RECT  1313.66 1773.56 1321.06 1785.74 ;
     RECT  1371.26 1758.86 1371.46 1786.16 ;
     RECT  1408.7 1767.88 1408.9 1786.78 ;
     RECT  2541.02 1774.16 2541.22 1788.02 ;
     RECT  1342.46 1783.22 1350.34 1788.68 ;
     RECT  2901.98 1766.4 2908.42 1788.86 ;
     RECT  1423.58 1771.88 1798.18 1788.88 ;
     RECT  2874.14 1780.68 2880.58 1789.7 ;
     RECT  2851.58 1782.78 2851.78 1789.92 ;
     RECT  2949.02 1769.34 2958.34 1790.76 ;
     RECT  2996.06 1773.54 2997.22 1791.18 ;
     RECT  2996.06 1791.18 3001.54 1791.6 ;
     RECT  1432.7 1788.88 1798.18 1793.5 ;
     RECT  2949.02 1790.76 2966.02 1794.54 ;
     RECT  2880.38 1789.7 2880.58 1794.74 ;
     RECT  2920.7 1794.54 2920.9 1795.8 ;
     RECT  2986.46 1791.6 3001.54 1796.22 ;
     RECT  2757.98 1780.68 2805.22 1797.48 ;
     RECT  2920.7 1795.8 2928.58 1797.9 ;
     RECT  2757.98 1797.48 2811.46 1799.16 ;
     RECT  2901.98 1788.86 2905.06 1799.16 ;
     RECT  2704.22 1761.78 2713.06 1800.42 ;
     RECT  2986.46 1796.22 3002.98 1800.62 ;
     RECT  2898.62 1799.16 2905.06 1800.84 ;
     RECT  2917.34 1797.9 2928.58 1801.26 ;
     RECT  2948.06 1794.54 2966.02 1801.26 ;
     RECT  2845.82 1789.92 2851.78 1803.36 ;
     RECT  2704.22 1800.42 2718.34 1804.62 ;
     RECT  2756.06 1799.16 2811.46 1804.82 ;
     RECT  1371.26 1786.16 1371.94 1805.06 ;
     RECT  2838.14 1803.36 2851.78 1805.88 ;
     RECT  2916.86 1801.26 2928.58 1805.88 ;
     RECT  2756.06 1804.82 2762.5 1806.3 ;
     RECT  2776.7 1804.82 2811.46 1806.5 ;
     RECT  2895.74 1800.84 2905.06 1806.72 ;
     RECT  2916.86 1805.88 2937.22 1806.72 ;
     RECT  2948.06 1801.26 2969.86 1806.72 ;
     RECT  2823.26 1803.36 2823.46 1807.14 ;
     RECT  2838.14 1805.88 2853.7 1807.14 ;
     RECT  2916.86 1806.72 2969.86 1807.76 ;
     RECT  1313.66 1785.74 1328.74 1808.42 ;
     RECT  1342.46 1788.68 1350.82 1808.42 ;
     RECT  918.14 1725.68 918.34 1809.04 ;
     RECT  2823.26 1807.14 2853.7 1810.08 ;
     RECT  2916.86 1807.76 2920.9 1810.7 ;
     RECT  2995.58 1800.62 3002.98 1810.7 ;
     RECT  2694.62 1804.62 2718.34 1810.92 ;
     RECT  2694.62 1810.92 2723.14 1811.34 ;
     RECT  2686.46 1811.34 2723.14 1811.96 ;
     RECT  2823.26 1810.08 2856.1 1812.6 ;
     RECT  2866.46 1810.5 2874.34 1812.6 ;
     RECT  2931.74 1807.76 2969.86 1812.6 ;
     RECT  1432.7 1793.5 1788.1 1812.62 ;
     RECT  2889.02 1806.72 2905.06 1813.02 ;
     RECT  2931.74 1812.6 2975.62 1813.22 ;
     RECT  2823.26 1812.6 2874.34 1813.86 ;
     RECT  2933.18 1813.22 2975.62 1814.06 ;
     RECT  2996.06 1810.7 3002.98 1814.06 ;
     RECT  1371.26 1805.06 1372.42 1816.4 ;
     RECT  1111.58 1714.34 1111.78 1816.6 ;
     RECT  2776.7 1806.5 2790.34 1817.64 ;
     RECT  2802.14 1806.5 2811.46 1817.64 ;
     RECT  2752.7 1806.3 2762.5 1818.48 ;
     RECT  2776.7 1817.64 2811.46 1818.48 ;
     RECT  2822.3 1813.86 2874.34 1818.48 ;
     RECT  1428.86 1812.62 1788.1 1819.12 ;
     RECT  2686.46 1811.96 2694.82 1819.52 ;
     RECT  2776.7 1818.48 2874.34 1819.74 ;
     RECT  2937.02 1814.06 2975.62 1819.94 ;
     RECT  2937.02 1819.94 2974.18 1820.36 ;
     RECT  2773.34 1819.74 2874.34 1820.78 ;
     RECT  2996.06 1814.06 3001.54 1820.78 ;
     RECT  3026.3 1807.14 3026.5 1820.78 ;
     RECT  1428.86 1819.12 1730.02 1821.22 ;
     RECT  2918.3 1810.7 2920.9 1821.84 ;
     RECT  2889.02 1813.02 2906.98 1822.04 ;
     RECT  1532.06 1821.22 1730.02 1822.06 ;
     RECT  1400.06 1787 1400.26 1822.28 ;
     RECT  1416.38 1818.92 1416.58 1822.28 ;
     RECT  2939.9 1820.36 2974.18 1822.46 ;
     RECT  2940.38 1822.46 2974.18 1823.3 ;
     RECT  1532.06 1822.06 1729.54 1825 ;
     RECT  2752.7 1818.48 2762.98 1825.62 ;
     RECT  2841.98 1820.78 2874.34 1826.24 ;
     RECT  2918.3 1821.84 2922.34 1826.46 ;
     RECT  1313.66 1808.42 1350.82 1826.48 ;
     RECT  1741.82 1819.12 1788.1 1826.68 ;
     RECT  3222 1757 3470 1827 ;
     RECT  2940.38 1823.3 2972.26 1827.5 ;
     RECT  1400.06 1822.28 1416.58 1828.16 ;
     RECT  1428.86 1821.22 1522.18 1828.16 ;
     RECT  2694.62 1819.52 2694.82 1828.34 ;
     RECT  2744.06 1825.62 2762.98 1828.34 ;
     RECT  2841.98 1826.24 2842.66 1829.18 ;
     RECT  2752.7 1828.34 2762.98 1830.02 ;
     RECT  2853.5 1826.24 2874.34 1830.66 ;
     RECT  2889.02 1822.04 2903.14 1830.66 ;
     RECT  2773.34 1820.78 2832.1 1830.86 ;
     RECT  2914.94 1826.46 2922.34 1830.86 ;
     RECT  2831.9 1830.86 2832.1 1834.64 ;
     RECT  1558.46 1825 1729.54 1834.66 ;
     RECT  2657.18 1811.34 2657.38 1835.48 ;
     RECT  2707.58 1811.96 2723.14 1836.32 ;
     RECT  2841.98 1829.18 2842.18 1836.32 ;
     RECT  -70 1767 178 1837 ;
     RECT  2853.5 1830.66 2903.14 1838.22 ;
     RECT  2914.94 1830.86 2921.38 1838.22 ;
     RECT  1558.46 1834.66 1718.98 1838.44 ;
     RECT  1559.9 1838.44 1718.98 1838.86 ;
     RECT  2708.54 1836.32 2723.14 1839.06 ;
     RECT  2940.38 1827.5 2944.9 1840.32 ;
     RECT  2954.78 1827.5 2972.26 1840.32 ;
     RECT  2940.38 1840.32 2972.26 1842 ;
     RECT  2853.5 1838.22 2921.38 1842.42 ;
     RECT  2940.38 1842 2974.18 1842.42 ;
     RECT  1400.06 1828.16 1522.18 1842.44 ;
     RECT  1398.14 1842.44 1522.18 1842.64 ;
     RECT  1741.82 1826.68 1782.34 1842.64 ;
     RECT  2708.54 1839.06 2723.62 1843.04 ;
     RECT  2940.38 1842.42 2981.38 1843.26 ;
     RECT  2852.06 1842.42 2921.38 1843.88 ;
     RECT  2773.34 1830.86 2821.54 1845.14 ;
     RECT  1559.9 1838.86 1711.78 1845.16 ;
     RECT  1708.7 1845.16 1711.78 1846.84 ;
     RECT  2839.58 1838.64 2840.26 1848.92 ;
     RECT  2914.94 1843.88 2921.38 1848.92 ;
     RECT  2919.74 1848.92 2921.38 1849.34 ;
     RECT  1532.06 1825 1548.58 1850.2 ;
     RECT  2752.7 1830.02 2762.5 1851.02 ;
     RECT  2940.38 1843.26 2985.22 1851.02 ;
     RECT  2708.54 1843.04 2714.02 1851.86 ;
     RECT  2708.54 1851.86 2712.1 1853.12 ;
     RECT  2812.7 1845.14 2821.54 1853.12 ;
     RECT  2756.06 1851.02 2762.5 1853.34 ;
     RECT  2773.34 1845.14 2802.34 1853.34 ;
     RECT  2940.38 1851.02 2978.98 1853.34 ;
     RECT  2919.74 1849.34 2920.9 1853.54 ;
     RECT  3040.7 1806.72 3040.9 1853.96 ;
     RECT  2852.06 1843.88 2903.62 1854.8 ;
     RECT  2920.7 1853.54 2920.9 1855.64 ;
     RECT  2708.54 1853.12 2708.74 1856.06 ;
     RECT  2937.5 1853.34 2978.98 1856.06 ;
     RECT  2756.06 1853.34 2802.34 1856.28 ;
     RECT  2812.7 1853.12 2812.9 1856.28 ;
     RECT  2874.14 1854.8 2903.62 1856.28 ;
     RECT  2756.06 1856.28 2812.9 1856.48 ;
     RECT  2852.06 1854.8 2862.34 1856.7 ;
     RECT  2874.14 1856.28 2907.46 1856.9 ;
     RECT  2943.74 1856.06 2978.98 1856.9 ;
     RECT  2874.14 1856.9 2877.7 1857.32 ;
     RECT  2968.7 1856.9 2978.98 1857.74 ;
     RECT  1532.54 1850.2 1548.58 1857.76 ;
     RECT  1711.58 1846.84 1711.78 1858.18 ;
     RECT  2731.1 1854.18 2731.3 1859.64 ;
     RECT  2893.34 1856.9 2907.46 1860.48 ;
     RECT  3009.02 1856.7 3009.22 1860.68 ;
     RECT  2893.34 1860.48 2907.94 1860.9 ;
     RECT  2893.34 1860.9 2909.38 1861.1 ;
     RECT  2729.18 1859.64 2731.3 1861.52 ;
     RECT  1386.14 1820.18 1386.34 1861.76 ;
     RECT  1398.14 1842.64 1403.62 1861.76 ;
     RECT  1416.38 1842.64 1522.18 1862.8 ;
     RECT  2845.82 1856.7 2862.34 1864.88 ;
     RECT  1416.38 1862.8 1422.82 1864.9 ;
     RECT  2824.22 1863 2824.42 1865.52 ;
     RECT  2900.54 1861.1 2909.38 1865.72 ;
     RECT  2943.74 1856.9 2958.82 1866.78 ;
     RECT  1559.9 1845.16 1697.86 1866.8 ;
     RECT  2933.66 1866.78 2958.82 1867.4 ;
     RECT  2823.26 1865.52 2824.42 1867.82 ;
     RECT  2845.82 1864.88 2861.86 1867.82 ;
     RECT  2845.82 1867.82 2847.94 1868.04 ;
     RECT  2823.26 1867.82 2823.46 1868.66 ;
     RECT  2943.74 1867.4 2958.82 1869.08 ;
     RECT  2901.02 1865.72 2909.38 1869.5 ;
     RECT  1743.26 1842.64 1782.34 1869.52 ;
     RECT  2859.74 1867.82 2861.86 1870.34 ;
     RECT  2973.98 1857.74 2978.98 1870.56 ;
     RECT  2729.18 1861.52 2729.38 1871.18 ;
     RECT  2756.06 1856.48 2807.62 1871.18 ;
     RECT  2971.58 1870.56 2978.98 1871.4 ;
     RECT  1364.06 1816.4 1372.42 1871.42 ;
     RECT  1386.14 1861.76 1403.62 1871.42 ;
     RECT  2901.02 1869.5 2907.46 1871.6 ;
     RECT  2971.1 1871.4 2978.98 1871.6 ;
     RECT  1532.54 1857.76 1547.14 1872.88 ;
     RECT  2843.42 1868.04 2847.94 1873.28 ;
     RECT  2756.06 1871.18 2764.42 1874.12 ;
     RECT  2877.5 1857.32 2877.7 1874.12 ;
     RECT  2946.62 1869.08 2958.82 1874.54 ;
     RECT  2971.1 1871.6 2978.5 1874.54 ;
     RECT  2971.1 1874.54 2973.22 1875.38 ;
     RECT  2513.66 1863.42 2513.86 1875.8 ;
     RECT  2971.58 1875.38 2973.22 1876.22 ;
     RECT  2091.26 1849.16 2091.46 1876.46 ;
     RECT  1744.22 1869.52 1782.34 1877.08 ;
     RECT  2971.58 1876.22 2971.78 1880 ;
     RECT  2776.7 1871.18 2807.62 1881.9 ;
     RECT  2776.7 1881.9 2812.9 1882.52 ;
     RECT  2845.82 1873.28 2847.94 1883.36 ;
     RECT  2845.82 1883.36 2846.02 1884.2 ;
     RECT  2946.62 1874.54 2958.34 1886.1 ;
     RECT  2781.5 1882.52 2812.9 1886.3 ;
     RECT  1534.94 1872.88 1547.14 1886.32 ;
     RECT  3092.06 1554.74 3092.26 1889.06 ;
     RECT  2996.06 1820.78 2997.22 1890.08 ;
     RECT  1434.62 1862.8 1522.18 1891.16 ;
     RECT  1534.94 1886.32 1544.74 1891.16 ;
     RECT  698.3 1745 698.5 1892.84 ;
     RECT  2756.06 1874.12 2761.06 1893.02 ;
     RECT  2943.26 1886.1 2958.34 1893.24 ;
     RECT  2859.74 1870.34 2859.94 1894.5 ;
     RECT  1434.62 1891.16 1544.74 1894.72 ;
     RECT  2856.86 1894.5 2859.94 1894.92 ;
     RECT  2901.98 1871.6 2907.46 1895.12 ;
     RECT  2357.66 1675.28 2358.34 1895.14 ;
     RECT  691.58 1892.84 698.5 1896.2 ;
     RECT  2782.46 1886.3 2812.9 1896.38 ;
     RECT  2891.42 1887.78 2891.62 1897.44 ;
     RECT  2901.98 1895.12 2902.18 1897.44 ;
     RECT  2372.06 1856.7 2372.26 1898.48 ;
     RECT  687.26 1896.2 698.5 1899.14 ;
     RECT  2856.86 1894.92 2861.86 1899.32 ;
     RECT  2791.1 1896.38 2812.9 1899.74 ;
     RECT  2857.82 1899.32 2861.86 1899.96 ;
     RECT  2358.14 1895.14 2358.34 1900.4 ;
     RECT  2565.5 1889.88 2565.7 1901.84 ;
     RECT  976.7 1774.6 1022.02 1902.7 ;
     RECT  3092.06 1889.06 3098.98 1903.76 ;
     RECT  1744.7 1877.08 1782.34 1904.38 ;
     RECT  2940.38 1893.24 2958.34 1905.84 ;
     RECT  2978.3 1893.66 2978.5 1905.84 ;
     RECT  2501.66 1905.86 2501.86 1906.28 ;
     RECT  2940.38 1905.84 2961.22 1906.68 ;
     RECT  2501.66 1906.28 2509.06 1907.1 ;
     RECT  2891.42 1897.44 2902.18 1907.52 ;
     RECT  2940.38 1906.68 2961.7 1907.52 ;
     RECT  2977.34 1905.84 2978.5 1907.52 ;
     RECT  1558.46 1866.8 1697.86 1907.96 ;
     RECT  2891.42 1907.52 2913.7 1908.36 ;
     RECT  2793.02 1899.74 2812.9 1909.2 ;
     RECT  2997.02 1890.08 2997.22 1909.2 ;
     RECT  2832.38 1907.1 2840.74 1909.62 ;
     RECT  2877.02 1906.52 2878.66 1909.62 ;
     RECT  2891.42 1908.36 2919.46 1909.62 ;
     RECT  1364.06 1871.42 1403.62 1910.26 ;
     RECT  2940.38 1907.52 2978.5 1910.88 ;
     RECT  2994.62 1909.2 2997.22 1910.88 ;
     RECT  2940.38 1910.88 2997.22 1911.3 ;
     RECT  1744.7 1904.38 1761.7 1911.52 ;
     RECT  2832.38 1909.62 2847.46 1911.72 ;
     RECT  2857.82 1899.96 2867.14 1911.72 ;
     RECT  3070.46 1898.72 3070.66 1911.74 ;
     RECT  3085.34 1903.76 3098.98 1911.74 ;
     RECT  2877.02 1909.62 2919.46 1912.98 ;
     RECT  2933.18 1911.3 2997.22 1912.98 ;
     RECT  682.94 1899.14 698.5 1914.26 ;
     RECT  2832.38 1911.72 2867.14 1914.66 ;
     RECT  2877.02 1912.98 2997.22 1914.66 ;
     RECT  681.5 1914.26 698.5 1915.1 ;
     RECT  2793.02 1909.2 2821.54 1916.76 ;
     RECT  2832.38 1914.66 2997.22 1916.76 ;
     RECT  2757.98 1893.02 2761.06 1916.96 ;
     RECT  976.7 1902.7 1010.5 1917.4 ;
     RECT  2793.02 1916.76 2997.22 1921.16 ;
     RECT  983.9 1917.4 1010.5 1921.6 ;
     RECT  681.5 1915.1 703.78 1922.24 ;
     RECT  994.46 1921.6 1010.5 1922.86 ;
     RECT  2463.26 1911.32 2463.46 1923.06 ;
     RECT  1021.82 1902.7 1022.02 1923.28 ;
     RECT  2699.9 1912.56 2700.1 1924.52 ;
     RECT  2501.66 1907.1 2517.22 1925.16 ;
     RECT  1434.62 1894.72 1538.98 1925.8 ;
     RECT  2358.14 1900.4 2358.82 1927.28 ;
     RECT  2371.1 1923.92 2371.3 1927.28 ;
     RECT  2454.14 1923.06 2463.46 1927.88 ;
     RECT  2821.34 1921.16 2997.22 1927.88 ;
     RECT  736.7 1837.82 736.9 1928.96 ;
     RECT  1422.62 1864.9 1422.82 1930 ;
     RECT  681.5 1922.24 704.26 1930.22 ;
     RECT  2757.98 1916.96 2758.66 1930.82 ;
     RECT  983.9 1921.6 984.1 1930.84 ;
     RECT  2793.02 1921.16 2810.02 1931.46 ;
     RECT  2821.34 1927.88 2981.86 1931.46 ;
     RECT  2793.02 1931.46 2981.86 1931.66 ;
     RECT  2757.98 1930.82 2758.18 1932.08 ;
     RECT  994.46 1922.86 1006.66 1932.52 ;
     RECT  1509.02 1925.8 1538.98 1933.16 ;
     RECT  1554.14 1907.96 1697.86 1933.16 ;
     RECT  2793.02 1931.66 2793.22 1935.86 ;
     RECT  2994.62 1927.88 2997.22 1935.86 ;
     RECT  722.78 1935.68 722.98 1936.1 ;
     RECT  736.7 1928.96 745.06 1936.1 ;
     RECT  2994.62 1935.86 2994.82 1936.28 ;
     RECT  722.78 1936.1 745.06 1936.52 ;
     RECT  997.82 1932.52 1006.66 1937.14 ;
     RECT  2686.46 1936.52 2688.1 1937.28 ;
     RECT  2629.82 1932.3 2630.02 1937.34 ;
     RECT  2640.38 1749.7 2640.58 1937.34 ;
     RECT  1434.62 1925.8 1498.66 1937.78 ;
     RECT  1509.02 1933.16 1697.86 1937.78 ;
     RECT  999.26 1937.14 1000.9 1938.4 ;
     RECT  2629.82 1937.34 2640.58 1938.62 ;
     RECT  2629.82 1938.62 2645.86 1938.82 ;
     RECT  2803.1 1931.66 2981.86 1939.22 ;
     RECT  2803.1 1939.22 2881.54 1939.64 ;
     RECT  2629.82 1938.82 2631.94 1939.86 ;
     RECT  1364.06 1910.26 1400.26 1940.3 ;
     RECT  2501.66 1925.16 2520.1 1940.48 ;
     RECT  2620.22 1939.86 2631.94 1940.48 ;
     RECT  1000.7 1938.4 1000.9 1940.5 ;
     RECT  1363.1 1940.3 1400.26 1940.72 ;
     RECT  2804.06 1939.64 2881.54 1942.16 ;
     RECT  2821.34 1942.16 2881.54 1942.58 ;
     RECT  2415.26 1942.4 2415.46 1942.82 ;
     RECT  2829.5 1942.58 2881.54 1943 ;
     RECT  2411.9 1942.82 2415.46 1943.24 ;
     RECT  2891.9 1939.22 2981.86 1943.64 ;
     RECT  2891.9 1943.64 2987.62 1943.84 ;
     RECT  2845.82 1943 2881.54 1944.26 ;
     RECT  2896.22 1943.84 2987.62 1944.26 ;
     RECT  2358.14 1927.28 2371.3 1944.5 ;
     RECT  2896.22 1944.26 2919.94 1945.52 ;
     RECT  2932.22 1944.26 2987.62 1946.16 ;
     RECT  2845.82 1944.26 2880.58 1946.78 ;
     RECT  2358.14 1944.5 2380.42 1947.86 ;
     RECT  2394.14 1947.02 2394.34 1947.86 ;
     RECT  2932.22 1946.16 2988.1 1948.26 ;
     RECT  1773.02 1904.38 1782.34 1948.28 ;
     RECT  680.54 1930.22 704.26 1948.7 ;
     RECT  2932.22 1948.26 2994.82 1948.88 ;
     RECT  1363.1 1940.72 1400.74 1949.12 ;
     RECT  2949.5 1948.88 2994.82 1949.72 ;
     RECT  2848.22 1946.78 2880.58 1950.14 ;
     RECT  2849.66 1950.14 2880.58 1950.56 ;
     RECT  2519.9 1940.48 2520.1 1950.98 ;
     RECT  3222 1827 3400 1951 ;
     RECT  2933.18 1948.88 2933.38 1951.82 ;
     RECT  722.3 1936.52 745.06 1952.9 ;
     RECT  2520.86 1952.9 2521.06 1953.04 ;
     RECT  2949.5 1949.72 2981.86 1953.08 ;
     RECT  2501.66 1940.48 2509.06 1953.1 ;
     RECT  2520.86 1953.04 2524.9 1953.24 ;
     RECT  680.54 1948.7 709.06 1953.32 ;
     RECT  721.82 1952.9 745.06 1953.32 ;
     RECT  2645.66 1938.82 2645.86 1953.74 ;
     RECT  2992.7 1949.72 2994.82 1953.92 ;
     RECT  2657.66 1936.52 2657.86 1953.94 ;
     RECT  2609.66 1749.4 2609.86 1954.58 ;
     RECT  2620.22 1940.48 2630.02 1954.76 ;
     RECT  2524.7 1953.24 2524.9 1954.78 ;
     RECT  669.02 1910.06 669.22 1955.42 ;
     RECT  2896.22 1945.52 2916.58 1955.6 ;
     RECT  2949.5 1953.08 2961.22 1955.6 ;
     RECT  2851.1 1950.56 2880.58 1956.02 ;
     RECT  2829.5 1943 2831.14 1956.44 ;
     RECT  2896.22 1955.6 2898.82 1956.86 ;
     RECT  2994.62 1953.92 2994.82 1956.86 ;
     RECT  2629.82 1954.76 2630.02 1957.7 ;
     RECT  2830.94 1956.44 2831.14 1957.7 ;
     RECT  2851.1 1956.02 2868.58 1957.7 ;
     RECT  2880.38 1956.02 2880.58 1957.7 ;
     RECT  2972.06 1953.08 2981.86 1957.7 ;
     RECT  2411.9 1943.24 2415.94 1957.92 ;
     RECT  1421.66 1947.44 1421.86 1958.36 ;
     RECT  2910.14 1955.6 2916.58 1959.8 ;
     RECT  2956.7 1955.6 2961.22 1959.8 ;
     RECT  2405.18 1957.92 2415.94 1960.08 ;
     RECT  2642.3 1953.74 2645.86 1960.08 ;
     RECT  668.54 1955.42 669.22 1960.88 ;
     RECT  680.54 1953.32 745.06 1960.88 ;
     RECT  0 1837 178 1961 ;
     RECT  3070.46 1911.74 3098.98 1962.14 ;
     RECT  2358.14 1947.86 2394.34 1962.98 ;
     RECT  1772.54 1948.28 1782.34 1964.86 ;
     RECT  2972.06 1957.7 2972.26 1965.26 ;
     RECT  1421.66 1958.36 1423.3 1965.5 ;
     RECT  1434.62 1937.78 1697.86 1965.5 ;
     RECT  2405.18 1960.08 2405.38 1965.68 ;
     RECT  2958.14 1959.8 2961.22 1965.68 ;
     RECT  1421.66 1965.5 1697.86 1965.7 ;
     RECT  2491.58 1949.1 2491.78 1968.42 ;
     RECT  2501.66 1953.1 2501.86 1968.42 ;
     RECT  2566.46 1957.5 2566.66 1969.68 ;
     RECT  2355.74 1962.98 2394.34 1970.74 ;
     RECT  2851.1 1957.7 2861.86 1973.88 ;
     RECT  2566.46 1969.68 2572.9 1974.5 ;
     RECT  2851.1 1973.88 2865.22 1974.92 ;
     RECT  2852.54 1974.92 2865.22 1975.76 ;
     RECT  2757.98 1969.26 2758.18 1976.4 ;
     RECT  1708.22 1864.7 1708.42 1976.84 ;
     RECT  2491.58 1968.42 2501.86 1979.54 ;
     RECT  1363.1 1949.12 1410.34 1979.98 ;
     RECT  2494.46 1979.54 2501.86 1980.8 ;
     RECT  2853.98 1975.76 2865.22 1980.8 ;
     RECT  2853.98 1980.8 2857.54 1982.06 ;
     RECT  668.54 1960.88 745.06 1982.3 ;
     RECT  2896.7 1956.86 2898.82 1983.32 ;
     RECT  2958.62 1965.68 2961.22 1983.32 ;
     RECT  2358.14 1970.74 2394.34 1985.66 ;
     RECT  2804.06 1942.16 2806.18 1986.68 ;
     RECT  2757.98 1976.4 2759.62 1988.36 ;
     RECT  1421.66 1965.7 1656.1 1990.48 ;
     RECT  2757.98 1988.36 2758.18 1992.56 ;
     RECT  2961.02 1983.32 2961.22 1992.98 ;
     RECT  1708.22 1976.84 1717.06 1993 ;
     RECT  1773.02 1964.86 1782.34 1993.64 ;
     RECT  2910.14 1959.8 2910.34 1995.92 ;
     RECT  2680.22 1961.7 2680.42 1996.34 ;
     RECT  2805.98 1986.68 2806.18 1996.76 ;
     RECT  2898.62 1983.32 2898.82 1998.86 ;
     RECT  2857.34 1982.06 2857.54 2003.9 ;
     RECT  2566.46 1974.5 2566.66 2004.32 ;
     RECT  668.06 1982.3 745.06 2005.4 ;
     RECT  2448.86 2007.76 2451.46 2008.34 ;
     RECT  2555.42 2007.92 2555.62 2008.34 ;
     RECT  3057.98 1935.26 3058.18 2008.34 ;
     RECT  3070.46 1962.14 3100.9 2008.34 ;
     RECT  1773.02 1993.64 1785.22 2008.96 ;
     RECT  2448.38 2008.34 2451.46 2010.24 ;
     RECT  1421.66 1990.48 1655.14 2010.44 ;
     RECT  1665.98 1965.7 1697.86 2010.44 ;
     RECT  1716.86 1993 1717.06 2012.12 ;
     RECT  1744.7 1911.52 1756.9 2013.8 ;
     RECT  2415.26 1960.08 2415.94 2016.1 ;
     RECT  2443.1 2015.9 2443.3 2016.32 ;
     RECT  1307.42 1826.48 1350.82 2016.475 ;
     RECT  2415.74 2016.1 2415.94 2016.52 ;
     RECT  2442.62 2016.32 2443.3 2016.74 ;
     RECT  2546.78 2008.34 2555.62 2016.88 ;
     RECT  2568.86 2016.74 2578.66 2016.88 ;
     RECT  2442.14 2016.74 2443.3 2017.16 ;
     RECT  2358.14 1985.66 2402.5 2017.36 ;
     RECT  2441.66 2017.16 2443.3 2017.58 ;
     RECT  2857.82 2008.32 2858.02 2018.82 ;
     RECT  2869.34 2016.72 2869.54 2018.82 ;
     RECT  2429.66 2016.74 2429.86 2019.16 ;
     RECT  2441.18 2017.58 2443.3 2019.16 ;
     RECT  2371.1 2017.36 2402.5 2019.88 ;
     RECT  2429.66 2019.16 2443.3 2019.88 ;
     RECT  2523.26 2020.1 2523.46 2020.52 ;
     RECT  3222 1951 3470 2021 ;
     RECT  2434.94 2019.88 2443.3 2021.56 ;
     RECT  2546.78 2016.88 2579.14 2021.64 ;
     RECT  2463.26 1927.88 2463.46 2021.98 ;
     RECT  2546.78 2021.64 2563.78 2021.98 ;
     RECT  2523.26 2020.52 2530.66 2022.62 ;
     RECT  2523.26 2022.62 2531.62 2023.04 ;
     RECT  2645.66 1960.08 2645.86 2023.04 ;
     RECT  2602.46 1954.58 2609.86 2023.24 ;
     RECT  2314.46 1668.56 2315.62 2027.02 ;
     RECT  2434.94 2021.56 2440.9 2027.02 ;
     RECT  2768.06 2022.6 2768.26 2027.84 ;
     RECT  1305.18 2016.475 1350.82 2027.875 ;
     RECT  2693.66 1999.92 2693.86 2030.36 ;
     RECT  1302.58 2027.875 1350.82 2030.6 ;
     RECT  -70 1961 178 2031 ;
     RECT  2638.46 2023.04 2645.86 2033.1 ;
     RECT  2824.22 1992.36 2824.42 2036.88 ;
     RECT  1302.58 2030.6 1351.3 2041.1 ;
     RECT  2857.82 2018.82 2869.54 2045.48 ;
     RECT  2857.82 2045.48 2863.3 2050.52 ;
     RECT  1421.66 2010.44 1697.86 2051.8 ;
     RECT  2546.78 2021.98 2563.3 2051.9 ;
     RECT  2573.66 2021.64 2579.14 2051.9 ;
     RECT  2602.46 2023.24 2602.66 2051.9 ;
     RECT  2380.22 2019.88 2402.5 2052.1 ;
     RECT  2516.06 2023.04 2531.62 2052.1 ;
     RECT  2602.46 2051.9 2605.06 2052.1 ;
     RECT  2824.22 2036.88 2824.9 2052.42 ;
     RECT  2632.22 2033.1 2645.86 2052.62 ;
     RECT  1422.14 2051.8 1697.86 2055.16 ;
     RECT  2810.3 2007.9 2810.5 2058.5 ;
     RECT  2501.66 1980.8 2501.86 2058.72 ;
     RECT  2821.34 2052.42 2824.9 2060.82 ;
     RECT  2863.1 2050.52 2863.3 2060.82 ;
     RECT  2696.06 2058.72 2696.26 2061.44 ;
     RECT  2946.62 2052.84 2946.82 2063.96 ;
     RECT  2863.1 2060.82 2868.58 2064.18 ;
     RECT  2382.62 2052.1 2402.5 2064.4 ;
     RECT  2382.62 2064.4 2386.66 2064.62 ;
     RECT  2483.9 2064.2 2484.1 2064.62 ;
     RECT  2381.66 2064.62 2386.66 2064.76 ;
     RECT  1364.06 1979.98 1410.34 2066.3 ;
     RECT  1422.14 2055.16 1693.06 2066.3 ;
     RECT  2472.86 2033.96 2473.06 2066.72 ;
     RECT  2815.58 2060.82 2824.9 2067.12 ;
     RECT  2863.1 2064.18 2872.9 2067.12 ;
     RECT  2358.14 2017.36 2359.3 2067.34 ;
     RECT  2863.1 2067.12 2875.3 2067.96 ;
     RECT  2815.58 2067.12 2826.34 2068.16 ;
     RECT  2863.1 2067.96 2880.1 2068.38 ;
     RECT  1713.98 2012.12 1717.06 2069.44 ;
     RECT  2378.3 2064.76 2386.66 2069.52 ;
     RECT  2483.9 2064.62 2484.58 2069.66 ;
     RECT  2382.14 2069.52 2386.66 2069.86 ;
     RECT  2467.58 2066.72 2473.06 2070.08 ;
     RECT  2483.9 2069.66 2491.3 2070.08 ;
     RECT  2359.1 2067.34 2359.3 2072.38 ;
     RECT  2718.62 2062.92 2718.82 2072.78 ;
     RECT  1364.06 2066.3 1693.06 2073.44 ;
     RECT  1364.06 2073.44 1697.86 2077.42 ;
     RECT  2861.18 2068.38 2880.1 2077.82 ;
     RECT  910.62 2072.98 910.82 2080.96 ;
     RECT  2937.5 2082.26 2937.7 2082.68 ;
     RECT  2937.02 2082.68 2937.7 2083 ;
     RECT  2861.18 2077.82 2874.34 2084.12 ;
     RECT  2934.62 2083 2937.7 2084.78 ;
     RECT  2861.18 2084.12 2872.9 2085.18 ;
     RECT  1773.02 2008.96 1782.34 2087.72 ;
     RECT  2658.14 2075.52 2658.34 2089.58 ;
     RECT  1364.06 2077.42 1378.66 2090.24 ;
     RECT  1390.46 2077.42 1697.86 2090.24 ;
     RECT  2501.66 2058.72 2506.18 2090.42 ;
     RECT  1300.22 2041.1 1351.3 2091.5 ;
     RECT  2519.9 2052.1 2531.62 2092.12 ;
     RECT  2546.78 2051.9 2582.02 2092.12 ;
     RECT  1300.22 2091.5 1353.7 2092.34 ;
     RECT  1364.06 2090.24 1697.86 2092.34 ;
     RECT  2467.58 2070.08 2491.3 2098 ;
     RECT  952.86 2078.44 953.06 2098.6 ;
     RECT  2638.46 2052.62 2645.86 2098.64 ;
     RECT  2934.62 2084.78 2941.06 2098.64 ;
     RECT  2604.86 2052.1 2605.06 2098.84 ;
     RECT  2483.9 2098 2491.3 2099.26 ;
     RECT  1773.02 2087.72 1787.62 2099.68 ;
     RECT  2467.58 2098 2473.06 2099.68 ;
     RECT  952.86 2098.6 953.54 2100.06 ;
     RECT  2467.58 2099.68 2467.78 2100.1 ;
     RECT  952.86 2100.06 953.06 2100.48 ;
     RECT  2484.38 2099.26 2491.3 2100.52 ;
     RECT  886.62 2045.68 886.82 2100.7 ;
     RECT  2491.1 2100.52 2491.3 2100.94 ;
     RECT  2816.06 2068.16 2826.34 2102.18 ;
     RECT  3057.98 2008.34 3100.9 2102.5 ;
     RECT  618.14 2069.24 618.34 2103.46 ;
     RECT  2400.86 2064.4 2402.5 2103.46 ;
     RECT  2442.62 2102.3 2446.18 2103.88 ;
     RECT  2402.3 2103.46 2402.5 2104.3 ;
     RECT  2858.78 2085.18 2872.9 2104.7 ;
     RECT  2519.9 2092.12 2582.02 2106.4 ;
     RECT  2382.62 2069.86 2386.66 2107.66 ;
     RECT  2519.9 2106.4 2535.94 2108.5 ;
     RECT  2860.22 2104.7 2863.3 2108.9 ;
     RECT  2452.7 2108.7 2452.9 2111.66 ;
     RECT  843.42 2109.1 843.62 2114.76 ;
     RECT  2860.22 2108.9 2860.9 2115.84 ;
     RECT  1300.22 2092.34 1697.86 2116.7 ;
     RECT  2546.78 2106.4 2582.02 2117.12 ;
     RECT  2546.78 2117.12 2588.26 2117.54 ;
     RECT  2519.9 2108.5 2534.98 2118.58 ;
     RECT  2519.9 2118.58 2520.1 2118.8 ;
     RECT  2519.42 2118.8 2520.1 2119.22 ;
     RECT  2501.66 2090.42 2502.34 2119.42 ;
     RECT  2616.86 2119.64 2617.06 2120.06 ;
     RECT  2616.86 2120.06 2625.7 2120.48 ;
     RECT  2517.5 2119.22 2520.1 2120.68 ;
     RECT  2616.86 2120.48 2628.1 2120.9 ;
     RECT  2502.14 2119.42 2502.34 2121.52 ;
     RECT  2546.78 2117.54 2596.42 2121.74 ;
     RECT  2609.66 2120.9 2628.1 2121.74 ;
     RECT  2517.5 2120.68 2519.62 2121.96 ;
     RECT  2858.78 2115.84 2860.9 2122.34 ;
     RECT  2546.78 2121.74 2628.1 2122.58 ;
     RECT  2638.46 2098.64 2646.34 2122.58 ;
     RECT  2530.46 2118.58 2534.98 2123.2 ;
     RECT  2546.78 2122.58 2646.34 2123.84 ;
     RECT  2663.9 2121.74 2664.1 2123.84 ;
     RECT  2440.22 2122.98 2440.42 2124.02 ;
     RECT  2544.86 2123.84 2646.34 2124.04 ;
     RECT  2378.78 2109.54 2378.98 2124.66 ;
     RECT  2378.78 2124.66 2384.26 2124.86 ;
     RECT  2646.14 2124.04 2646.34 2126.32 ;
     RECT  2656.22 2123.84 2664.1 2126.32 ;
     RECT  2544.86 2124.04 2631.46 2126.52 ;
     RECT  2858.78 2122.34 2860.42 2128.86 ;
     RECT  2816.06 2102.18 2824.42 2129.06 ;
     RECT  954.78 2125.9 954.98 2130.1 ;
     RECT  2920.7 2111.66 2920.9 2132.24 ;
     RECT  2932.22 2098.64 2941.06 2132.24 ;
     RECT  2877.98 2133.92 2878.18 2134.34 ;
     RECT  1299.26 2116.7 1697.86 2134.76 ;
     RECT  2877.98 2134.34 2882.02 2134.76 ;
     RECT  2877.5 2134.76 2882.02 2135.18 ;
     RECT  2877.5 2135.18 2882.98 2136.86 ;
     RECT  2877.5 2136.86 2887.3 2137.7 ;
     RECT  2850.14 2128.86 2860.42 2141.48 ;
     RECT  668.06 2005.4 752.74 2142.1 ;
     RECT  2920.7 2132.24 2941.06 2142.1 ;
     RECT  2934.62 2142.1 2941.06 2142.48 ;
     RECT  1299.26 2134.76 1702.66 2142.52 ;
     RECT  2920.7 2142.1 2923.3 2142.52 ;
     RECT  1166.46 2136.4 1166.66 2142.7 ;
     RECT  2920.7 2142.52 2920.9 2142.94 ;
     RECT  2718.62 2101.14 2718.82 2143.34 ;
     RECT  752.06 2142.1 752.74 2144.2 ;
     RECT  3222 2021 3400 2145 ;
     RECT  952.38 2130.1 954.98 2146.48 ;
     RECT  2850.14 2141.48 2867.14 2147.12 ;
     RECT  1740.38 2013.8 1756.9 2148.82 ;
     RECT  897.66 2093.56 897.86 2149 ;
     RECT  910.62 2080.96 914.66 2149 ;
     RECT  1153.02 2149 1154.18 2149.76 ;
     RECT  2824.22 2129.06 2824.42 2150.06 ;
     RECT  1299.26 2142.52 1378.66 2150.08 ;
     RECT  834.78 2137.66 834.98 2151.1 ;
     RECT  880.86 2100.7 886.82 2151.1 ;
     RECT  897.66 2149 914.66 2151.1 ;
     RECT  1165.02 2142.7 1166.66 2152.14 ;
     RECT  880.86 2151.1 914.66 2152.36 ;
     RECT  952.38 2146.48 955.46 2152.56 ;
     RECT  1125.66 2152.36 1125.86 2153.62 ;
     RECT  2742.62 1936.52 2742.82 2153.88 ;
     RECT  834.78 2151.1 839.78 2154.46 ;
     RECT  1165.02 2152.14 1165.22 2154.46 ;
     RECT  0 2031 178 2155 ;
     RECT  834.78 2154.46 847.46 2156.56 ;
     RECT  2384.06 2124.86 2384.26 2156.78 ;
     RECT  2850.14 2147.12 2850.34 2158.24 ;
     RECT  2865.5 2147.12 2867.14 2158.24 ;
     RECT  952.38 2152.56 954.98 2159.28 ;
     RECT  2452.7 2111.66 2457.22 2159.3 ;
     RECT  2850.14 2158.24 2867.14 2159.3 ;
     RECT  877.5 2152.36 914.66 2160.34 ;
     RECT  2646.14 2126.32 2664.1 2160.72 ;
     RECT  2940.86 2142.48 2941.06 2160.72 ;
     RECT  2530.46 2123.2 2530.66 2163.32 ;
     RECT  2437.34 2133.5 2437.54 2163.52 ;
     RECT  2544.86 2126.52 2545.06 2163.74 ;
     RECT  2555.42 2126.52 2631.46 2163.74 ;
     RECT  2646.14 2160.72 2646.34 2163.94 ;
     RECT  1027.26 2156.98 1027.46 2164.12 ;
     RECT  2732.54 2163.74 2732.74 2164.16 ;
     RECT  2656.22 2160.72 2664.1 2164.36 ;
     RECT  2544.86 2163.74 2631.46 2164.78 ;
     RECT  1125.66 2153.62 1132.1 2164.96 ;
     RECT  1163.1 2154.46 1165.22 2164.96 ;
     RECT  1125.18 2164.96 1132.1 2165.38 ;
     RECT  1142.46 2160.34 1142.66 2165.38 ;
     RECT  834.78 2156.56 858.02 2166.42 ;
     RECT  2544.86 2164.78 2625.7 2166.46 ;
     RECT  847.26 2166.42 856.1 2167.26 ;
     RECT  1160.7 2164.96 1165.22 2167.26 ;
     RECT  2663.9 2164.36 2664.1 2167.3 ;
     RECT  2877.5 2137.7 2890.66 2167.3 ;
     RECT  1027.26 2164.12 1031.3 2167.48 ;
     RECT  2857.34 2159.3 2867.14 2167.52 ;
     RECT  2877.5 2167.3 2879.62 2167.52 ;
     RECT  3057.98 2102.5 3099.46 2167.56 ;
     RECT  1160.7 2167.26 1163.3 2167.9 ;
     RECT  2544.86 2166.46 2624.74 2168.14 ;
     RECT  2808.86 2167.36 2810.02 2168.14 ;
     RECT  2890.46 2167.3 2890.66 2168.14 ;
     RECT  759.9 2151.1 760.1 2168.32 ;
     RECT  929.34 2133.88 929.54 2168.32 ;
     RECT  1125.18 2165.38 1142.66 2168.32 ;
     RECT  1153.02 2167.9 1163.3 2168.32 ;
     RECT  952.38 2159.28 952.58 2168.52 ;
     RECT  2544.86 2168.14 2563.3 2168.56 ;
     RECT  926.46 2168.32 929.54 2169.16 ;
     RECT  2580.86 2168.14 2624.74 2169.4 ;
     RECT  2624.06 2169.4 2624.74 2170.24 ;
     RECT  2580.86 2169.4 2609.86 2170.66 ;
     RECT  926.46 2169.16 933.38 2170.84 ;
     RECT  2441.66 2167.36 2444.26 2170.88 ;
     RECT  2523.26 2163.32 2530.66 2170.88 ;
     RECT  2581.82 2170.66 2609.86 2171.08 ;
     RECT  2521.82 2170.88 2530.66 2171.3 ;
     RECT  2544.86 2168.56 2547.94 2171.3 ;
     RECT  2624.06 2170.24 2624.26 2171.92 ;
     RECT  759.9 2168.32 769.22 2172.3 ;
     RECT  2559.74 2168.56 2563.3 2172.34 ;
     RECT  2857.34 2167.52 2879.62 2172.76 ;
     RECT  2732.06 2164.16 2732.74 2173.18 ;
     RECT  2857.34 2172.76 2858.98 2173.18 ;
     RECT  802.14 2152.78 802.34 2173.56 ;
     RECT  1125.18 2168.32 1163.3 2173.56 ;
     RECT  1390.46 2142.52 1702.66 2173.82 ;
     RECT  1713.98 2069.44 1714.18 2173.82 ;
     RECT  2691.26 2167.1 2691.46 2174.24 ;
     RECT  2441.66 2170.88 2444.74 2174.4 ;
     RECT  2588.06 2171.08 2609.86 2174.44 ;
     RECT  668.06 2142.1 736.9 2174.86 ;
     RECT  2588.06 2174.44 2602.66 2174.86 ;
     RECT  2735.9 2174.66 2736.1 2175.08 ;
     RECT  1131.9 2173.56 1163.3 2175.24 ;
     RECT  2602.46 2174.86 2602.66 2175.28 ;
     RECT  847.26 2167.26 847.46 2175.66 ;
     RECT  2691.26 2174.24 2692.9 2175.7 ;
     RECT  2588.06 2174.86 2588.26 2176.68 ;
     RECT  3207.26 1965.08 3207.46 2176.68 ;
     RECT  1025.82 2167.48 1031.3 2176.72 ;
     RECT  870.3 2160.34 914.66 2177.34 ;
     RECT  1752.86 2148.82 1756.9 2178.22 ;
     RECT  2874.62 2172.76 2879.62 2178.86 ;
     RECT  668.06 2174.86 731.62 2179.06 ;
     RECT  926.46 2170.84 937.22 2179.24 ;
     RECT  897.66 2177.34 914.66 2179.66 ;
     RECT  3057.98 2167.56 3073.06 2179.9 ;
     RECT  1390.46 2173.82 1714.18 2180.32 ;
     RECT  2454.62 2159.3 2457.22 2181.56 ;
     RECT  2858.78 2173.18 2858.98 2181.58 ;
     RECT  2874.62 2178.86 2880.1 2181.58 ;
     RECT  1025.34 2176.72 1031.3 2181.76 ;
     RECT  1002.78 2154.46 1002.98 2182.18 ;
     RECT  2819.42 2181.8 2819.62 2182.22 ;
     RECT  2723.9 2174.24 2724.1 2182.42 ;
     RECT  2735.9 2175.08 2736.58 2182.84 ;
     RECT  834.78 2166.42 834.98 2183.02 ;
     RECT  870.3 2177.34 886.82 2183.22 ;
     RECT  1131.9 2175.24 1160.9 2183.22 ;
     RECT  2832.38 2163.32 2832.58 2183.26 ;
     RECT  2818.94 2182.22 2819.62 2183.32 ;
     RECT  2874.62 2181.58 2879.14 2183.68 ;
     RECT  3084.86 2167.56 3099.46 2183.68 ;
     RECT  1142.46 2183.22 1160.9 2184.06 ;
     RECT  668.06 2179.06 731.14 2184.1 ;
     RECT  2878.94 2183.68 2879.14 2184.1 ;
     RECT  3085.82 2183.68 3099.46 2184.1 ;
     RECT  970.62 2152.78 970.82 2184.28 ;
     RECT  2815.1 2183.32 2819.62 2185.16 ;
     RECT  1025.34 2181.76 1038.02 2185.32 ;
     RECT  2814.14 2185.16 2819.62 2185.8 ;
     RECT  995.58 2182.18 1002.98 2186.16 ;
     RECT  1145.82 2184.06 1160.9 2187 ;
     RECT  882.78 2183.22 886.82 2187.22 ;
     RECT  897.66 2179.66 915.14 2187.22 ;
     RECT  997.98 2186.16 1002.98 2188.26 ;
     RECT  2819.42 2185.8 2819.62 2189.14 ;
     RECT  1421.66 2180.32 1714.18 2189.56 ;
     RECT  1131.9 2183.22 1132.1 2189.74 ;
     RECT  2736.38 2182.84 2736.58 2189.98 ;
     RECT  1126.14 2189.74 1132.1 2190.16 ;
     RECT  1027.26 2185.32 1038.02 2191.62 ;
     RECT  969.66 2184.28 970.82 2192.04 ;
     RECT  1027.26 2191.62 1031.3 2192.04 ;
     RECT  1028.22 2192.04 1031.3 2192.88 ;
     RECT  870.3 2183.22 870.5 2193.72 ;
     RECT  1390.46 2180.32 1411.3 2193.76 ;
     RECT  635.42 2012.12 635.62 2195.66 ;
     RECT  1172.7 2193.94 1172.9 2196.04 ;
     RECT  1145.82 2187 1153.22 2197.08 ;
     RECT  635.42 2195.66 638.98 2197.76 ;
     RECT  1170.78 2196.04 1172.9 2200.02 ;
     RECT  998.94 2188.26 1002.98 2200.44 ;
     RECT  1145.82 2197.08 1146.02 2200.86 ;
     RECT  2605.82 2184.3 2606.02 2200.88 ;
     RECT  834.78 2183.02 838.34 2201.5 ;
     RECT  863.1 2195.62 863.3 2201.5 ;
     RECT  882.78 2187.22 915.14 2201.5 ;
     RECT  925.5 2179.24 937.22 2201.5 ;
     RECT  956.7 2194.78 956.9 2201.5 ;
     RECT  1028.22 2192.88 1029.86 2201.7 ;
     RECT  1119.42 2190.16 1132.1 2201.7 ;
     RECT  769.02 2172.3 769.22 2202.34 ;
     RECT  834.78 2201.5 847.94 2202.34 ;
     RECT  1170.78 2200.02 1170.98 2202.54 ;
     RECT  2691.26 2175.7 2691.46 2203 ;
     RECT  2521.82 2171.3 2547.94 2204.04 ;
     RECT  3086.3 2184.1 3099.46 2204.04 ;
     RECT  816.06 2100.28 816.26 2205.28 ;
     RECT  827.1 2202.34 847.94 2205.28 ;
     RECT  1119.42 2201.7 1126.34 2205.9 ;
     RECT  859.26 2201.5 863.3 2208.22 ;
     RECT  859.26 2208.22 866.66 2208.64 ;
     RECT  879.9 2201.5 937.22 2208.64 ;
     RECT  766.14 2202.34 769.22 2209.9 ;
     RECT  2508.86 2164.16 2509.06 2210.88 ;
     RECT  2541.5 2204.04 2547.94 2211.82 ;
     RECT  2611.1 2201.94 2611.3 2212.22 ;
     RECT  2541.5 2211.82 2546.98 2212.24 ;
     RECT  2559.74 2172.34 2559.94 2212.66 ;
     RECT  2521.82 2204.04 2530.66 2213.08 ;
     RECT  3222 2145 3470 2215 ;
     RECT  2541.5 2212.24 2541.7 2215.6 ;
     RECT  2521.82 2213.08 2523.46 2216.02 ;
     RECT  859.26 2208.64 937.22 2216.2 ;
     RECT  2521.82 2216.02 2522.02 2216.44 ;
     RECT  859.26 2216.2 937.7 2216.82 ;
     RECT  816.06 2205.28 847.94 2217.24 ;
     RECT  998.94 2200.44 999.14 2217.24 ;
     RECT  1740.38 2148.82 1740.58 2217.5 ;
     RECT  1421.66 2189.56 1655.14 2217.7 ;
     RECT  2436.86 2197 2437.06 2217.72 ;
     RECT  3066.62 2179.9 3073.06 2217.72 ;
     RECT  956.7 2201.5 957.38 2217.88 ;
     RECT  1446.62 2217.7 1655.14 2219.8 ;
     RECT  1665.5 2189.56 1714.18 2220.64 ;
     RECT  1390.46 2193.76 1410.34 2220.86 ;
     RECT  1421.66 2217.7 1436.74 2220.86 ;
     RECT  2405.66 2220.86 2405.86 2224.64 ;
     RECT  2457.02 2181.56 2457.22 2224.84 ;
     RECT  2591.42 2224.36 2599.3 2224.84 ;
     RECT  -70 2155 178 2225 ;
     RECT  2405.18 2224.64 2405.86 2227.16 ;
     RECT  861.18 2216.82 937.7 2228.58 ;
     RECT  1773.02 2099.68 1782.34 2228.84 ;
     RECT  1765.82 2228.84 1782.34 2229.12 ;
     RECT  861.18 2228.58 886.34 2230.48 ;
     RECT  2405.18 2227.16 2412.58 2231.78 ;
     RECT  1390.46 2220.86 1436.74 2231.9 ;
     RECT  1446.62 2219.8 1504.42 2231.9 ;
     RECT  897.66 2228.58 937.7 2232.36 ;
     RECT  1515.74 2219.8 1655.14 2232.4 ;
     RECT  954.78 2217.88 957.38 2233.62 ;
     RECT  1390.46 2231.9 1504.42 2235.76 ;
     RECT  1629.02 2232.4 1655.14 2235.98 ;
     RECT  1665.98 2220.64 1714.18 2235.98 ;
     RECT  860.22 2230.48 886.34 2236.14 ;
     RECT  861.18 2236.14 886.34 2236.98 ;
     RECT  830.94 2217.24 847.94 2237.82 ;
     RECT  954.78 2233.62 956.9 2238.24 ;
     RECT  631.58 2197.76 638.98 2238.92 ;
     RECT  668.06 2184.1 730.18 2239.12 ;
     RECT  1421.66 2235.76 1504.42 2239.12 ;
     RECT  867.42 2236.98 886.34 2239.72 ;
     RECT  897.66 2232.36 929.54 2239.72 ;
     RECT  622.46 2238.92 638.98 2239.76 ;
     RECT  1299.26 2150.08 1353.7 2239.96 ;
     RECT  816.06 2217.24 818.18 2241.18 ;
     RECT  834.78 2237.82 847.94 2241.18 ;
     RECT  1629.02 2235.98 1714.18 2241.22 ;
     RECT  1797.98 1793.5 1798.18 2242.195 ;
     RECT  3087.26 2204.04 3099.46 2242.195 ;
     RECT  2405.18 2231.78 2415.94 2243.32 ;
     RECT  956.7 2238.24 956.9 2243.5 ;
     RECT  969.66 2192.04 969.86 2243.5 ;
     RECT  1544.06 2232.4 1618.18 2243.74 ;
     RECT  2562.62 2213.72 2562.82 2246.26 ;
     RECT  1422.14 2239.12 1504.42 2246.68 ;
     RECT  956.7 2243.5 969.86 2247.06 ;
     RECT  622.46 2239.76 639.94 2247.32 ;
     RECT  846.78 2241.18 846.98 2247.48 ;
     RECT  1793.18 2242.195 1798.18 2247.765 ;
     RECT  3087.26 2242.195 3106.82 2247.765 ;
     RECT  1739.9 2217.5 1740.58 2249.2 ;
     RECT  1515.74 2232.4 1530.82 2249.62 ;
     RECT  1629.02 2241.22 1702.66 2250.04 ;
     RECT  2314.46 2027.02 2314.66 2250.04 ;
     RECT  2390.3 2204.48 2390.5 2250.46 ;
     RECT  2405.18 2243.32 2412.58 2251.72 ;
     RECT  786.62 2026.4 786.82 2251.9 ;
     RECT  867.42 2239.72 929.54 2252.1 ;
     RECT  1515.74 2249.62 1518.34 2252.14 ;
     RECT  3087.26 2247.765 3104.22 2252.14 ;
     RECT  1652.06 2250.04 1702.66 2253.2 ;
     RECT  1713.98 2241.22 1714.18 2253.2 ;
     RECT  3066.62 2217.72 3071.14 2253.4 ;
     RECT  2404.7 2251.72 2412.58 2253.7 ;
     RECT  2405.18 2253.7 2412.58 2253.82 ;
     RECT  892.38 2252.1 929.54 2254 ;
     RECT  2405.18 2253.82 2405.86 2254.24 ;
     RECT  622.46 2247.32 640.42 2258.24 ;
     RECT  650.3 2138.12 650.5 2258.24 ;
     RECT  956.7 2247.06 960.26 2258.62 ;
     RECT  867.42 2252.1 880.1 2258.82 ;
     RECT  1795.78 2247.765 1798.18 2259.165 ;
     RECT  3099.26 2252.14 3104.22 2259.165 ;
     RECT  867.42 2258.82 879.62 2259.24 ;
     RECT  1119.42 2205.9 1119.62 2260.3 ;
     RECT  1422.62 2246.68 1504.42 2260.54 ;
     RECT  1517.18 2252.14 1518.34 2262.22 ;
     RECT  3066.62 2253.4 3066.82 2262.22 ;
     RECT  2405.66 2254.24 2405.86 2262.64 ;
     RECT  3087.26 2252.14 3087.46 2263.06 ;
     RECT  1499.9 2260.54 1504.42 2263.28 ;
     RECT  1773.02 2229.12 1782.34 2264.32 ;
     RECT  3099.26 2259.165 3099.46 2264.74 ;
     RECT  1263.26 2261.6 1263.46 2264.96 ;
     RECT  892.38 2254 936.74 2265.96 ;
     RECT  892.38 2265.96 929.54 2266.38 ;
     RECT  1824.38 1911.74 1824.58 2266.64 ;
     RECT  1773.02 2264.32 1781.86 2267.9 ;
     RECT  892.38 2266.38 929.06 2269.12 ;
     RECT  1299.26 2239.96 1351.3 2271.88 ;
     RECT  724.7 2239.12 730.18 2272.9 ;
     RECT  1544.06 2243.74 1544.26 2274.62 ;
     RECT  1556.06 2243.74 1618.18 2274.62 ;
     RECT  1422.62 2260.54 1489.06 2275.66 ;
     RECT  1541.18 2274.62 1618.18 2276.5 ;
     RECT  801.66 2256.94 801.86 2277.3 ;
     RECT  1499.9 2263.28 1505.86 2278.6 ;
     RECT  1119.42 2260.3 1127.3 2279.62 ;
     RECT  979.26 2272.06 979.46 2279.82 ;
     RECT  1541.18 2276.5 1562.02 2280.28 ;
     RECT  1299.26 2271.88 1300.42 2283.235 ;
     RECT  1310.78 2271.88 1351.3 2283.235 ;
     RECT  1740.38 2249.2 1740.58 2284.28 ;
     RECT  1541.18 2280.28 1559.14 2284.9 ;
     RECT  1764.86 2267.9 1781.86 2286.16 ;
     RECT  953.34 2258.62 960.26 2286.76 ;
     RECT  1428.86 2275.66 1489.06 2287.42 ;
     RECT  834.78 2241.18 834.98 2288.64 ;
     RECT  886.62 2269.12 929.06 2289.06 ;
     RECT  896.22 2289.06 929.06 2292 ;
     RECT  1117.98 2279.62 1127.3 2292 ;
     RECT  953.34 2286.76 962.18 2293.06 ;
     RECT  1117.98 2292 1124.9 2293.68 ;
     RECT  1504.22 2278.6 1505.86 2295.4 ;
     RECT  1797.98 2259.165 1798.18 2296.46 ;
     RECT  622.46 2258.24 650.5 2299.18 ;
     RECT  1299.26 2283.235 1351.3 2300.205 ;
     RECT  896.22 2292 927.14 2300.4 ;
     RECT  867.42 2259.24 875.78 2300.82 ;
     RECT  1227.26 2300.66 1227.46 2301.08 ;
     RECT  766.14 2209.9 771.14 2301.24 ;
     RECT  724.7 2272.9 732.26 2302.08 ;
     RECT  781.98 2251.9 786.82 2302.08 ;
     RECT  943.26 2293.48 943.46 2302.3 ;
     RECT  953.34 2293.06 964.1 2302.3 ;
     RECT  1954.46 1798.34 1954.66 2303.6 ;
     RECT  1450.46 2287.42 1489.06 2304.86 ;
     RECT  867.42 2300.82 867.62 2308.38 ;
     RECT  899.1 2300.4 927.14 2308.38 ;
     RECT  903.9 2308.38 927.14 2309.22 ;
     RECT  904.38 2309.22 927.14 2315.52 ;
     RECT  943.26 2302.3 964.1 2316.36 ;
     RECT  1119.42 2293.68 1124.9 2316.78 ;
     RECT  766.14 2301.24 770.18 2322.66 ;
     RECT  624.38 2299.18 650.5 2323.76 ;
     RECT  668.06 2239.12 714.82 2323.76 ;
     RECT  1299.26 2300.205 1300.42 2323.76 ;
     RECT  1310.78 2300.205 1351.3 2323.76 ;
     RECT  951.9 2316.36 964.1 2324.34 ;
     RECT  910.14 2315.52 927.14 2326.02 ;
     RECT  910.62 2326.02 927.14 2326.44 ;
     RECT  956.7 2324.34 964.1 2326.86 ;
     RECT  956.7 2326.86 961.22 2327.28 ;
     RECT  724.7 2302.08 730.18 2330.06 ;
     RECT  597.5 2317.88 597.7 2330.26 ;
     RECT  624.38 2323.76 714.82 2331.32 ;
     RECT  724.7 2330.06 736.9 2331.32 ;
     RECT  624.38 2331.32 736.9 2332.16 ;
     RECT  956.7 2327.28 960.26 2335.68 ;
     RECT  624.38 2332.16 742.66 2338.24 ;
     RECT  769.02 2322.66 770.18 2338.62 ;
     RECT  3222 2215 3400 2339 ;
     RECT  910.62 2326.44 915.62 2345.76 ;
     RECT  769.98 2338.62 770.18 2346.18 ;
     RECT  0 2225 178 2349 ;
     RECT  915.42 2345.76 915.62 2353.12 ;
     RECT  926.94 2326.44 927.14 2353.12 ;
     RECT  915.42 2353.12 927.14 2357.1 ;
     RECT  915.42 2357.1 921.38 2360.46 ;
     RECT  1752.86 2178.22 1754.02 2361.34 ;
     RECT  638.78 2338.24 742.66 2361.76 ;
     RECT  1629.02 2250.04 1638.82 2365.12 ;
     RECT  816.06 2241.18 816.26 2365.92 ;
     RECT  1652.06 2253.2 1714.18 2372.26 ;
     RECT  915.42 2360.46 915.62 2374.32 ;
     RECT  1364.06 2150.08 1378.66 2375.62 ;
     RECT  1371.26 2375.62 1378.66 2378.14 ;
     RECT  680.54 2361.76 742.66 2378.52 ;
     RECT  1629.02 2365.12 1637.38 2379.82 ;
     RECT  786.62 2302.08 786.82 2381.08 ;
     RECT  1299.26 2323.76 1351.3 2381.5 ;
     RECT  1328.06 2381.5 1351.3 2383.6 ;
     RECT  638.78 2361.76 669.22 2386.44 ;
     RECT  1220.06 2301.08 1227.46 2394.1 ;
     RECT  624.38 2338.24 624.58 2394.94 ;
     RECT  1256.06 2264.96 1263.46 2394.94 ;
     RECT  638.78 2386.44 650.5 2395.36 ;
     RECT  1263.26 2394.94 1263.46 2395.36 ;
     RECT  712.7 2378.52 742.66 2402.08 ;
     RECT  1220.06 2394.1 1220.26 2402.5 ;
     RECT  724.7 2402.08 742.66 2402.92 ;
     RECT  742.46 2402.92 742.66 2403.34 ;
     RECT  1299.26 2381.5 1315.78 2405.44 ;
     RECT  1572.86 2276.5 1618.18 2408.38 ;
     RECT  3222 2339 3470 2409 ;
     RECT  1594.46 2408.38 1618.18 2409.22 ;
     RECT  638.78 2395.36 640.42 2412.16 ;
     RECT  1299.26 2405.44 1308.1 2412.16 ;
     RECT  1572.86 2408.38 1580.74 2415.94 ;
     RECT  1504.22 2295.4 1504.42 2416.36 ;
     RECT  -70 2349 178 2419 ;
     RECT  680.54 2378.52 701.54 2419.1 ;
     RECT  712.7 2402.08 714.82 2419.1 ;
     RECT  650.3 2395.36 650.5 2422.66 ;
     RECT  1328.06 2383.6 1349.86 2429.38 ;
     RECT  1119.42 2316.78 1119.62 2433.96 ;
     RECT  1371.26 2378.14 1371.94 2434 ;
     RECT  680.54 2419.1 714.82 2448.28 ;
     RECT  1371.26 2434 1371.46 2456.26 ;
     RECT  1336.22 2429.38 1349.86 2457.1 ;
     RECT  1299.26 2412.16 1300.42 2459.62 ;
     RECT  1349.66 2457.1 1349.86 2468.86 ;
     RECT  1390.46 2235.76 1410.34 2479.36 ;
     RECT  1390.46 2479.36 1400.26 2487.76 ;
     RECT  1336.22 2457.1 1336.42 2494.7 ;
     RECT  668.06 2386.44 669.22 2507.5 ;
     RECT  1284.38 1567.76 1284.58 2509.18 ;
     RECT  956.7 2335.68 956.9 2512.08 ;
     RECT  638.78 2412.16 638.98 2516.32 ;
     RECT  668.06 2507.5 668.74 2520.94 ;
     RECT  681.02 2448.28 714.82 2525.14 ;
     RECT  1089.5 1925.6 1089.7 2529.76 ;
     RECT  3222 2409 3400 2533 ;
     RECT  668.06 2520.94 668.26 2537.74 ;
     RECT  681.98 2525.14 714.82 2541.94 ;
     RECT  0 2419 178 2543 ;
     RECT  724.7 2402.92 730.18 2543.2 ;
     RECT  681.98 2541.94 712.9 2545.3 ;
     RECT  1300.22 2459.62 1300.42 2547.715 ;
     RECT  724.7 2543.2 724.9 2549.08 ;
     RECT  708.86 2545.3 712.9 2552.86 ;
     RECT  1300.22 2547.715 1306.82 2553.285 ;
     RECT  681.98 2545.3 694.82 2553.7 ;
     RECT  1796.06 2296.46 1798.18 2555.8 ;
     RECT  682.46 2553.7 694.82 2556.22 ;
     RECT  712.7 2552.86 712.9 2558.32 ;
     RECT  683.42 2556.22 694.82 2559.115 ;
     RECT  683.42 2559.115 697.42 2564.685 ;
     RECT  1300.22 2553.285 1304.22 2564.685 ;
     RECT  683.42 2564.685 690.82 2565.88 ;
     RECT  690.62 2565.88 690.82 2573.02 ;
     RECT  3222 2533 3470 2603 ;
     RECT  -70 2543 178 2613 ;
     RECT  1654.94 2372.26 1714.18 2653.24 ;
     RECT  1629.02 2379.82 1630.18 2725.06 ;
     RECT  3222 2603 3400 2727 ;
     RECT  0 2613 178 2737 ;
     RECT  3222 2727 3470 2797 ;
     RECT  -70 2737 178 2807 ;
     RECT  2049.02 2193.14 2049.22 2868.92 ;
     RECT  2091.26 1876.46 2091.94 2876.06 ;
     RECT  1428.86 2287.42 1436.74 2876.26 ;
     RECT  1393.82 2487.76 1400.26 2883.62 ;
     RECT  1925.66 2298.98 1925.86 2890.76 ;
     RECT  1428.86 2876.26 1436.26 2890.96 ;
     RECT  1541.18 2284.9 1556.26 2895.16 ;
     RECT  1410.14 2479.36 1410.34 2898.1 ;
     RECT  1674.62 2653.24 1714.18 2901.88 ;
     RECT  1764.86 2286.16 1776.1 2904.82 ;
     RECT  1551.26 2895.16 1556.26 2907.76 ;
     RECT  1572.86 2415.94 1580.26 2907.76 ;
     RECT  1617.98 2409.22 1618.18 2907.76 ;
     RECT  1729.34 1834.66 1729.54 2909.02 ;
     RECT  1428.86 2890.96 1429.06 2911.54 ;
     RECT  1450.46 2304.86 1490.98 2911.54 ;
     RECT  2016.38 1752.98 2016.58 2912.18 ;
     RECT  1517.18 2262.22 1517.38 2912.6 ;
     RECT  1529.66 2249.62 1530.82 2912.6 ;
     RECT  1629.98 2725.06 1630.18 2912.6 ;
     RECT  1541.18 2895.16 1541.38 2915.12 ;
     RECT  1551.26 2907.76 1552.42 2915.12 ;
     RECT  1594.46 2409.22 1603.78 2915.12 ;
     RECT  1818.62 2266.64 1824.58 2915.12 ;
     RECT  1841.18 2259.92 1841.38 2915.12 ;
     RECT  1875.26 2883.62 1875.46 2915.12 ;
     RECT  1897.82 2343.5 1898.02 2915.12 ;
     RECT  1490.78 2911.54 1490.98 2915.54 ;
     RECT  1625.66 2912.6 1630.18 2915.54 ;
     RECT  1654.94 2653.24 1659.46 2915.54 ;
     RECT  1740.38 2284.28 1741.54 2915.54 ;
     RECT  1752.86 2361.34 1753.06 2915.54 ;
     RECT  1768.22 2904.82 1776.1 2915.54 ;
     RECT  1796.06 2555.8 1796.26 2915.54 ;
     RECT  1818.62 2915.12 1825.06 2915.54 ;
     RECT  1841.18 2915.12 1846.66 2915.54 ;
     RECT  1869.02 2915.12 1875.46 2915.54 ;
     RECT  1977.5 2027.24 1977.7 2915.54 ;
     RECT  1674.62 2901.88 1710.82 2915.74 ;
     RECT  1336.22 2494.7 1345.06 2917 ;
     RECT  1517.18 2912.6 1530.82 2917 ;
     RECT  1594.46 2915.12 1609.06 2917 ;
     RECT  1739.9 2915.54 1753.06 2917 ;
     RECT  1490.78 2915.54 1495.3 2917.22 ;
     RECT  1947.74 2303.6 1954.66 2917.22 ;
     RECT  1300.22 2564.685 1300.42 2919.32 ;
     RECT  3222 2797 3400 2921 ;
     RECT  0 2807 178 2931 ;
     RECT  1299.74 2919.32 1300.42 2942.155 ;
     RECT  1322.3 2437.16 1322.5 2942.155 ;
     RECT  1344.86 2917 1345.06 2942.155 ;
     RECT  1371.26 2918.9 1371.46 2942.155 ;
     RECT  1389.98 2883.62 1400.26 2942.155 ;
     RECT  1427.42 2916.8 1427.62 2942.155 ;
     RECT  1450.46 2911.54 1451.62 2942.155 ;
     RECT  1468.7 2911.54 1479.94 2942.155 ;
     RECT  1490.78 2917.22 1501.06 2942.155 ;
     RECT  1519.1 2917 1530.82 2942.155 ;
     RECT  1541.18 2915.12 1552.42 2942.155 ;
     RECT  1573.82 2907.76 1580.26 2942.155 ;
     RECT  1595.9 2917 1609.06 2942.155 ;
     RECT  1625.66 2915.54 1632.1 2942.155 ;
     RECT  1652.54 2915.54 1659.46 2942.155 ;
     RECT  1685.18 2915.74 1710.82 2942.155 ;
     RECT  1720.7 2919.32 1720.9 2942.155 ;
     RECT  1739.9 2917 1747.3 2942.155 ;
     RECT  1764.38 2915.54 1776.1 2942.155 ;
     RECT  1786.46 2915.54 1796.26 2942.155 ;
     RECT  1814.78 2915.54 1825.06 2942.155 ;
     RECT  1837.34 2915.54 1854.34 2942.155 ;
     RECT  1869.02 2915.54 1876.9 2942.155 ;
     RECT  1897.82 2915.12 1902.82 2942.155 ;
     RECT  1920.38 2890.76 1925.86 2942.155 ;
     RECT  1947.74 2917.22 1955.62 2942.155 ;
     RECT  1965.98 2915.54 1966.18 2942.155 ;
     RECT  1977.02 2915.54 1977.7 2942.155 ;
     RECT  2016.38 2912.18 2021.38 2942.155 ;
     RECT  2049.02 2868.92 2055.46 2942.155 ;
     RECT  2077.34 2307.38 2077.54 2942.155 ;
     RECT  2091.26 2876.06 2101.54 2942.155 ;
     RECT  1299.74 2942.155 1663.085 2947.725 ;
     RECT  1317.665 2947.725 1663.085 2953.555 ;
     RECT  1674.62 2915.74 1674.82 2953.555 ;
     RECT  1685.18 2942.155 1720.9 2953.555 ;
     RECT  1736.755 2942.155 2101.54 2953.555 ;
     RECT  1299.74 2947.725 1305.1 2959.125 ;
     RECT  1317.665 2953.555 1720.9 2959.125 ;
     RECT  1731.135 2953.555 2101.54 2959.125 ;
     RECT  1685.18 2959.125 1710.82 2959.3 ;
     RECT  3222 2921 3470 2991 ;
     RECT  -70 2931 178 3001 ;
     RECT  1344.86 2959.125 1345.06 3009.5 ;
     RECT  1814.78 2959.125 1825.06 3009.5 ;
     RECT  1965.98 2959.125 1966.18 3009.5 ;
     RECT  1299.74 2959.125 1300.42 3010.555 ;
     RECT  1322.3 2959.125 1322.5 3010.555 ;
     RECT  1344.38 3009.5 1345.06 3010.555 ;
     RECT  1371.26 2959.125 1371.46 3010.555 ;
     RECT  1389.98 2959.125 1400.26 3010.555 ;
     RECT  1427.42 2959.125 1427.62 3010.555 ;
     RECT  1450.46 2959.125 1451.62 3010.555 ;
     RECT  1468.7 2959.125 1479.94 3010.555 ;
     RECT  1490.78 2959.125 1501.06 3010.555 ;
     RECT  1519.1 2959.125 1530.82 3010.555 ;
     RECT  1541.18 2959.125 1552.42 3010.555 ;
     RECT  1573.82 2959.125 1580.26 3010.555 ;
     RECT  1595.9 2959.125 1609.06 3010.555 ;
     RECT  1625.66 2959.125 1632.1 3010.555 ;
     RECT  1652.54 2959.125 1659.46 3010.555 ;
     RECT  1685.18 2959.3 1690.18 3010.555 ;
     RECT  1700.54 2959.3 1710.82 3010.555 ;
     RECT  1720.7 2959.125 1720.9 3010.555 ;
     RECT  1739.9 2959.125 1747.3 3010.555 ;
     RECT  1764.38 2959.125 1775.62 3010.555 ;
     RECT  1786.46 2959.125 1796.26 3010.555 ;
     RECT  1814.3 3009.5 1825.06 3010.555 ;
     RECT  1837.34 2959.125 1854.34 3010.555 ;
     RECT  1869.02 2959.125 1876.9 3010.555 ;
     RECT  1897.82 2959.125 1902.82 3010.555 ;
     RECT  1920.38 2959.125 1925.86 3010.555 ;
     RECT  1947.74 2959.125 1955.62 3010.555 ;
     RECT  1965.5 3009.5 1966.18 3010.555 ;
     RECT  1977.02 2959.125 1977.7 3010.555 ;
     RECT  2016.38 2959.125 2021.38 3010.555 ;
     RECT  2049.02 2959.125 2055.46 3010.555 ;
     RECT  2077.34 2959.125 2077.54 3010.555 ;
     RECT  2091.26 2959.125 2101.54 3010.555 ;
     RECT  1299.74 3010.555 1663.085 3016.125 ;
     RECT  1317.665 3016.125 1663.085 3021.955 ;
     RECT  1674.62 2959.125 1674.82 3021.955 ;
     RECT  1685.18 3010.555 1720.9 3021.955 ;
     RECT  1736.755 3010.555 2101.54 3021.955 ;
     RECT  1299.74 3016.125 1305.1 3027.525 ;
     RECT  1317.665 3021.955 1720.9 3027.525 ;
     RECT  1731.135 3021.955 2101.54 3027.525 ;
     RECT  2091.26 3027.525 2101.54 3031.68 ;
     RECT  2092.7 3031.68 2101.54 3032.5 ;
     RECT  1764.38 3027.525 1776.1 3033.96 ;
     RECT  1367.9 3027.525 1371.46 3036.24 ;
     RECT  1674.62 3027.525 1674.82 3038.3 ;
     RECT  1685.18 3027.525 1690.18 3038.3 ;
     RECT  1739.9 3027.525 1747.3 3038.3 ;
     RECT  2077.34 3027.525 2077.54 3038.3 ;
     RECT  1674.62 3038.3 1690.18 3038.5 ;
     RECT  1764.86 3033.96 1776.1 3038.5 ;
     RECT  1897.82 3027.525 1902.82 3038.5 ;
     RECT  2077.34 3038.3 2079.94 3038.5 ;
     RECT  1299.74 3027.525 1300.42 3045.16 ;
     RECT  1344.38 3027.525 1344.58 3045.16 ;
     RECT  1977.02 3027.525 1977.7 3047.44 ;
     RECT  2112.38 3036.04 2112.58 3048.46 ;
     RECT  1299.74 3045.16 1301.38 3049.52 ;
     RECT  1965.5 3027.525 1965.7 3049.52 ;
     RECT  1977.02 3047.44 1980.58 3049.52 ;
     RECT  2079.74 3038.5 2079.94 3049.52 ;
     RECT  1322.3 3027.525 1332.1 3049.72 ;
     RECT  1344.38 3045.16 1353.7 3049.72 ;
     RECT  2016.38 3027.525 2021.38 3049.72 ;
     RECT  1573.82 3027.525 1580.26 3050.36 ;
     RECT  2016.38 3049.72 2032.9 3050.56 ;
     RECT  2093.66 3032.5 2101.54 3050.56 ;
     RECT  1367.9 3036.24 1368.1 3051.2 ;
     RECT  2093.18 3050.78 2093.38 3051.2 ;
     RECT  1367.9 3051.2 1375.3 3051.4 ;
     RECT  2016.38 3050.56 2031.46 3051.4 ;
     RECT  1720.7 3027.525 1720.9 3051.62 ;
     RECT  1353.5 3049.72 1353.7 3052 ;
     RECT  1427.42 3027.525 1427.62 3052 ;
     RECT  2078.3 3049.52 2079.94 3052 ;
     RECT  1675.58 3038.5 1690.18 3052.04 ;
     RECT  1353.5 3052 1356.1 3052.2 ;
     RECT  2078.3 3052 2080.9 3052.2 ;
     RECT  2108.54 3052 2108.74 3052.24 ;
     RECT  1450.46 3027.525 1451.62 3052.46 ;
     RECT  1468.7 3027.525 1479.94 3052.46 ;
     RECT  1490.78 3027.525 1501.06 3052.46 ;
     RECT  1625.66 3027.525 1632.1 3052.46 ;
     RECT  1652.54 3027.525 1659.46 3052.46 ;
     RECT  1674.14 3052.04 1690.18 3052.46 ;
     RECT  1700.54 3027.525 1710.34 3052.46 ;
     RECT  2080.7 3052.2 2080.9 3052.46 ;
     RECT  2092.7 3051.2 2093.38 3052.46 ;
     RECT  2080.7 3052.46 2093.38 3052.66 ;
     RECT  1423.1 3052 1427.62 3052.88 ;
     RECT  1445.18 3052.46 1451.62 3052.88 ;
     RECT  1652.54 3052.46 1660.42 3052.88 ;
     RECT  1739.9 3038.3 1747.78 3052.88 ;
     RECT  1786.46 3027.525 1796.26 3052.88 ;
     RECT  1837.34 3027.525 1854.34 3052.88 ;
     RECT  1869.02 3027.525 1876.9 3052.88 ;
     RECT  1898.3 3038.5 1902.82 3052.88 ;
     RECT  1322.3 3049.72 1327.78 3053.08 ;
     RECT  1423.1 3052.88 1451.62 3053.08 ;
     RECT  1519.1 3027.525 1530.82 3053.08 ;
     RECT  1541.18 3027.525 1552.42 3053.08 ;
     RECT  1736.06 3052.88 1747.78 3053.08 ;
     RECT  1814.3 3027.525 1825.06 3053.08 ;
     RECT  1868.06 3052.88 1876.9 3053.08 ;
     RECT  1965.5 3049.52 1980.58 3053.08 ;
     RECT  1299.74 3049.52 1306.66 3053.3 ;
     RECT  1322.3 3053.08 1325.86 3053.3 ;
     RECT  1428.86 3053.08 1451.62 3053.3 ;
     RECT  1541.66 3053.08 1552.42 3053.3 ;
     RECT  1573.82 3050.36 1581.22 3053.3 ;
     RECT  1595.9 3027.525 1609.06 3053.3 ;
     RECT  1625.66 3052.46 1636.42 3053.3 ;
     RECT  1652.06 3052.88 1660.42 3053.3 ;
     RECT  1674.14 3052.46 1710.34 3053.3 ;
     RECT  1736.06 3053.08 1747.3 3053.3 ;
     RECT  1764.86 3038.5 1775.62 3053.3 ;
     RECT  1785.5 3052.88 1796.26 3053.3 ;
     RECT  1837.34 3052.88 1854.82 3053.3 ;
     RECT  1898.3 3052.88 1903.3 3053.3 ;
     RECT  1920.38 3027.525 1925.86 3053.3 ;
     RECT  1947.74 3027.525 1955.62 3053.3 ;
     RECT  1299.74 3053.3 1325.86 3053.5 ;
     RECT  1355.9 3052.2 1356.1 3053.5 ;
     RECT  1367.9 3051.4 1368.1 3053.5 ;
     RECT  1389.98 3027.525 1400.26 3053.5 ;
     RECT  1468.7 3052.46 1480.9 3053.5 ;
     RECT  1869.98 3053.08 1876.9 3053.5 ;
     RECT  1943.9 3053.3 1955.62 3053.5 ;
     RECT  1965.98 3053.08 1980.58 3053.5 ;
     RECT  2016.38 3051.4 2021.38 3053.5 ;
     RECT  2049.02 3027.525 2055.46 3053.5 ;
     RECT  1299.74 3053.5 1312.9 3058.84 ;
     RECT  1390.94 3053.5 1400.26 3059.04 ;
     RECT  1428.86 3053.3 1452.1 3060.1 ;
     RECT  1836.38 3053.3 1854.82 3060.1 ;
     RECT  1965.98 3053.5 1977.7 3060.1 ;
     RECT  1299.26 3058.84 1312.9 3060.22 ;
     RECT  1288.22 3036.04 1288.42 3063.58 ;
     RECT  1305.5 3060.22 1312.9 3065.88 ;
     RECT  1305.5 3065.88 1306.66 3066.1 ;
     RECT  1295.42 3065.68 1295.62 3066.94 ;
     RECT  1674.14 3053.3 1710.82 3067.1 ;
     RECT  1720.7 3051.62 1721.86 3067.1 ;
     RECT  2087.9 3052.66 2093.38 3067.96 ;
     RECT  2087.9 3067.96 2099.62 3073.66 ;
     RECT  1300.22 3072.52 1300.42 3074.08 ;
     RECT  1325.66 3053.5 1325.86 3076.675 ;
     RECT  1393.82 3059.04 1400.26 3076.675 ;
     RECT  1428.86 3060.1 1429.54 3076.675 ;
     RECT  1440.38 3060.1 1452.1 3076.675 ;
     RECT  1468.7 3053.5 1479.94 3076.675 ;
     RECT  1490.78 3052.46 1502.5 3076.675 ;
     RECT  1519.1 3053.08 1530.34 3076.675 ;
     RECT  1541.66 3053.3 1553.38 3076.675 ;
     RECT  1569.98 3053.3 1581.22 3076.675 ;
     RECT  1592.54 3053.3 1636.42 3076.675 ;
     RECT  1648.7 3053.3 1660.42 3076.675 ;
     RECT  1735.1 3053.3 1747.3 3076.675 ;
     RECT  1764.38 3053.3 1775.62 3076.675 ;
     RECT  1785.5 3053.3 1798.18 3076.675 ;
     RECT  1814.78 3053.08 1825.06 3076.675 ;
     RECT  1836.38 3060.1 1854.34 3076.675 ;
     RECT  1869.98 3053.5 1875.46 3076.675 ;
     RECT  1893.5 3053.3 1904.26 3076.675 ;
     RECT  1916.06 3053.3 1927.3 3076.675 ;
     RECT  1943.9 3053.5 1955.14 3076.675 ;
     RECT  1966.46 3060.1 1977.7 3076.675 ;
     RECT  2016.38 3053.5 2016.58 3076.675 ;
     RECT  2050.46 3053.5 2050.66 3076.675 ;
     RECT  2087.9 3073.66 2098.98 3076.675 ;
     RECT  1300.86 3076.675 1663.085 3082.245 ;
     RECT  1735.1 3076.675 2098.98 3082.245 ;
     RECT  1317.665 3082.245 1663.085 3088.075 ;
     RECT  1674.14 3067.1 1721.86 3088.075 ;
     RECT  1735.1 3082.245 2082.175 3088.075 ;
     RECT  1303.46 3082.245 1305.1 3093.645 ;
     RECT  1317.665 3088.075 2082.175 3093.645 ;
     RECT  2094.74 3082.245 2096.38 3093.645 ;
     RECT  1490.78 3093.645 1502.5 3110.3 ;
     RECT  1592.54 3093.645 1636.42 3110.5 ;
     RECT  1541.66 3093.645 1550.98 3111.28 ;
     RECT  3222 2991 3400 3115 ;
     RECT  1592.54 3110.5 1635.94 3116.04 ;
     RECT  1592.54 3116.04 1610.5 3117.7 ;
     RECT  0 3001 178 3125 ;
     RECT  1620.38 3116.04 1635.94 3132.1 ;
     RECT  1393.82 3093.645 1400.26 3145.075 ;
     RECT  1428.86 3093.645 1429.54 3145.075 ;
     RECT  1440.38 3093.645 1452.1 3145.075 ;
     RECT  1468.7 3093.645 1479.94 3145.075 ;
     RECT  1490.3 3110.3 1502.5 3145.075 ;
     RECT  1519.1 3093.645 1530.34 3145.075 ;
     RECT  1541.66 3111.28 1554.34 3145.075 ;
     RECT  1569.98 3093.645 1581.22 3145.075 ;
     RECT  1592.54 3117.7 1609.54 3145.075 ;
     RECT  1620.38 3132.1 1634.5 3145.075 ;
     RECT  1648.22 3093.645 1659.94 3145.075 ;
     RECT  1735.1 3093.645 1747.3 3145.075 ;
     RECT  1764.38 3093.645 1775.62 3145.075 ;
     RECT  1785.5 3093.645 1798.18 3145.075 ;
     RECT  1814.78 3093.645 1825.06 3145.075 ;
     RECT  1836.38 3093.645 1854.34 3145.075 ;
     RECT  1869.98 3093.645 1875.46 3145.075 ;
     RECT  1893.5 3093.645 1903.3 3145.075 ;
     RECT  1916.06 3093.645 1927.3 3145.075 ;
     RECT  1943.9 3093.645 1955.14 3145.075 ;
     RECT  1966.46 3093.645 1977.7 3145.075 ;
     RECT  2016.38 3093.645 2016.58 3145.075 ;
     RECT  1300.86 3145.075 1663.085 3150.645 ;
     RECT  1735.1 3145.075 2098.98 3150.645 ;
     RECT  1317.665 3150.645 1663.085 3156.475 ;
     RECT  1674.14 3093.645 1721.86 3156.475 ;
     RECT  1735.1 3150.645 2082.175 3156.475 ;
     RECT  1303.46 3150.645 1305.1 3162.045 ;
     RECT  1317.665 3156.475 2082.175 3162.045 ;
     RECT  2094.74 3150.645 2096.38 3162.045 ;
     RECT  1620.38 3162.045 1635.46 3168.1 ;
     RECT  1468.7 3162.045 1479.94 3183.7 ;
     RECT  1490.3 3162.045 1502.5 3183.7 ;
     RECT  1519.1 3162.045 1530.34 3183.7 ;
     RECT  1620.38 3168.1 1632.1 3183.7 ;
     RECT  1648.22 3162.045 1659.94 3183.7 ;
     RECT  1674.14 3162.045 1721.86 3183.7 ;
     RECT  1785.5 3162.045 1798.18 3183.7 ;
     RECT  1869.98 3162.045 1875.46 3183.7 ;
     RECT  1943.9 3162.045 1955.14 3183.7 ;
     RECT  1652.54 3183.7 1659.94 3184.12 ;
     RECT  1869.98 3183.7 1874.98 3184.12 ;
     RECT  3222 3115 3470 3185 ;
     RECT  1428.86 3162.045 1429.54 3187.06 ;
     RECT  1569.98 3162.045 1581.22 3187.06 ;
     RECT  1836.38 3162.045 1854.34 3187.06 ;
     RECT  1429.34 3187.06 1429.54 3187.48 ;
     RECT  1440.38 3162.045 1452.1 3187.48 ;
     RECT  1468.7 3183.7 1478.98 3187.48 ;
     RECT  1490.3 3183.7 1501.54 3187.48 ;
     RECT  1523.9 3183.7 1529.86 3187.48 ;
     RECT  1541.66 3162.045 1552.42 3187.48 ;
     RECT  1569.98 3187.06 1580.26 3187.48 ;
     RECT  1592.54 3162.045 1609.54 3187.48 ;
     RECT  1620.38 3183.7 1631.14 3187.48 ;
     RECT  1653.5 3184.12 1659.94 3187.48 ;
     RECT  1674.14 3183.7 1690.18 3187.48 ;
     RECT  1700.06 3183.7 1720.9 3187.48 ;
     RECT  1735.1 3162.045 1747.3 3187.48 ;
     RECT  1764.38 3162.045 1775.62 3187.48 ;
     RECT  1785.5 3183.7 1797.22 3187.48 ;
     RECT  1814.78 3162.045 1825.06 3187.48 ;
     RECT  1836.38 3187.06 1836.58 3187.48 ;
     RECT  1847.42 3187.06 1854.34 3187.48 ;
     RECT  1870.94 3184.12 1874.98 3187.48 ;
     RECT  1893.5 3162.045 1903.3 3187.48 ;
     RECT  1916.06 3162.045 1927.3 3187.48 ;
     RECT  1943.9 3183.7 1954.66 3187.48 ;
     RECT  1966.46 3162.045 1977.7 3187.48 ;
     RECT  1495.1 3187.48 1500.58 3187.9 ;
     RECT  1546.94 3187.48 1547.14 3187.9 ;
     RECT  1495.1 3187.9 1495.3 3188.32 ;
     RECT  1472.54 3187.48 1472.74 3189.16 ;
     RECT  1674.14 3187.48 1675.78 3190 ;
     RECT  1689.98 3187.48 1690.18 3191.26 ;
     RECT  1653.5 3187.48 1653.7 3191.68 ;
     RECT  1746.14 3187.48 1746.82 3191.68 ;
     RECT  1674.14 3190 1674.34 3192.1 ;
     RECT  1700.54 3187.48 1709.86 3192.1 ;
     RECT  1971.74 3187.48 1977.7 3192.1 ;
     RECT  1700.54 3192.1 1705.54 3192.52 ;
     RECT  -70 3125 178 3195 ;
     RECT  1705.34 3192.52 1705.54 3195.04 ;
     RECT  1746.62 3191.68 1746.82 3195.04 ;
     RECT  1579.1 3187.48 1580.26 3197.14 ;
     RECT  1773.5 3187.48 1775.62 3197.14 ;
     RECT  1954.46 3187.48 1954.66 3197.14 ;
     RECT  1450.46 3187.48 1450.66 3203.44 ;
     RECT  1393.82 3162.045 1400.26 3203.86 ;
     RECT  1775.42 3197.14 1775.62 3211.1 ;
     RECT  1775.42 3211.1 1776.1 3211.3 ;
     RECT  0 3195 178 3220 ;
     RECT  3222 3185 3400 3220 ;
     RECT  0 3220 180 3222 ;
     RECT  1393.82 3203.86 1394.02 3222 ;
     RECT  1579.1 3197.14 1579.3 3222 ;
     RECT  1629.98 3187.48 1630.18 3222 ;
     RECT  1775.9 3211.3 1776.1 3222 ;
     RECT  1824.38 3187.48 1824.58 3222 ;
     RECT  1977.5 3192.1 1977.7 3222 ;
     RECT  2016.38 3162.045 2016.58 3222 ;
     RECT  2365.34 2135.18 2365.54 3222 ;
     RECT  3220 3220 3400 3222 ;
     RECT  0 3222 3400 3400 ;
     RECT  215 3400 285 3470 ;
     RECT  409 3400 479 3470 ;
     RECT  603 3400 673 3470 ;
     RECT  797 3400 867 3470 ;
     RECT  991 3400 1061 3470 ;
     RECT  1185 3400 1255 3470 ;
     RECT  1379 3400 1449 3470 ;
     RECT  1573 3400 1643 3470 ;
     RECT  1767 3400 1837 3470 ;
     RECT  1961 3400 2031 3470 ;
     RECT  2155 3400 2225 3470 ;
     RECT  2349 3400 2419 3470 ;
     RECT  2543 3400 2613 3470 ;
     RECT  2737 3400 2807 3470 ;
     RECT  2931 3400 3001 3470 ;
     RECT  3125 3400 3195 3470 ;
    LAYER TopMetal1 ;
     RECT  -70 215 0 285 ;
     RECT  -70 409 0 479 ;
     RECT  -70 603 0 673 ;
     RECT  -70 797 0 867 ;
     RECT  -70 991 0 1061 ;
     RECT  -70 1185 0 1255 ;
     RECT  -70 1379 0 1449 ;
     RECT  -70 1573 0 1643 ;
     RECT  -70 1767 0 1837 ;
     RECT  -70 1961 0 2031 ;
     RECT  -70 2155 0 2225 ;
     RECT  -70 2349 0 2419 ;
     RECT  -70 2543 0 2613 ;
     RECT  -70 2737 0 2807 ;
     RECT  -70 2931 0 3001 ;
     RECT  -70 3125 0 3195 ;
     RECT  0 0 178 3400 ;
     RECT  178 0 205 212 ;
     RECT  178 3188 215 3400 ;
     RECT  205 -70 275 212 ;
     RECT  215 3188 285 3470 ;
     RECT  275 0 399 212 ;
     RECT  285 3188 409 3400 ;
     RECT  399 -70 469 212 ;
     RECT  409 3188 479 3470 ;
     RECT  469 0 593 212 ;
     RECT  479 3188 603 3400 ;
     RECT  593 -70 663 212 ;
     RECT  603 3188 673 3470 ;
     RECT  693 2016.26 695.6 2022.26 ;
     RECT  693 2283.02 695.6 2289.02 ;
     RECT  693 2547.5 695.6 2553.5 ;
     RECT  699.5 2200.84 716.98 2202.48 ;
     RECT  699.5 2089.12 717.94 2090.76 ;
     RECT  657.74 2385.52 737.9 2387.16 ;
     RECT  663 0 787 212 ;
     RECT  673 3188 797 3400 ;
     RECT  787 -70 857 212 ;
     RECT  797 3188 867 3470 ;
     RECT  857 0 981 212 ;
     RECT  867 3188 991 3400 ;
     RECT  993 616.34 995.6 622.34 ;
     RECT  993 782.78 995.6 788.78 ;
     RECT  993 946.94 995.6 952.94 ;
     RECT  995.6 782.78 999.98 800.18 ;
     RECT  999.98 782.78 1023.7 827.64 ;
     RECT  981 -70 1051 212 ;
     RECT  991 3188 1061 3470 ;
     RECT  1051 0 1175 212 ;
     RECT  1061 3188 1185 3400 ;
     RECT  1175 -70 1245 212 ;
     RECT  1185 3188 1255 3470 ;
     RECT  1287.5 3035.32 1294.7 3036.96 ;
     RECT  1294.7 3035.32 1299.5 3066.6 ;
     RECT  1299.5 3035.32 1300.68 3073.44 ;
     RECT  1255 3188 1300.68 3400 ;
     RECT  1300.68 2941.94 1303.28 2947.94 ;
     RECT  1300.68 3010.34 1303.28 3082.46 ;
     RECT  695.6 2016.26 1304.4 2033.66 ;
     RECT  695.6 2283.02 1304.4 2300.42 ;
     RECT  695.6 2547.5 1304.4 2564.9 ;
     RECT  1304.4 2016.26 1307 2022.26 ;
     RECT  1304.4 2283.02 1307 2289.02 ;
     RECT  1304.4 2547.5 1307 2553.5 ;
     RECT  737.9 2378.68 1315.06 2387.16 ;
     RECT  1315.06 2378.68 1339.06 2380.32 ;
     RECT  1245 0 1369 212 ;
     RECT  1300.68 3144.86 1379 3400 ;
     RECT  995.6 616.34 1404.4 633.74 ;
     RECT  1023.7 782.78 1404.4 800.18 ;
     RECT  995.6 946.94 1404.4 964.34 ;
     RECT  1404.4 616.34 1407 622.34 ;
     RECT  1404.4 782.78 1407 788.78 ;
     RECT  1404.4 946.94 1407 952.94 ;
     RECT  1303.28 3010.34 1424.02 3093.86 ;
     RECT  1369 -70 1439 212 ;
     RECT  1379 3144.86 1449 3470 ;
     RECT  1439 0 1563 212 ;
     RECT  1449 3144.86 1573 3400 ;
     RECT  1580.78 1991.08 1588.46 1992.72 ;
     RECT  1424.02 3076.46 1607.66 3093.86 ;
     RECT  1573 3144.86 1607.66 3470 ;
     RECT  1607.66 3076.46 1614.1 3470 ;
     RECT  1563 -70 1633 212 ;
     RECT  1614.1 3144.86 1643 3470 ;
     RECT  1614.1 3076.46 1706.54 3093.86 ;
     RECT  1643 3144.86 1706.54 3400 ;
     RECT  1424.02 3010.34 1708.46 3027.74 ;
     RECT  1706.54 3076.46 1708.46 3400 ;
     RECT  1708.46 3010.34 1710.58 3400 ;
     RECT  1710.58 3010.34 1720.66 3093.86 ;
     RECT  1633 0 1757 212 ;
     RECT  1504.94 2196.28 1765.1 2197.92 ;
     RECT  1710.58 3144.86 1767 3400 ;
     RECT  1683.98 1446.16 1788.14 1447.8 ;
     RECT  1765.1 2196.28 1791 2229.84 ;
     RECT  1791 1017.62 1795.6 1023.62 ;
     RECT  1791 1628.66 1795.6 1634.66 ;
     RECT  1791 2196.28 1795.6 2247.98 ;
     RECT  1757 -70 1827 212 ;
     RECT  1767 3144.86 1837 3470 ;
     RECT  1827 0 1951 212 ;
     RECT  1837 3144.86 1961 3400 ;
     RECT  1720.66 3010.34 1979.66 3027.74 ;
     RECT  1720.66 3076.46 1979.66 3093.86 ;
     RECT  1951 -70 2021 212 ;
     RECT  1961 3144.86 2031 3470 ;
     RECT  1303.28 2941.94 2096.56 2959.34 ;
     RECT  1979.66 3010.34 2096.56 3093.86 ;
     RECT  2096.56 2941.94 2099.16 2947.94 ;
     RECT  2096.56 3010.34 2099.16 3082.46 ;
     RECT  2031 3144.86 2099.16 3400 ;
     RECT  2099.16 3035.32 2100.34 3068.88 ;
     RECT  2100.34 3035.32 2109.46 3052.92 ;
     RECT  2109.46 3035.32 2113.3 3036.96 ;
     RECT  2021 0 2145 212 ;
     RECT  2099.16 3188 2155 3400 ;
     RECT  2145 -70 2215 212 ;
     RECT  2155 3188 2225 3470 ;
     RECT  2215 0 2339 212 ;
     RECT  2225 3188 2349 3400 ;
     RECT  2339 -70 2409 212 ;
     RECT  1588.46 1991.08 2411.18 2001.84 ;
     RECT  2349 3188 2419 3470 ;
     RECT  1795.6 2196.28 2437.78 2259.38 ;
     RECT  2437.78 2216.8 2508.14 2259.38 ;
     RECT  2409 0 2533 212 ;
     RECT  2508.14 2209.96 2537.9 2259.38 ;
     RECT  2419 3188 2543 3400 ;
     RECT  2546.06 2125.6 2564.3 2127.24 ;
     RECT  2564.3 2118.76 2573.9 2127.24 ;
     RECT  2537.9 2203.12 2573.9 2259.38 ;
     RECT  2573.9 2118.76 2574.58 2259.38 ;
     RECT  2533 -70 2603 212 ;
     RECT  2543 3188 2613 3470 ;
     RECT  1788.14 1446.16 2630.54 1466.04 ;
     RECT  2411.18 1959.16 2643.22 2001.84 ;
     RECT  2574.58 2125.6 2650.42 2259.38 ;
     RECT  2630.54 1409.68 2708.02 1466.04 ;
     RECT  2603 0 2727 212 ;
     RECT  2708.02 1409.68 2736.34 1459.2 ;
     RECT  2613 3188 2737 3400 ;
     RECT  2650.42 2159.8 2741.9 2259.38 ;
     RECT  2736.34 1409.68 2782.7 1454.64 ;
     RECT  2727 -70 2797 212 ;
     RECT  2737 3188 2807 3470 ;
     RECT  2741.9 2152.96 2866.42 2259.38 ;
     RECT  2797 0 2921 212 ;
     RECT  2807 3188 2931 3400 ;
     RECT  2866.42 2159.8 2941.78 2259.38 ;
     RECT  2921 -70 2991 212 ;
     RECT  2931 3188 3001 3470 ;
     RECT  2782.7 1409.68 3074.26 1466.04 ;
     RECT  2941.78 2166.64 3078.58 2259.38 ;
     RECT  3078.58 2175.76 3094.9 2259.38 ;
     RECT  3074.26 1453 3095.86 1466.04 ;
     RECT  2643.22 1991.08 3100.66 2001.84 ;
     RECT  3095.86 1453 3101.14 1459.2 ;
     RECT  1795.6 1017.62 3104.4 1035.02 ;
     RECT  1795.6 1628.66 3104.4 1646.06 ;
     RECT  3094.9 2241.98 3104.4 2259.38 ;
     RECT  3104.4 1017.62 3107 1023.62 ;
     RECT  3104.4 1628.66 3107 1634.66 ;
     RECT  3104.4 2241.98 3107 2247.98 ;
     RECT  2991 0 3115 212 ;
     RECT  3001 3188 3125 3400 ;
     RECT  3115 -70 3185 212 ;
     RECT  3125 3188 3195 3470 ;
     RECT  3185 0 3222 212 ;
     RECT  3101.14 1453 3222 1454.64 ;
     RECT  3094.9 2175.76 3222 2177.4 ;
     RECT  3195 3188 3222 3400 ;
     RECT  3222 0 3400 3400 ;
     RECT  3400 205 3470 275 ;
     RECT  3400 399 3470 469 ;
     RECT  3400 593 3470 663 ;
     RECT  3400 787 3470 857 ;
     RECT  3400 981 3470 1051 ;
     RECT  3400 1175 3470 1245 ;
     RECT  3400 1369 3470 1439 ;
     RECT  3400 1563 3470 1633 ;
     RECT  3400 1757 3470 1827 ;
     RECT  3400 1951 3470 2021 ;
     RECT  3400 2145 3470 2215 ;
     RECT  3400 2339 3470 2409 ;
     RECT  3400 2533 3470 2603 ;
     RECT  3400 2727 3470 2797 ;
     RECT  3400 2921 3470 2991 ;
     RECT  3400 3115 3470 3185 ;
    LAYER TopMetal2 ;
     RECT  205 -70 275 0 ;
     RECT  399 -70 469 0 ;
     RECT  593 -70 663 0 ;
     RECT  787 -70 857 0 ;
     RECT  981 -70 1051 0 ;
     RECT  1175 -70 1245 0 ;
     RECT  1369 -70 1439 0 ;
     RECT  1563 -70 1633 0 ;
     RECT  1757 -70 1827 0 ;
     RECT  1951 -70 2021 0 ;
     RECT  2145 -70 2215 0 ;
     RECT  2339 -70 2409 0 ;
     RECT  2533 -70 2603 0 ;
     RECT  2727 -70 2797 0 ;
     RECT  2921 -70 2991 0 ;
     RECT  3115 -70 3185 0 ;
     RECT  0 0 280 8.5 ;
     RECT  394 0 474 8.5 ;
     RECT  588 0 668 8.5 ;
     RECT  782 0 862 8.5 ;
     RECT  976 0 1056 8.5 ;
     RECT  1170 0 1250 8.5 ;
     RECT  1364 0 1444 8.5 ;
     RECT  1558 0 1638 8.5 ;
     RECT  1752 0 1832 8.5 ;
     RECT  1946 0 2026 8.5 ;
     RECT  2140 0 2220 8.5 ;
     RECT  2334 0 2414 8.5 ;
     RECT  2528 0 2608 8.5 ;
     RECT  2722 0 2802 8.5 ;
     RECT  2916 0 2996 8.5 ;
     RECT  3110 0 3400 8.5 ;
     RECT  0 8.5 3400 205 ;
     RECT  0 205 3470 212 ;
     RECT  0 212 212 215 ;
     RECT  3188 212 3470 275 ;
     RECT  3188 275 3400 280 ;
     RECT  -70 215 212 285 ;
     RECT  0 285 212 290 ;
     RECT  3188 280 3391.5 394 ;
     RECT  3188 394 3400 399 ;
     RECT  8.5 290 212 404 ;
     RECT  0 404 212 409 ;
     RECT  3188 399 3470 469 ;
     RECT  3188 469 3400 474 ;
     RECT  -70 409 212 479 ;
     RECT  0 479 212 484 ;
     RECT  3188 474 3391.5 588 ;
     RECT  3188 588 3400 593 ;
     RECT  8.5 484 212 598 ;
     RECT  0 598 212 603 ;
     RECT  1111 212 1117 616.34 ;
     RECT  1383 616.34 1389 627.74 ;
     RECT  3188 593 3470 663 ;
     RECT  3188 663 3400 668 ;
     RECT  -70 603 212 673 ;
     RECT  0 673 212 678 ;
     RECT  3188 668 3391.5 782 ;
     RECT  3188 782 3400 787 ;
     RECT  8.5 678 212 792 ;
     RECT  0 792 212 797 ;
     RECT  3188 787 3470 857 ;
     RECT  3188 857 3400 862 ;
     RECT  -70 797 212 867 ;
     RECT  0 867 212 872 ;
     RECT  3188 862 3391.5 976 ;
     RECT  3188 976 3400 981 ;
     RECT  8.5 872 212 986 ;
     RECT  0 986 212 991 ;
     RECT  1927 212 1933 1017.62 ;
     RECT  2539 212 2545 1017.62 ;
     RECT  2743 212 2749 1017.62 ;
     RECT  3015 1017.62 3021 1029.02 ;
     RECT  3188 981 3470 1051 ;
     RECT  3188 1051 3400 1056 ;
     RECT  -70 991 212 1061 ;
     RECT  0 1061 212 1066 ;
     RECT  3188 1056 3391.5 1170 ;
     RECT  3188 1170 3400 1175 ;
     RECT  8.5 1066 212 1180 ;
     RECT  0 1180 212 1185 ;
     RECT  3188 1175 3470 1245 ;
     RECT  3188 1245 3400 1250 ;
     RECT  -70 1185 212 1255 ;
     RECT  0 1255 212 1260 ;
     RECT  3188 1250 3391.5 1364 ;
     RECT  3188 1364 3400 1369 ;
     RECT  8.5 1260 212 1374 ;
     RECT  0 1374 212 1379 ;
     RECT  3188 1369 3470 1439 ;
     RECT  3188 1439 3400 1444 ;
     RECT  -70 1379 212 1449 ;
     RECT  0 1449 212 1454 ;
     RECT  3188 1444 3391.5 1558 ;
     RECT  3188 1558 3400 1563 ;
     RECT  8.5 1454 212 1568 ;
     RECT  0 1568 212 1573 ;
     RECT  3188 1563 3470 1633 ;
     RECT  3188 1633 3400 1638 ;
     RECT  -70 1573 212 1643 ;
     RECT  0 1643 212 1648 ;
     RECT  3188 1638 3391.5 1752 ;
     RECT  3188 1752 3400 1757 ;
     RECT  8.5 1648 212 1762 ;
     RECT  0 1762 212 1767 ;
     RECT  3188 1757 3470 1827 ;
     RECT  3188 1827 3400 1832 ;
     RECT  -70 1767 212 1837 ;
     RECT  0 1837 212 1842 ;
     RECT  3188 1832 3391.5 1946 ;
     RECT  3188 1946 3400 1951 ;
     RECT  8.5 1842 212 1956 ;
     RECT  0 1956 212 1961 ;
     RECT  3188 1951 3470 2021 ;
     RECT  3188 2021 3400 2026 ;
     RECT  771 212 777 2027.66 ;
     RECT  -70 1961 212 2031 ;
     RECT  0 2031 212 2036 ;
     RECT  3188 2026 3391.5 2140 ;
     RECT  3188 2140 3400 2145 ;
     RECT  8.5 2036 212 2150 ;
     RECT  0 2150 212 2155 ;
     RECT  3188 2145 3470 2215 ;
     RECT  3188 2215 3400 2220 ;
     RECT  -70 2155 212 2225 ;
     RECT  0 2225 212 2230 ;
     RECT  2131 212 2205 2247.98 ;
     RECT  2743 1017.62 2817 2247.98 ;
     RECT  2947 1029.02 3021 2247.98 ;
     RECT  3188 2220 3391.5 2334 ;
     RECT  3188 2334 3400 2339 ;
     RECT  8.5 2230 212 2344 ;
     RECT  0 2344 212 2349 ;
     RECT  3188 2339 3470 2409 ;
     RECT  3188 2409 3400 2414 ;
     RECT  -70 2349 212 2419 ;
     RECT  0 2419 212 2424 ;
     RECT  3188 2414 3391.5 2528 ;
     RECT  3188 2528 3400 2533 ;
     RECT  8.5 2424 212 2538 ;
     RECT  0 2538 212 2543 ;
     RECT  703 2027.66 777 2564.9 ;
     RECT  907 212 981 2564.9 ;
     RECT  3188 2533 3470 2603 ;
     RECT  3188 2603 3400 2608 ;
     RECT  -70 2543 212 2613 ;
     RECT  0 2613 212 2618 ;
     RECT  3188 2608 3391.5 2722 ;
     RECT  3188 2722 3400 2727 ;
     RECT  8.5 2618 212 2732 ;
     RECT  0 2732 212 2737 ;
     RECT  3188 2727 3470 2797 ;
     RECT  3188 2797 3400 2802 ;
     RECT  -70 2737 212 2807 ;
     RECT  0 2807 212 2812 ;
     RECT  3188 2802 3391.5 2916 ;
     RECT  3188 2916 3400 2921 ;
     RECT  8.5 2812 212 2926 ;
     RECT  0 2926 212 2931 ;
     RECT  1587 2941.94 1593 2953.34 ;
     RECT  1791 1017.62 1797 2953.34 ;
     RECT  3188 2921 3470 2991 ;
     RECT  3188 2991 3400 2996 ;
     RECT  -70 2931 212 3001 ;
     RECT  0 3001 212 3006 ;
     RECT  3188 2996 3391.5 3110 ;
     RECT  3188 3110 3400 3115 ;
     RECT  8.5 3006 212 3120 ;
     RECT  0 3120 212 3125 ;
     RECT  3188 3115 3470 3185 ;
     RECT  -70 3125 212 3188 ;
     RECT  771 2564.9 777 3188 ;
     RECT  975 2564.9 981 3188 ;
     RECT  1111 616.34 1185 3188 ;
     RECT  1315 627.74 1389 3188 ;
     RECT  1519 2953.34 1593 3188 ;
     RECT  1723 2953.34 1797 3188 ;
     RECT  1927 1017.62 2001 3188 ;
     RECT  2131 2247.98 2137 3188 ;
     RECT  2335 212 2409 3188 ;
     RECT  2539 1017.62 2613 3188 ;
     RECT  2743 2247.98 2749 3188 ;
     RECT  2947 2247.98 2953 3188 ;
     RECT  3188 3185 3400 3188 ;
     RECT  -70 3188 3400 3195 ;
     RECT  0 3195 3400 3391.5 ;
     RECT  0 3391.5 290 3400 ;
     RECT  404 3391.5 484 3400 ;
     RECT  598 3391.5 678 3400 ;
     RECT  792 3391.5 872 3400 ;
     RECT  986 3391.5 1066 3400 ;
     RECT  1180 3391.5 1260 3400 ;
     RECT  1374 3391.5 1454 3400 ;
     RECT  1568 3391.5 1648 3400 ;
     RECT  1762 3391.5 1842 3400 ;
     RECT  1956 3391.5 2036 3400 ;
     RECT  2150 3391.5 2230 3400 ;
     RECT  2344 3391.5 2424 3400 ;
     RECT  2538 3391.5 2618 3400 ;
     RECT  2732 3391.5 2812 3400 ;
     RECT  2926 3391.5 3006 3400 ;
     RECT  3120 3391.5 3400 3400 ;
     RECT  215 3400 285 3470 ;
     RECT  409 3400 479 3470 ;
     RECT  603 3400 673 3470 ;
     RECT  797 3400 867 3470 ;
     RECT  991 3400 1061 3470 ;
     RECT  1185 3400 1255 3470 ;
     RECT  1379 3400 1449 3470 ;
     RECT  1573 3400 1643 3470 ;
     RECT  1767 3400 1837 3470 ;
     RECT  1961 3400 2031 3470 ;
     RECT  2155 3400 2225 3470 ;
     RECT  2349 3400 2419 3470 ;
     RECT  2543 3400 2613 3470 ;
     RECT  2737 3400 2807 3470 ;
     RECT  2931 3400 3001 3470 ;
     RECT  3125 3400 3195 3470 ;
  END
END croc_chip
END LIBRARY
