VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO dmi_jtag
  FOREIGN dmi_jtag 0 0 ;
  CLASS BLOCK ;
  SIZE 600 BY 574.56 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VDDIO
    USE POWER ;
    DIRECTION INOUT ;
  END VDDIO
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN VSSIO
    USE GROUND ;
    DIRECTION INOUT ;
  END VSSIO
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 353.12 0.72 353.32 ;
    END
  END clk_i
  PIN dmi_req_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 242.24 600 242.44 ;
    END
  END dmi_req_o_0_
  PIN dmi_req_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 300.2 600 300.4 ;
    END
  END dmi_req_o_10_
  PIN dmi_req_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 297.68 600 297.88 ;
    END
  END dmi_req_o_11_
  PIN dmi_req_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 312.8 600 313 ;
    END
  END dmi_req_o_12_
  PIN dmi_req_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 355.64 600 355.84 ;
    END
  END dmi_req_o_13_
  PIN dmi_req_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 302.72 600 302.92 ;
    END
  END dmi_req_o_14_
  PIN dmi_req_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 290.12 600 290.32 ;
    END
  END dmi_req_o_15_
  PIN dmi_req_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 295.16 600 295.36 ;
    END
  END dmi_req_o_16_
  PIN dmi_req_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 345.56 600 345.76 ;
    END
  END dmi_req_o_17_
  PIN dmi_req_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 332.96 600 333.16 ;
    END
  END dmi_req_o_18_
  PIN dmi_req_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 282.56 600 282.76 ;
    END
  END dmi_req_o_19_
  PIN dmi_req_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 280.04 600 280.24 ;
    END
  END dmi_req_o_1_
  PIN dmi_req_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 277.52 600 277.72 ;
    END
  END dmi_req_o_20_
  PIN dmi_req_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 307.76 600 307.96 ;
    END
  END dmi_req_o_21_
  PIN dmi_req_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 335.48 600 335.68 ;
    END
  END dmi_req_o_22_
  PIN dmi_req_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 272.48 600 272.68 ;
    END
  END dmi_req_o_23_
  PIN dmi_req_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 269.96 600 270.16 ;
    END
  END dmi_req_o_24_
  PIN dmi_req_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 310.28 600 310.48 ;
    END
  END dmi_req_o_25_
  PIN dmi_req_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 267.44 600 267.64 ;
    END
  END dmi_req_o_26_
  PIN dmi_req_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 317.84 600 318.04 ;
    END
  END dmi_req_o_27_
  PIN dmi_req_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 338 600 338.2 ;
    END
  END dmi_req_o_28_
  PIN dmi_req_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 348.08 600 348.28 ;
    END
  END dmi_req_o_29_
  PIN dmi_req_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 285.08 600 285.28 ;
    END
  END dmi_req_o_2_
  PIN dmi_req_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 259.88 600 260.08 ;
    END
  END dmi_req_o_30_
  PIN dmi_req_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 275 600 275.2 ;
    END
  END dmi_req_o_31_
  PIN dmi_req_o_32_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 315.32 600 315.52 ;
    END
  END dmi_req_o_32_
  PIN dmi_req_o_33_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 353.12 600 353.32 ;
    END
  END dmi_req_o_33_
  PIN dmi_req_o_34_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 254.84 600 255.04 ;
    END
  END dmi_req_o_34_
  PIN dmi_req_o_35_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 264.92 600 265.12 ;
    END
  END dmi_req_o_35_
  PIN dmi_req_o_36_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 340.52 600 340.72 ;
    END
  END dmi_req_o_36_
  PIN dmi_req_o_37_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 292.64 600 292.84 ;
    END
  END dmi_req_o_37_
  PIN dmi_req_o_38_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 252.32 600 252.52 ;
    END
  END dmi_req_o_38_
  PIN dmi_req_o_39_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 320.36 600 320.56 ;
    END
  END dmi_req_o_39_
  PIN dmi_req_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 322.88 600 323.08 ;
    END
  END dmi_req_o_3_
  PIN dmi_req_o_40_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 325.4 600 325.6 ;
    END
  END dmi_req_o_40_
  PIN dmi_req_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 247.28 600 247.48 ;
    END
  END dmi_req_o_4_
  PIN dmi_req_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 262.4 600 262.6 ;
    END
  END dmi_req_o_5_
  PIN dmi_req_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 330.44 600 330.64 ;
    END
  END dmi_req_o_6_
  PIN dmi_req_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 350.6 600 350.8 ;
    END
  END dmi_req_o_7_
  PIN dmi_req_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 244.76 600 244.96 ;
    END
  END dmi_req_o_8_
  PIN dmi_req_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 305.24 600 305.44 ;
    END
  END dmi_req_o_9_
  PIN dmi_req_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 272.48 0.72 272.68 ;
    END
  END dmi_req_ready_i
  PIN dmi_req_valid_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 343.04 600 343.24 ;
    END
  END dmi_req_valid_o
  PIN dmi_resp_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 302.72 0.72 302.92 ;
    END
  END dmi_resp_i_0_
  PIN dmi_resp_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 257.36 0.72 257.56 ;
    END
  END dmi_resp_i_10_
  PIN dmi_resp_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 287.6 0.72 287.8 ;
    END
  END dmi_resp_i_11_
  PIN dmi_resp_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 307.76 0.72 307.96 ;
    END
  END dmi_resp_i_12_
  PIN dmi_resp_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 247.28 0.72 247.48 ;
    END
  END dmi_resp_i_13_
  PIN dmi_resp_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 295.16 0.72 295.36 ;
    END
  END dmi_resp_i_14_
  PIN dmi_resp_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 312.8 0.72 313 ;
    END
  END dmi_resp_i_15_
  PIN dmi_resp_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 315.32 0.72 315.52 ;
    END
  END dmi_resp_i_16_
  PIN dmi_resp_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 317.84 0.72 318.04 ;
    END
  END dmi_resp_i_17_
  PIN dmi_resp_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 267.44 0.72 267.64 ;
    END
  END dmi_resp_i_18_
  PIN dmi_resp_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 277.52 0.72 277.72 ;
    END
  END dmi_resp_i_19_
  PIN dmi_resp_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 297.68 0.72 297.88 ;
    END
  END dmi_resp_i_1_
  PIN dmi_resp_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 325.4 0.72 325.6 ;
    END
  END dmi_resp_i_20_
  PIN dmi_resp_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 290.12 0.72 290.32 ;
    END
  END dmi_resp_i_21_
  PIN dmi_resp_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 264.92 0.72 265.12 ;
    END
  END dmi_resp_i_22_
  PIN dmi_resp_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 330.44 0.72 330.64 ;
    END
  END dmi_resp_i_23_
  PIN dmi_resp_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 332.96 0.72 333.16 ;
    END
  END dmi_resp_i_24_
  PIN dmi_resp_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 254.84 0.72 255.04 ;
    END
  END dmi_resp_i_25_
  PIN dmi_resp_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 320.36 0.72 320.56 ;
    END
  END dmi_resp_i_26_
  PIN dmi_resp_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 338 0.72 338.2 ;
    END
  END dmi_resp_i_27_
  PIN dmi_resp_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 327.92 0.72 328.12 ;
    END
  END dmi_resp_i_28_
  PIN dmi_resp_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 285.08 0.72 285.28 ;
    END
  END dmi_resp_i_29_
  PIN dmi_resp_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 262.4 0.72 262.6 ;
    END
  END dmi_resp_i_2_
  PIN dmi_resp_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 249.8 0.72 250 ;
    END
  END dmi_resp_i_30_
  PIN dmi_resp_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 310.28 0.72 310.48 ;
    END
  END dmi_resp_i_31_
  PIN dmi_resp_i_32_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 282.56 0.72 282.76 ;
    END
  END dmi_resp_i_32_
  PIN dmi_resp_i_33_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 340.52 0.72 340.72 ;
    END
  END dmi_resp_i_33_
  PIN dmi_resp_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 300.2 0.72 300.4 ;
    END
  END dmi_resp_i_3_
  PIN dmi_resp_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 343.04 0.72 343.24 ;
    END
  END dmi_resp_i_4_
  PIN dmi_resp_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 280.04 0.72 280.24 ;
    END
  END dmi_resp_i_5_
  PIN dmi_resp_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 322.88 0.72 323.08 ;
    END
  END dmi_resp_i_6_
  PIN dmi_resp_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 259.88 0.72 260.08 ;
    END
  END dmi_resp_i_7_
  PIN dmi_resp_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 305.24 0.72 305.44 ;
    END
  END dmi_resp_i_8_
  PIN dmi_resp_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 252.32 0.72 252.52 ;
    END
  END dmi_resp_i_9_
  PIN dmi_resp_ready_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 257.36 600 257.56 ;
    END
  END dmi_resp_ready_o
  PIN dmi_resp_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 345.56 0.72 345.76 ;
    END
  END dmi_resp_valid_i
  PIN dmi_rst_no
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 287.6 600 287.8 ;
    END
  END dmi_rst_no
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 275 0.72 275.2 ;
    END
  END rst_ni
  PIN tck_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 348.08 0.72 348.28 ;
    END
  END tck_i
  PIN td_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 269.96 0.72 270.16 ;
    END
  END td_i
  PIN td_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 249.8 600 250 ;
    END
  END td_o
  PIN tdo_oe_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 327.92 600 328.12 ;
    END
  END tdo_oe_o
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 350.6 0.72 350.8 ;
    END
  END testmode_i
  PIN tms_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 292.64 0.72 292.84 ;
    END
  END tms_i
  PIN trst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 335.48 0.72 335.68 ;
    END
  END trst_ni
  OBS
    LAYER Metal1 ;
     RECT  25.44 26.24 574.56 237.64 ;
     RECT  25.44 237.64 575.12 239.32 ;
     RECT  25.44 239.32 575.6 251.5 ;
     RECT  25.44 251.5 576.08 255.02 ;
     RECT  12.4 259.9 12.56 262.58 ;
     RECT  598.96 256.12 599.12 263.68 ;
     RECT  595.12 263.68 599.12 270.14 ;
     RECT  7.12 275.02 7.28 283.16 ;
     RECT  25.44 255.02 575.6 285.1 ;
     RECT  24.88 285.1 575.6 286.52 ;
     RECT  598.96 270.14 599.12 305.42 ;
     RECT  25.44 286.52 575.6 310.72 ;
     RECT  24.88 310.72 575.6 312.82 ;
     RECT  23.92 312.82 575.6 316.76 ;
     RECT  25.44 316.76 575.6 319.7 ;
     RECT  25.44 319.7 575.12 334.82 ;
     RECT  25.44 334.82 574.56 345.58 ;
     RECT  25.44 345.58 575.12 348.1 ;
     RECT  25.44 348.1 575.6 357.5 ;
     RECT  25.44 357.5 575.12 365.06 ;
     RECT  25.44 365.06 574.56 574.78 ;
    LAYER Metal2 ;
     RECT  0.38 255.26 0.48 262.18 ;
     RECT  0.38 277.94 0.48 287.38 ;
     RECT  0.38 298.94 0.48 330.22 ;
     RECT  0.38 345.98 0.48 352.9 ;
     RECT  0.48 247.28 1.06 353.32 ;
     RECT  1.06 247.28 7.3 350.8 ;
     RECT  7.3 277.94 27.26 348.28 ;
     RECT  7.3 247.28 28.7 267.64 ;
     RECT  27.26 277.1 28.7 348.28 ;
     RECT  28.7 247.28 32.26 348.28 ;
     RECT  32.26 247.28 32.74 338.2 ;
     RECT  32.26 346.82 86.98 348.28 ;
     RECT  32.74 249.8 98.5 338.2 ;
     RECT  86.98 346.82 115.1 347.02 ;
     RECT  98.5 249.8 115.3 336.1 ;
     RECT  115.1 346.82 115.3 347.86 ;
     RECT  115.3 249.8 116.74 334.84 ;
     RECT  116.74 251.48 124.9 334.84 ;
     RECT  124.9 251.9 138.82 334.84 ;
     RECT  138.82 254.42 143.675 334.84 ;
     RECT  115.3 347.66 143.675 347.86 ;
     RECT  143.675 254.42 146.02 347.86 ;
     RECT  146.02 255.26 154.94 347.86 ;
     RECT  155.305 376.625 155.8 376.855 ;
     RECT  154.94 254.84 156.46 347.86 ;
     RECT  156.46 255.26 158.02 347.86 ;
     RECT  158.02 257.78 158.3 347.86 ;
     RECT  158.3 257.78 161.1 350.38 ;
     RECT  161.1 257.78 161.875 352.9 ;
     RECT  155.8 375.79 163.1 376.855 ;
     RECT  163.1 375.38 163.78 381.46 ;
     RECT  161.875 257.78 165.02 353.74 ;
     RECT  163.78 381.26 167.785 381.46 ;
     RECT  171.74 209.9 172.22 212.62 ;
     RECT  171.74 221.24 172.22 222.7 ;
     RECT  172.22 209.9 172.64 222.7 ;
     RECT  172.64 209.865 173.66 222.7 ;
     RECT  173.66 209.48 174.14 228.58 ;
     RECT  165.02 257.78 174.62 356.68 ;
     RECT  174.14 206.54 175.04 236.98 ;
     RECT  167.785 381.26 175.235 384.415 ;
     RECT  174.62 247.28 176.94 356.68 ;
     RECT  175.04 205.53 178.46 236.98 ;
     RECT  176.94 247.28 178.46 357.52 ;
     RECT  175.235 381.26 179.42 384.4 ;
     RECT  178.46 205.53 179.9 357.52 ;
     RECT  179.9 205.53 180.86 360.04 ;
     RECT  180.86 205.53 181.34 365.08 ;
     RECT  179.42 377.9 181.34 384.4 ;
     RECT  181.34 205.53 184.22 384.4 ;
     RECT  184.22 202.34 184.42 384.4 ;
     RECT  184.42 202.34 185.12 360.04 ;
     RECT  185.12 202.305 185.38 360.04 ;
     RECT  184.42 371.18 185.66 384.4 ;
     RECT  185.38 273.74 185.86 360.04 ;
     RECT  185.38 202.305 186.14 263.86 ;
     RECT  185.86 273.74 186.34 357.94 ;
     RECT  185.66 371.18 190.885 384.82 ;
     RECT  190.885 371.18 191.9 387.76 ;
     RECT  186.34 274.16 192.58 357.94 ;
     RECT  186.14 201.92 193.34 263.86 ;
     RECT  193.34 201.5 194.3 263.86 ;
     RECT  192.58 274.58 194.3 357.94 ;
     RECT  191.9 371.18 194.3 388.6 ;
     RECT  194.3 201.5 198.14 265.54 ;
     RECT  198.14 201.08 198.34 265.54 ;
     RECT  198.34 201.92 200.26 265.54 ;
     RECT  194.3 274.58 200.74 388.6 ;
     RECT  200.26 206.12 203.42 265.54 ;
     RECT  200.74 274.58 203.42 387.76 ;
     RECT  203.42 206.12 204.58 387.76 ;
     RECT  204.58 213.09 206.605 387.76 ;
     RECT  206.605 213.09 210.325 384.15 ;
     RECT  210.325 213.26 213.22 384.15 ;
     RECT  213.22 213.68 217.525 384.15 ;
     RECT  217.525 213.68 220.9 382.72 ;
     RECT  220.9 213.68 221.61 380.62 ;
     RECT  221.61 213.68 221.86 380.54 ;
     RECT  221.86 213.68 222.56 338.79 ;
     RECT  221.86 349.34 223.05 380.54 ;
     RECT  223.05 352.28 228.4 380.54 ;
     RECT  222.56 213.09 230.005 338.79 ;
     RECT  228.4 352.28 231.21 380.045 ;
     RECT  230.005 213.26 232.22 338.79 ;
     RECT  231.21 352.28 232.22 378.1 ;
     RECT  232.22 213.26 240.1 378.1 ;
     RECT  240.1 217.04 249.22 378.1 ;
     RECT  249.22 217.04 249.34 373.48 ;
     RECT  249.34 217.04 252.86 372.64 ;
     RECT  252.86 206.54 253.06 372.64 ;
     RECT  253.06 206.54 253.76 358.36 ;
     RECT  253.06 367.4 254.5 372.64 ;
     RECT  253.76 205.53 255.26 358.36 ;
     RECT  255.26 198.98 256.16 358.36 ;
     RECT  256.16 197.97 263.9 358.36 ;
     RECT  263.9 197.72 268.9 358.36 ;
     RECT  268.9 198.56 275.14 358.36 ;
     RECT  275.14 198.56 275.62 353.32 ;
     RECT  275.62 198.56 276.58 349.12 ;
     RECT  276.58 198.56 278.06 345.76 ;
     RECT  278.06 198.14 279.46 345.76 ;
     RECT  279.46 198.14 279.68 339.04 ;
     RECT  279.68 197.97 281.13 339.04 ;
     RECT  281.13 197.97 287.125 323.92 ;
     RECT  287.125 201.08 287.62 323.92 ;
     RECT  254.5 370.76 287.9 370.96 ;
     RECT  287.9 370.76 288.1 372.22 ;
     RECT  287.62 201.5 289.06 323.92 ;
     RECT  281.13 335.48 289.06 339.04 ;
     RECT  289.06 336.32 289.34 339.04 ;
     RECT  288.86 348.5 289.34 348.7 ;
     RECT  289.34 336.32 290.5 349.96 ;
     RECT  289.06 202.34 295.285 323.92 ;
     RECT  295.285 204.44 296.94 323.92 ;
     RECT  296.94 204.44 297.5 327.7 ;
     RECT  290.5 336.32 297.5 348.7 ;
     RECT  297.5 204.44 298.66 348.7 ;
     RECT  298.66 205.53 311.125 348.7 ;
     RECT  311.125 209.48 311.14 348.7 ;
     RECT  311.14 209.9 315.445 348.7 ;
     RECT  315.445 233.42 315.94 348.7 ;
     RECT  315.94 240.98 316.42 348.7 ;
     RECT  316.42 242.66 316.7 348.7 ;
     RECT  288.1 372.02 316.7 372.22 ;
     RECT  315.445 209.9 316.885 223.96 ;
     RECT  316.7 372.02 316.9 372.64 ;
     RECT  316.885 210.74 318.82 223.96 ;
     RECT  318.82 210.74 319.78 216.4 ;
     RECT  319.78 210.74 321.22 213.88 ;
     RECT  316.7 242.66 332.74 349.12 ;
     RECT  332.74 243.08 338.5 349.12 ;
     RECT  338.5 243.5 346.41 349.12 ;
     RECT  316.9 372.44 354.62 372.64 ;
     RECT  354.14 391.34 355.04 392.38 ;
     RECT  355.04 391.305 356.06 392.38 ;
     RECT  356.06 390.92 357.02 392.38 ;
     RECT  354.62 372.44 359.42 373.48 ;
     RECT  359.42 365.3 359.9 373.48 ;
     RECT  359.9 365.3 361.075 375.16 ;
     RECT  357.02 388.4 361.34 392.38 ;
     RECT  361.34 387.98 362.24 392.38 ;
     RECT  361.075 364.46 365.66 375.16 ;
     RECT  362.24 386.97 365.66 392.38 ;
     RECT  346.41 244.76 366.62 349.12 ;
     RECT  366.62 244.76 367.58 352.9 ;
     RECT  365.66 364.46 367.58 392.38 ;
     RECT  367.58 244.76 380.54 392.38 ;
     RECT  380.54 244.76 380.795 394.9 ;
     RECT  380.795 244.76 382.46 398.68 ;
     RECT  382.46 244.76 388.7 399.94 ;
     RECT  388.7 244.76 394.885 402.88 ;
     RECT  394.885 244.76 395.62 403.3 ;
     RECT  395.62 244.76 397.06 402.88 ;
     RECT  397.06 244.76 402.82 402.04 ;
     RECT  402.82 244.76 415.58 399.94 ;
     RECT  415.58 244.76 416.54 401.2 ;
     RECT  416.54 244.76 427.1 402.88 ;
     RECT  427.1 244.76 432.86 404.56 ;
     RECT  432.86 244.76 438.14 406.66 ;
     RECT  438.14 244.76 445.82 410.44 ;
     RECT  445.82 244.76 452.26 410.86 ;
     RECT  452.26 244.76 454.66 407.92 ;
     RECT  454.66 244.76 461.86 407.08 ;
     RECT  461.86 244.76 468.58 406.24 ;
     RECT  468.58 244.76 468.86 398.68 ;
     RECT  468.86 244.34 470.5 398.68 ;
     RECT  470.5 244.34 473.18 397.84 ;
     RECT  473.18 242.66 473.38 397.84 ;
     RECT  473.38 242.66 480.58 388.6 ;
     RECT  480.58 242.66 482.5 388.18 ;
     RECT  482.5 367.82 483.94 388.18 ;
     RECT  482.5 242.66 485.18 357.52 ;
     RECT  483.94 367.82 485.86 378.94 ;
     RECT  485.18 241.82 491.42 357.52 ;
     RECT  491.42 241.82 492.58 357.94 ;
     RECT  492.58 241.82 496.45 357.135 ;
     RECT  496.45 241.82 503.605 357.1 ;
     RECT  503.605 241.82 503.62 356.26 ;
     RECT  503.62 241.82 505.34 294.52 ;
     RECT  503.62 303.14 506.98 356.26 ;
     RECT  506.98 303.14 518.3 355.84 ;
     RECT  505.34 239.72 519.66 294.52 ;
     RECT  518.3 303.14 519.66 357.94 ;
     RECT  519.66 239.72 523.58 357.94 ;
     RECT  523.58 238.46 525.5 357.94 ;
     RECT  485.86 367.82 525.5 368.44 ;
     RECT  525.5 238.46 525.7 368.44 ;
     RECT  483.94 387.98 536.26 388.18 ;
     RECT  525.7 238.46 536.74 368.02 ;
     RECT  536.74 238.46 549.02 360.46 ;
     RECT  549.02 238.46 552.86 360.88 ;
     RECT  552.86 238.46 556.22 364.66 ;
     RECT  556.22 238.46 558.14 365.92 ;
     RECT  558.14 236.36 558.34 365.92 ;
     RECT  558.34 237.62 558.82 365.92 ;
     RECT  558.82 237.62 575.14 365.08 ;
     RECT  575.14 239.3 575.62 357.52 ;
     RECT  575.62 239.72 599.52 355.84 ;
     RECT  599.52 239.72 599.62 247.06 ;
     RECT  599.52 260.3 599.62 262.18 ;
     RECT  599.52 275.42 599.62 286.54 ;
     RECT  599.52 298.1 599.62 315.1 ;
     RECT  599.52 325.82 599.62 350.38 ;
    LAYER Metal3 ;
     RECT  261.5 198.14 269.38 198.56 ;
     RECT  280.7 198.14 280.9 198.56 ;
     RECT  260.54 198.56 280.9 199.4 ;
     RECT  193.34 201.5 193.54 201.92 ;
     RECT  191.42 201.92 200.26 202.34 ;
     RECT  190.46 202.34 200.26 203.18 ;
     RECT  260.54 199.4 290.5 203.18 ;
     RECT  187.1 203.18 200.26 206.12 ;
     RECT  260.54 203.18 298.66 206.12 ;
     RECT  309.5 205.7 309.7 206.12 ;
     RECT  257.66 206.12 309.7 206.96 ;
     RECT  176.06 206.12 200.26 209.48 ;
     RECT  213.02 213.26 213.22 213.68 ;
     RECT  231.26 213.26 235.3 213.68 ;
     RECT  257.66 206.96 314.5 213.88 ;
     RECT  173.66 209.48 200.26 214.1 ;
     RECT  173.66 214.1 203.14 214.52 ;
     RECT  213.02 213.68 238.66 214.52 ;
     RECT  173.66 214.52 238.66 217.04 ;
     RECT  173.66 217.04 241.06 217.24 ;
     RECT  257.66 213.88 311.14 217.24 ;
     RECT  257.66 217.24 310.18 217.46 ;
     RECT  176.06 217.24 241.06 218.3 ;
     RECT  252.38 217.46 310.18 224.38 ;
     RECT  295.1 224.38 310.18 227.74 ;
     RECT  176.06 218.3 242.02 228.8 ;
     RECT  252.38 224.38 282.82 228.8 ;
     RECT  176.06 228.8 282.82 236.14 ;
     RECT  186.62 236.14 282.82 236.36 ;
     RECT  565.34 235.52 567.46 236.36 ;
     RECT  537.02 238.88 537.22 239.3 ;
     RECT  295.58 227.74 310.18 239.72 ;
     RECT  507.26 239.3 507.46 239.72 ;
     RECT  506.78 239.72 507.46 240.14 ;
     RECT  528.38 239.3 537.22 240.14 ;
     RECT  556.7 236.36 567.46 240.34 ;
     RECT  506.3 240.14 507.46 240.56 ;
     RECT  294.62 239.72 310.18 240.98 ;
     RECT  186.62 236.36 284.26 242.66 ;
     RECT  186.62 242.66 284.74 243.08 ;
     RECT  294.62 240.98 316.42 243.08 ;
     RECT  497.66 240.56 514.18 243.08 ;
     RECT  335.9 242.66 336.1 243.5 ;
     RECT  477.98 240.56 478.18 243.7 ;
     RECT  186.62 243.08 316.42 244.34 ;
     RECT  186.62 244.34 324.58 246.86 ;
     RECT  335.9 243.5 338.5 246.86 ;
     RECT  186.62 246.86 338.5 247.06 ;
     RECT  349.82 243.92 350.02 247.28 ;
     RECT  497.66 243.08 515.62 247.28 ;
     RECT  527.9 240.14 545.86 247.28 ;
     RECT  349.82 247.28 355.3 247.7 ;
     RECT  349.82 247.7 359.14 248.12 ;
     RECT  369.98 247.28 370.18 248.12 ;
     RECT  490.46 247.28 545.86 250.64 ;
     RECT  176.06 236.14 176.26 251.06 ;
     RECT  186.62 247.06 199.78 251.06 ;
     RECT  469.34 246.44 470.5 251.06 ;
     RECT  176.06 251.06 199.78 251.26 ;
     RECT  44.54 248.12 44.74 251.48 ;
     RECT  209.66 247.06 338.5 251.48 ;
     RECT  349.82 248.12 370.18 251.48 ;
     RECT  381.5 251.06 381.7 251.48 ;
     RECT  456.38 250.64 456.58 251.48 ;
     RECT  468.38 251.06 470.5 251.48 ;
     RECT  481.34 250.64 546.34 251.48 ;
     RECT  556.7 240.34 566.98 251.48 ;
     RECT  481.34 251.48 566.98 251.68 ;
     RECT  133.34 250.64 135.46 251.9 ;
     RECT  33.98 251.48 44.74 252.32 ;
     RECT  32.06 252.32 44.74 254.42 ;
     RECT  121.82 251.48 122.02 254.42 ;
     RECT  133.34 251.9 138.82 254.42 ;
     RECT  31.1 254.42 44.74 254.84 ;
     RECT  121.82 254.42 143.62 254.84 ;
     RECT  209.66 251.48 388.9 254.84 ;
     RECT  456.38 251.48 470.5 254.84 ;
     RECT  481.34 251.68 566.5 254.84 ;
     RECT  91.58 254.84 91.78 255.68 ;
     RECT  121.82 254.84 157.06 255.68 ;
     RECT  30.62 254.84 44.74 256.1 ;
     RECT  209.66 254.84 396.1 256.1 ;
     RECT  121.82 255.68 164.26 257.36 ;
     RECT  176.06 251.26 197.38 257.36 ;
     RECT  91.58 255.68 100.42 257.78 ;
     RECT  209.66 256.1 400.42 258.2 ;
     RECT  436.22 257.78 436.42 258.62 ;
     RECT  121.82 257.36 197.38 258.82 ;
     RECT  453.98 254.84 566.5 258.82 ;
     RECT  453.98 258.82 513.22 259.24 ;
     RECT  209.66 258.2 402.34 259.46 ;
     RECT  430.46 258.62 436.42 259.46 ;
     RECT  30.62 256.1 53.86 259.66 ;
     RECT  453.98 259.24 508.9 259.66 ;
     RECT  31.1 259.66 53.86 260.08 ;
     RECT  121.82 258.82 183.94 261.56 ;
     RECT  121.34 261.56 183.94 262.4 ;
     RECT  430.46 259.46 443.62 262.4 ;
     RECT  118.94 262.4 183.94 262.6 ;
     RECT  427.58 262.4 443.62 265.34 ;
     RECT  453.98 259.66 507.94 265.34 ;
     RECT  194.3 258.82 197.38 265.54 ;
     RECT  31.58 260.08 53.86 265.76 ;
     RECT  91.58 257.78 108.1 266.6 ;
     RECT  209.66 259.46 411.94 266.6 ;
     RECT  427.58 265.34 507.94 266.6 ;
     RECT  209.66 266.6 412.9 266.8 ;
     RECT  90.62 266.6 109.06 267.02 ;
     RECT  118.94 262.6 179.62 267.02 ;
     RECT  211.1 266.8 412.9 267.02 ;
     RECT  424.7 266.6 507.94 267.02 ;
     RECT  523.1 258.82 566.5 267.02 ;
     RECT  90.62 267.02 179.62 267.44 ;
     RECT  211.1 267.02 507.94 268.48 ;
     RECT  213.98 268.48 507.94 269.96 ;
     RECT  523.1 267.02 566.98 269.96 ;
     RECT  31.58 265.76 60.1 270.58 ;
     RECT  86.3 267.44 179.62 270.58 ;
     RECT  86.3 270.58 148.9 271 ;
     RECT  213.98 269.96 566.98 273.1 ;
     RECT  160.22 270.58 179.62 273.74 ;
     RECT  31.58 270.58 55.78 274.16 ;
     RECT  160.22 273.74 186.34 276.26 ;
     RECT  86.78 271 148.9 277.72 ;
     RECT  160.22 276.26 191.62 278.36 ;
     RECT  219.26 273.1 566.98 278.56 ;
     RECT  160.22 278.36 200.74 278.78 ;
     RECT  28.7 274.16 55.78 280.88 ;
     RECT  143.42 277.72 148.9 280.88 ;
     RECT  160.22 278.78 203.62 280.88 ;
     RECT  28.7 280.88 58.18 281.5 ;
     RECT  30.14 281.5 58.18 282.14 ;
     RECT  86.78 277.72 132.58 282.14 ;
     RECT  519.26 278.56 566.98 282.34 ;
     RECT  143.42 280.88 203.62 282.56 ;
     RECT  143.42 282.56 205.54 284.86 ;
     RECT  143.42 284.86 203.62 285.7 ;
     RECT  84.86 282.14 132.58 285.92 ;
     RECT  219.26 278.56 509.38 286.34 ;
     RECT  30.14 282.14 60.1 288.02 ;
     RECT  537.02 282.34 566.98 288.44 ;
     RECT  519.26 282.34 526.66 289.06 ;
     RECT  30.14 288.02 63.94 289.28 ;
     RECT  81.02 285.92 132.58 289.28 ;
     RECT  143.42 285.7 202.66 289.28 ;
     RECT  216.86 286.34 509.38 289.28 ;
     RECT  519.26 289.06 525.22 289.28 ;
     RECT  30.14 289.28 202.66 289.48 ;
     RECT  537.02 288.44 569.38 292.42 ;
     RECT  216.86 289.28 525.22 292.84 ;
     RECT  472.7 292.84 507.94 293.26 ;
     RECT  537.5 292.42 569.38 293.26 ;
     RECT  518.78 292.84 525.22 293.68 ;
     RECT  30.14 289.48 120.58 293.9 ;
     RECT  489.5 293.26 507.94 294.1 ;
     RECT  490.46 294.1 507.94 294.52 ;
     RECT  472.7 293.26 478.18 294.94 ;
     RECT  216.86 292.84 456.58 296 ;
     RECT  151.1 289.48 202.66 296.42 ;
     RECT  151.1 296.42 203.14 296.62 ;
     RECT  179.9 296.62 203.14 296.84 ;
     RECT  216.38 296 456.58 297.26 ;
     RECT  179.9 296.84 203.62 297.68 ;
     RECT  151.1 296.62 169.06 297.88 ;
     RECT  179.9 297.68 204.1 299.36 ;
     RECT  215.42 297.26 456.58 299.36 ;
     RECT  29.18 293.9 120.58 299.78 ;
     RECT  132.86 289.48 138.82 299.78 ;
     RECT  151.1 297.88 168.58 299.78 ;
     RECT  519.74 293.68 525.22 303.56 ;
     RECT  179.9 299.36 456.58 303.98 ;
     RECT  475.1 294.94 478.18 303.98 ;
     RECT  490.94 294.52 507.94 303.98 ;
     RECT  519.74 303.56 527.14 303.98 ;
     RECT  179.9 303.98 457.06 304.4 ;
     RECT  490.94 303.98 527.14 304.4 ;
     RECT  537.5 293.26 567.46 304.4 ;
     RECT  29.18 299.78 168.58 304.82 ;
     RECT  179.9 304.4 464.26 304.82 ;
     RECT  475.1 303.98 478.66 304.82 ;
     RECT  488.54 304.4 527.14 304.82 ;
     RECT  179.9 304.82 527.14 307.76 ;
     RECT  537.02 304.4 567.46 307.76 ;
     RECT  179.9 307.76 567.46 308.38 ;
     RECT  28.22 304.82 168.58 308.6 ;
     RECT  179.9 308.38 490.18 308.6 ;
     RECT  28.22 308.6 490.18 311.74 ;
     RECT  28.22 311.74 169.06 313 ;
     RECT  28.22 313 131.14 313.42 ;
     RECT  179.9 311.74 490.18 314.26 ;
     RECT  183.26 314.26 490.18 315.52 ;
     RECT  29.18 313.42 131.14 315.94 ;
     RECT  500.06 308.38 538.18 315.94 ;
     RECT  185.18 315.52 440.26 316.78 ;
     RECT  500.06 315.94 509.38 316.78 ;
     RECT  521.66 315.94 538.18 318.68 ;
     RECT  549.5 308.38 567.46 318.68 ;
     RECT  521.66 318.68 568.42 319.72 ;
     RECT  555.26 319.72 568.42 320.14 ;
     RECT  74.78 315.94 131.14 322.24 ;
     RECT  185.18 316.78 438.82 322.24 ;
     RECT  0.86 272.48 1.06 322.88 ;
     RECT  75.26 322.24 131.14 322.88 ;
     RECT  143.9 313 169.06 322.88 ;
     RECT  29.18 315.94 63.94 323.08 ;
     RECT  291.74 322.24 438.82 323.08 ;
     RECT  453.5 315.52 490.18 323.5 ;
     RECT  475.58 323.5 490.18 323.92 ;
     RECT  75.26 322.88 169.06 326.66 ;
     RECT  297.5 323.08 438.82 326.66 ;
     RECT  453.5 323.5 464.74 326.66 ;
     RECT  501.5 316.78 509.38 326.66 ;
     RECT  75.26 326.66 174.82 326.86 ;
     RECT  29.18 323.08 57.22 327.28 ;
     RECT  567.26 320.14 568.42 327.28 ;
     RECT  51.26 327.28 51.46 327.7 ;
     RECT  75.26 326.86 75.46 327.7 ;
     RECT  85.82 326.86 131.14 327.7 ;
     RECT  297.5 326.66 464.74 327.7 ;
     RECT  85.82 327.7 122.5 328.12 ;
     RECT  598.46 327.08 598.66 328.12 ;
     RECT  297.5 327.7 391.78 328.54 ;
     RECT  86.78 328.12 122.5 329.38 ;
     RECT  144.38 326.86 174.82 329.6 ;
     RECT  185.18 322.24 280.42 329.6 ;
     RECT  86.78 329.38 114.82 329.8 ;
     RECT  555.26 320.14 557.38 330.02 ;
     RECT  29.18 327.28 41.38 330.64 ;
     RECT  86.78 329.8 105.22 330.64 ;
     RECT  86.78 330.64 88.9 331.06 ;
     RECT  300.38 328.54 391.78 331.06 ;
     RECT  489.02 323.92 490.18 331.28 ;
     RECT  501.02 326.66 509.38 331.28 ;
     RECT  521.66 319.72 544.42 331.28 ;
     RECT  555.26 330.02 566.02 331.28 ;
     RECT  30.14 330.64 41.38 331.48 ;
     RECT  98.78 330.64 101.38 331.48 ;
     RECT  300.38 331.06 383.62 333.58 ;
     RECT  475.58 323.92 478.66 333.8 ;
     RECT  489.02 331.28 566.02 333.8 ;
     RECT  336.86 333.58 383.62 334.42 ;
     RECT  475.58 333.8 566.02 334.42 ;
     RECT  403.1 327.7 464.74 334.64 ;
     RECT  475.58 334.42 496.42 334.64 ;
     RECT  99.26 331.48 101.38 334.84 ;
     RECT  144.38 329.6 280.42 334.84 ;
     RECT  300.38 333.58 326.98 334.84 ;
     RECT  336.86 334.42 351.94 334.84 ;
     RECT  555.74 334.42 566.02 337.16 ;
     RECT  362.3 334.42 383.62 337.36 ;
     RECT  338.78 334.84 351.94 337.78 ;
     RECT  300.38 334.84 313.06 338.2 ;
     RECT  338.78 337.78 347.14 338.2 ;
     RECT  373.34 337.36 383.62 338.2 ;
     RECT  403.1 334.64 496.42 338.2 ;
     RECT  300.38 338.2 307.78 338.62 ;
     RECT  340.22 338.2 347.14 338.62 ;
     RECT  555.74 337.16 566.98 338.84 ;
     RECT  30.14 331.48 32.26 340.72 ;
     RECT  305.66 338.62 307.78 341.14 ;
     RECT  346.94 338.62 347.14 341.14 ;
     RECT  403.1 338.2 465.7 341.36 ;
     RECT  144.38 334.84 224.26 341.98 ;
     RECT  307.58 341.14 307.78 341.98 ;
     RECT  555.74 338.84 567.46 341.98 ;
     RECT  400.22 341.36 465.7 342.2 ;
     RECT  0.38 322.88 1.06 342.4 ;
     RECT  395.9 342.2 465.7 342.62 ;
     RECT  381.98 338.2 383.62 343.04 ;
     RECT  395.42 342.62 465.7 343.04 ;
     RECT  32.06 340.72 32.26 343.24 ;
     RECT  153.98 341.98 224.26 344.5 ;
     RECT  156.86 344.5 224.26 345.14 ;
     RECT  235.58 334.84 280.42 345.14 ;
     RECT  475.58 338.2 496.42 346.18 ;
     RECT  156.86 345.14 280.42 346.6 ;
     RECT  156.86 346.6 277.06 347.02 ;
     RECT  475.58 346.18 479.62 347.02 ;
     RECT  86.78 331.06 86.98 348.28 ;
     RECT  477.98 347.02 479.62 348.7 ;
     RECT  381.98 343.04 465.7 348.92 ;
     RECT  489.5 346.18 496.42 348.92 ;
     RECT  507.26 334.42 545.38 348.92 ;
     RECT  489.5 348.92 545.38 349.34 ;
     RECT  555.74 341.98 566.98 349.34 ;
     RECT  156.86 347.02 206.5 349.54 ;
     RECT  381.02 348.92 465.7 349.76 ;
     RECT  489.5 349.34 566.98 349.96 ;
     RECT  380.54 349.76 465.7 350.18 ;
     RECT  158.3 349.54 206.5 350.38 ;
     RECT  216.86 347.02 277.06 350.8 ;
     RECT  216.86 350.8 275.62 351.22 ;
     RECT  380.54 350.18 466.66 352.48 ;
     RECT  531.74 349.96 566.98 352.48 ;
     RECT  0.38 342.4 0.58 352.9 ;
     RECT  161.18 350.38 206.5 352.9 ;
     RECT  216.86 351.22 264.58 352.9 ;
     RECT  478.94 348.7 479.62 352.9 ;
     RECT  216.86 352.9 264.1 353.32 ;
     RECT  274.94 351.22 275.62 353.32 ;
     RECT  161.18 352.9 166.66 354.16 ;
     RECT  489.5 349.96 516.58 354.16 ;
     RECT  489.5 354.16 504.1 355.84 ;
     RECT  161.18 354.16 165.22 356.68 ;
     RECT  216.86 353.32 263.14 356.68 ;
     RECT  177.02 352.9 206.5 356.9 ;
     RECT  177.02 356.9 206.98 357.32 ;
     RECT  216.86 356.68 256.42 357.32 ;
     RECT  177.02 357.32 256.42 357.52 ;
     RECT  489.5 355.84 500.26 357.52 ;
     RECT  542.3 352.48 566.98 357.52 ;
     RECT  179.9 357.52 256.42 357.94 ;
     RECT  491.42 357.52 500.26 357.94 ;
     RECT  274.94 353.32 275.14 358.36 ;
     RECT  366.62 352.7 366.82 359.84 ;
     RECT  179.9 357.94 253.06 360.04 ;
     RECT  478.94 352.9 479.14 360.26 ;
     RECT  531.74 352.48 531.94 360.46 ;
     RECT  366.62 359.84 368.26 360.68 ;
     RECT  380.54 352.48 463.3 360.68 ;
     RECT  192.86 360.04 253.06 360.88 ;
     RECT  549.02 357.52 566.98 360.88 ;
     RECT  500.06 357.94 500.26 361.72 ;
     RECT  552.86 360.88 566.98 361.72 ;
     RECT  195.26 360.88 253.06 364.24 ;
     RECT  552.86 361.72 566.5 364.24 ;
     RECT  552.86 364.24 563.14 364.66 ;
     RECT  473.66 360.26 479.14 364.88 ;
     RECT  556.22 364.66 563.14 365.08 ;
     RECT  558.14 365.08 563.14 365.5 ;
     RECT  233.66 364.24 253.06 367.18 ;
     RECT  473.66 364.88 481.54 367.82 ;
     RECT  366.62 360.68 463.3 368.02 ;
     RECT  367.58 368.02 463.3 368.24 ;
     RECT  473.66 367.82 482.5 368.24 ;
     RECT  195.26 364.24 223.3 371.6 ;
     RECT  181.82 360.04 182.02 372.44 ;
     RECT  193.34 371.6 223.3 372.44 ;
     RECT  367.58 368.24 482.5 373.9 ;
     RECT  181.82 372.44 223.3 375.8 ;
     RECT  233.66 367.18 249.22 375.8 ;
     RECT  181.82 375.8 249.22 376.42 ;
     RECT  161.18 356.68 163.3 376.84 ;
     RECT  249.02 376.42 249.22 378.1 ;
     RECT  368.06 373.9 482.5 378.94 ;
     RECT  181.82 376.42 234.82 379.78 ;
     RECT  416.06 378.94 482.5 379.78 ;
     RECT  220.22 379.78 234.82 380.2 ;
     RECT  163.1 376.84 163.3 381.46 ;
     RECT  368.06 378.94 406.18 383.14 ;
     RECT  416.54 379.78 482.5 383.14 ;
     RECT  368.06 383.14 371.14 383.56 ;
     RECT  381.02 383.14 406.18 383.56 ;
     RECT  181.82 379.78 210.34 383.98 ;
     RECT  181.82 383.98 205.06 384.4 ;
     RECT  368.06 383.56 368.74 387.34 ;
     RECT  416.54 383.14 482.02 387.34 ;
     RECT  191.42 384.4 205.06 387.76 ;
     RECT  368.54 387.34 368.74 387.76 ;
     RECT  416.54 387.34 481.06 387.76 ;
     RECT  191.9 387.76 192.58 388.18 ;
     RECT  192.38 388.18 192.58 388.6 ;
     RECT  416.54 387.76 477.22 388.6 ;
     RECT  388.7 383.56 406.18 388.82 ;
     RECT  388.7 388.82 406.66 390.5 ;
     RECT  416.54 388.6 471.46 390.5 ;
     RECT  388.7 390.5 471.46 394.9 ;
     RECT  390.62 394.9 471.46 398.26 ;
     RECT  390.62 398.26 401.38 398.68 ;
     RECT  414.62 398.26 471.46 398.68 ;
     RECT  414.62 398.68 468.58 399.1 ;
     RECT  415.58 399.1 468.58 401.2 ;
     RECT  394.94 398.68 397.06 401.62 ;
     RECT  395.42 401.62 397.06 402.88 ;
     RECT  416.54 401.2 468.58 402.88 ;
     RECT  395.42 402.88 395.62 403.3 ;
     RECT  427.1 402.88 468.58 404.56 ;
     RECT  432.86 404.56 468.58 406.24 ;
     RECT  432.86 406.24 449.86 406.66 ;
     RECT  461.66 406.24 461.86 407.08 ;
     RECT  438.14 406.66 449.86 410.02 ;
     RECT  438.14 410.02 446.5 410.44 ;
     RECT  446.3 410.44 446.5 410.86 ;
    LAYER Metal4 ;
     RECT  0.86 342.2 7.1 342.4 ;
     RECT  50.3 311.12 60.58 311.32 ;
     RECT  7.1 342.2 86.78 350.8 ;
     RECT  101.18 281.72 121.34 281.92 ;
     RECT  126.62 299.78 160.22 299.98 ;
     RECT  121.34 281.72 160.7 285.28 ;
     RECT  3.26 269.96 163.58 270.16 ;
     RECT  160.7 281.72 163.58 289.48 ;
     RECT  163.58 269.96 166.18 289.48 ;
     RECT  107.9 259.04 168.38 259.24 ;
     RECT  168.38 257.36 176.54 259.24 ;
     RECT  160.22 299.78 182.3 300.82 ;
     RECT  176.06 239.72 183.46 239.92 ;
     RECT  166.18 269.96 184.7 270.58 ;
     RECT  166.18 281.72 184.7 289.48 ;
     RECT  182.3 299.78 184.7 301.24 ;
     RECT  156.38 311.96 184.7 312.16 ;
     RECT  184.7 299.78 185.18 312.16 ;
     RECT  0.38 322.88 185.18 323.08 ;
     RECT  185.18 299.78 186.62 323.08 ;
     RECT  184.7 269.96 188.54 289.48 ;
     RECT  186.62 299.78 188.54 323.5 ;
     RECT  188.54 269.96 190.66 323.5 ;
     RECT  176.54 254.84 193.54 259.24 ;
     RECT  189.98 372.44 194.98 372.64 ;
     RECT  86.78 334.22 195.74 350.8 ;
     RECT  194.3 360.68 195.74 360.88 ;
     RECT  187.1 209.48 196.42 209.68 ;
     RECT  195.74 334.22 200.54 360.88 ;
     RECT  200.54 333.8 200.74 360.88 ;
     RECT  200.74 360.68 201.22 360.88 ;
     RECT  192.86 223.34 201.7 223.54 ;
     RECT  200.74 333.8 203.14 350.8 ;
     RECT  183.26 384.2 203.14 384.4 ;
     RECT  205.34 367.4 207.46 367.6 ;
     RECT  204.86 232.16 209.38 232.36 ;
     RECT  193.54 257.36 214.94 259.24 ;
     RECT  190.66 269.96 214.94 323.08 ;
     RECT  201.98 243.92 218.78 244.12 ;
     RECT  218.78 236.36 218.98 244.12 ;
     RECT  203.14 334.22 219.26 350.8 ;
     RECT  214.94 257.36 222.62 323.08 ;
     RECT  219.26 334.22 224.74 353.32 ;
     RECT  222.62 254.84 234.14 323.08 ;
     RECT  234.62 375.8 235.1 376 ;
     RECT  234.14 254.84 237.22 323.92 ;
     RECT  224.74 334.22 239.9 350.8 ;
     RECT  239.9 334.22 241.34 351.22 ;
     RECT  237.22 257.36 241.54 323.92 ;
     RECT  235.58 221.24 242.02 221.44 ;
     RECT  235.1 372.44 242.98 376 ;
     RECT  241.54 257.36 244.9 323.5 ;
     RECT  218.98 236.36 246.82 236.56 ;
     RECT  242.98 375.8 247.78 376 ;
     RECT  241.34 334.22 248.26 353.32 ;
     RECT  244.9 257.36 249.98 323.08 ;
     RECT  249.98 252.32 252.1 323.08 ;
     RECT  248.26 334.22 266.98 351.22 ;
     RECT  252.1 257.36 271.3 323.08 ;
     RECT  270.14 239.72 275.42 239.92 ;
     RECT  275.42 236.36 275.62 239.92 ;
     RECT  266.3 206.54 276.86 206.74 ;
     RECT  266.98 334.22 277.06 350.8 ;
     RECT  276.86 206.54 278.02 210.1 ;
     RECT  278.02 209.48 281.38 210.1 ;
     RECT  281.38 209.9 281.86 210.1 ;
     RECT  271.3 257.36 283.1 257.56 ;
     RECT  271.3 266.18 283.1 323.08 ;
     RECT  283.1 257.36 283.3 323.08 ;
     RECT  275.62 236.36 284.26 236.56 ;
     RECT  283.3 295.58 284.54 323.08 ;
     RECT  277.06 334.22 284.54 342.4 ;
     RECT  283.3 257.36 295.3 284.44 ;
     RECT  295.3 266.18 301.82 284.44 ;
     RECT  295.3 257.36 304.22 257.56 ;
     RECT  301.82 266.18 304.22 285.28 ;
     RECT  302.3 215.78 305.66 215.98 ;
     RECT  284.54 295.58 306.82 342.4 ;
     RECT  305.66 213.68 307.78 215.98 ;
     RECT  307.78 213.68 309.22 214.3 ;
     RECT  309.22 214.1 310.66 214.3 ;
     RECT  304.22 257.36 312.86 285.28 ;
     RECT  312.86 254 317.18 285.28 ;
     RECT  306.82 295.58 322.18 327.28 ;
     RECT  317.18 254 324.38 285.7 ;
     RECT  322.18 326.66 326.78 327.28 ;
     RECT  306.82 342.2 326.78 342.4 ;
     RECT  324.38 251.48 327.94 285.7 ;
     RECT  327.94 251.48 337.54 285.28 ;
     RECT  322.18 295.58 339.74 315.94 ;
     RECT  339.74 295.58 344.74 316.78 ;
     RECT  337.54 251.48 345.7 259.24 ;
     RECT  337.54 269.96 350.3 285.28 ;
     RECT  344.74 295.58 350.3 315.52 ;
     RECT  345.7 254.42 355.1 259.24 ;
     RECT  355.1 251.48 362.78 259.24 ;
     RECT  350.3 269.96 362.78 315.52 ;
     RECT  362.78 251.48 370.46 315.52 ;
     RECT  370.46 251.48 371.14 315.94 ;
     RECT  370.94 367.82 375.74 368.02 ;
     RECT  371.14 257.36 376.42 315.94 ;
     RECT  375.74 367.82 381.7 368.44 ;
     RECT  376.42 257.36 385.06 315.52 ;
     RECT  384.38 353.54 385.82 360.88 ;
     RECT  385.06 257.36 393.5 289.9 ;
     RECT  385.06 300.2 393.5 315.52 ;
     RECT  393.5 257.36 395.14 315.52 ;
     RECT  392.54 398.48 397.54 398.68 ;
     RECT  385.82 351.86 398.78 360.88 ;
     RECT  398.78 351.86 400.22 367.18 ;
     RECT  326.78 326.66 400.7 342.4 ;
     RECT  400.22 351.86 400.7 368.44 ;
     RECT  395.14 257.36 403.3 289.9 ;
     RECT  400.7 326.66 403.3 368.44 ;
     RECT  403.3 326.66 404.26 367.18 ;
     RECT  403.3 270.8 405.5 289.9 ;
     RECT  395.14 300.62 405.5 315.52 ;
     RECT  406.46 392.18 407.42 392.38 ;
     RECT  404.26 326.66 407.62 360.46 ;
     RECT  407.62 326.66 408.1 357.1 ;
     RECT  408.1 326.66 410.5 356.68 ;
     RECT  410.5 326.66 411.46 346.18 ;
     RECT  410.5 356.48 411.46 356.68 ;
     RECT  411.46 326.66 411.94 345.76 ;
     RECT  407.42 392.18 417.02 394.9 ;
     RECT  417.02 392.18 417.5 402.46 ;
     RECT  417.5 390.08 420.1 402.46 ;
     RECT  406.46 375.8 423.46 376 ;
     RECT  420.1 390.08 423.46 399.94 ;
     RECT  405.5 270.8 425.38 315.52 ;
     RECT  425.38 274.16 426.82 315.52 ;
     RECT  426.62 360.26 428.74 360.46 ;
     RECT  429.02 361.1 429.5 361.72 ;
     RECT  426.82 274.16 432.1 274.78 ;
     RECT  429.5 361.1 433.54 364.66 ;
     RECT  423.46 394.7 433.82 399.94 ;
     RECT  433.54 361.1 434.02 361.72 ;
     RECT  434.02 361.1 434.98 361.3 ;
     RECT  426.82 288.86 436.42 315.52 ;
     RECT  432.1 274.58 438.14 274.78 ;
     RECT  436.42 288.86 442.18 293.26 ;
     RECT  433.82 394.28 442.94 399.94 ;
     RECT  411.94 326.66 444.58 342.4 ;
     RECT  442.18 288.86 446.98 292.42 ;
     RECT  438.14 274.58 448.42 277.72 ;
     RECT  442.94 387.56 449.86 399.94 ;
     RECT  449.86 390.92 450.34 399.94 ;
     RECT  446.98 288.86 450.82 289.9 ;
     RECT  446.78 357.74 452.74 357.94 ;
     RECT  448.42 274.58 453.5 274.78 ;
     RECT  450.34 394.28 453.7 399.94 ;
     RECT  453.5 273.74 454.66 274.78 ;
     RECT  453.7 394.28 458.78 399.1 ;
     RECT  458.78 387.56 460.9 399.1 ;
     RECT  454.66 274.58 463.78 274.78 ;
     RECT  436.42 304.82 464.06 315.52 ;
     RECT  444.58 326.66 464.06 338.2 ;
     RECT  460.9 393.44 465.22 399.1 ;
     RECT  464.06 304.82 468.1 338.2 ;
     RECT  465.22 394.7 468.58 398.68 ;
     RECT  468.1 311.96 469.06 338.2 ;
     RECT  468.58 395.54 469.54 398.68 ;
     RECT  446.3 375.8 472.22 376 ;
     RECT  469.54 398.48 472.42 398.68 ;
     RECT  472.22 375.8 475.3 380.2 ;
     RECT  475.3 380 481.06 380.2 ;
     RECT  450.82 289.7 488.26 289.9 ;
     RECT  489.5 349.76 494.5 349.96 ;
     RECT  488.06 266.18 494.98 266.38 ;
     RECT  469.06 326.66 501.22 338.2 ;
     RECT  469.06 311.96 502.18 315.52 ;
     RECT  502.18 311.96 507.46 312.16 ;
     RECT  501.22 327.08 508.9 338.2 ;
     RECT  508.9 327.08 512.26 334.84 ;
     RECT  556.22 285.08 561.22 285.28 ;
     RECT  403.3 257.36 590.5 257.56 ;
     RECT  512.26 327.08 598.66 327.28 ;
    LAYER Metal5 ;
     RECT  403.58 356.06 403.78 365.08 ;
  END
END dmi_jtag
END LIBRARY
