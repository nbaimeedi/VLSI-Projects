VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO dm_top
  FOREIGN dm_top 0 0 ;
  CLASS BLOCK ;
  SIZE 600 BY 580.12 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VDDIO
    USE POWER ;
    DIRECTION INOUT ;
  END VDDIO
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN VSSIO
    USE GROUND ;
    DIRECTION INOUT ;
  END VSSIO
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 529.52 0.72 529.72 ;
    END
  END clk_i
  PIN debug_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 476.6 600 476.8 ;
    END
  END debug_req_o
  PIN dmactive_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 388.4 600 388.6 ;
    END
  END dmactive_o
  PIN dmi_req_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 300.2 0.72 300.4 ;
    END
  END dmi_req_i_0_
  PIN dmi_req_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 123.8 0.72 124 ;
    END
  END dmi_req_i_10_
  PIN dmi_req_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 297.68 0.72 297.88 ;
    END
  END dmi_req_i_11_
  PIN dmi_req_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 184.28 0.72 184.48 ;
    END
  END dmi_req_i_12_
  PIN dmi_req_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 307.76 0.72 307.96 ;
    END
  END dmi_req_i_13_
  PIN dmi_req_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 310.28 0.72 310.48 ;
    END
  END dmi_req_i_14_
  PIN dmi_req_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 262.4 0.72 262.6 ;
    END
  END dmi_req_i_15_
  PIN dmi_req_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 312.8 0.72 313 ;
    END
  END dmi_req_i_16_
  PIN dmi_req_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 181.76 0.72 181.96 ;
    END
  END dmi_req_i_17_
  PIN dmi_req_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 317.84 0.72 318.04 ;
    END
  END dmi_req_i_18_
  PIN dmi_req_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 292.64 0.72 292.84 ;
    END
  END dmi_req_i_19_
  PIN dmi_req_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 242.24 0.72 242.44 ;
    END
  END dmi_req_i_1_
  PIN dmi_req_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 121.28 0.72 121.48 ;
    END
  END dmi_req_i_20_
  PIN dmi_req_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 179.24 0.72 179.44 ;
    END
  END dmi_req_i_21_
  PIN dmi_req_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 290.12 0.72 290.32 ;
    END
  END dmi_req_i_22_
  PIN dmi_req_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 327.92 0.72 328.12 ;
    END
  END dmi_req_i_23_
  PIN dmi_req_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 330.44 0.72 330.64 ;
    END
  END dmi_req_i_24_
  PIN dmi_req_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 332.96 0.72 333.16 ;
    END
  END dmi_req_i_25_
  PIN dmi_req_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 176.72 0.72 176.92 ;
    END
  END dmi_req_i_26_
  PIN dmi_req_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 335.48 0.72 335.68 ;
    END
  END dmi_req_i_27_
  PIN dmi_req_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 338 0.72 338.2 ;
    END
  END dmi_req_i_28_
  PIN dmi_req_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 340.52 0.72 340.72 ;
    END
  END dmi_req_i_29_
  PIN dmi_req_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 285.08 0.72 285.28 ;
    END
  END dmi_req_i_2_
  PIN dmi_req_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 174.2 0.72 174.4 ;
    END
  END dmi_req_i_30_
  PIN dmi_req_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 118.76 0.72 118.96 ;
    END
  END dmi_req_i_31_
  PIN dmi_req_i_32_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 348.08 0.72 348.28 ;
    END
  END dmi_req_i_32_
  PIN dmi_req_i_33_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 282.56 0.72 282.76 ;
    END
  END dmi_req_i_33_
  PIN dmi_req_i_34_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 350.6 0.72 350.8 ;
    END
  END dmi_req_i_34_
  PIN dmi_req_i_35_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 171.68 0.72 171.88 ;
    END
  END dmi_req_i_35_
  PIN dmi_req_i_36_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 355.64 0.72 355.84 ;
    END
  END dmi_req_i_36_
  PIN dmi_req_i_37_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 93.56 0.72 93.76 ;
    END
  END dmi_req_i_37_
  PIN dmi_req_i_38_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 358.16 0.72 358.36 ;
    END
  END dmi_req_i_38_
  PIN dmi_req_i_39_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 154.04 0.72 154.24 ;
    END
  END dmi_req_i_39_
  PIN dmi_req_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 169.16 0.72 169.36 ;
    END
  END dmi_req_i_3_
  PIN dmi_req_i_40_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 116.24 0.72 116.44 ;
    END
  END dmi_req_i_40_
  PIN dmi_req_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 365.72 0.72 365.92 ;
    END
  END dmi_req_i_4_
  PIN dmi_req_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 368.24 0.72 368.44 ;
    END
  END dmi_req_i_5_
  PIN dmi_req_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 370.76 0.72 370.96 ;
    END
  END dmi_req_i_6_
  PIN dmi_req_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 166.64 0.72 166.84 ;
    END
  END dmi_req_i_7_
  PIN dmi_req_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 373.28 0.72 373.48 ;
    END
  END dmi_req_i_8_
  PIN dmi_req_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 375.8 0.72 376 ;
    END
  END dmi_req_i_9_
  PIN dmi_req_ready_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 436.28 600 436.48 ;
    END
  END dmi_req_ready_o
  PIN dmi_req_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 378.32 0.72 378.52 ;
    END
  END dmi_req_valid_i
  PIN dmi_resp_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 295.16 600 295.36 ;
    END
  END dmi_resp_o_0_
  PIN dmi_resp_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 292.64 600 292.84 ;
    END
  END dmi_resp_o_10_
  PIN dmi_resp_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 315.32 600 315.52 ;
    END
  END dmi_resp_o_11_
  PIN dmi_resp_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 390.92 600 391.12 ;
    END
  END dmi_resp_o_12_
  PIN dmi_resp_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 287.6 600 287.8 ;
    END
  END dmi_resp_o_13_
  PIN dmi_resp_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 343.04 600 343.24 ;
    END
  END dmi_resp_o_14_
  PIN dmi_resp_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 305.24 600 305.44 ;
    END
  END dmi_resp_o_15_
  PIN dmi_resp_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 282.56 600 282.76 ;
    END
  END dmi_resp_o_16_
  PIN dmi_resp_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 393.44 600 393.64 ;
    END
  END dmi_resp_o_17_
  PIN dmi_resp_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 277.52 600 277.72 ;
    END
  END dmi_resp_o_18_
  PIN dmi_resp_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 438.8 600 439 ;
    END
  END dmi_resp_o_19_
  PIN dmi_resp_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 275 600 275.2 ;
    END
  END dmi_resp_o_1_
  PIN dmi_resp_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 300.2 600 300.4 ;
    END
  END dmi_resp_o_20_
  PIN dmi_resp_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 395.96 600 396.16 ;
    END
  END dmi_resp_o_21_
  PIN dmi_resp_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 310.28 600 310.48 ;
    END
  END dmi_resp_o_22_
  PIN dmi_resp_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 267.44 600 267.64 ;
    END
  END dmi_resp_o_23_
  PIN dmi_resp_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 264.92 600 265.12 ;
    END
  END dmi_resp_o_24_
  PIN dmi_resp_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 262.4 600 262.6 ;
    END
  END dmi_resp_o_25_
  PIN dmi_resp_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 398.48 600 398.68 ;
    END
  END dmi_resp_o_26_
  PIN dmi_resp_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 441.32 600 441.52 ;
    END
  END dmi_resp_o_27_
  PIN dmi_resp_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 257.36 600 257.56 ;
    END
  END dmi_resp_o_28_
  PIN dmi_resp_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 254.84 600 255.04 ;
    END
  END dmi_resp_o_29_
  PIN dmi_resp_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 348.08 600 348.28 ;
    END
  END dmi_resp_o_2_
  PIN dmi_resp_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 401 600 401.2 ;
    END
  END dmi_resp_o_30_
  PIN dmi_resp_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 249.8 600 250 ;
    END
  END dmi_resp_o_31_
  PIN dmi_resp_o_32_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 247.28 600 247.48 ;
    END
  END dmi_resp_o_32_
  PIN dmi_resp_o_33_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 317.84 600 318.04 ;
    END
  END dmi_resp_o_33_
  PIN dmi_resp_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 443.84 600 444.04 ;
    END
  END dmi_resp_o_3_
  PIN dmi_resp_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 403.52 600 403.72 ;
    END
  END dmi_resp_o_4_
  PIN dmi_resp_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 239.72 600 239.92 ;
    END
  END dmi_resp_o_5_
  PIN dmi_resp_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 320.36 600 320.56 ;
    END
  END dmi_resp_o_6_
  PIN dmi_resp_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 237.2 600 237.4 ;
    END
  END dmi_resp_o_7_
  PIN dmi_resp_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 234.68 600 234.88 ;
    END
  END dmi_resp_o_8_
  PIN dmi_resp_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 406.04 600 406.24 ;
    END
  END dmi_resp_o_9_
  PIN dmi_resp_ready_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 272.48 0.72 272.68 ;
    END
  END dmi_resp_ready_i
  PIN dmi_resp_valid_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 461.48 600 461.68 ;
    END
  END dmi_resp_valid_o
  PIN dmi_rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 164.12 0.72 164.32 ;
    END
  END dmi_rst_ni
  PIN hartinfo_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 113.72 0.72 113.92 ;
    END
  END hartinfo_i_0_
  PIN hartinfo_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 385.88 0.72 386.08 ;
    END
  END hartinfo_i_10_
  PIN hartinfo_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 269.96 0.72 270.16 ;
    END
  END hartinfo_i_11_
  PIN hartinfo_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 388.4 0.72 388.6 ;
    END
  END hartinfo_i_12_
  PIN hartinfo_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 161.6 0.72 161.8 ;
    END
  END hartinfo_i_13_
  PIN hartinfo_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 267.44 0.72 267.64 ;
    END
  END hartinfo_i_14_
  PIN hartinfo_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 264.92 0.72 265.12 ;
    END
  END hartinfo_i_15_
  PIN hartinfo_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 395.96 0.72 396.16 ;
    END
  END hartinfo_i_16_
  PIN hartinfo_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 398.48 0.72 398.68 ;
    END
  END hartinfo_i_17_
  PIN hartinfo_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 159.08 0.72 159.28 ;
    END
  END hartinfo_i_18_
  PIN hartinfo_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 91.04 0.72 91.24 ;
    END
  END hartinfo_i_19_
  PIN hartinfo_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 403.52 0.72 403.72 ;
    END
  END hartinfo_i_1_
  PIN hartinfo_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 406.04 0.72 406.24 ;
    END
  END hartinfo_i_20_
  PIN hartinfo_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 408.56 0.72 408.76 ;
    END
  END hartinfo_i_21_
  PIN hartinfo_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 156.56 0.72 156.76 ;
    END
  END hartinfo_i_22_
  PIN hartinfo_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 411.08 0.72 411.28 ;
    END
  END hartinfo_i_23_
  PIN hartinfo_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 413.6 0.72 413.8 ;
    END
  END hartinfo_i_24_
  PIN hartinfo_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 416.12 0.72 416.32 ;
    END
  END hartinfo_i_25_
  PIN hartinfo_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 111.2 0.72 111.4 ;
    END
  END hartinfo_i_26_
  PIN hartinfo_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 418.64 0.72 418.84 ;
    END
  END hartinfo_i_27_
  PIN hartinfo_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 80.96 0.72 81.16 ;
    END
  END hartinfo_i_28_
  PIN hartinfo_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 423.68 0.72 423.88 ;
    END
  END hartinfo_i_29_
  PIN hartinfo_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 232.16 0.72 232.36 ;
    END
  END hartinfo_i_2_
  PIN hartinfo_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 426.2 0.72 426.4 ;
    END
  END hartinfo_i_30_
  PIN hartinfo_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 302.72 0.72 302.92 ;
    END
  END hartinfo_i_31_
  PIN hartinfo_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 151.52 0.72 151.72 ;
    END
  END hartinfo_i_3_
  PIN hartinfo_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 254.84 0.72 255.04 ;
    END
  END hartinfo_i_4_
  PIN hartinfo_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 433.76 0.72 433.96 ;
    END
  END hartinfo_i_5_
  PIN hartinfo_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 360.68 0.72 360.88 ;
    END
  END hartinfo_i_6_
  PIN hartinfo_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 275 0.72 275.2 ;
    END
  END hartinfo_i_7_
  PIN hartinfo_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 149 0.72 149.2 ;
    END
  END hartinfo_i_8_
  PIN hartinfo_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 441.32 0.72 441.52 ;
    END
  END hartinfo_i_9_
  PIN master_add_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 345.56 600 345.76 ;
    END
  END master_add_o_0_
  PIN master_add_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 227.12 600 227.32 ;
    END
  END master_add_o_10_
  PIN master_add_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 224.6 600 224.8 ;
    END
  END master_add_o_11_
  PIN master_add_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 408.56 600 408.76 ;
    END
  END master_add_o_12_
  PIN master_add_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 222.08 600 222.28 ;
    END
  END master_add_o_13_
  PIN master_add_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 219.56 600 219.76 ;
    END
  END master_add_o_14_
  PIN master_add_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 244.76 600 244.96 ;
    END
  END master_add_o_15_
  PIN master_add_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 327.92 600 328.12 ;
    END
  END master_add_o_16_
  PIN master_add_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 411.08 600 411.28 ;
    END
  END master_add_o_17_
  PIN master_add_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 212 600 212.2 ;
    END
  END master_add_o_18_
  PIN master_add_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 209.48 600 209.68 ;
    END
  END master_add_o_19_
  PIN master_add_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 330.44 600 330.64 ;
    END
  END master_add_o_1_
  PIN master_add_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 446.36 600 446.56 ;
    END
  END master_add_o_20_
  PIN master_add_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 413.6 600 413.8 ;
    END
  END master_add_o_21_
  PIN master_add_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 204.44 600 204.64 ;
    END
  END master_add_o_22_
  PIN master_add_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 332.96 600 333.16 ;
    END
  END master_add_o_23_
  PIN master_add_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 199.4 600 199.6 ;
    END
  END master_add_o_24_
  PIN master_add_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 302.72 600 302.92 ;
    END
  END master_add_o_25_
  PIN master_add_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 416.12 600 416.32 ;
    END
  END master_add_o_26_
  PIN master_add_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 335.48 600 335.68 ;
    END
  END master_add_o_27_
  PIN master_add_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 191.84 600 192.04 ;
    END
  END master_add_o_28_
  PIN master_add_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 338 600 338.2 ;
    END
  END master_add_o_29_
  PIN master_add_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 259.88 600 260.08 ;
    END
  END master_add_o_2_
  PIN master_add_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 448.88 600 449.08 ;
    END
  END master_add_o_30_
  PIN master_add_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 312.8 600 313 ;
    END
  END master_add_o_31_
  PIN master_add_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 418.64 600 418.84 ;
    END
  END master_add_o_3_
  PIN master_add_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 181.76 600 181.96 ;
    END
  END master_add_o_4_
  PIN master_add_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 340.52 600 340.72 ;
    END
  END master_add_o_5_
  PIN master_add_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 206.96 600 207.16 ;
    END
  END master_add_o_6_
  PIN master_add_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 176.72 600 176.92 ;
    END
  END master_add_o_7_
  PIN master_add_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 464 600 464.2 ;
    END
  END master_add_o_8_
  PIN master_add_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 360.68 600 360.88 ;
    END
  END master_add_o_9_
  PIN master_be_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 174.2 600 174.4 ;
    END
  END master_be_o_0_
  PIN master_be_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 297.68 600 297.88 ;
    END
  END master_be_o_1_
  PIN master_be_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 171.68 600 171.88 ;
    END
  END master_be_o_2_
  PIN master_be_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 421.16 600 421.36 ;
    END
  END master_be_o_3_
  PIN master_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 443.84 0.72 444.04 ;
    END
  END master_gnt_i
  PIN master_r_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 446.36 0.72 446.56 ;
    END
  END master_r_err_i
  PIN master_r_other_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 249.8 0.72 250 ;
    END
  END master_r_other_err_i
  PIN master_r_rdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 108.68 0.72 108.88 ;
    END
  END master_r_rdata_i_0_
  PIN master_r_rdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 451.4 0.72 451.6 ;
    END
  END master_r_rdata_i_10_
  PIN master_r_rdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 224.6 0.72 224.8 ;
    END
  END master_r_rdata_i_11_
  PIN master_r_rdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 247.28 0.72 247.48 ;
    END
  END master_r_rdata_i_12_
  PIN master_r_rdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 322.88 0.72 323.08 ;
    END
  END master_r_rdata_i_13_
  PIN master_r_rdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 458.96 0.72 459.16 ;
    END
  END master_r_rdata_i_14_
  PIN master_r_rdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 146.48 0.72 146.68 ;
    END
  END master_r_rdata_i_15_
  PIN master_r_rdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 244.76 0.72 244.96 ;
    END
  END master_r_rdata_i_16_
  PIN master_r_rdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 431.24 0.72 431.44 ;
    END
  END master_r_rdata_i_17_
  PIN master_r_rdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 277.52 0.72 277.72 ;
    END
  END master_r_rdata_i_18_
  PIN master_r_rdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 421.16 0.72 421.36 ;
    END
  END master_r_rdata_i_19_
  PIN master_r_rdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 88.52 0.72 88.72 ;
    END
  END master_r_rdata_i_1_
  PIN master_r_rdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 464 0.72 464.2 ;
    END
  END master_r_rdata_i_20_
  PIN master_r_rdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 453.92 0.72 454.12 ;
    END
  END master_r_rdata_i_21_
  PIN master_r_rdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 106.16 0.72 106.36 ;
    END
  END master_r_rdata_i_22_
  PIN master_r_rdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 239.72 0.72 239.92 ;
    END
  END master_r_rdata_i_23_
  PIN master_r_rdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 401 0.72 401.2 ;
    END
  END master_r_rdata_i_24_
  PIN master_r_rdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 438.8 0.72 439 ;
    END
  END master_r_rdata_i_25_
  PIN master_r_rdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 143.96 0.72 144.16 ;
    END
  END master_r_rdata_i_26_
  PIN master_r_rdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 237.2 0.72 237.4 ;
    END
  END master_r_rdata_i_27_
  PIN master_r_rdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 471.56 0.72 471.76 ;
    END
  END master_r_rdata_i_28_
  PIN master_r_rdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 380.84 0.72 381.04 ;
    END
  END master_r_rdata_i_29_
  PIN master_r_rdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 103.64 0.72 103.84 ;
    END
  END master_r_rdata_i_2_
  PIN master_r_rdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 234.68 0.72 234.88 ;
    END
  END master_r_rdata_i_30_
  PIN master_r_rdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 476.6 0.72 476.8 ;
    END
  END master_r_rdata_i_31_
  PIN master_r_rdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 363.2 0.72 363.4 ;
    END
  END master_r_rdata_i_3_
  PIN master_r_rdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 479.12 0.72 479.32 ;
    END
  END master_r_rdata_i_4_
  PIN master_r_rdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 141.44 0.72 141.64 ;
    END
  END master_r_rdata_i_5_
  PIN master_r_rdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 353.12 0.72 353.32 ;
    END
  END master_r_rdata_i_6_
  PIN master_r_rdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 466.52 0.72 466.72 ;
    END
  END master_r_rdata_i_7_
  PIN master_r_rdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 343.04 0.72 343.24 ;
    END
  END master_r_rdata_i_8_
  PIN master_r_rdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 229.64 0.72 229.84 ;
    END
  END master_r_rdata_i_9_
  PIN master_r_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 280.04 0.72 280.24 ;
    END
  END master_r_valid_i
  PIN master_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 214.52 600 214.72 ;
    END
  END master_req_o
  PIN master_wdata_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 169.16 600 169.36 ;
    END
  END master_wdata_o_0_
  PIN master_wdata_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 474.08 600 474.28 ;
    END
  END master_wdata_o_10_
  PIN master_wdata_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 451.4 600 451.6 ;
    END
  END master_wdata_o_11_
  PIN master_wdata_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 232.16 600 232.36 ;
    END
  END master_wdata_o_12_
  PIN master_wdata_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 164.12 600 164.32 ;
    END
  END master_wdata_o_13_
  PIN master_wdata_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 242.24 600 242.44 ;
    END
  END master_wdata_o_14_
  PIN master_wdata_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 350.6 600 350.8 ;
    END
  END master_wdata_o_15_
  PIN master_wdata_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 161.6 600 161.8 ;
    END
  END master_wdata_o_16_
  PIN master_wdata_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 252.32 600 252.52 ;
    END
  END master_wdata_o_17_
  PIN master_wdata_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 307.76 600 307.96 ;
    END
  END master_wdata_o_18_
  PIN master_wdata_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 353.12 600 353.32 ;
    END
  END master_wdata_o_19_
  PIN master_wdata_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 423.68 600 423.88 ;
    END
  END master_wdata_o_1_
  PIN master_wdata_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 269.96 600 270.16 ;
    END
  END master_wdata_o_20_
  PIN master_wdata_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 189.32 600 189.52 ;
    END
  END master_wdata_o_21_
  PIN master_wdata_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 355.64 600 355.84 ;
    END
  END master_wdata_o_22_
  PIN master_wdata_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 280.04 600 280.24 ;
    END
  END master_wdata_o_23_
  PIN master_wdata_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 166.64 600 166.84 ;
    END
  END master_wdata_o_24_
  PIN master_wdata_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 471.56 600 471.76 ;
    END
  END master_wdata_o_25_
  PIN master_wdata_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 358.16 600 358.36 ;
    END
  END master_wdata_o_26_
  PIN master_wdata_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 196.88 600 197.08 ;
    END
  END master_wdata_o_27_
  PIN master_wdata_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 453.92 600 454.12 ;
    END
  END master_wdata_o_28_
  PIN master_wdata_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 184.28 600 184.48 ;
    END
  END master_wdata_o_29_
  PIN master_wdata_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 426.2 600 426.4 ;
    END
  END master_wdata_o_2_
  PIN master_wdata_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 179.24 600 179.44 ;
    END
  END master_wdata_o_30_
  PIN master_wdata_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 466.52 600 466.72 ;
    END
  END master_wdata_o_31_
  PIN master_wdata_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 149 600 149.2 ;
    END
  END master_wdata_o_3_
  PIN master_wdata_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 363.2 600 363.4 ;
    END
  END master_wdata_o_4_
  PIN master_wdata_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 146.48 600 146.68 ;
    END
  END master_wdata_o_5_
  PIN master_wdata_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 143.96 600 144.16 ;
    END
  END master_wdata_o_6_
  PIN master_wdata_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 141.44 600 141.64 ;
    END
  END master_wdata_o_7_
  PIN master_wdata_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 365.72 600 365.92 ;
    END
  END master_wdata_o_8_
  PIN master_wdata_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 380.84 600 381.04 ;
    END
  END master_wdata_o_9_
  PIN master_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 229.64 600 229.84 ;
    END
  END master_we_o
  PIN ndmreset_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 486.68 0.72 486.88 ;
    END
  END ndmreset_ack_i
  PIN ndmreset_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 428.72 600 428.92 ;
    END
  END ndmreset_o
  PIN next_dm_addr_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 325.4 0.72 325.6 ;
    END
  END next_dm_addr_i_0_
  PIN next_dm_addr_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 227.12 0.72 227.32 ;
    END
  END next_dm_addr_i_10_
  PIN next_dm_addr_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 461.48 0.72 461.68 ;
    END
  END next_dm_addr_i_11_
  PIN next_dm_addr_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 315.32 0.72 315.52 ;
    END
  END next_dm_addr_i_12_
  PIN next_dm_addr_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 86 0.72 86.2 ;
    END
  END next_dm_addr_i_13_
  PIN next_dm_addr_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 138.92 0.72 139.12 ;
    END
  END next_dm_addr_i_14_
  PIN next_dm_addr_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 305.24 0.72 305.44 ;
    END
  END next_dm_addr_i_15_
  PIN next_dm_addr_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 491.72 0.72 491.92 ;
    END
  END next_dm_addr_i_16_
  PIN next_dm_addr_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 494.24 0.72 494.44 ;
    END
  END next_dm_addr_i_17_
  PIN next_dm_addr_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 222.08 0.72 222.28 ;
    END
  END next_dm_addr_i_18_
  PIN next_dm_addr_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 496.76 0.72 496.96 ;
    END
  END next_dm_addr_i_19_
  PIN next_dm_addr_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 456.44 0.72 456.64 ;
    END
  END next_dm_addr_i_1_
  PIN next_dm_addr_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 212 0.72 212.2 ;
    END
  END next_dm_addr_i_20_
  PIN next_dm_addr_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 219.56 0.72 219.76 ;
    END
  END next_dm_addr_i_21_
  PIN next_dm_addr_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 199.4 0.72 199.6 ;
    END
  END next_dm_addr_i_22_
  PIN next_dm_addr_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 393.44 0.72 393.64 ;
    END
  END next_dm_addr_i_23_
  PIN next_dm_addr_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 136.4 0.72 136.6 ;
    END
  END next_dm_addr_i_24_
  PIN next_dm_addr_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 217.04 0.72 217.24 ;
    END
  END next_dm_addr_i_25_
  PIN next_dm_addr_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 499.28 0.72 499.48 ;
    END
  END next_dm_addr_i_26_
  PIN next_dm_addr_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 390.92 0.72 391.12 ;
    END
  END next_dm_addr_i_27_
  PIN next_dm_addr_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 501.8 0.72 502 ;
    END
  END next_dm_addr_i_28_
  PIN next_dm_addr_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 214.52 0.72 214.72 ;
    END
  END next_dm_addr_i_29_
  PIN next_dm_addr_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 101.12 0.72 101.32 ;
    END
  END next_dm_addr_i_2_
  PIN next_dm_addr_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 252.32 0.72 252.52 ;
    END
  END next_dm_addr_i_30_
  PIN next_dm_addr_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 504.32 0.72 504.52 ;
    END
  END next_dm_addr_i_31_
  PIN next_dm_addr_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 186.8 0.72 187 ;
    END
  END next_dm_addr_i_3_
  PIN next_dm_addr_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 133.88 0.72 134.08 ;
    END
  END next_dm_addr_i_4_
  PIN next_dm_addr_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 287.6 0.72 287.8 ;
    END
  END next_dm_addr_i_5_
  PIN next_dm_addr_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 320.36 0.72 320.56 ;
    END
  END next_dm_addr_i_6_
  PIN next_dm_addr_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 209.48 0.72 209.68 ;
    END
  END next_dm_addr_i_7_
  PIN next_dm_addr_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 78.44 0.72 78.64 ;
    END
  END next_dm_addr_i_8_
  PIN next_dm_addr_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 481.64 0.72 481.84 ;
    END
  END next_dm_addr_i_9_
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 474.08 0.72 474.28 ;
    END
  END rst_ni
  PIN slave_addr_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 206.96 0.72 207.16 ;
    END
  END slave_addr_i_0_
  PIN slave_addr_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 257.36 0.72 257.56 ;
    END
  END slave_addr_i_10_
  PIN slave_addr_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 506.84 0.72 507.04 ;
    END
  END slave_addr_i_11_
  PIN slave_addr_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 579.92 0.72 580.12 ;
    END
  END slave_addr_i_12_
  PIN slave_addr_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 577.4 0.72 577.6 ;
    END
  END slave_addr_i_13_
  PIN slave_addr_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 574.88 0.72 575.08 ;
    END
  END slave_addr_i_14_
  PIN slave_addr_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 572.36 0.72 572.56 ;
    END
  END slave_addr_i_15_
  PIN slave_addr_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 569.84 0.72 570.04 ;
    END
  END slave_addr_i_16_
  PIN slave_addr_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 567.32 0.72 567.52 ;
    END
  END slave_addr_i_17_
  PIN slave_addr_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 564.8 0.72 565 ;
    END
  END slave_addr_i_18_
  PIN slave_addr_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 562.28 0.72 562.48 ;
    END
  END slave_addr_i_19_
  PIN slave_addr_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 131.36 0.72 131.56 ;
    END
  END slave_addr_i_1_
  PIN slave_addr_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 559.76 0.72 559.96 ;
    END
  END slave_addr_i_20_
  PIN slave_addr_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 557.24 0.72 557.44 ;
    END
  END slave_addr_i_21_
  PIN slave_addr_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 554.72 0.72 554.92 ;
    END
  END slave_addr_i_22_
  PIN slave_addr_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 552.2 0.72 552.4 ;
    END
  END slave_addr_i_23_
  PIN slave_addr_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 549.68 0.72 549.88 ;
    END
  END slave_addr_i_24_
  PIN slave_addr_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 547.16 0.72 547.36 ;
    END
  END slave_addr_i_25_
  PIN slave_addr_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 544.64 0.72 544.84 ;
    END
  END slave_addr_i_26_
  PIN slave_addr_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 542.12 0.72 542.32 ;
    END
  END slave_addr_i_27_
  PIN slave_addr_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 539.6 0.72 539.8 ;
    END
  END slave_addr_i_28_
  PIN slave_addr_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 537.08 0.72 537.28 ;
    END
  END slave_addr_i_29_
  PIN slave_addr_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 204.44 0.72 204.64 ;
    END
  END slave_addr_i_2_
  PIN slave_addr_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 534.56 0.72 534.76 ;
    END
  END slave_addr_i_30_
  PIN slave_addr_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 532.04 0.72 532.24 ;
    END
  END slave_addr_i_31_
  PIN slave_addr_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 345.56 0.72 345.76 ;
    END
  END slave_addr_i_3_
  PIN slave_addr_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 514.4 0.72 514.6 ;
    END
  END slave_addr_i_4_
  PIN slave_addr_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 516.92 0.72 517.12 ;
    END
  END slave_addr_i_5_
  PIN slave_addr_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 201.92 0.72 202.12 ;
    END
  END slave_addr_i_6_
  PIN slave_addr_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 511.88 0.72 512.08 ;
    END
  END slave_addr_i_7_
  PIN slave_addr_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 448.88 0.72 449.08 ;
    END
  END slave_addr_i_8_
  PIN slave_addr_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 519.44 0.72 519.64 ;
    END
  END slave_addr_i_9_
  PIN slave_be_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 128.84 0.72 129.04 ;
    END
  END slave_be_i_0_
  PIN slave_be_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 383.36 0.72 383.56 ;
    END
  END slave_be_i_1_
  PIN slave_be_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 484.16 0.72 484.36 ;
    END
  END slave_be_i_2_
  PIN slave_be_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 428.72 0.72 428.92 ;
    END
  END slave_be_i_3_
  PIN slave_rdata_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 368.24 600 368.44 ;
    END
  END slave_rdata_o_0_
  PIN slave_rdata_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 138.92 600 139.12 ;
    END
  END slave_rdata_o_10_
  PIN slave_rdata_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 154.04 600 154.24 ;
    END
  END slave_rdata_o_11_
  PIN slave_rdata_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 133.88 600 134.08 ;
    END
  END slave_rdata_o_12_
  PIN slave_rdata_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 370.76 600 370.96 ;
    END
  END slave_rdata_o_13_
  PIN slave_rdata_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 285.08 600 285.28 ;
    END
  END slave_rdata_o_14_
  PIN slave_rdata_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 322.88 600 323.08 ;
    END
  END slave_rdata_o_15_
  PIN slave_rdata_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 131.36 600 131.56 ;
    END
  END slave_rdata_o_16_
  PIN slave_rdata_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 373.28 600 373.48 ;
    END
  END slave_rdata_o_17_
  PIN slave_rdata_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 431.24 600 431.44 ;
    END
  END slave_rdata_o_18_
  PIN slave_rdata_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 272.48 600 272.68 ;
    END
  END slave_rdata_o_19_
  PIN slave_rdata_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 456.44 600 456.64 ;
    END
  END slave_rdata_o_1_
  PIN slave_rdata_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 375.8 600 376 ;
    END
  END slave_rdata_o_20_
  PIN slave_rdata_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 186.8 600 187 ;
    END
  END slave_rdata_o_21_
  PIN slave_rdata_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 128.84 600 129.04 ;
    END
  END slave_rdata_o_22_
  PIN slave_rdata_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 126.32 600 126.52 ;
    END
  END slave_rdata_o_23_
  PIN slave_rdata_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 378.32 600 378.52 ;
    END
  END slave_rdata_o_24_
  PIN slave_rdata_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 156.56 600 156.76 ;
    END
  END slave_rdata_o_25_
  PIN slave_rdata_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 194.36 600 194.56 ;
    END
  END slave_rdata_o_26_
  PIN slave_rdata_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 217.04 600 217.24 ;
    END
  END slave_rdata_o_27_
  PIN slave_rdata_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 433.76 600 433.96 ;
    END
  END slave_rdata_o_28_
  PIN slave_rdata_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 290.12 600 290.32 ;
    END
  END slave_rdata_o_29_
  PIN slave_rdata_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 469.04 600 469.24 ;
    END
  END slave_rdata_o_2_
  PIN slave_rdata_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 136.4 600 136.6 ;
    END
  END slave_rdata_o_30_
  PIN slave_rdata_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 383.36 600 383.56 ;
    END
  END slave_rdata_o_31_
  PIN slave_rdata_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 151.52 600 151.72 ;
    END
  END slave_rdata_o_3_
  PIN slave_rdata_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 159.08 600 159.28 ;
    END
  END slave_rdata_o_4_
  PIN slave_rdata_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 458.96 600 459.16 ;
    END
  END slave_rdata_o_5_
  PIN slave_rdata_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 385.88 600 386.08 ;
    END
  END slave_rdata_o_6_
  PIN slave_rdata_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 123.8 600 124 ;
    END
  END slave_rdata_o_7_
  PIN slave_rdata_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 201.92 600 202.12 ;
    END
  END slave_rdata_o_8_
  PIN slave_rdata_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  599.28 325.4 600 325.6 ;
    END
  END slave_rdata_o_9_
  PIN slave_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 196.88 0.72 197.08 ;
    END
  END slave_req_i
  PIN slave_wdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 98.6 0.72 98.8 ;
    END
  END slave_wdata_i_0_
  PIN slave_wdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 259.88 0.72 260.08 ;
    END
  END slave_wdata_i_10_
  PIN slave_wdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 469.04 0.72 469.24 ;
    END
  END slave_wdata_i_11_
  PIN slave_wdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 194.36 0.72 194.56 ;
    END
  END slave_wdata_i_12_
  PIN slave_wdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 126.32 0.72 126.52 ;
    END
  END slave_wdata_i_13_
  PIN slave_wdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 295.16 0.72 295.36 ;
    END
  END slave_wdata_i_14_
  PIN slave_wdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 521.96 0.72 522.16 ;
    END
  END slave_wdata_i_15_
  PIN slave_wdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 191.84 0.72 192.04 ;
    END
  END slave_wdata_i_16_
  PIN slave_wdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 524.48 0.72 524.68 ;
    END
  END slave_wdata_i_17_
  PIN slave_wdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 509.36 0.72 509.56 ;
    END
  END slave_wdata_i_18_
  PIN slave_wdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 83.48 0.72 83.68 ;
    END
  END slave_wdata_i_19_
  PIN slave_wdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 189.32 0.72 189.52 ;
    END
  END slave_wdata_i_1_
  PIN slave_wdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 436.28 0.72 436.48 ;
    END
  END slave_wdata_i_20_
  PIN slave_wdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 527 0.72 527.2 ;
    END
  END slave_wdata_i_21_
  PIN slave_wdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 489.2 0.72 489.4 ;
    END
  END slave_wdata_i_22_
  PIN slave_wdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 96.08 0.72 96.28 ;
    END
  END slave_wdata_i_23_
  PIN slave_wdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 33.08 0.72 33.28 ;
    END
  END slave_wdata_i_24_
  PIN slave_wdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 63.32 0.72 63.52 ;
    END
  END slave_wdata_i_25_
  PIN slave_wdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 40.64 0.72 40.84 ;
    END
  END slave_wdata_i_26_
  PIN slave_wdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 48.2 0.72 48.4 ;
    END
  END slave_wdata_i_27_
  PIN slave_wdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 65.84 0.72 66.04 ;
    END
  END slave_wdata_i_28_
  PIN slave_wdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 50.72 0.72 50.92 ;
    END
  END slave_wdata_i_29_
  PIN slave_wdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 73.4 0.72 73.6 ;
    END
  END slave_wdata_i_2_
  PIN slave_wdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 58.28 0.72 58.48 ;
    END
  END slave_wdata_i_30_
  PIN slave_wdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 35.6 0.72 35.8 ;
    END
  END slave_wdata_i_31_
  PIN slave_wdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 38.12 0.72 38.32 ;
    END
  END slave_wdata_i_3_
  PIN slave_wdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 70.88 0.72 71.08 ;
    END
  END slave_wdata_i_4_
  PIN slave_wdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 45.68 0.72 45.88 ;
    END
  END slave_wdata_i_5_
  PIN slave_wdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 75.92 0.72 76.12 ;
    END
  END slave_wdata_i_6_
  PIN slave_wdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 53.24 0.72 53.44 ;
    END
  END slave_wdata_i_7_
  PIN slave_wdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 60.8 0.72 61 ;
    END
  END slave_wdata_i_8_
  PIN slave_wdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 43.16 0.72 43.36 ;
    END
  END slave_wdata_i_9_
  PIN slave_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 68.36 0.72 68.56 ;
    END
  END slave_we_i
  PIN testmode_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 30.56 0.72 30.76 ;
    END
  END testmode_i
  PIN unavailable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 55.76 0.72 55.96 ;
    END
  END unavailable_i
  OBS
    LAYER Metal1 ;
     RECT  0.88 65.86 1.04 88.54 ;
     RECT  20.16 22.46 579.84 88.54 ;
     RECT  598.96 176.74 599.12 181.78 ;
     RECT  598 181.78 599.12 189.34 ;
     RECT  0.88 88.54 579.84 204.2 ;
     RECT  595.6 189.34 599.12 205.04 ;
     RECT  597.04 205.04 599.12 219.58 ;
     RECT  594.16 219.58 599.12 222.1 ;
     RECT  1.36 204.2 579.84 225.04 ;
     RECT  593.68 222.1 599.12 227.14 ;
     RECT  590.32 227.14 599.12 242 ;
     RECT  593.68 242 599.12 249.14 ;
     RECT  596.08 249.14 599.12 256.28 ;
     RECT  596.08 256.28 598.64 263.42 ;
     RECT  597.04 263.42 598.64 283.16 ;
     RECT  597.04 283.16 597.2 335.92 ;
     RECT  597.04 335.92 597.68 343.48 ;
     RECT  597.04 343.48 598.64 360.86 ;
     RECT  597.04 360.86 598.16 363.22 ;
     RECT  589.84 363.22 598.16 364.64 ;
     RECT  597.04 364.64 598.16 366.32 ;
     RECT  0.4 225.04 579.84 370.52 ;
     RECT  597.52 366.32 598.16 377.5 ;
     RECT  0.4 370.52 2.48 391.78 ;
     RECT  0.4 391.78 4.88 392.2 ;
     RECT  0.4 392.2 6.32 393.46 ;
     RECT  0.4 393.46 7.28 406.22 ;
     RECT  597.52 377.5 599.6 413.36 ;
     RECT  0.4 406.22 6.8 416.3 ;
     RECT  0.4 416.3 4.88 423.86 ;
     RECT  597.52 413.36 599.12 436.46 ;
     RECT  597.52 436.46 598.64 446.54 ;
     RECT  0.4 423.86 2.48 461.66 ;
     RECT  597.52 446.54 597.68 461.66 ;
     RECT  17.68 370.52 579.84 479.3 ;
     RECT  0.4 461.66 2 481.82 ;
     RECT  0.4 481.82 1.52 504.5 ;
     RECT  0.4 504.5 1.04 522.14 ;
     RECT  0.4 522.14 0.56 529.28 ;
     RECT  20.16 479.3 579.84 578.56 ;
    LAYER Metal2 ;
     RECT  0.38 94.4 0.48 95.86 ;
     RECT  0.38 126.74 0.48 128.62 ;
     RECT  0.38 144.38 0.48 146.26 ;
     RECT  0.38 182.18 0.48 184.06 ;
     RECT  0.38 232.58 0.48 232.78 ;
     RECT  0.38 295.58 0.48 297.46 ;
     RECT  0.38 338.84 0.48 355.42 ;
     RECT  0.38 376.22 0.48 377.26 ;
     RECT  0.38 471.98 0.48 473.86 ;
     RECT  0.38 529.1 0.48 529.3 ;
     RECT  0.48 33.08 1.06 529.72 ;
     RECT  1.06 33.08 3.46 527.2 ;
     RECT  3.46 86 4.42 255.04 ;
     RECT  3.46 264.92 4.42 527.2 ;
     RECT  4.42 391.76 6.34 527.2 ;
     RECT  4.42 264.92 6.82 381.04 ;
     RECT  6.34 416.12 6.82 527.2 ;
     RECT  4.42 86 7.3 224.8 ;
     RECT  4.42 234.68 7.3 255.04 ;
     RECT  6.82 264.92 7.3 282.76 ;
     RECT  6.82 291.38 7.3 381.04 ;
     RECT  6.34 391.76 7.3 406.24 ;
     RECT  7.3 88.52 10.66 108.88 ;
     RECT  6.82 421.16 10.66 527.2 ;
     RECT  10.66 94.4 11.14 108.88 ;
     RECT  7.3 234.68 11.62 247.48 ;
     RECT  7.3 141.44 12.1 146.68 ;
     RECT  7.3 277.52 13.06 280.24 ;
     RECT  11.14 94.4 14.5 106.36 ;
     RECT  7.3 291.38 17.66 345.34 ;
     RECT  7.3 354.38 17.66 381.04 ;
     RECT  14.5 94.82 17.86 106.36 ;
     RECT  10.66 421.16 17.86 479.32 ;
     RECT  7.3 174.2 19.58 192.04 ;
     RECT  7.3 204.02 19.58 204.64 ;
     RECT  7.3 216.62 19.58 224.8 ;
     RECT  17.86 421.16 20.26 476.8 ;
     RECT  19.58 163.7 20.74 195.4 ;
     RECT  11.62 234.68 20.905 244.96 ;
     RECT  13.06 280.04 20.905 280.24 ;
     RECT  17.66 291.38 21.22 381.04 ;
     RECT  7.3 121.28 21.385 129.04 ;
     RECT  20.905 261.965 21.4 262.195 ;
     RECT  12.1 146.06 21.98 146.68 ;
     RECT  20.74 163.7 21.98 194.98 ;
     RECT  19.58 204.02 21.98 224.8 ;
     RECT  20.905 234.68 21.98 252.115 ;
     RECT  21.385 121.28 22.46 131.155 ;
     RECT  21.98 141.44 22.46 146.68 ;
     RECT  17.86 106.16 22.94 106.36 ;
     RECT  22.46 119.6 22.94 131.155 ;
     RECT  22.46 141.44 22.94 150.88 ;
     RECT  21.98 159.92 22.94 194.98 ;
     RECT  20.26 466.52 23.14 476.8 ;
     RECT  21.98 204.02 23.42 252.115 ;
     RECT  21.4 261.965 23.42 263.03 ;
     RECT  7.3 391.76 23.62 401.2 ;
     RECT  20.905 280.04 24.38 282.355 ;
     RECT  21.22 291.38 24.38 377.68 ;
     RECT  23.42 204.02 24.86 263.03 ;
     RECT  24.38 278.36 24.86 377.68 ;
     RECT  17.86 94.82 25.705 95.44 ;
     RECT  23.14 469.04 26.02 476.8 ;
     RECT  20.26 421.16 27.94 456.64 ;
     RECT  22.94 106.16 29.18 194.98 ;
     RECT  24.86 204.02 29.18 377.68 ;
     RECT  26.02 469.04 29.86 472.18 ;
     RECT  29.18 106.16 33.5 377.68 ;
     RECT  25.705 88.085 33.98 95.44 ;
     RECT  33.5 105.32 33.98 377.68 ;
     RECT  33.865 72.965 34.36 73.195 ;
     RECT  27.94 426.2 35.62 456.64 ;
     RECT  3.46 33.08 35.9 63.52 ;
     RECT  33.98 88.085 37.34 377.68 ;
     RECT  34.36 72.965 37.82 74.03 ;
     RECT  37.82 72.965 38.3 76.54 ;
     RECT  37.34 85.16 38.3 377.68 ;
     RECT  35.9 33.08 39.145 63.94 ;
     RECT  38.3 72.965 39.145 377.68 ;
     RECT  39.145 33.08 41.66 377.68 ;
     RECT  41.66 33.08 91.1 378.1 ;
     RECT  35.62 436.28 102.82 456.64 ;
     RECT  10.66 489.2 105.22 527.2 ;
     RECT  91.1 33.08 107.14 378.52 ;
     RECT  107.14 35.6 114.14 378.52 ;
     RECT  23.62 391.76 115.1 394.06 ;
     RECT  114.14 35.6 117.5 379.78 ;
     RECT  117.5 35.6 118.46 380.62 ;
     RECT  118.46 35.6 124.7 381.04 ;
     RECT  115.1 390.5 124.7 394.06 ;
     RECT  105.22 489.2 128.26 524.68 ;
     RECT  124.7 35.6 133.54 394.06 ;
     RECT  133.54 54.5 139.3 394.06 ;
     RECT  139.3 54.92 142.645 394.06 ;
     RECT  128.26 496.76 142.66 524.68 ;
     RECT  142.66 516.92 145.54 524.68 ;
     RECT  142.645 55.76 146.02 394.06 ;
     RECT  29.86 469.04 154.66 469.24 ;
     RECT  133.54 35.6 158.02 43.36 ;
     RECT  142.66 496.76 158.02 507.04 ;
     RECT  146.02 56.18 159.69 394.06 ;
     RECT  159.69 56.18 165.5 381.04 ;
     RECT  158.02 38.12 166.94 43.36 ;
     RECT  165.5 51.98 166.94 381.04 ;
     RECT  158.02 496.76 170.98 496.96 ;
     RECT  166.94 38.12 173.66 381.04 ;
     RECT  159.69 390.5 173.66 394.06 ;
     RECT  173.66 38.12 194.5 394.06 ;
     RECT  194.5 38.12 199.78 43.36 ;
     RECT  102.82 441.32 205.54 456.64 ;
     RECT  194.5 51.98 215.295 394.06 ;
     RECT  215.295 51.14 216.86 394.06 ;
     RECT  216.86 50.72 218.02 394.06 ;
     RECT  218.02 50.72 218.72 388.6 ;
     RECT  199.78 38.12 220.42 38.32 ;
     RECT  205.54 443.84 220.42 456.64 ;
     RECT  218.72 50.55 220.585 388.6 ;
     RECT  220.585 47.765 221.08 388.6 ;
     RECT  221.08 46.93 223.58 388.6 ;
     RECT  35.62 426.2 223.78 426.4 ;
     RECT  223.58 43.58 225.22 388.6 ;
     RECT  225.22 46.52 227.42 388.6 ;
     RECT  227.42 46.52 228.82 390.28 ;
     RECT  228.82 46.52 229.34 391.33 ;
     RECT  229.34 46.52 229.82 391.54 ;
     RECT  229.82 46.52 244.9 392.38 ;
     RECT  145.54 516.92 248.26 519.64 ;
     RECT  158.02 506.84 250.66 507.04 ;
     RECT  220.42 443.84 254.5 449.08 ;
     RECT  244.9 46.52 258.34 391.54 ;
     RECT  258.34 46.94 261.02 391.54 ;
     RECT  261.02 46.94 262.18 394.48 ;
     RECT  248.26 516.92 262.66 517.12 ;
     RECT  262.18 51.14 263.42 394.48 ;
     RECT  263.42 51.14 265.06 395.74 ;
     RECT  265.06 54.92 271.285 395.74 ;
     RECT  271.285 55.76 273.02 395.74 ;
     RECT  273.02 55.76 273.43 399.1 ;
     RECT  273.43 55.76 274.66 395.74 ;
     RECT  274.66 58.11 275.125 395.74 ;
     RECT  275.125 59.54 278.5 395.74 ;
     RECT  278.5 65.67 284.74 395.74 ;
     RECT  284.74 65.67 286.18 395.32 ;
     RECT  286.18 65.67 286.645 394.9 ;
     RECT  286.645 65.84 288.1 394.9 ;
     RECT  288.1 68.78 289.06 394.9 ;
     RECT  289.06 72.14 290.02 394.9 ;
     RECT  290.02 72.14 293.38 391.54 ;
     RECT  293.38 77.17 295.685 391.54 ;
     RECT  295.685 77.18 296.74 391.54 ;
     RECT  296.74 77.18 302.02 391.12 ;
     RECT  302.02 82.22 302.405 391.12 ;
     RECT  302.405 103.47 302.485 391.12 ;
     RECT  302.485 104.9 302.965 391.12 ;
     RECT  302.405 82.22 305.365 93.09 ;
     RECT  302.965 104.9 307.3 388.6 ;
     RECT  305.365 82.22 307.78 91.66 ;
     RECT  307.78 91.46 308.74 91.66 ;
     RECT  307.3 104.9 308.74 115.18 ;
     RECT  308.74 104.9 309.22 105.1 ;
     RECT  308.74 114.56 309.22 114.76 ;
     RECT  307.3 125.06 311.42 388.6 ;
     RECT  311.42 125.06 316.42 392.38 ;
     RECT  316.42 125.06 320.74 391.54 ;
     RECT  320.74 125.06 320.98 390.7 ;
     RECT  320.98 125.06 327.94 388.6 ;
     RECT  327.94 125.06 331.78 384.82 ;
     RECT  331.78 125.06 333.7 383.99 ;
     RECT  333.7 126.74 341.285 383.99 ;
     RECT  254.5 443.84 346.66 446.56 ;
     RECT  341.285 126.74 351.46 380.62 ;
     RECT  351.46 130.52 351.925 380.62 ;
     RECT  351.925 130.94 361.82 380.62 ;
     RECT  361.82 130.1 366.62 380.62 ;
     RECT  366.62 130.1 374.5 381.04 ;
     RECT  374.5 132.62 386.78 381.04 ;
     RECT  386.78 130.52 387.26 381.04 ;
     RECT  387.26 130.1 387.46 381.04 ;
     RECT  387.46 132.62 393.7 381.04 ;
     RECT  393.7 133.46 395.9 381.04 ;
     RECT  346.66 443.84 413.86 444.04 ;
     RECT  412.22 471.56 418.46 471.76 ;
     RECT  419.42 123.8 423.74 124 ;
     RECT  395.9 133.46 423.74 381.46 ;
     RECT  418.46 466.52 425.66 471.76 ;
     RECT  423.74 123.8 429.02 381.46 ;
     RECT  422.78 453.92 429.02 454.12 ;
     RECT  429.02 123.8 429.22 382.72 ;
     RECT  246.62 428.72 430.46 428.92 ;
     RECT  429.22 123.8 434.5 381.04 ;
     RECT  429.02 451.4 434.78 454.12 ;
     RECT  434.5 123.8 447.74 379.36 ;
     RECT  447.74 123.8 451.58 381.46 ;
     RECT  451.58 123.8 453.5 382.72 ;
     RECT  453.5 123.8 453.98 386.5 ;
     RECT  434.78 451.4 454.94 456.64 ;
     RECT  425.66 466.52 454.94 474.28 ;
     RECT  453.98 123.8 457.34 387.34 ;
     RECT  457.34 123.8 459.26 390.28 ;
     RECT  430.46 421.16 459.74 428.92 ;
     RECT  459.26 123.8 472.22 392.38 ;
     RECT  472.22 123.8 472.9 394.06 ;
     RECT  472.9 159.08 474.14 394.06 ;
     RECT  474.14 159.08 474.33 396.16 ;
     RECT  472.9 123.8 474.34 149.62 ;
     RECT  474.34 143.96 474.82 149.62 ;
     RECT  474.82 143.96 475.3 145 ;
     RECT  474.33 159.08 475.3 214.72 ;
     RECT  475.3 172.1 476.26 202.12 ;
     RECT  476.26 201.92 476.98 202.12 ;
     RECT  476.26 172.1 477.22 173.14 ;
     RECT  475.3 159.08 478.18 159.7 ;
     RECT  476.26 183.02 478.18 190.78 ;
     RECT  472.22 441.32 488.06 441.52 ;
     RECT  454.94 451.4 488.06 474.28 ;
     RECT  459.74 421.16 488.54 431.44 ;
     RECT  488.06 441.32 488.54 474.28 ;
     RECT  474.33 229.64 490.94 396.16 ;
     RECT  475.3 214.52 503.9 214.72 ;
     RECT  490.94 229.64 510.62 403.72 ;
     RECT  510.62 229.64 514.66 406.24 ;
     RECT  514.66 353.96 518.02 406.24 ;
     RECT  503.9 214.52 518.3 216.82 ;
     RECT  514.66 229.64 524.54 344.5 ;
     RECT  524.54 229.64 524.74 348.28 ;
     RECT  478.18 185.54 528.86 185.74 ;
     RECT  478.18 159.08 536.06 159.28 ;
     RECT  518.02 362.78 542.02 406.24 ;
     RECT  474.34 123.8 590.3 134.08 ;
     RECT  500.06 146.48 590.3 146.68 ;
     RECT  536.06 159.08 590.3 166.84 ;
     RECT  528.86 185.54 590.3 192.04 ;
     RECT  528.86 204.86 590.3 205.06 ;
     RECT  518.3 214.52 590.3 217.24 ;
     RECT  524.74 229.64 590.3 320.56 ;
     RECT  524.74 329.18 590.3 348.28 ;
     RECT  542.02 364.04 590.3 406.24 ;
     RECT  590.3 123.8 593.66 217.24 ;
     RECT  590.3 227.12 593.66 348.28 ;
     RECT  593.66 123.8 594.62 348.28 ;
     RECT  590.3 358.16 594.62 406.24 ;
     RECT  488.54 421.16 596.06 474.28 ;
     RECT  594.62 123.8 597.5 406.24 ;
     RECT  596.06 416.12 597.5 474.28 ;
     RECT  597.5 123.8 598.94 474.28 ;
     RECT  598.94 123.8 599.52 476.8 ;
     RECT  599.52 185.54 599.62 186.58 ;
     RECT  599.52 247.7 599.62 249.58 ;
     RECT  599.52 262.82 599.62 264.7 ;
     RECT  599.52 290.54 599.62 292.42 ;
     RECT  599.52 329.18 599.62 330.22 ;
     RECT  599.52 340.94 599.62 342.82 ;
     RECT  599.52 364.04 599.62 365.5 ;
     RECT  599.52 382.1 599.62 383.14 ;
     RECT  599.52 413.18 599.62 413.38 ;
    LAYER Metal3 ;
     RECT  220.22 38.12 220.42 43.58 ;
     RECT  220.22 43.58 225.22 46.52 ;
     RECT  253.82 46.52 254.02 46.94 ;
     RECT  220.22 46.52 230.02 50.3 ;
     RECT  106.94 33.08 107.14 50.72 ;
     RECT  220.22 50.3 231.46 50.72 ;
     RECT  186.62 50.72 186.82 51.14 ;
     RECT  157.82 35.6 158.02 51.56 ;
     RECT  168.86 50.72 169.06 51.56 ;
     RECT  253.82 46.94 262.18 51.56 ;
     RECT  215.9 50.72 237.7 53.24 ;
     RECT  249.5 51.56 262.18 53.24 ;
     RECT  182.3 51.14 187.78 54.08 ;
     RECT  199.58 43.16 199.78 54.08 ;
     RECT  133.34 48.2 133.54 54.5 ;
     RECT  157.82 51.56 169.06 54.5 ;
     RECT  182.3 54.08 199.78 54.5 ;
     RECT  103.1 50.72 107.14 54.92 ;
     RECT  119.9 40.64 120.1 54.92 ;
     RECT  133.34 54.5 139.3 54.92 ;
     RECT  157.82 54.5 169.54 54.92 ;
     RECT  181.34 54.5 199.78 54.92 ;
     RECT  215.9 53.24 262.18 54.92 ;
     RECT  133.34 54.92 142.66 55.76 ;
     RECT  103.1 54.92 120.1 58.28 ;
     RECT  133.34 55.76 143.62 58.28 ;
     RECT  92.54 58.28 120.1 58.7 ;
     RECT  129.98 58.28 143.62 58.7 ;
     RECT  157.82 54.92 203.14 58.7 ;
     RECT  215.9 54.92 267.94 59.12 ;
     RECT  156.38 58.7 203.62 59.54 ;
     RECT  214.94 59.12 267.94 59.54 ;
     RECT  92.54 58.7 143.62 62.06 ;
     RECT  65.18 62.06 66.34 62.48 ;
     RECT  91.1 62.06 143.62 62.48 ;
     RECT  61.82 62.48 69.22 63.32 ;
     RECT  91.1 62.48 144.1 63.32 ;
     RECT  61.82 63.32 144.1 63.94 ;
     RECT  156.38 59.54 273.22 65 ;
     RECT  44.06 61.64 44.26 65.84 ;
     RECT  61.82 63.94 76.42 65.84 ;
     RECT  89.18 63.94 144.1 65.84 ;
     RECT  156.38 65 275.14 65.84 ;
     RECT  89.18 65.84 275.14 66.68 ;
     RECT  89.18 66.68 276.1 67.1 ;
     RECT  287.9 65.84 288.1 67.1 ;
     RECT  89.18 67.1 290.02 68.36 ;
     RECT  44.06 65.84 76.42 73.82 ;
     RECT  44.06 73.82 77.86 74.66 ;
     RECT  44.06 74.66 78.34 75.92 ;
     RECT  89.18 68.36 292.9 75.92 ;
     RECT  0.86 65.84 1.06 77.18 ;
     RECT  44.06 75.92 292.9 77.18 ;
     RECT  44.06 77.18 298.66 78.44 ;
     RECT  41.18 78.44 298.66 80.96 ;
     RECT  41.18 80.96 301.54 84.74 ;
     RECT  40.7 84.74 301.54 86 ;
     RECT  38.3 86 301.54 86.84 ;
     RECT  38.3 86.84 302.98 88.1 ;
     RECT  29.66 88.1 302.98 89.36 ;
     RECT  28.7 89.36 302.98 96.7 ;
     RECT  28.7 96.7 301.54 114.56 ;
     RECT  25.34 114.56 301.54 119.38 ;
     RECT  28.7 119.38 301.54 122.32 ;
     RECT  28.7 122.32 297.7 122.74 ;
     RECT  30.62 122.74 297.7 124.84 ;
     RECT  0.86 77.18 6.34 126.74 ;
     RECT  308.54 122.54 309.22 127.16 ;
     RECT  320.06 125.06 320.26 127.16 ;
     RECT  308.54 127.16 320.26 130.1 ;
     RECT  335.9 127.58 336.1 130.1 ;
     RECT  352.22 126.74 352.42 130.1 ;
     RECT  362.3 129.68 362.5 130.1 ;
     RECT  308.54 130.1 336.1 130.52 ;
     RECT  352.22 130.1 362.5 130.52 ;
     RECT  386.3 130.1 386.5 130.52 ;
     RECT  386.3 130.52 386.98 131.36 ;
     RECT  308.54 130.52 362.5 133.88 ;
     RECT  386.3 131.36 387.46 133.88 ;
     RECT  386.3 133.88 393.22 134.3 ;
     RECT  380.06 134.3 393.22 135.14 ;
     RECT  405.98 134.3 406.18 135.14 ;
     RECT  30.62 124.84 297.22 135.56 ;
     RECT  308.54 133.88 363.46 135.56 ;
     RECT  374.3 135.14 393.22 135.56 ;
     RECT  30.62 135.56 363.46 136.82 ;
     RECT  373.82 135.56 393.22 136.82 ;
     RECT  405.5 135.14 406.18 136.82 ;
     RECT  417.02 136.4 417.22 136.82 ;
     RECT  30.62 136.82 393.22 137.66 ;
     RECT  405.5 136.82 417.22 137.66 ;
     RECT  431.9 137.24 432.1 137.66 ;
     RECT  25.82 137.66 393.22 138.08 ;
     RECT  405.5 137.66 432.58 138.08 ;
     RECT  442.46 137.66 442.66 138.08 ;
     RECT  453.02 138.5 453.22 139.34 ;
     RECT  474.62 131.36 474.82 139.76 ;
     RECT  452.54 139.34 453.22 141.44 ;
     RECT  452.54 141.44 454.18 141.86 ;
     RECT  466.46 139.76 474.82 141.86 ;
     RECT  25.82 138.08 442.66 142.7 ;
     RECT  452.54 141.86 474.82 142.7 ;
     RECT  25.82 142.7 474.82 148.78 ;
     RECT  593.18 149.84 593.38 150.68 ;
     RECT  25.82 148.78 474.34 156.56 ;
     RECT  593.18 150.68 594.82 156.56 ;
     RECT  593.18 156.56 598.66 157.6 ;
     RECT  23.42 156.56 474.34 164.96 ;
     RECT  593.18 157.6 593.38 167.48 ;
     RECT  23.42 164.96 474.82 167.9 ;
     RECT  23.42 167.9 475.78 172.1 ;
     RECT  23.42 172.1 477.22 174.82 ;
     RECT  23.42 174.82 476.74 175.66 ;
     RECT  0.86 126.74 10.66 176.92 ;
     RECT  23.42 175.66 475.3 179.66 ;
     RECT  22.46 179.66 475.3 186.38 ;
     RECT  536.06 166.64 536.26 191.84 ;
     RECT  22.46 186.38 476.26 194.98 ;
     RECT  593.18 167.48 599.14 202.12 ;
     RECT  23.9 194.98 476.26 205.28 ;
     RECT  23.42 205.28 476.26 205.9 ;
     RECT  23.42 205.9 473.86 210.1 ;
     RECT  23.9 210.1 469.54 212.2 ;
     RECT  0.86 176.92 6.34 214.52 ;
     RECT  528.86 191.84 536.26 217.04 ;
     RECT  0.86 214.52 7.3 219.98 ;
     RECT  23.9 212.2 467.62 222.08 ;
     RECT  23.9 222.08 468.1 222.28 ;
     RECT  23.9 222.28 467.62 228.16 ;
     RECT  0.86 219.98 10.66 232.58 ;
     RECT  23.9 228.16 351.94 234.68 ;
     RECT  362.3 228.16 467.62 237.5 ;
     RECT  22.94 234.68 351.94 238.04 ;
     RECT  362.3 237.5 468.58 238.04 ;
     RECT  22.94 238.04 468.58 241.18 ;
     RECT  0.38 232.58 10.66 244.76 ;
     RECT  22.94 241.18 383.62 244.76 ;
     RECT  393.5 241.18 468.58 247.28 ;
     RECT  393.5 247.28 475.3 248.54 ;
     RECT  0.38 244.76 383.62 251.9 ;
     RECT  393.5 248.54 482.98 251.9 ;
     RECT  0.38 251.9 482.98 252.32 ;
     RECT  0.38 252.32 486.34 255.88 ;
     RECT  593.18 202.12 598.66 256.1 ;
     RECT  0.86 255.88 486.34 258.62 ;
     RECT  0.86 258.62 489.22 263.86 ;
     RECT  0.86 263.86 475.3 270.16 ;
     RECT  485.66 263.86 489.22 273.32 ;
     RECT  0.86 270.16 474.34 273.52 ;
     RECT  485.66 273.32 492.1 278.78 ;
     RECT  484.7 278.78 492.1 282.56 ;
     RECT  0.86 273.52 473.86 284.66 ;
     RECT  484.7 282.56 495.94 284.66 ;
     RECT  505.82 262.4 506.02 285.08 ;
     RECT  505.82 285.08 511.3 286.34 ;
     RECT  528.86 217.04 543.46 286.34 ;
     RECT  0.86 284.66 495.94 286.76 ;
     RECT  505.82 286.34 543.46 286.76 ;
     RECT  0.86 286.76 543.46 293.06 ;
     RECT  568.7 300.2 568.9 307.12 ;
     RECT  0.38 293.06 543.46 310.9 ;
     RECT  0.38 310.9 512.26 312.16 ;
     RECT  528.86 310.9 543.46 313.84 ;
     RECT  593.18 256.1 599.14 319.52 ;
     RECT  0.38 312.16 509.86 324.14 ;
     RECT  0.38 324.14 517.54 327.08 ;
     RECT  0.38 327.08 518.02 331.06 ;
     RECT  118.94 331.06 518.02 333.8 ;
     RECT  118.94 333.8 521.38 334.42 ;
     RECT  120.38 334.42 521.38 338.2 ;
     RECT  536.06 313.84 543.46 338.62 ;
     RECT  120.38 338.2 519.94 339.04 ;
     RECT  0.38 331.06 109.06 345.56 ;
     RECT  120.38 339.04 511.3 345.56 ;
     RECT  590.78 319.52 599.14 345.76 ;
     RECT  592.22 345.76 599.14 346.18 ;
     RECT  0.38 345.56 511.3 350.6 ;
     RECT  0.38 350.6 518.02 357.1 ;
     RECT  0.38 357.1 508.42 360.04 ;
     RECT  399.74 360.04 508.42 364.24 ;
     RECT  592.7 346.18 599.14 364.66 ;
     RECT  0.38 360.04 388.9 365.92 ;
     RECT  0.38 365.92 387.94 366.34 ;
     RECT  453.5 364.24 508.42 369.5 ;
     RECT  399.74 364.24 439.78 369.7 ;
     RECT  402.62 369.7 439.78 371.8 ;
     RECT  404.06 371.8 439.78 372.22 ;
     RECT  453.5 369.5 509.38 372.22 ;
     RECT  0.38 366.34 378.82 373.9 ;
     RECT  0.38 373.9 55.78 375.58 ;
     RECT  543.26 338.62 543.46 376 ;
     RECT  55.58 375.58 55.78 376.42 ;
     RECT  66.62 373.9 378.82 376.42 ;
     RECT  66.62 376.42 66.82 376.84 ;
     RECT  454.94 372.22 509.38 376.84 ;
     RECT  77.18 376.42 77.38 377.26 ;
     RECT  91.1 376.42 378.82 377.26 ;
     RECT  0.38 375.58 41.86 378.1 ;
     RECT  404.54 372.22 439.78 378.1 ;
     RECT  91.1 377.26 366.82 378.52 ;
     RECT  102.62 378.52 366.82 379.36 ;
     RECT  404.54 378.1 434.98 379.78 ;
     RECT  117.98 379.36 366.82 380.2 ;
     RECT  117.98 380.2 346.66 380.62 ;
     RECT  366.62 380.2 366.82 381.04 ;
     RECT  124.7 380.62 346.66 383.14 ;
     RECT  124.7 383.14 331.78 383.98 ;
     RECT  341.66 383.14 346.66 383.98 ;
     RECT  124.7 383.98 158.5 384.4 ;
     RECT  171.26 383.98 320.74 384.4 ;
     RECT  171.26 384.4 176.26 384.82 ;
     RECT  187.1 384.4 320.74 384.82 ;
     RECT  330.62 383.98 331.78 384.82 ;
     RECT  191.9 384.82 320.74 385.24 ;
     RECT  198.14 385.24 320.74 386.5 ;
     RECT  330.62 384.82 330.82 386.5 ;
     RECT  198.14 386.5 296.26 386.92 ;
     RECT  205.34 386.92 296.26 387.76 ;
     RECT  454.94 376.84 507.94 387.76 ;
     RECT  0.38 378.1 32.26 388.9 ;
     RECT  306.14 386.5 320.74 390.28 ;
     RECT  243.74 387.76 296.26 391.33 ;
     RECT  205.34 387.76 230.02 391.54 ;
     RECT  244.7 391.33 296.26 391.54 ;
     RECT  311.42 390.28 320.74 391.54 ;
     RECT  470.3 387.76 493.54 391.54 ;
     RECT  487.1 391.54 491.14 391.96 ;
     RECT  244.7 391.54 289.54 392.38 ;
     RECT  311.42 391.54 311.62 392.38 ;
     RECT  205.34 391.54 210.34 393.22 ;
     RECT  246.62 392.38 289.54 394.48 ;
     RECT  273.98 394.48 284.74 394.9 ;
     RECT  273.98 394.9 278.98 395.74 ;
     RECT  474.14 391.54 474.34 396.16 ;
     RECT  273.98 395.74 275.14 398.68 ;
     RECT  274.46 398.68 274.66 399.1 ;
     RECT  507.74 387.76 507.94 401.2 ;
     RECT  488.54 391.96 491.14 403.72 ;
     RECT  171.26 384.82 171.46 417.5 ;
     RECT  220.7 391.54 223.78 417.5 ;
     RECT  488.54 403.72 488.74 417.5 ;
     RECT  128.06 384.4 158.5 417.7 ;
     RECT  170.78 417.5 171.46 417.7 ;
     RECT  488.06 417.5 488.74 417.7 ;
     RECT  413.66 379.78 434.98 421.36 ;
     RECT  220.22 417.5 223.78 426.4 ;
     RECT  246.62 394.48 262.66 428.92 ;
     RECT  454.94 387.76 459.94 431.44 ;
     RECT  102.62 379.36 105.7 436.48 ;
     RECT  0.86 388.9 32.26 439 ;
     RECT  205.34 393.22 205.54 441.52 ;
     RECT  413.66 421.36 422.98 444.04 ;
     RECT  488.06 417.7 488.26 444.04 ;
     RECT  346.46 383.98 346.66 446.56 ;
     RECT  248.06 428.92 262.66 449.08 ;
     RECT  418.46 444.04 422.98 454.12 ;
     RECT  220.22 426.4 220.42 456.64 ;
     RECT  434.78 421.36 434.98 456.64 ;
     RECT  454.94 431.44 455.14 459.16 ;
     RECT  0.86 439 26.02 464.2 ;
     RECT  418.46 454.12 418.66 466.72 ;
     RECT  128.06 417.7 158.02 469.24 ;
     RECT  593.18 364.66 599.14 469.24 ;
     RECT  25.82 464.2 26.02 476.8 ;
     RECT  598.94 469.24 599.14 476.8 ;
     RECT  0.86 464.2 10.66 484.36 ;
     RECT  0.86 484.36 5.86 486.88 ;
     RECT  128.06 469.24 145.54 489.4 ;
     RECT  105.5 436.48 105.7 489.5 ;
     RECT  105.02 489.5 105.7 489.7 ;
     RECT  1.34 486.88 5.86 491.92 ;
     RECT  5.66 491.92 5.86 494.44 ;
     RECT  170.78 417.7 170.98 496.96 ;
     RECT  155.42 469.24 158.02 499.48 ;
     RECT  157.82 499.48 158.02 502 ;
     RECT  248.06 449.08 250.66 507.04 ;
     RECT  134.3 489.4 145.54 509.56 ;
     RECT  134.3 509.56 134.5 514.6 ;
     RECT  262.46 449.08 262.66 517.12 ;
     RECT  248.06 507.04 248.26 519.64 ;
     RECT  145.34 509.56 145.54 524.68 ;
     RECT  105.02 489.7 105.22 527.2 ;
    LAYER Metal4 ;
     RECT  0.38 225.02 0.86 225.22 ;
     RECT  0.38 293.06 0.86 293.26 ;
     RECT  0.38 322.88 0.86 323.92 ;
     RECT  0.38 255.68 1.34 255.88 ;
     RECT  0.86 293.06 1.34 296.2 ;
     RECT  1.34 284.66 1.82 296.2 ;
     RECT  1.34 305.24 1.82 305.44 ;
     RECT  1.34 433.76 2.02 433.96 ;
     RECT  0.86 218.3 2.3 225.22 ;
     RECT  1.82 274.16 2.3 274.36 ;
     RECT  0.86 65.84 3.26 66.04 ;
     RECT  1.34 255.68 4.22 262.6 ;
     RECT  2.3 274.16 4.22 274.78 ;
     RECT  3.26 202.34 5.66 202.54 ;
     RECT  0.86 322.88 5.66 328.12 ;
     RECT  3.26 60.8 7.1 83.68 ;
     RECT  2.78 130.1 7.1 130.3 ;
     RECT  3.74 172.52 7.1 172.72 ;
     RECT  5.66 197.3 7.1 202.54 ;
     RECT  2.3 218.3 7.1 232.36 ;
     RECT  4.22 255.68 7.1 274.78 ;
     RECT  1.82 284.66 7.1 305.44 ;
     RECT  5.66 316.16 7.1 328.12 ;
     RECT  3.26 373.28 7.1 373.48 ;
     RECT  7.1 60.8 14.3 101.32 ;
     RECT  7.1 350.6 22.94 350.8 ;
     RECT  7.1 186.8 23.42 232.36 ;
     RECT  7.1 242.24 23.42 328.12 ;
     RECT  22.94 350.6 24.86 353.74 ;
     RECT  7.1 365.72 24.86 373.48 ;
     RECT  23.42 186.8 28.22 328.12 ;
     RECT  7.1 340.94 36.86 341.14 ;
     RECT  24.86 350.6 36.86 373.48 ;
     RECT  7.1 149 37.34 172.72 ;
     RECT  28.22 186.8 37.34 329.8 ;
     RECT  14.3 60.8 40.22 102.16 ;
     RECT  7.1 111.2 40.22 118.96 ;
     RECT  37.34 149 43.1 329.8 ;
     RECT  36.86 340.94 43.1 373.48 ;
     RECT  40.22 60.8 56.06 118.96 ;
     RECT  7.1 130.1 57.5 139.12 ;
     RECT  43.1 149 57.5 373.48 ;
     RECT  56.06 60.8 61.82 119.38 ;
     RECT  57.5 130.1 61.82 373.48 ;
     RECT  61.82 60.8 87.26 373.48 ;
     RECT  87.26 60.8 96.38 376.42 ;
     RECT  96.38 60.8 129.5 378.52 ;
     RECT  129.5 60.8 148.22 379.36 ;
     RECT  148.22 60.8 161.18 380.2 ;
     RECT  161.18 58.28 176.06 380.2 ;
     RECT  176.06 54.92 181.34 380.2 ;
     RECT  181.34 54.5 183.46 380.2 ;
     RECT  3.26 45.68 186.82 45.88 ;
     RECT  183.46 54.92 197.86 380.2 ;
     RECT  197.86 59.54 209.66 380.2 ;
     RECT  209.66 59.54 215.9 387.76 ;
     RECT  215.9 58.28 216.1 387.76 ;
     RECT  216.1 58.7 225.98 387.76 ;
     RECT  225.98 50.72 231.94 387.76 ;
     RECT  231.94 50.72 237.7 111.82 ;
     RECT  237.7 58.7 240.38 111.82 ;
     RECT  231.94 121.7 240.38 387.76 ;
     RECT  240.38 58.7 245.38 387.76 ;
     RECT  245.38 119.18 246.34 387.76 ;
     RECT  245.38 58.7 248.74 105.1 ;
     RECT  246.34 119.18 248.74 380.2 ;
     RECT  248.74 122.54 254.98 380.2 ;
     RECT  3.26 511.88 256.9 512.08 ;
     RECT  248.74 59.12 258.34 105.1 ;
     RECT  258.34 66.68 261.7 105.1 ;
     RECT  254.98 122.54 263.62 129.04 ;
     RECT  261.7 84.32 264.1 105.1 ;
     RECT  258.62 54.92 267.94 55.12 ;
     RECT  254.98 137.66 268.22 380.2 ;
     RECT  268.22 137.66 268.42 387.76 ;
     RECT  261.7 66.68 269.38 70.24 ;
     RECT  269.38 68.36 271.3 70.24 ;
     RECT  268.42 137.66 272.26 223.96 ;
     RECT  264.1 85.16 273.7 105.1 ;
     RECT  268.42 232.58 273.98 387.76 ;
     RECT  273.7 85.16 278.78 99.22 ;
     RECT  273.98 232.58 279.46 391.54 ;
     RECT  272.26 137.66 280.7 223.12 ;
     RECT  279.46 232.58 280.7 380.2 ;
     RECT  278.78 84.74 286.18 99.22 ;
     RECT  284.06 113.3 287.62 114.34 ;
     RECT  280.7 137.66 288.1 380.2 ;
     RECT  263.62 122.96 290.98 129.04 ;
     RECT  286.18 85.16 291.94 99.22 ;
     RECT  279.46 391.34 291.94 391.54 ;
     RECT  290.98 122.96 292.22 126.52 ;
     RECT  292.22 119.6 292.42 126.52 ;
     RECT  271.3 68.36 292.9 68.56 ;
     RECT  292.42 119.6 294.82 119.8 ;
     RECT  291.94 85.16 295.3 92.5 ;
     RECT  295.3 91.88 296.26 92.5 ;
     RECT  288.1 137.66 296.54 223.96 ;
     RECT  288.1 232.58 296.54 380.2 ;
     RECT  296.54 137.66 302.3 380.2 ;
     RECT  302.3 137.66 318.82 386.08 ;
     RECT  318.82 137.66 322.66 383.98 ;
     RECT  322.66 137.66 341.86 380.62 ;
     RECT  341.86 137.66 350.98 380.2 ;
     RECT  350.98 137.66 351.46 221.86 ;
     RECT  351.46 137.66 352.9 216.82 ;
     RECT  350.98 232.16 352.9 380.2 ;
     RECT  352.9 137.66 354.14 161.38 ;
     RECT  354.14 133.88 363.46 161.38 ;
     RECT  363.46 137.66 366.34 161.38 ;
     RECT  366.34 154.46 379.58 161.38 ;
     RECT  352.9 170.42 379.58 216.82 ;
     RECT  352.9 232.16 380.26 379.78 ;
     RECT  379.58 154.46 381.22 221.44 ;
     RECT  381.22 170.42 381.7 221.44 ;
     RECT  381.7 187.22 382.18 221.44 ;
     RECT  366.34 137.66 384.1 143.74 ;
     RECT  381.22 154.46 388.9 161.38 ;
     RECT  381.7 170.42 388.9 176.08 ;
     RECT  382.18 187.22 389.86 197.08 ;
     RECT  388.9 175.88 392.74 176.08 ;
     RECT  389.86 192.26 395.9 197.08 ;
     RECT  382.18 206.96 396.1 221.44 ;
     RECT  396.1 221.24 397.06 221.44 ;
     RECT  396.1 206.96 398.02 212.2 ;
     RECT  380.26 236.36 399.94 379.78 ;
     RECT  395.9 192.26 402.34 198.34 ;
     RECT  402.34 192.26 403.1 194.56 ;
     RECT  398.02 209.06 403.3 212.2 ;
     RECT  403.1 186.8 403.58 194.56 ;
     RECT  403.58 183.44 403.78 194.56 ;
     RECT  399.94 238.88 404.74 379.78 ;
     RECT  403.78 183.44 406.18 187.42 ;
     RECT  404.74 238.88 408.58 377.26 ;
     RECT  384.1 140.18 409.34 143.74 ;
     RECT  408.58 239.3 409.54 377.26 ;
     RECT  409.34 140.18 409.82 145.84 ;
     RECT  409.54 239.3 412.42 376.84 ;
     RECT  409.82 140.18 413.38 147.1 ;
     RECT  403.3 209.48 413.66 212.2 ;
     RECT  412.42 244.34 414.34 376.84 ;
     RECT  388.9 161.18 414.62 161.38 ;
     RECT  414.62 157.4 415.1 161.38 ;
     RECT  406.18 183.44 416.06 183.64 ;
     RECT  415.1 157.4 416.54 167.68 ;
     RECT  416.06 183.44 417.02 191.62 ;
     RECT  413.38 140.18 417.98 145.84 ;
     RECT  416.54 157.4 420.86 173.98 ;
     RECT  417.02 183.44 420.86 194.56 ;
     RECT  420.86 157.4 421.34 194.56 ;
     RECT  421.34 157.4 421.82 195.82 ;
     RECT  413.66 209.48 421.82 213.04 ;
     RECT  414.34 244.34 423.26 376.42 ;
     RECT  417.98 138.92 423.74 145.84 ;
     RECT  421.82 157.4 423.74 213.04 ;
     RECT  423.26 242.24 428.06 376.42 ;
     RECT  423.74 138.92 429.02 213.46 ;
     RECT  428.06 235.94 431.14 376.42 ;
     RECT  431.14 239.3 434.5 376.42 ;
     RECT  434.5 269.54 435.94 376.42 ;
     RECT  434.5 239.3 438.82 260.5 ;
     RECT  429.02 138.92 450.14 217.24 ;
     RECT  438.82 252.32 453.7 260.5 ;
     RECT  435.94 271.64 455.42 376.42 ;
     RECT  455.42 269.54 456.58 376.42 ;
     RECT  450.14 138.92 457.54 218.08 ;
     RECT  457.54 138.92 466.46 217.24 ;
     RECT  453.7 252.32 468.38 258.82 ;
     RECT  456.58 273.32 468.38 376.42 ;
     RECT  468.38 252.32 470.98 376.42 ;
     RECT  470.98 269.96 471.46 376.42 ;
     RECT  466.46 136.4 474.34 217.24 ;
     RECT  471.46 269.96 475.3 292.84 ;
     RECT  474.34 194.36 476.26 217.24 ;
     RECT  476.26 194.36 476.74 202.12 ;
     RECT  470.98 252.32 489.22 258.82 ;
     RECT  475.3 273.32 489.22 292.84 ;
     RECT  489.22 273.32 492.1 292.42 ;
     RECT  492.1 273.74 497.66 292.42 ;
     RECT  471.46 304.82 497.66 376.42 ;
     RECT  497.66 273.74 501.22 376.42 ;
     RECT  489.22 252.32 505.82 256.3 ;
     RECT  501.22 273.74 506.5 298.72 ;
     RECT  506.5 273.74 506.98 292.42 ;
     RECT  476.74 194.36 518.3 195.82 ;
     RECT  501.22 308.18 529.06 376.42 ;
     RECT  529.06 319.1 536.26 376.42 ;
     RECT  476.26 212 543.46 217.24 ;
     RECT  505.82 252.32 554.5 262.6 ;
     RECT  474.34 136.4 590.5 184.48 ;
     RECT  518.3 194.36 590.5 197.08 ;
     RECT  543.46 212 590.5 212.2 ;
     RECT  438.82 239.3 590.5 242.44 ;
     RECT  554.5 252.32 590.5 256.3 ;
     RECT  506.98 273.74 590.5 291.58 ;
     RECT  536.26 319.1 590.5 334.42 ;
     RECT  419.42 433.76 590.5 433.96 ;
     RECT  590.5 319.1 590.98 319.72 ;
     RECT  536.26 345.56 592.7 376.42 ;
     RECT  592.7 344.3 592.9 376.42 ;
     RECT  590.5 149.84 593.38 157.6 ;
     RECT  592.9 370.76 593.86 376.42 ;
     RECT  590.5 285.5 594.34 291.58 ;
     RECT  593.38 150.68 594.82 157.6 ;
     RECT  590.5 329.6 594.82 334.42 ;
     RECT  590.5 273.74 595.3 273.94 ;
     RECT  592.9 344.3 595.3 360.04 ;
     RECT  593.86 375.38 595.3 376.42 ;
     RECT  529.06 308.18 595.78 308.38 ;
     RECT  590.5 239.3 596.26 239.5 ;
     RECT  594.82 330.44 596.26 334.42 ;
     RECT  595.3 359.84 596.26 360.04 ;
     RECT  590.98 319.1 596.74 319.3 ;
     RECT  594.34 287.6 597.22 291.58 ;
     RECT  596.26 334.22 597.22 334.42 ;
     RECT  597.22 287.6 597.7 287.8 ;
     RECT  590.5 255.68 598.18 256.3 ;
     RECT  594.82 157.4 598.66 157.6 ;
     RECT  595.3 376.22 598.66 376.42 ;
     RECT  595.3 344.3 598.94 346.18 ;
     RECT  590.5 167.48 599.14 167.68 ;
     RECT  598.18 256.1 599.14 256.3 ;
     RECT  598.94 343.88 599.14 346.18 ;
    LAYER Metal5 ;
     RECT  210.62 72.98 210.82 80.96 ;
     RECT  252.86 78.44 253.06 98.6 ;
     RECT  252.86 98.6 253.54 100.06 ;
     RECT  252.86 100.06 253.06 100.48 ;
     RECT  186.62 45.68 186.82 100.7 ;
     RECT  143.42 109.1 143.62 114.76 ;
     RECT  254.78 125.9 254.98 130.1 ;
     RECT  466.46 136.4 466.66 142.7 ;
     RECT  252.38 130.1 254.98 146.48 ;
     RECT  197.66 93.56 197.86 149 ;
     RECT  210.62 80.96 214.66 149 ;
     RECT  453.02 149 454.18 149.76 ;
     RECT  134.78 137.66 134.98 151.1 ;
     RECT  180.86 100.7 186.82 151.1 ;
     RECT  197.66 149 214.66 151.1 ;
     RECT  465.02 142.7 466.66 152.14 ;
     RECT  180.86 151.1 214.66 152.36 ;
     RECT  252.38 146.48 255.46 152.56 ;
     RECT  425.66 152.36 425.86 153.62 ;
     RECT  134.78 151.1 139.78 154.46 ;
     RECT  465.02 152.14 465.22 154.46 ;
     RECT  134.78 154.46 147.46 156.56 ;
     RECT  252.38 152.56 254.98 159.28 ;
     RECT  177.5 152.36 214.66 160.34 ;
     RECT  327.26 156.98 327.46 164.12 ;
     RECT  425.66 153.62 432.1 164.96 ;
     RECT  463.1 154.46 465.22 164.96 ;
     RECT  425.18 164.96 432.1 165.38 ;
     RECT  442.46 160.34 442.66 165.38 ;
     RECT  134.78 156.56 158.02 166.42 ;
     RECT  147.26 166.42 156.1 167.26 ;
     RECT  460.7 164.96 465.22 167.26 ;
     RECT  327.26 164.12 331.3 167.48 ;
     RECT  460.7 167.26 463.3 167.9 ;
     RECT  59.9 151.1 60.1 168.32 ;
     RECT  229.34 133.88 229.54 168.32 ;
     RECT  425.18 165.38 442.66 168.32 ;
     RECT  453.02 167.9 463.3 168.32 ;
     RECT  252.38 159.28 252.58 168.52 ;
     RECT  226.46 168.32 229.54 169.16 ;
     RECT  226.46 169.16 233.38 170.84 ;
     RECT  59.9 168.32 69.22 172.3 ;
     RECT  102.14 152.78 102.34 173.56 ;
     RECT  425.18 168.32 463.3 173.56 ;
     RECT  431.9 173.56 463.3 175.24 ;
     RECT  147.26 167.26 147.46 175.66 ;
     RECT  325.82 167.48 331.3 176.72 ;
     RECT  170.3 160.34 214.66 177.34 ;
     RECT  226.46 170.84 237.22 179.24 ;
     RECT  197.66 177.34 214.66 179.66 ;
     RECT  325.34 176.72 331.3 181.76 ;
     RECT  302.78 154.46 302.98 182.18 ;
     RECT  134.78 166.42 134.98 183.02 ;
     RECT  170.3 177.34 186.82 183.22 ;
     RECT  431.9 175.24 460.9 183.22 ;
     RECT  442.46 183.22 460.9 184.06 ;
     RECT  270.62 152.78 270.82 184.28 ;
     RECT  325.34 181.76 338.02 185.32 ;
     RECT  295.58 182.18 302.98 186.16 ;
     RECT  445.82 184.06 460.9 187 ;
     RECT  182.78 183.22 186.82 187.22 ;
     RECT  197.66 179.66 215.14 187.22 ;
     RECT  297.98 186.16 302.98 188.26 ;
     RECT  431.9 183.22 432.1 189.74 ;
     RECT  426.14 189.74 432.1 190.16 ;
     RECT  327.26 185.32 338.02 191.62 ;
     RECT  269.66 184.28 270.82 192.04 ;
     RECT  327.26 191.62 331.3 192.04 ;
     RECT  328.22 192.04 331.3 192.88 ;
     RECT  170.3 183.22 170.5 193.72 ;
     RECT  472.7 193.94 472.9 196.04 ;
     RECT  445.82 187 453.22 197.08 ;
     RECT  470.78 196.04 472.9 200.02 ;
     RECT  298.94 188.26 302.98 200.44 ;
     RECT  445.82 197.08 446.02 200.86 ;
     RECT  134.78 183.02 138.34 201.5 ;
     RECT  163.1 195.62 163.3 201.5 ;
     RECT  182.78 187.22 215.14 201.5 ;
     RECT  225.5 179.24 237.22 201.5 ;
     RECT  256.7 194.78 256.9 201.5 ;
     RECT  328.22 192.88 329.86 201.7 ;
     RECT  419.42 190.16 432.1 201.7 ;
     RECT  69.02 172.3 69.22 202.34 ;
     RECT  134.78 201.5 147.94 202.34 ;
     RECT  470.78 200.02 470.98 202.54 ;
     RECT  116.06 100.28 116.26 205.28 ;
     RECT  127.1 202.34 147.94 205.28 ;
     RECT  419.42 201.7 426.34 205.9 ;
     RECT  159.26 201.5 163.3 208.22 ;
     RECT  159.26 208.22 166.66 208.64 ;
     RECT  179.9 201.5 237.22 208.64 ;
     RECT  66.14 202.34 69.22 209.9 ;
     RECT  159.26 208.64 237.22 216.2 ;
     RECT  159.26 216.2 237.7 216.82 ;
     RECT  116.06 205.28 147.94 217.24 ;
     RECT  298.94 200.44 299.14 217.24 ;
     RECT  256.7 201.5 257.38 217.88 ;
     RECT  161.18 216.82 237.7 228.58 ;
     RECT  161.18 228.58 186.34 230.48 ;
     RECT  197.66 228.58 237.7 232.36 ;
     RECT  254.78 217.88 257.38 233.62 ;
     RECT  160.22 230.48 186.34 236.14 ;
     RECT  161.18 236.14 186.34 236.98 ;
     RECT  130.94 217.24 147.94 237.82 ;
     RECT  254.78 233.62 256.9 238.24 ;
     RECT  167.42 236.98 186.34 239.72 ;
     RECT  197.66 232.36 229.54 239.72 ;
     RECT  116.06 217.24 118.18 241.18 ;
     RECT  134.78 237.82 147.94 241.18 ;
     RECT  256.7 238.24 256.9 243.5 ;
     RECT  269.66 192.04 269.86 243.5 ;
     RECT  256.7 243.5 269.86 247.06 ;
     RECT  146.78 241.18 146.98 247.48 ;
     RECT  167.42 239.72 229.54 252.1 ;
     RECT  192.38 252.1 229.54 254 ;
     RECT  256.7 247.06 260.26 258.62 ;
     RECT  167.42 252.1 180.1 258.82 ;
     RECT  167.42 258.82 179.62 259.24 ;
     RECT  419.42 205.9 419.62 260.3 ;
     RECT  0.86 218.3 1.06 262.4 ;
     RECT  192.38 254 236.74 265.96 ;
     RECT  192.38 265.96 229.54 266.38 ;
     RECT  192.38 266.38 229.06 269.12 ;
     RECT  101.66 256.94 101.86 277.3 ;
     RECT  419.42 260.3 427.3 279.62 ;
     RECT  279.26 272.06 279.46 279.82 ;
     RECT  253.34 258.62 260.26 286.76 ;
     RECT  134.78 241.18 134.98 288.64 ;
     RECT  186.62 269.12 229.06 289.06 ;
     RECT  196.22 289.06 229.06 292 ;
     RECT  417.98 279.62 427.3 292 ;
     RECT  253.34 286.76 262.18 293.06 ;
     RECT  417.98 292 424.9 293.68 ;
     RECT  196.22 292 227.14 300.4 ;
     RECT  167.42 259.24 175.78 300.82 ;
     RECT  66.14 209.9 71.14 301.24 ;
     RECT  32.06 272.9 32.26 302.08 ;
     RECT  81.98 251.9 82.18 302.08 ;
     RECT  243.26 293.48 243.46 302.3 ;
     RECT  253.34 293.06 264.1 302.3 ;
     RECT  167.42 300.82 167.62 308.38 ;
     RECT  199.1 300.4 227.14 308.38 ;
     RECT  203.9 308.38 227.14 309.22 ;
     RECT  204.38 309.22 227.14 315.52 ;
     RECT  243.26 302.3 264.1 316.36 ;
     RECT  419.42 293.68 424.9 316.78 ;
     RECT  66.14 301.24 70.18 322.66 ;
     RECT  251.9 316.36 264.1 324.34 ;
     RECT  210.14 315.52 227.14 326.02 ;
     RECT  210.62 326.02 227.14 326.44 ;
     RECT  256.7 324.34 264.1 326.86 ;
     RECT  256.7 326.86 261.22 327.28 ;
     RECT  256.7 327.28 260.26 335.68 ;
     RECT  69.02 322.66 70.18 338.62 ;
     RECT  0.86 262.4 1.54 340.94 ;
     RECT  210.62 326.44 215.62 345.76 ;
     RECT  69.98 338.62 70.18 346.18 ;
     RECT  215.42 345.76 215.62 353.12 ;
     RECT  226.94 326.44 227.14 353.12 ;
     RECT  215.42 353.12 227.14 357.1 ;
     RECT  215.42 357.1 221.38 360.46 ;
     RECT  116.06 241.18 116.26 365.92 ;
     RECT  215.42 360.46 215.62 374.32 ;
     RECT  0.86 340.94 7.3 378.52 ;
     RECT  0.86 378.52 1.54 383.56 ;
     RECT  1.34 383.56 1.54 433.96 ;
     RECT  419.42 316.78 419.62 433.96 ;
     RECT  256.7 335.68 256.9 512.08 ;
  END
END dm_top
END LIBRARY
