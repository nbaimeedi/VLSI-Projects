VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO cve2_core
  FOREIGN cve2_core 0 0 ;
  CLASS BLOCK ;
  SIZE 815 BY 895.12 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN VDDIO
    USE POWER ;
    DIRECTION INOUT ;
  END VDDIO
  PIN VSSIO
    USE GROUND ;
    DIRECTION INOUT ;
  END VSSIO
  PIN crash_dump_o_64_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 17.96 815 18.16 ;
    END
  END crash_dump_o_64_
  PIN data_addr_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 20.48 815 20.68 ;
    END
  END data_addr_o_0_
  PIN data_addr_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 23 815 23.2 ;
    END
  END data_addr_o_1_
  PIN instr_addr_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 25.52 815 25.72 ;
    END
  END instr_addr_o_0_
  PIN instr_addr_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 28.04 815 28.24 ;
    END
  END instr_addr_o_1_
  PIN boot_addr_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 894.92 0.72 895.12 ;
    END
  END boot_addr_i_0_
  PIN boot_addr_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 768.92 0.72 769.12 ;
    END
  END boot_addr_i_10_
  PIN boot_addr_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 456.44 0.72 456.64 ;
    END
  END boot_addr_i_11_
  PIN boot_addr_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 458.96 0.72 459.16 ;
    END
  END boot_addr_i_12_
  PIN boot_addr_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 461.48 0.72 461.68 ;
    END
  END boot_addr_i_13_
  PIN boot_addr_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 464 0.72 464.2 ;
    END
  END boot_addr_i_14_
  PIN boot_addr_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 453.92 0.72 454.12 ;
    END
  END boot_addr_i_15_
  PIN boot_addr_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 466.52 0.72 466.72 ;
    END
  END boot_addr_i_16_
  PIN boot_addr_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 469.04 0.72 469.24 ;
    END
  END boot_addr_i_17_
  PIN boot_addr_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 471.56 0.72 471.76 ;
    END
  END boot_addr_i_18_
  PIN boot_addr_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 451.4 0.72 451.6 ;
    END
  END boot_addr_i_19_
  PIN boot_addr_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 892.4 0.72 892.6 ;
    END
  END boot_addr_i_1_
  PIN boot_addr_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 474.08 0.72 474.28 ;
    END
  END boot_addr_i_20_
  PIN boot_addr_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 476.6 0.72 476.8 ;
    END
  END boot_addr_i_21_
  PIN boot_addr_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 479.12 0.72 479.32 ;
    END
  END boot_addr_i_22_
  PIN boot_addr_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 448.88 0.72 449.08 ;
    END
  END boot_addr_i_23_
  PIN boot_addr_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 481.64 0.72 481.84 ;
    END
  END boot_addr_i_24_
  PIN boot_addr_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 484.16 0.72 484.36 ;
    END
  END boot_addr_i_25_
  PIN boot_addr_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 486.68 0.72 486.88 ;
    END
  END boot_addr_i_26_
  PIN boot_addr_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 446.36 0.72 446.56 ;
    END
  END boot_addr_i_27_
  PIN boot_addr_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 489.2 0.72 489.4 ;
    END
  END boot_addr_i_28_
  PIN boot_addr_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 491.72 0.72 491.92 ;
    END
  END boot_addr_i_29_
  PIN boot_addr_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 889.88 0.72 890.08 ;
    END
  END boot_addr_i_2_
  PIN boot_addr_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 494.24 0.72 494.44 ;
    END
  END boot_addr_i_30_
  PIN boot_addr_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 443.84 0.72 444.04 ;
    END
  END boot_addr_i_31_
  PIN boot_addr_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 887.36 0.72 887.56 ;
    END
  END boot_addr_i_3_
  PIN boot_addr_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 884.84 0.72 885.04 ;
    END
  END boot_addr_i_4_
  PIN boot_addr_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 882.32 0.72 882.52 ;
    END
  END boot_addr_i_5_
  PIN boot_addr_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 879.8 0.72 880 ;
    END
  END boot_addr_i_6_
  PIN boot_addr_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 877.28 0.72 877.48 ;
    END
  END boot_addr_i_7_
  PIN boot_addr_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 496.76 0.72 496.96 ;
    END
  END boot_addr_i_8_
  PIN boot_addr_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 499.28 0.72 499.48 ;
    END
  END boot_addr_i_9_
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 501.8 0.72 502 ;
    END
  END clk_i
  PIN core_busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 30.56 815 30.76 ;
    END
  END core_busy_o
  PIN crash_dump_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 33.08 815 33.28 ;
    END
  END crash_dump_o_0_
  PIN crash_dump_o_100_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 35.6 815 35.8 ;
    END
  END crash_dump_o_100_
  PIN crash_dump_o_101_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 38.12 815 38.32 ;
    END
  END crash_dump_o_101_
  PIN crash_dump_o_102_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 40.64 815 40.84 ;
    END
  END crash_dump_o_102_
  PIN crash_dump_o_103_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 43.16 815 43.36 ;
    END
  END crash_dump_o_103_
  PIN crash_dump_o_104_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 45.68 815 45.88 ;
    END
  END crash_dump_o_104_
  PIN crash_dump_o_105_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 48.2 815 48.4 ;
    END
  END crash_dump_o_105_
  PIN crash_dump_o_106_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 50.72 815 50.92 ;
    END
  END crash_dump_o_106_
  PIN crash_dump_o_107_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 53.24 815 53.44 ;
    END
  END crash_dump_o_107_
  PIN crash_dump_o_108_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 55.76 815 55.96 ;
    END
  END crash_dump_o_108_
  PIN crash_dump_o_109_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 58.28 815 58.48 ;
    END
  END crash_dump_o_109_
  PIN crash_dump_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 60.8 815 61 ;
    END
  END crash_dump_o_10_
  PIN crash_dump_o_110_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 63.32 815 63.52 ;
    END
  END crash_dump_o_110_
  PIN crash_dump_o_111_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 65.84 815 66.04 ;
    END
  END crash_dump_o_111_
  PIN crash_dump_o_112_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 68.36 815 68.56 ;
    END
  END crash_dump_o_112_
  PIN crash_dump_o_113_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 70.88 815 71.08 ;
    END
  END crash_dump_o_113_
  PIN crash_dump_o_114_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 73.4 815 73.6 ;
    END
  END crash_dump_o_114_
  PIN crash_dump_o_115_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 75.92 815 76.12 ;
    END
  END crash_dump_o_115_
  PIN crash_dump_o_116_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 78.44 815 78.64 ;
    END
  END crash_dump_o_116_
  PIN crash_dump_o_117_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 80.96 815 81.16 ;
    END
  END crash_dump_o_117_
  PIN crash_dump_o_118_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 83.48 815 83.68 ;
    END
  END crash_dump_o_118_
  PIN crash_dump_o_119_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 86 815 86.2 ;
    END
  END crash_dump_o_119_
  PIN crash_dump_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 88.52 815 88.72 ;
    END
  END crash_dump_o_11_
  PIN crash_dump_o_120_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 91.04 815 91.24 ;
    END
  END crash_dump_o_120_
  PIN crash_dump_o_121_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 93.56 815 93.76 ;
    END
  END crash_dump_o_121_
  PIN crash_dump_o_122_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 96.08 815 96.28 ;
    END
  END crash_dump_o_122_
  PIN crash_dump_o_123_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 98.6 815 98.8 ;
    END
  END crash_dump_o_123_
  PIN crash_dump_o_124_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 101.12 815 101.32 ;
    END
  END crash_dump_o_124_
  PIN crash_dump_o_125_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 103.64 815 103.84 ;
    END
  END crash_dump_o_125_
  PIN crash_dump_o_126_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 106.16 815 106.36 ;
    END
  END crash_dump_o_126_
  PIN crash_dump_o_127_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 108.68 815 108.88 ;
    END
  END crash_dump_o_127_
  PIN crash_dump_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 111.2 815 111.4 ;
    END
  END crash_dump_o_12_
  PIN crash_dump_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 113.72 815 113.92 ;
    END
  END crash_dump_o_13_
  PIN crash_dump_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 116.24 815 116.44 ;
    END
  END crash_dump_o_14_
  PIN crash_dump_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 118.76 815 118.96 ;
    END
  END crash_dump_o_15_
  PIN crash_dump_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 121.28 815 121.48 ;
    END
  END crash_dump_o_16_
  PIN crash_dump_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 123.8 815 124 ;
    END
  END crash_dump_o_17_
  PIN crash_dump_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 126.32 815 126.52 ;
    END
  END crash_dump_o_18_
  PIN crash_dump_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 128.84 815 129.04 ;
    END
  END crash_dump_o_19_
  PIN crash_dump_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 131.36 815 131.56 ;
    END
  END crash_dump_o_1_
  PIN crash_dump_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 133.88 815 134.08 ;
    END
  END crash_dump_o_20_
  PIN crash_dump_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 136.4 815 136.6 ;
    END
  END crash_dump_o_21_
  PIN crash_dump_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 138.92 815 139.12 ;
    END
  END crash_dump_o_22_
  PIN crash_dump_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 141.44 815 141.64 ;
    END
  END crash_dump_o_23_
  PIN crash_dump_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 143.96 815 144.16 ;
    END
  END crash_dump_o_24_
  PIN crash_dump_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 146.48 815 146.68 ;
    END
  END crash_dump_o_25_
  PIN crash_dump_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 149 815 149.2 ;
    END
  END crash_dump_o_26_
  PIN crash_dump_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 151.52 815 151.72 ;
    END
  END crash_dump_o_27_
  PIN crash_dump_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 154.04 815 154.24 ;
    END
  END crash_dump_o_28_
  PIN crash_dump_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 156.56 815 156.76 ;
    END
  END crash_dump_o_29_
  PIN crash_dump_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 159.08 815 159.28 ;
    END
  END crash_dump_o_2_
  PIN crash_dump_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 161.6 815 161.8 ;
    END
  END crash_dump_o_30_
  PIN crash_dump_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 164.12 815 164.32 ;
    END
  END crash_dump_o_31_
  PIN crash_dump_o_32_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 166.64 815 166.84 ;
    END
  END crash_dump_o_32_
  PIN crash_dump_o_33_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 169.16 815 169.36 ;
    END
  END crash_dump_o_33_
  PIN crash_dump_o_34_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 171.68 815 171.88 ;
    END
  END crash_dump_o_34_
  PIN crash_dump_o_35_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 174.2 815 174.4 ;
    END
  END crash_dump_o_35_
  PIN crash_dump_o_36_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 176.72 815 176.92 ;
    END
  END crash_dump_o_36_
  PIN crash_dump_o_37_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 179.24 815 179.44 ;
    END
  END crash_dump_o_37_
  PIN crash_dump_o_38_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 181.76 815 181.96 ;
    END
  END crash_dump_o_38_
  PIN crash_dump_o_39_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 184.28 815 184.48 ;
    END
  END crash_dump_o_39_
  PIN crash_dump_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 186.8 815 187 ;
    END
  END crash_dump_o_3_
  PIN crash_dump_o_40_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 189.32 815 189.52 ;
    END
  END crash_dump_o_40_
  PIN crash_dump_o_41_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 191.84 815 192.04 ;
    END
  END crash_dump_o_41_
  PIN crash_dump_o_42_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 194.36 815 194.56 ;
    END
  END crash_dump_o_42_
  PIN crash_dump_o_43_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 196.88 815 197.08 ;
    END
  END crash_dump_o_43_
  PIN crash_dump_o_44_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 199.4 815 199.6 ;
    END
  END crash_dump_o_44_
  PIN crash_dump_o_45_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 201.92 815 202.12 ;
    END
  END crash_dump_o_45_
  PIN crash_dump_o_46_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 204.44 815 204.64 ;
    END
  END crash_dump_o_46_
  PIN crash_dump_o_47_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 206.96 815 207.16 ;
    END
  END crash_dump_o_47_
  PIN crash_dump_o_48_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 209.48 815 209.68 ;
    END
  END crash_dump_o_48_
  PIN crash_dump_o_49_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 212 815 212.2 ;
    END
  END crash_dump_o_49_
  PIN crash_dump_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 214.52 815 214.72 ;
    END
  END crash_dump_o_4_
  PIN crash_dump_o_50_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 217.04 815 217.24 ;
    END
  END crash_dump_o_50_
  PIN crash_dump_o_51_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 219.56 815 219.76 ;
    END
  END crash_dump_o_51_
  PIN crash_dump_o_52_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 222.08 815 222.28 ;
    END
  END crash_dump_o_52_
  PIN crash_dump_o_53_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 224.6 815 224.8 ;
    END
  END crash_dump_o_53_
  PIN crash_dump_o_54_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 227.12 815 227.32 ;
    END
  END crash_dump_o_54_
  PIN crash_dump_o_55_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 229.64 815 229.84 ;
    END
  END crash_dump_o_55_
  PIN crash_dump_o_56_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 232.16 815 232.36 ;
    END
  END crash_dump_o_56_
  PIN crash_dump_o_57_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 234.68 815 234.88 ;
    END
  END crash_dump_o_57_
  PIN crash_dump_o_58_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 237.2 815 237.4 ;
    END
  END crash_dump_o_58_
  PIN crash_dump_o_59_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 239.72 815 239.92 ;
    END
  END crash_dump_o_59_
  PIN crash_dump_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 242.24 815 242.44 ;
    END
  END crash_dump_o_5_
  PIN crash_dump_o_60_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 244.76 815 244.96 ;
    END
  END crash_dump_o_60_
  PIN crash_dump_o_61_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 247.28 815 247.48 ;
    END
  END crash_dump_o_61_
  PIN crash_dump_o_62_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 249.8 815 250 ;
    END
  END crash_dump_o_62_
  PIN crash_dump_o_63_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 252.32 815 252.52 ;
    END
  END crash_dump_o_63_
  PIN crash_dump_o_65_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 254.84 815 255.04 ;
    END
  END crash_dump_o_65_
  PIN crash_dump_o_66_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 257.36 815 257.56 ;
    END
  END crash_dump_o_66_
  PIN crash_dump_o_67_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 259.88 815 260.08 ;
    END
  END crash_dump_o_67_
  PIN crash_dump_o_68_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 262.4 815 262.6 ;
    END
  END crash_dump_o_68_
  PIN crash_dump_o_69_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 264.92 815 265.12 ;
    END
  END crash_dump_o_69_
  PIN crash_dump_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 267.44 815 267.64 ;
    END
  END crash_dump_o_6_
  PIN crash_dump_o_70_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 269.96 815 270.16 ;
    END
  END crash_dump_o_70_
  PIN crash_dump_o_71_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 272.48 815 272.68 ;
    END
  END crash_dump_o_71_
  PIN crash_dump_o_72_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 275 815 275.2 ;
    END
  END crash_dump_o_72_
  PIN crash_dump_o_73_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 277.52 815 277.72 ;
    END
  END crash_dump_o_73_
  PIN crash_dump_o_74_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 280.04 815 280.24 ;
    END
  END crash_dump_o_74_
  PIN crash_dump_o_75_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 282.56 815 282.76 ;
    END
  END crash_dump_o_75_
  PIN crash_dump_o_76_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 285.08 815 285.28 ;
    END
  END crash_dump_o_76_
  PIN crash_dump_o_77_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 287.6 815 287.8 ;
    END
  END crash_dump_o_77_
  PIN crash_dump_o_78_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 290.12 815 290.32 ;
    END
  END crash_dump_o_78_
  PIN crash_dump_o_79_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 292.64 815 292.84 ;
    END
  END crash_dump_o_79_
  PIN crash_dump_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 295.16 815 295.36 ;
    END
  END crash_dump_o_7_
  PIN crash_dump_o_80_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 297.68 815 297.88 ;
    END
  END crash_dump_o_80_
  PIN crash_dump_o_81_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 300.2 815 300.4 ;
    END
  END crash_dump_o_81_
  PIN crash_dump_o_82_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 302.72 815 302.92 ;
    END
  END crash_dump_o_82_
  PIN crash_dump_o_83_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 305.24 815 305.44 ;
    END
  END crash_dump_o_83_
  PIN crash_dump_o_84_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 307.76 815 307.96 ;
    END
  END crash_dump_o_84_
  PIN crash_dump_o_85_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 310.28 815 310.48 ;
    END
  END crash_dump_o_85_
  PIN crash_dump_o_86_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 312.8 815 313 ;
    END
  END crash_dump_o_86_
  PIN crash_dump_o_87_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 315.32 815 315.52 ;
    END
  END crash_dump_o_87_
  PIN crash_dump_o_88_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 317.84 815 318.04 ;
    END
  END crash_dump_o_88_
  PIN crash_dump_o_89_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 320.36 815 320.56 ;
    END
  END crash_dump_o_89_
  PIN crash_dump_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 322.88 815 323.08 ;
    END
  END crash_dump_o_8_
  PIN crash_dump_o_90_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 325.4 815 325.6 ;
    END
  END crash_dump_o_90_
  PIN crash_dump_o_91_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 327.92 815 328.12 ;
    END
  END crash_dump_o_91_
  PIN crash_dump_o_92_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 330.44 815 330.64 ;
    END
  END crash_dump_o_92_
  PIN crash_dump_o_93_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 332.96 815 333.16 ;
    END
  END crash_dump_o_93_
  PIN crash_dump_o_94_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 335.48 815 335.68 ;
    END
  END crash_dump_o_94_
  PIN crash_dump_o_95_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 338 815 338.2 ;
    END
  END crash_dump_o_95_
  PIN crash_dump_o_96_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 340.52 815 340.72 ;
    END
  END crash_dump_o_96_
  PIN crash_dump_o_97_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 343.04 815 343.24 ;
    END
  END crash_dump_o_97_
  PIN crash_dump_o_98_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 345.56 815 345.76 ;
    END
  END crash_dump_o_98_
  PIN crash_dump_o_99_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 348.08 815 348.28 ;
    END
  END crash_dump_o_99_
  PIN crash_dump_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 350.6 815 350.8 ;
    END
  END crash_dump_o_9_
  PIN data_addr_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 353.12 815 353.32 ;
    END
  END data_addr_o_10_
  PIN data_addr_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 355.64 815 355.84 ;
    END
  END data_addr_o_11_
  PIN data_addr_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 358.16 815 358.36 ;
    END
  END data_addr_o_12_
  PIN data_addr_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 360.68 815 360.88 ;
    END
  END data_addr_o_13_
  PIN data_addr_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 363.2 815 363.4 ;
    END
  END data_addr_o_14_
  PIN data_addr_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 365.72 815 365.92 ;
    END
  END data_addr_o_15_
  PIN data_addr_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 368.24 815 368.44 ;
    END
  END data_addr_o_16_
  PIN data_addr_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 370.76 815 370.96 ;
    END
  END data_addr_o_17_
  PIN data_addr_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 373.28 815 373.48 ;
    END
  END data_addr_o_18_
  PIN data_addr_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 375.8 815 376 ;
    END
  END data_addr_o_19_
  PIN data_addr_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 378.32 815 378.52 ;
    END
  END data_addr_o_20_
  PIN data_addr_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 380.84 815 381.04 ;
    END
  END data_addr_o_21_
  PIN data_addr_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 383.36 815 383.56 ;
    END
  END data_addr_o_22_
  PIN data_addr_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 385.88 815 386.08 ;
    END
  END data_addr_o_23_
  PIN data_addr_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 388.4 815 388.6 ;
    END
  END data_addr_o_24_
  PIN data_addr_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 390.92 815 391.12 ;
    END
  END data_addr_o_25_
  PIN data_addr_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 393.44 815 393.64 ;
    END
  END data_addr_o_26_
  PIN data_addr_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 395.96 815 396.16 ;
    END
  END data_addr_o_27_
  PIN data_addr_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 398.48 815 398.68 ;
    END
  END data_addr_o_28_
  PIN data_addr_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 401 815 401.2 ;
    END
  END data_addr_o_29_
  PIN data_addr_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 403.52 815 403.72 ;
    END
  END data_addr_o_2_
  PIN data_addr_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 406.04 815 406.24 ;
    END
  END data_addr_o_30_
  PIN data_addr_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 408.56 815 408.76 ;
    END
  END data_addr_o_31_
  PIN data_addr_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 411.08 815 411.28 ;
    END
  END data_addr_o_3_
  PIN data_addr_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 413.6 815 413.8 ;
    END
  END data_addr_o_4_
  PIN data_addr_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 416.12 815 416.32 ;
    END
  END data_addr_o_5_
  PIN data_addr_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 418.64 815 418.84 ;
    END
  END data_addr_o_6_
  PIN data_addr_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 421.16 815 421.36 ;
    END
  END data_addr_o_7_
  PIN data_addr_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 423.68 815 423.88 ;
    END
  END data_addr_o_8_
  PIN data_addr_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 426.2 815 426.4 ;
    END
  END data_addr_o_9_
  PIN data_be_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 428.72 815 428.92 ;
    END
  END data_be_o_0_
  PIN data_be_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 431.24 815 431.44 ;
    END
  END data_be_o_1_
  PIN data_be_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 433.76 815 433.96 ;
    END
  END data_be_o_2_
  PIN data_be_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 436.28 815 436.48 ;
    END
  END data_be_o_3_
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 441.32 0.72 441.52 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 504.32 0.72 504.52 ;
    END
  END data_gnt_i
  PIN data_rdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 506.84 0.72 507.04 ;
    END
  END data_rdata_i_0_
  PIN data_rdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 509.36 0.72 509.56 ;
    END
  END data_rdata_i_10_
  PIN data_rdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 438.8 0.72 439 ;
    END
  END data_rdata_i_11_
  PIN data_rdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 511.88 0.72 512.08 ;
    END
  END data_rdata_i_12_
  PIN data_rdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 514.4 0.72 514.6 ;
    END
  END data_rdata_i_13_
  PIN data_rdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 516.92 0.72 517.12 ;
    END
  END data_rdata_i_14_
  PIN data_rdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 436.28 0.72 436.48 ;
    END
  END data_rdata_i_15_
  PIN data_rdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 519.44 0.72 519.64 ;
    END
  END data_rdata_i_16_
  PIN data_rdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 521.96 0.72 522.16 ;
    END
  END data_rdata_i_17_
  PIN data_rdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 524.48 0.72 524.68 ;
    END
  END data_rdata_i_18_
  PIN data_rdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 433.76 0.72 433.96 ;
    END
  END data_rdata_i_19_
  PIN data_rdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 527 0.72 527.2 ;
    END
  END data_rdata_i_1_
  PIN data_rdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 529.52 0.72 529.72 ;
    END
  END data_rdata_i_20_
  PIN data_rdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 532.04 0.72 532.24 ;
    END
  END data_rdata_i_21_
  PIN data_rdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 431.24 0.72 431.44 ;
    END
  END data_rdata_i_22_
  PIN data_rdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 534.56 0.72 534.76 ;
    END
  END data_rdata_i_23_
  PIN data_rdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 537.08 0.72 537.28 ;
    END
  END data_rdata_i_24_
  PIN data_rdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 539.6 0.72 539.8 ;
    END
  END data_rdata_i_25_
  PIN data_rdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 428.72 0.72 428.92 ;
    END
  END data_rdata_i_26_
  PIN data_rdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 542.12 0.72 542.32 ;
    END
  END data_rdata_i_27_
  PIN data_rdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 544.64 0.72 544.84 ;
    END
  END data_rdata_i_28_
  PIN data_rdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 547.16 0.72 547.36 ;
    END
  END data_rdata_i_29_
  PIN data_rdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 426.2 0.72 426.4 ;
    END
  END data_rdata_i_2_
  PIN data_rdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 549.68 0.72 549.88 ;
    END
  END data_rdata_i_30_
  PIN data_rdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 552.2 0.72 552.4 ;
    END
  END data_rdata_i_31_
  PIN data_rdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 554.72 0.72 554.92 ;
    END
  END data_rdata_i_3_
  PIN data_rdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 423.68 0.72 423.88 ;
    END
  END data_rdata_i_4_
  PIN data_rdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 557.24 0.72 557.44 ;
    END
  END data_rdata_i_5_
  PIN data_rdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 559.76 0.72 559.96 ;
    END
  END data_rdata_i_6_
  PIN data_rdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 562.28 0.72 562.48 ;
    END
  END data_rdata_i_7_
  PIN data_rdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 421.16 0.72 421.36 ;
    END
  END data_rdata_i_8_
  PIN data_rdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 564.8 0.72 565 ;
    END
  END data_rdata_i_9_
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 438.8 815 439 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 567.32 0.72 567.52 ;
    END
  END data_rvalid_i
  PIN data_wdata_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 441.32 815 441.52 ;
    END
  END data_wdata_o_0_
  PIN data_wdata_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 443.84 815 444.04 ;
    END
  END data_wdata_o_10_
  PIN data_wdata_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 446.36 815 446.56 ;
    END
  END data_wdata_o_11_
  PIN data_wdata_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 448.88 815 449.08 ;
    END
  END data_wdata_o_12_
  PIN data_wdata_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 451.4 815 451.6 ;
    END
  END data_wdata_o_13_
  PIN data_wdata_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 453.92 815 454.12 ;
    END
  END data_wdata_o_14_
  PIN data_wdata_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 456.44 815 456.64 ;
    END
  END data_wdata_o_15_
  PIN data_wdata_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 458.96 815 459.16 ;
    END
  END data_wdata_o_16_
  PIN data_wdata_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 461.48 815 461.68 ;
    END
  END data_wdata_o_17_
  PIN data_wdata_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 464 815 464.2 ;
    END
  END data_wdata_o_18_
  PIN data_wdata_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 466.52 815 466.72 ;
    END
  END data_wdata_o_19_
  PIN data_wdata_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 469.04 815 469.24 ;
    END
  END data_wdata_o_1_
  PIN data_wdata_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 471.56 815 471.76 ;
    END
  END data_wdata_o_20_
  PIN data_wdata_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 474.08 815 474.28 ;
    END
  END data_wdata_o_21_
  PIN data_wdata_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 476.6 815 476.8 ;
    END
  END data_wdata_o_22_
  PIN data_wdata_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 479.12 815 479.32 ;
    END
  END data_wdata_o_23_
  PIN data_wdata_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 481.64 815 481.84 ;
    END
  END data_wdata_o_24_
  PIN data_wdata_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 484.16 815 484.36 ;
    END
  END data_wdata_o_25_
  PIN data_wdata_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 486.68 815 486.88 ;
    END
  END data_wdata_o_26_
  PIN data_wdata_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 489.2 815 489.4 ;
    END
  END data_wdata_o_27_
  PIN data_wdata_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 491.72 815 491.92 ;
    END
  END data_wdata_o_28_
  PIN data_wdata_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 494.24 815 494.44 ;
    END
  END data_wdata_o_29_
  PIN data_wdata_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 496.76 815 496.96 ;
    END
  END data_wdata_o_2_
  PIN data_wdata_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 499.28 815 499.48 ;
    END
  END data_wdata_o_30_
  PIN data_wdata_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 501.8 815 502 ;
    END
  END data_wdata_o_31_
  PIN data_wdata_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 504.32 815 504.52 ;
    END
  END data_wdata_o_3_
  PIN data_wdata_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 506.84 815 507.04 ;
    END
  END data_wdata_o_4_
  PIN data_wdata_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 509.36 815 509.56 ;
    END
  END data_wdata_o_5_
  PIN data_wdata_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 511.88 815 512.08 ;
    END
  END data_wdata_o_6_
  PIN data_wdata_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 514.4 815 514.6 ;
    END
  END data_wdata_o_7_
  PIN data_wdata_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 516.92 815 517.12 ;
    END
  END data_wdata_o_8_
  PIN data_wdata_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 519.44 815 519.64 ;
    END
  END data_wdata_o_9_
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 602.6 815 602.8 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 569.84 0.72 570.04 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 418.64 0.72 418.84 ;
    END
  END fetch_enable_i
  PIN hart_id_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 572.36 0.72 572.56 ;
    END
  END hart_id_i_0_
  PIN hart_id_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 574.88 0.72 575.08 ;
    END
  END hart_id_i_10_
  PIN hart_id_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 577.4 0.72 577.6 ;
    END
  END hart_id_i_11_
  PIN hart_id_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 416.12 0.72 416.32 ;
    END
  END hart_id_i_12_
  PIN hart_id_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 579.92 0.72 580.12 ;
    END
  END hart_id_i_13_
  PIN hart_id_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 582.44 0.72 582.64 ;
    END
  END hart_id_i_14_
  PIN hart_id_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 584.96 0.72 585.16 ;
    END
  END hart_id_i_15_
  PIN hart_id_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 413.6 0.72 413.8 ;
    END
  END hart_id_i_16_
  PIN hart_id_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 587.48 0.72 587.68 ;
    END
  END hart_id_i_17_
  PIN hart_id_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 590 0.72 590.2 ;
    END
  END hart_id_i_18_
  PIN hart_id_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 592.52 0.72 592.72 ;
    END
  END hart_id_i_19_
  PIN hart_id_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 411.08 0.72 411.28 ;
    END
  END hart_id_i_1_
  PIN hart_id_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 595.04 0.72 595.24 ;
    END
  END hart_id_i_20_
  PIN hart_id_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 597.56 0.72 597.76 ;
    END
  END hart_id_i_21_
  PIN hart_id_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 600.08 0.72 600.28 ;
    END
  END hart_id_i_22_
  PIN hart_id_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 408.56 0.72 408.76 ;
    END
  END hart_id_i_23_
  PIN hart_id_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 602.6 0.72 602.8 ;
    END
  END hart_id_i_24_
  PIN hart_id_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 605.12 0.72 605.32 ;
    END
  END hart_id_i_25_
  PIN hart_id_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 607.64 0.72 607.84 ;
    END
  END hart_id_i_26_
  PIN hart_id_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 406.04 0.72 406.24 ;
    END
  END hart_id_i_27_
  PIN hart_id_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 610.16 0.72 610.36 ;
    END
  END hart_id_i_28_
  PIN hart_id_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 612.68 0.72 612.88 ;
    END
  END hart_id_i_29_
  PIN hart_id_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 615.2 0.72 615.4 ;
    END
  END hart_id_i_2_
  PIN hart_id_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 403.52 0.72 403.72 ;
    END
  END hart_id_i_30_
  PIN hart_id_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 617.72 0.72 617.92 ;
    END
  END hart_id_i_31_
  PIN hart_id_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 620.24 0.72 620.44 ;
    END
  END hart_id_i_3_
  PIN hart_id_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 622.76 0.72 622.96 ;
    END
  END hart_id_i_4_
  PIN hart_id_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 401 0.72 401.2 ;
    END
  END hart_id_i_5_
  PIN hart_id_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 625.28 0.72 625.48 ;
    END
  END hart_id_i_6_
  PIN hart_id_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 627.8 0.72 628 ;
    END
  END hart_id_i_7_
  PIN hart_id_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 630.32 0.72 630.52 ;
    END
  END hart_id_i_8_
  PIN hart_id_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 398.48 0.72 398.68 ;
    END
  END hart_id_i_9_
  PIN instr_addr_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 587.48 815 587.68 ;
    END
  END instr_addr_o_10_
  PIN instr_addr_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 532.04 815 532.24 ;
    END
  END instr_addr_o_11_
  PIN instr_addr_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 554.72 815 554.92 ;
    END
  END instr_addr_o_12_
  PIN instr_addr_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 600.08 815 600.28 ;
    END
  END instr_addr_o_13_
  PIN instr_addr_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 590 815 590.2 ;
    END
  END instr_addr_o_14_
  PIN instr_addr_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 524.48 815 524.68 ;
    END
  END instr_addr_o_15_
  PIN instr_addr_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 567.32 815 567.52 ;
    END
  END instr_addr_o_16_
  PIN instr_addr_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 552.2 815 552.4 ;
    END
  END instr_addr_o_17_
  PIN instr_addr_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 592.52 815 592.72 ;
    END
  END instr_addr_o_18_
  PIN instr_addr_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 569.84 815 570.04 ;
    END
  END instr_addr_o_19_
  PIN instr_addr_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 534.56 815 534.76 ;
    END
  END instr_addr_o_20_
  PIN instr_addr_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 597.56 815 597.76 ;
    END
  END instr_addr_o_21_
  PIN instr_addr_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 572.36 815 572.56 ;
    END
  END instr_addr_o_22_
  PIN instr_addr_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 557.24 815 557.44 ;
    END
  END instr_addr_o_23_
  PIN instr_addr_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 539.6 815 539.8 ;
    END
  END instr_addr_o_24_
  PIN instr_addr_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 574.88 815 575.08 ;
    END
  END instr_addr_o_25_
  PIN instr_addr_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 564.8 815 565 ;
    END
  END instr_addr_o_26_
  PIN instr_addr_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 529.52 815 529.72 ;
    END
  END instr_addr_o_27_
  PIN instr_addr_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 577.4 815 577.6 ;
    END
  END instr_addr_o_28_
  PIN instr_addr_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 562.28 815 562.48 ;
    END
  END instr_addr_o_29_
  PIN instr_addr_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 547.16 815 547.36 ;
    END
  END instr_addr_o_2_
  PIN instr_addr_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 579.92 815 580.12 ;
    END
  END instr_addr_o_30_
  PIN instr_addr_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 549.68 815 549.88 ;
    END
  END instr_addr_o_31_
  PIN instr_addr_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 527 815 527.2 ;
    END
  END instr_addr_o_3_
  PIN instr_addr_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 582.44 815 582.64 ;
    END
  END instr_addr_o_4_
  PIN instr_addr_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 537.08 815 537.28 ;
    END
  END instr_addr_o_5_
  PIN instr_addr_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 595.04 815 595.24 ;
    END
  END instr_addr_o_6_
  PIN instr_addr_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 542.12 815 542.32 ;
    END
  END instr_addr_o_7_
  PIN instr_addr_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 584.96 815 585.16 ;
    END
  END instr_addr_o_8_
  PIN instr_addr_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 521.96 815 522.16 ;
    END
  END instr_addr_o_9_
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 632.84 0.72 633.04 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 635.36 0.72 635.56 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 637.88 0.72 638.08 ;
    END
  END instr_rdata_i_0_
  PIN instr_rdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 395.96 0.72 396.16 ;
    END
  END instr_rdata_i_10_
  PIN instr_rdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 640.4 0.72 640.6 ;
    END
  END instr_rdata_i_11_
  PIN instr_rdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 642.92 0.72 643.12 ;
    END
  END instr_rdata_i_12_
  PIN instr_rdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 645.44 0.72 645.64 ;
    END
  END instr_rdata_i_13_
  PIN instr_rdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 393.44 0.72 393.64 ;
    END
  END instr_rdata_i_14_
  PIN instr_rdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 647.96 0.72 648.16 ;
    END
  END instr_rdata_i_15_
  PIN instr_rdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 650.48 0.72 650.68 ;
    END
  END instr_rdata_i_16_
  PIN instr_rdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 653 0.72 653.2 ;
    END
  END instr_rdata_i_17_
  PIN instr_rdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 655.52 0.72 655.72 ;
    END
  END instr_rdata_i_18_
  PIN instr_rdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 658.04 0.72 658.24 ;
    END
  END instr_rdata_i_19_
  PIN instr_rdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 660.56 0.72 660.76 ;
    END
  END instr_rdata_i_1_
  PIN instr_rdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 663.08 0.72 663.28 ;
    END
  END instr_rdata_i_20_
  PIN instr_rdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 665.6 0.72 665.8 ;
    END
  END instr_rdata_i_21_
  PIN instr_rdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 668.12 0.72 668.32 ;
    END
  END instr_rdata_i_22_
  PIN instr_rdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 670.64 0.72 670.84 ;
    END
  END instr_rdata_i_23_
  PIN instr_rdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 673.16 0.72 673.36 ;
    END
  END instr_rdata_i_24_
  PIN instr_rdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 675.68 0.72 675.88 ;
    END
  END instr_rdata_i_25_
  PIN instr_rdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 678.2 0.72 678.4 ;
    END
  END instr_rdata_i_26_
  PIN instr_rdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 680.72 0.72 680.92 ;
    END
  END instr_rdata_i_27_
  PIN instr_rdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 683.24 0.72 683.44 ;
    END
  END instr_rdata_i_28_
  PIN instr_rdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 685.76 0.72 685.96 ;
    END
  END instr_rdata_i_29_
  PIN instr_rdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 688.28 0.72 688.48 ;
    END
  END instr_rdata_i_2_
  PIN instr_rdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 690.8 0.72 691 ;
    END
  END instr_rdata_i_30_
  PIN instr_rdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 693.32 0.72 693.52 ;
    END
  END instr_rdata_i_31_
  PIN instr_rdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 695.84 0.72 696.04 ;
    END
  END instr_rdata_i_3_
  PIN instr_rdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 698.36 0.72 698.56 ;
    END
  END instr_rdata_i_4_
  PIN instr_rdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 700.88 0.72 701.08 ;
    END
  END instr_rdata_i_5_
  PIN instr_rdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 703.4 0.72 703.6 ;
    END
  END instr_rdata_i_6_
  PIN instr_rdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 705.92 0.72 706.12 ;
    END
  END instr_rdata_i_7_
  PIN instr_rdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 708.44 0.72 708.64 ;
    END
  END instr_rdata_i_8_
  PIN instr_rdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 710.96 0.72 711.16 ;
    END
  END instr_rdata_i_9_
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 559.76 815 559.96 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 713.48 0.72 713.68 ;
    END
  END instr_rvalid_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 716 0.72 716.2 ;
    END
  END irq_external_i
  PIN irq_fast_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 718.52 0.72 718.72 ;
    END
  END irq_fast_i_0_
  PIN irq_fast_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 721.04 0.72 721.24 ;
    END
  END irq_fast_i_10_
  PIN irq_fast_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 723.56 0.72 723.76 ;
    END
  END irq_fast_i_11_
  PIN irq_fast_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 726.08 0.72 726.28 ;
    END
  END irq_fast_i_12_
  PIN irq_fast_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 728.6 0.72 728.8 ;
    END
  END irq_fast_i_13_
  PIN irq_fast_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 731.12 0.72 731.32 ;
    END
  END irq_fast_i_14_
  PIN irq_fast_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 733.64 0.72 733.84 ;
    END
  END irq_fast_i_15_
  PIN irq_fast_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 736.16 0.72 736.36 ;
    END
  END irq_fast_i_1_
  PIN irq_fast_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 738.68 0.72 738.88 ;
    END
  END irq_fast_i_2_
  PIN irq_fast_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 741.2 0.72 741.4 ;
    END
  END irq_fast_i_3_
  PIN irq_fast_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 743.72 0.72 743.92 ;
    END
  END irq_fast_i_4_
  PIN irq_fast_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 746.24 0.72 746.44 ;
    END
  END irq_fast_i_5_
  PIN irq_fast_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 748.76 0.72 748.96 ;
    END
  END irq_fast_i_6_
  PIN irq_fast_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 751.28 0.72 751.48 ;
    END
  END irq_fast_i_7_
  PIN irq_fast_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 753.8 0.72 754 ;
    END
  END irq_fast_i_8_
  PIN irq_fast_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 756.32 0.72 756.52 ;
    END
  END irq_fast_i_9_
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 758.84 0.72 759.04 ;
    END
  END irq_nm_i
  PIN irq_pending_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  814.28 544.64 815 544.84 ;
    END
  END irq_pending_o
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 761.36 0.72 761.56 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 763.88 0.72 764.08 ;
    END
  END irq_timer_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 766.4 0.72 766.6 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 874.76 0.72 874.96 ;
    END
  END test_en_i
  OBS
    LAYER Metal1 ;
     RECT  789.52 17.98 789.68 20.5 ;
     RECT  789.04 20.5 789.68 23.02 ;
     RECT  781.84 23.02 789.68 26.24 ;
     RECT  25.44 26.24 789.68 30.58 ;
     RECT  25.44 30.58 795.44 35.62 ;
     RECT  25.44 35.62 799.28 38.14 ;
     RECT  810.64 33.1 810.8 38.14 ;
     RECT  25.44 38.14 810.8 39.56 ;
     RECT  25.44 39.56 802.64 50.74 ;
     RECT  25.44 50.74 803.12 51.16 ;
     RECT  813.52 40.66 813.68 51.16 ;
     RECT  25.44 51.16 813.68 58.3 ;
     RECT  25.44 58.3 814.16 111.64 ;
     RECT  25.44 111.64 814.64 144.56 ;
     RECT  25.44 144.56 814.16 193.28 ;
     RECT  25.44 193.28 813.68 207.82 ;
     RECT  24.88 207.82 813.68 214.54 ;
     RECT  18.16 214.54 813.68 217.06 ;
     RECT  18.16 217.06 814.16 232.6 ;
     RECT  18.16 232.6 814.64 233.6 ;
     RECT  1.84 193.12 2 242.26 ;
     RECT  18.16 233.6 797.36 252.34 ;
     RECT  807.28 233.6 814.64 252.34 ;
     RECT  1.84 242.26 3.44 254.44 ;
     RECT  18.16 252.34 814.64 254.44 ;
     RECT  1.84 254.44 814.64 270.98 ;
     RECT  1.84 270.98 813.68 271.82 ;
     RECT  806.32 271.82 813.68 273.92 ;
     RECT  807.28 273.92 813.68 276.02 ;
     RECT  1.84 271.82 795.44 282.16 ;
     RECT  807.28 276.02 812.24 292.66 ;
     RECT  806.32 292.66 812.24 298.54 ;
     RECT  806.32 298.54 812.72 306.1 ;
     RECT  806.32 306.1 814.16 309.62 ;
     RECT  807.28 309.62 814.16 310.46 ;
     RECT  807.28 310.46 812.72 323.74 ;
     RECT  806.32 323.74 812.72 325 ;
     RECT  806.32 325 814.16 330.62 ;
     RECT  806.8 330.62 814.16 333.14 ;
     RECT  806.8 333.14 813.68 338.18 ;
     RECT  812.08 338.18 813.68 356.08 ;
     RECT  809.2 356.08 813.68 367.12 ;
     RECT  809.2 367.12 814.16 388.58 ;
     RECT  0.4 282.16 795.44 405.8 ;
     RECT  812.56 388.58 814.16 416.3 ;
     RECT  812.56 416.3 812.72 426.38 ;
     RECT  0.4 405.8 791.6 440.66 ;
     RECT  0.4 440.66 791.12 451.42 ;
     RECT  810.16 441.34 810.32 458.98 ;
     RECT  809.2 458.98 810.32 460.82 ;
     RECT  0.4 451.42 799.28 462.08 ;
     RECT  809.2 460.82 809.36 469.06 ;
     RECT  0.4 462.08 792.56 475.36 ;
     RECT  802.48 469.06 809.36 475.36 ;
     RECT  0.4 475.36 809.36 484.76 ;
     RECT  0.4 484.76 807.92 486.86 ;
     RECT  802 486.86 807.92 496.94 ;
     RECT  802.48 496.94 807.92 501.56 ;
     RECT  0.4 486.86 792.08 507.44 ;
     RECT  802.48 501.56 802.64 520.46 ;
     RECT  0.4 507.44 791.6 522.56 ;
     RECT  0.4 522.56 791.12 539.62 ;
     RECT  0.4 539.62 795.44 570.86 ;
     RECT  0.4 570.86 791.6 584.98 ;
     RECT  0.4 584.98 792.56 587.66 ;
     RECT  17.68 587.66 792.56 605.3 ;
     RECT  0.4 587.66 6.32 610.34 ;
     RECT  17.68 605.3 790.64 613.28 ;
     RECT  17.68 613.28 790.16 617.06 ;
     RECT  17.68 617.06 789.6 642.1 ;
     RECT  0.4 610.34 4.88 643.36 ;
     RECT  14.8 642.1 789.6 643.36 ;
     RECT  0.4 643.36 789.6 643.52 ;
     RECT  0.4 643.52 4.88 725.84 ;
     RECT  0.88 725.84 4.88 736.34 ;
     RECT  0.88 736.34 3.92 743.9 ;
     RECT  1.36 743.9 3.92 748.94 ;
     RECT  2.8 748.94 3.92 753.98 ;
     RECT  3.76 753.98 3.92 759.02 ;
     RECT  17.68 643.52 789.6 769.1 ;
     RECT  25.44 769.1 789.6 888.52 ;
    LAYER Metal2 ;
     RECT  0.38 400.58 0.48 400.78 ;
     RECT  0.38 412.34 0.48 413.38 ;
     RECT  0.38 505.16 0.48 506.62 ;
     RECT  0.38 522.38 0.48 529.3 ;
     RECT  0.38 540.02 0.48 543.58 ;
     RECT  0.38 578.66 0.48 579.7 ;
     RECT  0.38 638.3 0.48 645.22 ;
     RECT  0.38 671.06 0.48 672.52 ;
     RECT  0.38 707.18 0.48 708.22 ;
     RECT  0.38 723.14 0.48 725.86 ;
     RECT  0.48 393.44 1.06 769.12 ;
     RECT  0.86 309.02 1.34 309.22 ;
     RECT  1.06 731.12 1.54 769.12 ;
     RECT  1.54 731.12 2.02 741.4 ;
     RECT  0.38 282.14 2.3 282.34 ;
     RECT  1.06 393.44 2.5 721.24 ;
     RECT  2.5 393.44 3.46 713.68 ;
     RECT  2.02 733.64 3.94 741.4 ;
     RECT  1.54 751.28 3.94 769.12 ;
     RECT  3.46 630.32 4.42 675.88 ;
     RECT  3.94 736.16 4.42 741.4 ;
     RECT  2.78 339.68 4.7 339.88 ;
     RECT  4.42 736.16 4.9 736.36 ;
     RECT  3.94 751.28 4.9 751.48 ;
     RECT  4.22 261.56 5.18 261.76 ;
     RECT  5.18 261.56 5.66 264.7 ;
     RECT  3.46 393.44 5.86 617.92 ;
     RECT  2.3 282.14 6.14 290.74 ;
     RECT  5.86 406.04 6.34 617.92 ;
     RECT  3.94 761.36 6.34 769.12 ;
     RECT  5.86 393.44 7.3 396.16 ;
     RECT  6.34 406.04 7.3 602.8 ;
     RECT  6.34 612.68 7.3 617.92 ;
     RECT  4.42 632.84 7.3 675.88 ;
     RECT  3.46 690.8 7.3 713.68 ;
     RECT  5.66 261.56 10.46 272.26 ;
     RECT  4.7 339.68 10.94 343.66 ;
     RECT  7.3 411.08 11.14 600.28 ;
     RECT  11.14 411.08 11.62 597.76 ;
     RECT  11.62 411.08 14.02 582.64 ;
     RECT  7.3 395.96 14.3 396.16 ;
     RECT  6.14 282.14 14.5 294.52 ;
     RECT  14.3 395.96 14.5 397 ;
     RECT  14.02 411.08 14.5 565 ;
     RECT  6.34 766.4 17.86 769.12 ;
     RECT  14.02 574.88 18.34 582.64 ;
     RECT  14.5 411.08 18.82 564.16 ;
     RECT  11.62 592.52 18.82 597.76 ;
     RECT  10.94 331.7 19.1 343.66 ;
     RECT  1.34 309.02 24.38 313.84 ;
     RECT  19.1 324.98 24.38 343.66 ;
     RECT  18.14 214.52 24.86 214.72 ;
     RECT  18.82 592.52 25.06 592.72 ;
     RECT  17.86 766.4 26.78 766.6 ;
     RECT  26.78 765.56 26.98 766.6 ;
     RECT  7.3 692.9 28.7 713.68 ;
     RECT  7.3 637.88 29.18 675.88 ;
     RECT  18.82 412.34 29.66 564.16 ;
     RECT  24.86 207.8 30.14 214.72 ;
     RECT  29.66 179.66 30.56 182.38 ;
     RECT  30.14 206.54 30.62 214.72 ;
     RECT  30.14 227.96 30.62 231.94 ;
     RECT  1.82 193.1 31.1 193.3 ;
     RECT  29.66 412.34 31.1 569.2 ;
     RECT  18.34 578.24 31.1 578.44 ;
     RECT  30.56 179.625 31.58 182.38 ;
     RECT  3.26 242.24 31.58 242.44 ;
     RECT  10.46 254.42 31.58 272.26 ;
     RECT  24.38 309.02 31.58 343.66 ;
     RECT  31.58 179.24 32 182.38 ;
     RECT  31.1 191.42 32 193.3 ;
     RECT  30.62 206.54 32 231.94 ;
     RECT  29.18 629.48 32.06 675.88 ;
     RECT  32 179.24 33.02 193.3 ;
     RECT  31.58 242.24 33.5 274.78 ;
     RECT  14.5 283.4 33.5 294.52 ;
     RECT  32 205.53 34.46 232.95 ;
     RECT  33.5 242.24 34.46 294.52 ;
     RECT  32.06 628.22 35.14 675.88 ;
     RECT  33.02 178.82 35.42 193.3 ;
     RECT  34.46 205.53 35.42 294.52 ;
     RECT  31.58 304.4 35.42 343.66 ;
     RECT  23.9 358.58 35.42 358.78 ;
     RECT  35.42 178.82 35.9 343.66 ;
     RECT  35.14 629.48 35.9 675.88 ;
     RECT  28.7 691.22 35.9 713.68 ;
     RECT  35.42 358.58 36.1 367.6 ;
     RECT  3.74 377.06 36.86 377.26 ;
     RECT  35.9 629.48 37.54 676.72 ;
     RECT  35.9 178.82 37.82 345.34 ;
     RECT  36.86 374.96 37.82 377.26 ;
     RECT  35.9 387.56 37.82 387.76 ;
     RECT  37.82 178.82 38.3 345.76 ;
     RECT  38.3 171.68 38.78 345.76 ;
     RECT  38.78 170.84 39.26 345.76 ;
     RECT  31.1 412.34 39.26 578.44 ;
     RECT  39.26 167.9 40.22 345.76 ;
     RECT  39.26 412.34 40.7 584.74 ;
     RECT  40.22 167.9 43.1 346.6 ;
     RECT  36.1 358.58 43.1 358.78 ;
     RECT  37.82 374.96 43.58 387.76 ;
     RECT  14.5 396.8 43.58 397 ;
     RECT  43.1 610.58 44 613.3 ;
     RECT  43.1 167.9 44.06 358.78 ;
     RECT  44 610.545 44.06 613.3 ;
     RECT  43.58 374.96 45.5 397 ;
     RECT  44.06 164.54 45.98 358.78 ;
     RECT  45.5 372.86 45.98 397 ;
     RECT  44.06 607.22 46.46 613.3 ;
     RECT  45.98 164.54 47.36 397 ;
     RECT  46.46 607.22 47.9 614.56 ;
     RECT  47.36 164.505 48.38 397 ;
     RECT  47.9 607.22 48.38 614.98 ;
     RECT  37.54 635.36 48.38 676.72 ;
     RECT  48.38 629.48 48.86 676.72 ;
     RECT  48.38 607.22 49.28 617.5 ;
     RECT  48.38 164.12 50.3 397 ;
     RECT  49.28 607.22 50.3 618.51 ;
     RECT  48.86 628.22 50.3 676.72 ;
     RECT  50.3 164.12 50.78 398.68 ;
     RECT  40.7 412.34 50.78 597.34 ;
     RECT  50.3 607.22 52.22 676.72 ;
     RECT  50.78 164.12 52.42 597.34 ;
     RECT  52.42 428.72 52.7 597.34 ;
     RECT  52.22 606.38 52.7 676.72 ;
     RECT  52.42 164.12 55.1 420.1 ;
     RECT  35.9 691.22 57.5 714.1 ;
     RECT  57.5 690.8 57.98 714.1 ;
     RECT  52.7 428.72 58.46 676.72 ;
     RECT  57.98 688.28 58.46 714.1 ;
     RECT  55.1 163.7 66.14 420.1 ;
     RECT  58.46 428.72 66.14 714.1 ;
     RECT  66.14 163.7 69.98 714.1 ;
     RECT  69.98 156.14 79.58 714.1 ;
     RECT  79.58 153.62 83.42 714.1 ;
     RECT  83.42 152.78 83.9 716.2 ;
     RECT  83.9 151.94 94.46 716.2 ;
     RECT  94.46 151.94 96.38 716.62 ;
     RECT  96.38 146.06 96.8 716.62 ;
     RECT  96.8 146.06 97.28 716.79 ;
     RECT  97.28 145.05 100.22 716.79 ;
     RECT  100.22 145.05 101.12 727.54 ;
     RECT  101.12 145.05 102.14 727.575 ;
     RECT  102.14 145.05 105.02 728.38 ;
     RECT  105.02 144.8 112.9 728.38 ;
     RECT  112.9 145.64 113.86 728.38 ;
     RECT  113.86 146.06 114.82 728.38 ;
     RECT  114.82 146.06 121.045 727.54 ;
     RECT  121.045 146.06 123.2 726.7 ;
     RECT  123.2 145.05 124.42 726.7 ;
     RECT  124.42 145.05 125.86 725.02 ;
     RECT  125.86 145.05 136.22 724.6 ;
     RECT  136.22 144.8 139.1 727.12 ;
     RECT  139.1 142.7 141.02 727.12 ;
     RECT  141.02 141.44 141.22 727.12 ;
     RECT  141.22 141.86 142.46 727.12 ;
     RECT  142.46 141.86 144.58 727.96 ;
     RECT  144.58 141.86 149.66 727.12 ;
     RECT  149.66 138.5 151.52 727.12 ;
     RECT  151.52 137.49 157.54 727.12 ;
     RECT  157.54 137.49 158.965 726.7 ;
     RECT  158.965 137.66 172.22 726.7 ;
     RECT  172.22 134.3 173.12 728.8 ;
     RECT  173.12 134.265 174.14 728.8 ;
     RECT  174.14 133.88 180.38 728.8 ;
     RECT  180.38 133.46 181.54 728.8 ;
     RECT  181.54 133.46 183.46 727.96 ;
     RECT  183.46 133.46 186.805 727.54 ;
     RECT  186.805 133.46 187.1 726.7 ;
     RECT  187.1 130.94 190.18 726.7 ;
     RECT  190.18 130.94 190.46 724.615 ;
     RECT  190.46 130.52 196.7 724.615 ;
     RECT  196.7 123.38 198.56 724.615 ;
     RECT  198.56 122.37 199.1 724.615 ;
     RECT  199.1 115.82 201.5 724.615 ;
     RECT  201.5 114.56 204.515 724.615 ;
     RECT  204.515 114.56 204.965 723.78 ;
     RECT  209.66 104.06 210.14 104.26 ;
     RECT  204.965 114.56 210.14 721.24 ;
     RECT  210.14 104.06 210.56 721.24 ;
     RECT  210.56 104.025 214.18 721.24 ;
     RECT  214.18 104.025 216.1 714.1 ;
     RECT  216.1 104.025 218.3 713.68 ;
     RECT  218.3 101.12 220.22 713.68 ;
     RECT  220.22 96.08 222.14 713.68 ;
     RECT  222.14 91.46 224.48 713.68 ;
     RECT  224.48 88.905 225.5 713.68 ;
     RECT  220.22 77.6 228.38 77.8 ;
     RECT  225.5 88.52 228.38 713.68 ;
     RECT  228.38 76.76 235.78 713.68 ;
     RECT  235.78 77.18 251.9 713.68 ;
     RECT  251.9 77.18 262.46 714.52 ;
     RECT  262.46 77.18 264.32 715.78 ;
     RECT  264.32 77.18 270.14 716.79 ;
     RECT  270.14 76.76 270.62 716.79 ;
     RECT  270.62 76.76 271.1 719.98 ;
     RECT  271.1 76.76 271.3 723.34 ;
     RECT  271.3 77.01 275.9 723.34 ;
     RECT  275.9 77.01 276.38 724.18 ;
     RECT  276.38 77.01 277.34 725.02 ;
     RECT  277.34 77.01 278.02 727.96 ;
     RECT  278.02 77.01 279.445 727.12 ;
     RECT  279.445 77.18 285.22 727.12 ;
     RECT  285.22 80.96 287.62 727.12 ;
     RECT  287.62 81.38 289.06 727.12 ;
     RECT  289.06 84.32 290.02 727.12 ;
     RECT  30.62 764.3 290.98 764.5 ;
     RECT  290.02 86.42 291.26 727.12 ;
     RECT  291.26 86.42 294.62 735.52 ;
     RECT  294.62 86.42 296.48 736.36 ;
     RECT  296.48 86.42 300.1 739.47 ;
     RECT  300.1 86.42 300.775 158.86 ;
     RECT  300.775 85.58 301.555 158.86 ;
     RECT  300.1 167.48 303.925 739.47 ;
     RECT  301.555 84.74 309.98 158.86 ;
     RECT  303.925 167.48 309.98 739.3 ;
     RECT  309.98 84.74 310.375 739.3 ;
     RECT  310.375 78.02 311.155 739.3 ;
     RECT  311.155 77.18 311.42 739.3 ;
     RECT  311.42 74.24 312.38 739.3 ;
     RECT  312.38 73.4 313.28 739.3 ;
     RECT  313.28 73.4 322.46 739.47 ;
     RECT  322.46 70.46 323.36 739.47 ;
     RECT  323.36 69.45 326.3 739.47 ;
     RECT  326.3 69.45 331.1 739.72 ;
     RECT  331.1 65 337.82 739.72 ;
     RECT  337.82 58.28 340.22 739.72 ;
     RECT  340.22 57.86 348.1 739.72 ;
     RECT  348.1 57.86 354.82 736.36 ;
     RECT  354.82 60.8 360.1 736.36 ;
     RECT  360.1 60.8 363.97 735.135 ;
     RECT  363.97 60.8 380.48 735.1 ;
     RECT  380.48 60.8 380.77 735.135 ;
     RECT  386.3 51.14 387.2 52.18 ;
     RECT  387.2 51.105 388.22 52.18 ;
     RECT  380.77 60.8 388.22 735.1 ;
     RECT  388.22 51.105 389.18 735.1 ;
     RECT  389.18 50.3 394.66 735.1 ;
     RECT  394.66 50.3 395.9 732.16 ;
     RECT  395.9 48.2 396.1 732.16 ;
     RECT  396.1 48.2 397.34 731.91 ;
     RECT  397.34 43.58 401.18 731.91 ;
     RECT  401.18 43.16 403.1 731.91 ;
     RECT  403.1 41.06 404 731.91 ;
     RECT  404 39.21 404.06 731.91 ;
     RECT  404.06 38.54 404.245 731.91 ;
     RECT  404.245 38.54 408.86 731.32 ;
     RECT  408.86 29.3 410.5 731.32 ;
     RECT  410.5 29.3 417.5 730.9 ;
     RECT  417.5 27.2 421.54 730.9 ;
     RECT  421.54 27.2 422.02 726.28 ;
     RECT  422.02 28.04 423.94 726.28 ;
     RECT  423.94 28.04 427.78 714.52 ;
     RECT  427.78 698.78 428.74 714.52 ;
     RECT  428.74 708.43 429.125 714.52 ;
     RECT  429.125 708.44 429.7 714.52 ;
     RECT  423.94 726.08 429.7 726.28 ;
     RECT  427.78 28.04 432.1 685.12 ;
     RECT  428.74 698.78 433.06 699.4 ;
     RECT  432.1 28.04 434.5 681.34 ;
     RECT  434.5 33.08 434.98 681.34 ;
     RECT  434.98 34.34 436.9 678.82 ;
     RECT  433.06 698.78 439.78 698.98 ;
     RECT  436.9 34.34 441.22 677.56 ;
     RECT  441.22 34.34 445.54 676.3 ;
     RECT  445.54 34.34 451.78 672.1 ;
     RECT  451.78 34.34 460.42 671.68 ;
     RECT  460.42 36.02 460.9 671.68 ;
     RECT  460.9 39.21 462.34 671.68 ;
     RECT  462.34 39.21 467.14 666.64 ;
     RECT  467.14 39.21 467.62 651.52 ;
     RECT  467.14 666.44 467.62 666.64 ;
     RECT  467.62 39.21 468.34 625.9 ;
     RECT  468.34 39.21 468.565 625.48 ;
     RECT  467.62 635.78 468.58 651.52 ;
     RECT  468.58 635.78 469.06 642.7 ;
     RECT  468.565 40.64 469.075 625.48 ;
     RECT  469.06 636.2 470.98 642.7 ;
     RECT  469.075 40.64 471.94 620.86 ;
     RECT  471.94 46.1 472.9 620.86 ;
     RECT  472.9 46.77 475.285 620.86 ;
     RECT  429.7 714.32 477.7 714.52 ;
     RECT  470.98 642.5 480.38 642.7 ;
     RECT  475.285 47.78 482.3 620.86 ;
     RECT  480.38 635.78 483.26 642.7 ;
     RECT  483.26 635.78 484.7 643.96 ;
     RECT  484.7 635.78 485.18 644.8 ;
     RECT  482.3 47.78 485.42 622.12 ;
     RECT  485.18 635.78 485.42 648.16 ;
     RECT  485.42 47.78 485.66 648.16 ;
     RECT  485.66 47.78 486.14 649 ;
     RECT  485.18 670.22 486.14 670.84 ;
     RECT  486.14 668.12 486.62 672.1 ;
     RECT  486.62 668.12 487.1 675.46 ;
     RECT  487.1 668.12 487.58 676.72 ;
     RECT  486.14 47.78 489.02 655.72 ;
     RECT  489.02 47.78 489.5 656.14 ;
     RECT  487.58 668.12 489.5 682.18 ;
     RECT  489.5 47.78 489.98 685.96 ;
     RECT  489.5 715.58 491.42 715.78 ;
     RECT  490.46 728.18 491.42 728.38 ;
     RECT  489.98 696.26 491.9 696.46 ;
     RECT  491.9 696.26 493.34 697.72 ;
     RECT  489.98 47.78 493.82 686.8 ;
     RECT  493.34 696.26 493.82 701.5 ;
     RECT  493.82 47.78 494.78 701.5 ;
     RECT  494.78 47.78 496.7 705.28 ;
     RECT  491.42 715.58 496.7 728.38 ;
     RECT  496.7 47.78 497.38 728.38 ;
     RECT  497.38 51.98 498.62 728.38 ;
     RECT  498.62 51.98 501.82 729.22 ;
     RECT  501.82 51.98 503.9 732.16 ;
     RECT  503.9 51.98 506.3 736.78 ;
     RECT  506.3 51.98 506.78 737.2 ;
     RECT  506.78 51.98 508.22 738.88 ;
     RECT  508.22 51.98 510.14 746.44 ;
     RECT  510.14 51.98 511.58 750.64 ;
     RECT  511.58 51.98 512.54 751.48 ;
     RECT  512.06 760.94 512.54 761.56 ;
     RECT  512.54 51.98 512.78 761.56 ;
     RECT  512.78 51.98 513.5 762.82 ;
     RECT  513.5 51.98 517.34 764.5 ;
     RECT  517.34 51.98 518.3 766.18 ;
     RECT  518.3 51.98 522.62 766.6 ;
     RECT  522.62 51.98 528.86 768.7 ;
     RECT  528.86 51.98 529.34 769.96 ;
     RECT  529.34 51.98 533.18 776.26 ;
     RECT  533.18 51.98 534.505 776.68 ;
     RECT  534.505 46.505 537.98 776.68 ;
     RECT  537.98 46.505 540.825 777.1 ;
     RECT  540.825 46.505 541.34 780.46 ;
     RECT  541.34 46.505 543.74 788.44 ;
     RECT  543.74 46.505 546.62 791.38 ;
     RECT  546.62 46.505 549.925 794.74 ;
     RECT  549.925 46.505 553.06 796 ;
     RECT  553.06 46.505 562.46 795.58 ;
     RECT  562.46 46.505 566.435 798.1 ;
     RECT  566.435 47.34 566.885 798.1 ;
     RECT  566.885 47.36 567.46 798.1 ;
     RECT  567.46 50.875 568.17 798.1 ;
     RECT  568.17 51.98 570.14 798.1 ;
     RECT  569.18 807.14 570.14 807.34 ;
     RECT  570.14 51.98 577.1 807.34 ;
     RECT  577.1 51.98 577.34 808.18 ;
     RECT  559.58 834.44 579.74 834.64 ;
     RECT  577.82 818.48 580.585 818.68 ;
     RECT  580.585 818.48 580.7 822.04 ;
     RECT  577.34 51.98 581.9 809.86 ;
     RECT  580.7 818.48 581.9 823.3 ;
     RECT  581.9 51.98 583.58 823.3 ;
     RECT  583.58 51.98 590.02 824.98 ;
     RECT  590.02 51.98 590.3 52.18 ;
     RECT  590.3 51.14 590.5 52.18 ;
     RECT  590.02 62.48 592.22 824.98 ;
     RECT  592.22 62.48 592.42 825.82 ;
     RECT  592.42 71.72 592.7 825.82 ;
     RECT  579.74 834.44 592.7 835.9 ;
     RECT  592.7 71.72 597.98 835.9 ;
     RECT  597.98 71.72 600.58 836.74 ;
     RECT  600.58 71.72 609.465 836.32 ;
     RECT  609.465 71.72 612.86 837.58 ;
     RECT  612.86 71.72 614.78 840.52 ;
     RECT  614.78 71.72 615.74 841.36 ;
     RECT  615.74 71.72 619.1 841.78 ;
     RECT  619.1 71.3 623.42 841.78 ;
     RECT  623.42 71.3 626.78 842.2 ;
     RECT  626.78 71.3 629.38 844.72 ;
     RECT  629.38 71.3 638.98 841.78 ;
     RECT  638.98 833.6 642.82 833.8 ;
     RECT  638.98 71.3 648.1 823.3 ;
     RECT  648.1 105.32 657.22 823.3 ;
     RECT  657.22 105.32 657.7 822.04 ;
     RECT  657.7 802.1 660.58 822.04 ;
     RECT  660.58 802.1 662.02 821.62 ;
     RECT  662.02 815.54 662.5 821.62 ;
     RECT  662.02 802.1 663.94 802.3 ;
     RECT  648.1 71.3 669.5 96.28 ;
     RECT  657.7 105.32 686.98 792.22 ;
     RECT  686.98 792.02 691.3 792.22 ;
     RECT  686.98 105.32 692.26 780.04 ;
     RECT  669.5 71.3 695.9 96.7 ;
     RECT  692.26 105.32 695.9 777.52 ;
     RECT  695.9 71.3 697.54 777.52 ;
     RECT  662.5 815.54 701.38 815.74 ;
     RECT  697.54 115.4 705.7 777.52 ;
     RECT  705.7 755.9 708.58 776.68 ;
     RECT  708.58 755.9 709.06 774.16 ;
     RECT  709.06 773.12 709.54 774.16 ;
     RECT  709.54 773.12 710.02 773.74 ;
     RECT  710.02 773.12 710.98 773.32 ;
     RECT  705.7 115.4 711.46 746.02 ;
     RECT  709.06 760.52 711.46 760.72 ;
     RECT  711.46 124.22 712.42 746.02 ;
     RECT  712.42 124.22 712.9 730.9 ;
     RECT  712.42 745.82 712.9 746.02 ;
     RECT  712.9 124.22 714.835 729.22 ;
     RECT  714.835 671.48 715.3 729.22 ;
     RECT  715.3 671.48 718.18 727.12 ;
     RECT  718.18 671.9 718.66 727.12 ;
     RECT  718.66 671.9 719.14 724.18 ;
     RECT  719.14 716.21 719.38 724.18 ;
     RECT  714.835 124.22 719.62 662.86 ;
     RECT  719.14 671.9 719.62 706.12 ;
     RECT  719.38 716.84 719.62 724.18 ;
     RECT  719.62 125.06 720.1 662.86 ;
     RECT  719.62 677.36 720.1 706.12 ;
     RECT  719.62 716.84 720.34 719.56 ;
     RECT  720.1 125.06 720.58 653.2 ;
     RECT  720.58 125.06 721.54 652.36 ;
     RECT  720.1 677.36 721.54 705.28 ;
     RECT  721.54 621.92 722.02 652.36 ;
     RECT  720.1 662.66 722.02 662.86 ;
     RECT  721.54 701.72 722.5 705.28 ;
     RECT  721.54 125.06 723.46 613.3 ;
     RECT  721.54 677.36 723.46 692.68 ;
     RECT  722.02 621.92 724.66 651.94 ;
     RECT  724.66 621.92 724.9 627.58 ;
     RECT  724.66 637.04 724.9 651.94 ;
     RECT  723.46 692.48 724.9 692.68 ;
     RECT  724.9 637.04 725.38 637.24 ;
     RECT  723.46 681.14 725.38 681.34 ;
     RECT  724.9 622.76 725.62 627.58 ;
     RECT  724.9 648.38 725.86 651.94 ;
     RECT  720.34 719.36 725.86 719.56 ;
     RECT  725.62 627.38 727.3 627.58 ;
     RECT  725.86 651.74 727.3 651.94 ;
     RECT  723.46 125.06 735.74 603.39 ;
     RECT  723.46 612.68 735.74 613.3 ;
     RECT  735.74 125.06 737.6 614.14 ;
     RECT  737.6 125.06 738.62 614.175 ;
     RECT  738.62 125.06 739.58 614.56 ;
     RECT  739.58 125.06 740.48 621.7 ;
     RECT  740.48 125.06 741.02 621.735 ;
     RECT  741.02 125.06 741.7 622.12 ;
     RECT  741.7 125.06 745.06 621.7 ;
     RECT  745.06 164.96 755.84 621.7 ;
     RECT  755.84 164.96 756.38 621.735 ;
     RECT  651.26 39.38 759.26 39.58 ;
     RECT  590.5 51.14 759.26 51.34 ;
     RECT  756.38 164.96 768.38 622.12 ;
     RECT  768.38 164.96 775.78 625.9 ;
     RECT  775.78 164.96 781.045 621.7 ;
     RECT  745.06 125.06 781.34 156.34 ;
     RECT  781.045 164.96 781.34 620.86 ;
     RECT  759.26 39.38 781.82 51.34 ;
     RECT  781.34 125.06 784.42 620.86 ;
     RECT  781.82 23 785.66 23.2 ;
     RECT  781.82 33.08 785.66 51.34 ;
     RECT  784.42 125.06 785.845 618.51 ;
     RECT  697.54 71.3 788.06 105.52 ;
     RECT  785.66 23 789.02 51.34 ;
     RECT  785.845 125.06 789.22 617.08 ;
     RECT  789.02 20.48 789.5 51.34 ;
     RECT  789.5 17.96 789.7 51.34 ;
     RECT  789.22 125.06 790.18 414.22 ;
     RECT  789.22 423.26 790.18 617.08 ;
     RECT  790.18 125.06 790.66 345.76 ;
     RECT  790.18 423.68 790.66 613.3 ;
     RECT  790.66 423.68 791.62 612.04 ;
     RECT  790.66 125.06 792.1 342.4 ;
     RECT  790.18 354.8 792.58 414.22 ;
     RECT  791.62 443.84 792.58 612.04 ;
     RECT  792.1 340.52 793.54 342.4 ;
     RECT  789.7 17.96 799.1 30.76 ;
     RECT  789.7 39.38 799.1 51.34 ;
     RECT  791.62 423.68 801.5 433.96 ;
     RECT  792.58 443.84 801.5 602.38 ;
     RECT  801.5 423.68 802.46 602.38 ;
     RECT  592.42 62.48 803.42 62.68 ;
     RECT  788.06 71.3 803.42 106.36 ;
     RECT  711.46 115.4 806.3 115.6 ;
     RECT  792.1 125.06 806.3 330.22 ;
     RECT  793.54 340.52 806.3 340.72 ;
     RECT  792.58 354.8 806.3 413.8 ;
     RECT  802.46 423.68 806.3 602.8 ;
     RECT  792.58 611.84 806.5 612.04 ;
     RECT  799.1 17.96 806.78 51.34 ;
     RECT  803.42 62.48 806.78 106.36 ;
     RECT  806.3 115.4 806.78 330.64 ;
     RECT  806.3 340.52 806.78 343.24 ;
     RECT  806.78 17.96 807.74 106.36 ;
     RECT  806.78 115.4 807.74 343.24 ;
     RECT  807.74 17.96 811.1 343.24 ;
     RECT  806.3 354.8 811.1 602.8 ;
     RECT  811.1 17.96 814.56 602.8 ;
     RECT  814.56 25.94 814.66 27.4 ;
     RECT  814.56 48.62 814.66 50.5 ;
     RECT  814.56 61.22 814.66 62.68 ;
     RECT  814.56 111.62 814.66 111.82 ;
     RECT  814.56 125.06 814.66 126.1 ;
     RECT  814.56 144.38 814.66 144.58 ;
     RECT  814.56 154.46 814.66 163.9 ;
     RECT  814.56 185.54 814.66 186.58 ;
     RECT  814.56 232.58 814.66 247.06 ;
     RECT  814.56 277.94 814.66 297.46 ;
     RECT  814.56 306.5 814.66 315.1 ;
     RECT  814.56 353.54 814.66 375.58 ;
     RECT  814.56 391.34 814.66 393.22 ;
     RECT  814.56 406.46 814.66 407.92 ;
     RECT  814.56 449.3 814.66 450.76 ;
     RECT  814.56 464.42 814.66 466.3 ;
     RECT  814.56 498.02 814.66 499.06 ;
     RECT  814.56 520.7 814.66 524.26 ;
     RECT  814.56 534.98 814.66 602.38 ;
    LAYER Metal3 ;
     RECT  421.82 27.2 422.02 28.04 ;
     RECT  421.82 28.04 422.98 28.88 ;
     RECT  434.3 28.04 434.5 28.88 ;
     RECT  421.82 28.88 434.5 31.82 ;
     RECT  417.02 31.82 434.5 32.24 ;
     RECT  412.22 32.24 434.5 34.34 ;
     RECT  412.22 34.34 439.78 35.6 ;
     RECT  412.22 35.6 448.9 36.02 ;
     RECT  411.26 36.02 450.34 38.54 ;
     RECT  460.7 36.02 460.9 38.54 ;
     RECT  411.26 38.54 460.9 39.38 ;
     RECT  404.06 39.38 460.9 39.8 ;
     RECT  404.06 39.8 462.34 40.22 ;
     RECT  810.62 43.16 810.82 45.68 ;
     RECT  403.1 40.22 468.58 46.94 ;
     RECT  403.1 46.94 472.9 47.36 ;
     RECT  400.22 47.36 472.9 48.2 ;
     RECT  542.3 47.78 542.5 48.2 ;
     RECT  395.9 48.2 472.9 50.3 ;
     RECT  539.42 48.2 548.26 50.3 ;
     RECT  395.9 50.3 474.34 50.72 ;
     RECT  538.94 50.3 548.26 51.14 ;
     RECT  561.5 50.72 561.7 51.14 ;
     RECT  388.22 50.72 479.62 51.56 ;
     RECT  497.18 47.78 497.38 54.5 ;
     RECT  538.94 51.14 561.7 54.92 ;
     RECT  388.22 51.56 480.1 55.34 ;
     RECT  489.98 54.5 497.38 55.34 ;
     RECT  340.7 57.86 340.9 58.28 ;
     RECT  388.22 55.34 497.38 58.28 ;
     RECT  538.94 54.92 569.86 58.28 ;
     RECT  528.86 51.98 529.06 58.7 ;
     RECT  538.94 58.28 571.3 58.7 ;
     RECT  337.82 58.28 340.9 59.54 ;
     RECT  528.86 58.7 577.06 59.54 ;
     RECT  354.62 57.86 354.82 60.8 ;
     RECT  524.54 59.54 577.06 60.8 ;
     RECT  589.82 58.7 590.02 60.8 ;
     RECT  524.54 60.8 590.02 62.06 ;
     RECT  517.34 62.06 590.98 64.9 ;
     RECT  337.82 59.54 341.38 65 ;
     RECT  331.1 65 341.38 65.84 ;
     RECT  354.62 60.8 362.5 65.84 ;
     RECT  377.18 65.42 377.38 65.84 ;
     RECT  388.22 58.28 498.82 65.84 ;
     RECT  517.34 64.9 590.5 65.84 ;
     RECT  331.1 65.84 500.74 66.26 ;
     RECT  331.1 66.26 504.58 67.94 ;
     RECT  331.1 67.94 506.02 69.2 ;
     RECT  331.1 69.2 506.98 69.62 ;
     RECT  325.82 69.62 506.98 70.04 ;
     RECT  325.34 70.04 506.98 70.88 ;
     RECT  516.86 65.84 590.5 70.88 ;
     RECT  802.46 45.68 810.82 72.14 ;
     RECT  242.3 76.76 242.5 77.18 ;
     RECT  240.38 77.18 242.5 77.6 ;
     RECT  273.02 77.6 273.22 78.02 ;
     RECT  268.7 78.02 273.22 78.44 ;
     RECT  285.02 77.18 285.22 78.44 ;
     RECT  315.26 73.4 315.46 78.44 ;
     RECT  325.34 70.88 590.5 78.44 ;
     RECT  237.5 77.6 250.18 80.96 ;
     RECT  268.7 78.44 285.22 80.96 ;
     RECT  315.26 78.44 590.5 80.96 ;
     RECT  268.7 80.96 287.62 81.38 ;
     RECT  621.02 80.96 621.22 81.38 ;
     RECT  621.02 81.38 629.38 81.8 ;
     RECT  231.26 80.96 252.1 82.22 ;
     RECT  268.7 81.38 289.06 82.22 ;
     RECT  620.54 81.8 629.38 83.06 ;
     RECT  315.26 80.96 594.82 84.32 ;
     RECT  614.3 83.06 629.38 84.32 ;
     RECT  315.26 84.32 595.78 85.16 ;
     RECT  613.34 84.32 630.34 85.16 ;
     RECT  302.78 84.74 302.98 85.58 ;
     RECT  315.26 85.16 630.82 85.58 ;
     RECT  231.26 82.22 289.06 86.42 ;
     RECT  302.78 85.58 630.82 86.42 ;
     RECT  231.26 86.42 630.82 88.52 ;
     RECT  228.38 88.52 630.82 88.94 ;
     RECT  223.58 88.94 630.82 91.46 ;
     RECT  222.14 91.46 630.82 96.08 ;
     RECT  222.14 96.08 633.7 100.7 ;
     RECT  222.14 100.7 637.06 101.12 ;
     RECT  218.3 101.12 637.06 103.64 ;
     RECT  773.66 91.04 773.86 103.64 ;
     RECT  211.58 103.64 637.06 108.26 ;
     RECT  802.46 72.14 813.22 108.68 ;
     RECT  210.14 108.26 637.06 111.2 ;
     RECT  210.14 111.2 641.38 114.56 ;
     RECT  210.14 114.56 643.3 114.98 ;
     RECT  209.18 114.98 643.3 115.4 ;
     RECT  205.82 115.4 643.3 120.02 ;
     RECT  201.02 120.02 643.3 122.96 ;
     RECT  721.82 78.86 722.02 126.74 ;
     RECT  201.02 122.96 647.14 130.52 ;
     RECT  195.74 130.52 647.14 130.94 ;
     RECT  187.1 130.94 647.14 136.4 ;
     RECT  175.58 133.88 175.78 136.82 ;
     RECT  175.58 136.82 176.26 137.66 ;
     RECT  167.9 137.66 176.26 138.08 ;
     RECT  155.42 138.08 176.26 138.5 ;
     RECT  187.1 136.4 656.74 138.5 ;
     RECT  139.58 141.44 141.7 142.7 ;
     RECT  139.1 142.7 141.7 143.96 ;
     RECT  155.42 138.5 656.74 143.96 ;
     RECT  139.1 143.96 656.74 144.8 ;
     RECT  100.7 145.22 100.9 145.64 ;
     RECT  97.82 145.64 122.5 146.48 ;
     RECT  136.22 144.8 656.74 146.48 ;
     RECT  97.82 146.48 656.74 149 ;
     RECT  97.82 149 664.42 149.42 ;
     RECT  96.38 149.42 664.42 152.98 ;
     RECT  96.38 152.98 100.9 153.2 ;
     RECT  79.58 153.62 79.78 156.56 ;
     RECT  76.7 156.56 79.78 157.82 ;
     RECT  76.7 157.82 84.1 158.66 ;
     RECT  93.98 153.2 100.9 158.66 ;
     RECT  111.26 152.98 664.42 160.76 ;
     RECT  740.06 160.34 740.26 161.18 ;
     RECT  111.26 160.76 671.14 161.6 ;
     RECT  684.38 160.76 684.58 161.6 ;
     RECT  734.3 161.18 740.26 162.02 ;
     RECT  76.7 158.66 100.9 163.28 ;
     RECT  111.26 161.6 673.06 163.28 ;
     RECT  76.7 163.28 673.06 163.7 ;
     RECT  683.9 161.6 684.58 163.7 ;
     RECT  695.9 101.12 696.1 163.7 ;
     RECT  55.1 163.7 55.3 164.12 ;
     RECT  55.1 164.12 64.9 164.54 ;
     RECT  76.7 163.7 696.1 164.54 ;
     RECT  734.3 162.02 742.66 164.54 ;
     RECT  766.46 103.64 773.86 165.5 ;
     RECT  75.74 164.54 696.1 167.68 ;
     RECT  54.62 164.54 64.9 167.9 ;
     RECT  39.26 167.9 39.46 168.32 ;
     RECT  54.62 167.9 65.86 168.32 ;
     RECT  39.26 168.32 65.86 169.16 ;
     RECT  39.26 169.16 69.22 173.56 ;
     RECT  79.1 167.68 696.1 176.3 ;
     RECT  716.06 126.74 722.02 178.82 ;
     RECT  39.26 173.56 66.82 179.24 ;
     RECT  734.3 164.54 745.06 179.24 ;
     RECT  79.1 176.3 697.06 179.66 ;
     RECT  712.22 178.82 722.02 179.66 ;
     RECT  734.3 179.24 751.3 179.66 ;
     RECT  77.66 179.66 697.06 180.5 ;
     RECT  709.34 179.66 722.02 180.5 ;
     RECT  33.02 179.24 66.82 183.44 ;
     RECT  77.66 180.5 722.02 183.44 ;
     RECT  734.3 179.66 755.14 183.44 ;
     RECT  18.62 179.66 18.82 183.86 ;
     RECT  33.02 183.44 755.14 183.86 ;
     RECT  765.98 165.5 773.86 183.86 ;
     RECT  788.06 106.16 788.26 183.86 ;
     RECT  33.02 183.86 773.86 186.8 ;
     RECT  783.74 183.86 788.26 186.8 ;
     RECT  33.02 186.8 788.74 191.2 ;
     RECT  37.34 191.2 788.74 192.88 ;
     RECT  802.46 108.68 813.7 201.92 ;
     RECT  37.34 192.88 788.26 202.12 ;
     RECT  37.34 202.12 130.18 206.74 ;
     RECT  39.26 206.74 130.18 213.68 ;
     RECT  142.94 202.12 788.26 213.68 ;
     RECT  802.46 201.92 814.18 213.88 ;
     RECT  10.46 183.86 18.82 223.76 ;
     RECT  39.26 213.68 788.26 225.02 ;
     RECT  810.14 213.88 814.18 232.36 ;
     RECT  35.9 225.02 788.26 235.94 ;
     RECT  35.9 235.94 788.74 236.56 ;
     RECT  810.62 232.36 814.18 242.44 ;
     RECT  35.9 236.56 788.26 244.12 ;
     RECT  4.7 223.76 18.82 244.76 ;
     RECT  811.1 242.44 814.18 246.64 ;
     RECT  811.1 246.64 813.7 248.32 ;
     RECT  35.9 244.12 787.3 251.48 ;
     RECT  35.42 251.48 787.3 251.68 ;
     RECT  811.1 248.32 813.22 252.74 ;
     RECT  806.3 252.74 813.22 255.04 ;
     RECT  35.42 251.68 784.9 257.14 ;
     RECT  35.42 257.14 783.46 266.8 ;
     RECT  4.7 244.76 25.06 269.12 ;
     RECT  37.34 266.8 783.46 287.6 ;
     RECT  37.34 287.6 788.74 289.48 ;
     RECT  811.1 255.04 813.22 298.94 ;
     RECT  38.3 289.48 788.74 300.62 ;
     RECT  36.86 300.62 788.74 302.3 ;
     RECT  36.86 302.3 791.62 303.34 ;
     RECT  0.86 269.12 25.06 303.98 ;
     RECT  806.3 298.94 813.22 305.44 ;
     RECT  38.3 303.34 791.62 316.7 ;
     RECT  36.38 316.7 791.62 327.28 ;
     RECT  0.86 303.98 25.54 336.74 ;
     RECT  36.38 327.28 783.46 336.74 ;
     RECT  0.86 336.74 783.46 338 ;
     RECT  0.86 338 785.86 342.4 ;
     RECT  811.1 305.44 813.22 345.76 ;
     RECT  0.86 342.4 783.46 346.6 ;
     RECT  811.1 345.76 811.3 350.8 ;
     RECT  43.1 346.6 783.46 360.68 ;
     RECT  0.86 346.6 32.74 366.56 ;
     RECT  43.1 360.68 783.94 366.56 ;
     RECT  0.86 366.56 783.94 367.6 ;
     RECT  43.1 367.6 783.94 383.36 ;
     RECT  795.26 373.7 795.46 383.36 ;
     RECT  807.26 356.9 807.46 383.56 ;
     RECT  43.1 383.36 795.46 387.76 ;
     RECT  43.58 387.76 783.94 394.06 ;
     RECT  50.3 394.06 783.94 398.68 ;
     RECT  53.66 398.68 783.94 399.52 ;
     RECT  54.62 399.52 783.94 406.04 ;
     RECT  54.62 406.04 785.38 408.98 ;
     RECT  795.26 387.76 795.46 408.98 ;
     RECT  806.3 420.32 806.5 421.36 ;
     RECT  54.62 408.98 795.46 423.68 ;
     RECT  0.86 367.6 32.74 426.2 ;
     RECT  52.22 423.68 795.46 429.98 ;
     RECT  50.78 429.98 795.46 431.24 ;
     RECT  0.86 426.2 35.62 436.28 ;
     RECT  50.78 431.24 802.66 436.28 ;
     RECT  0.86 436.28 802.66 456.44 ;
     RECT  0.86 456.44 810.82 499.9 ;
     RECT  0.86 499.9 802.66 507.04 ;
     RECT  0.86 507.04 799.3 521.12 ;
     RECT  0.86 521.12 802.66 526.16 ;
     RECT  0.86 526.16 806.5 526.78 ;
     RECT  795.26 526.78 806.5 537.28 ;
     RECT  795.26 537.28 802.66 544.84 ;
     RECT  0.86 526.78 785.38 549.26 ;
     RECT  0.38 549.26 785.38 565.42 ;
     RECT  0.38 565.42 43.78 575.08 ;
     RECT  53.66 565.42 785.38 577.4 ;
     RECT  0.38 575.08 12.58 577.6 ;
     RECT  24.86 575.08 43.78 579.28 ;
     RECT  41.18 579.28 43.78 580.34 ;
     RECT  53.66 577.4 786.34 580.34 ;
     RECT  41.18 580.34 786.34 582.44 ;
     RECT  802.46 544.84 802.66 587.48 ;
     RECT  0.38 577.6 11.62 590.2 ;
     RECT  24.86 579.28 29.38 592.72 ;
     RECT  0.38 590.2 11.14 594.4 ;
     RECT  41.18 582.44 792.58 594.82 ;
     RECT  44.06 594.82 792.58 598.18 ;
     RECT  0.86 594.4 11.14 600.28 ;
     RECT  47.42 598.18 792.58 600.7 ;
     RECT  0.86 600.28 7.3 602.8 ;
     RECT  47.42 600.7 730.66 602.8 ;
     RECT  802.46 587.48 806.5 602.8 ;
     RECT  47.42 602.8 729.7 603.22 ;
     RECT  47.42 603.22 722.5 610.78 ;
     RECT  741.98 600.7 792.58 611.62 ;
     RECT  806.3 602.8 806.5 612.04 ;
     RECT  741.98 611.62 782.98 613.52 ;
     RECT  0.86 602.8 6.34 617.3 ;
     RECT  0.86 617.3 7.3 617.92 ;
     RECT  48.86 610.78 722.5 618.34 ;
     RECT  740.54 613.52 782.98 618.34 ;
     RECT  740.54 618.34 780.1 619.18 ;
     RECT  0.86 617.92 6.34 619.4 ;
     RECT  48.86 618.34 477.22 620.86 ;
     RECT  751.58 619.18 780.1 620.86 ;
     RECT  740.54 619.18 741.22 621.7 ;
     RECT  754.94 620.86 780.1 621.7 ;
     RECT  489.5 618.34 722.5 621.92 ;
     RECT  741.02 621.7 741.22 622.12 ;
     RECT  756.38 621.7 756.58 622.12 ;
     RECT  489.5 621.92 723.94 622.54 ;
     RECT  696.38 622.54 723.94 622.76 ;
     RECT  489.5 622.54 685.54 622.96 ;
     RECT  771.26 621.7 780.1 625.06 ;
     RECT  775.58 625.06 780.1 625.9 ;
     RECT  489.5 622.96 685.06 629.06 ;
     RECT  488.06 629.06 685.06 629.48 ;
     RECT  28.7 592.72 29.38 629.68 ;
     RECT  0.38 619.4 6.34 632.42 ;
     RECT  487.1 629.48 685.06 632.84 ;
     RECT  696.38 622.76 725.38 632.84 ;
     RECT  0.38 632.42 7.3 633.04 ;
     RECT  487.1 632.84 726.34 633.88 ;
     RECT  779.9 625.9 780.1 633.88 ;
     RECT  48.86 620.86 469.06 635.98 ;
     RECT  487.1 633.88 725.38 637.04 ;
     RECT  483.26 637.04 725.38 637.24 ;
     RECT  483.26 637.24 723.94 643.96 ;
     RECT  48.86 635.98 468.58 644.38 ;
     RECT  48.86 644.38 311.62 644.8 ;
     RECT  0.38 633.04 6.34 647.96 ;
     RECT  486.62 643.96 723.94 649 ;
     RECT  486.62 649 722.02 649.84 ;
     RECT  50.3 644.8 311.62 651.1 ;
     RECT  486.62 649.84 721.54 651.1 ;
     RECT  321.98 644.38 468.1 651.52 ;
     RECT  489.5 651.1 721.54 652.36 ;
     RECT  50.78 651.1 311.62 654.46 ;
     RECT  489.5 652.36 719.14 654.88 ;
     RECT  321.98 651.52 466.18 655.52 ;
     RECT  321.5 655.52 466.18 656.98 ;
     RECT  489.5 654.88 716.26 658.66 ;
     RECT  51.26 654.46 311.62 659.72 ;
     RECT  321.5 656.98 462.34 659.72 ;
     RECT  490.46 658.66 716.26 660.76 ;
     RECT  0.38 647.96 7.3 663.7 ;
     RECT  51.26 659.72 462.34 667.48 ;
     RECT  55.58 667.48 462.34 667.9 ;
     RECT  57.5 667.9 462.34 670 ;
     RECT  490.46 660.76 713.38 670.64 ;
     RECT  489.98 670.64 713.38 671.48 ;
     RECT  57.5 670 451.78 671.68 ;
     RECT  462.14 670 462.34 671.68 ;
     RECT  489.98 671.48 717.22 671.9 ;
     RECT  57.5 671.68 445.54 674.2 ;
     RECT  489.98 671.9 718.66 674.84 ;
     RECT  63.74 674.2 445.54 675.04 ;
     RECT  65.18 675.04 445.54 676.3 ;
     RECT  65.18 676.3 441.22 676.72 ;
     RECT  487.1 674.84 718.66 676.72 ;
     RECT  65.66 676.72 441.22 677.56 ;
     RECT  489.5 676.72 718.66 677.98 ;
     RECT  65.66 677.56 439.78 680.08 ;
     RECT  489.98 677.98 718.66 682.4 ;
     RECT  489.98 682.4 719.14 685.76 ;
     RECT  489.98 685.76 719.62 686.8 ;
     RECT  65.66 680.08 419.62 688.7 ;
     RECT  65.18 688.7 419.62 690.16 ;
     RECT  28.7 629.68 28.9 691.42 ;
     RECT  490.46 686.8 719.62 692.68 ;
     RECT  259.58 690.16 419.62 693.1 ;
     RECT  66.62 690.16 249.7 693.94 ;
     RECT  248.06 693.94 249.7 694.36 ;
     RECT  261.02 693.1 419.62 694.36 ;
     RECT  66.62 693.94 238.18 696.46 ;
     RECT  66.62 696.46 230.5 697.3 ;
     RECT  249.5 694.36 249.7 697.3 ;
     RECT  490.46 692.68 718.66 697.72 ;
     RECT  432.86 680.08 439.78 698.98 ;
     RECT  432.86 698.98 433.06 699.4 ;
     RECT  66.62 697.3 230.02 700.46 ;
     RECT  66.14 700.46 230.02 701.08 ;
     RECT  263.9 694.36 419.62 701.08 ;
     RECT  72.38 701.08 220.9 701.5 ;
     RECT  74.78 701.5 220.9 704.02 ;
     RECT  693.98 697.72 718.66 705.08 ;
     RECT  267.26 701.08 419.62 705.7 ;
     RECT  490.46 697.72 683.14 705.7 ;
     RECT  74.78 704.02 216.58 707.8 ;
     RECT  494.3 705.7 683.14 707.8 ;
     RECT  74.78 707.8 212.74 708.64 ;
     RECT  693.98 705.08 719.14 710.12 ;
     RECT  83.42 708.64 212.74 711.58 ;
     RECT  499.1 707.8 683.14 712.64 ;
     RECT  693.5 710.12 719.14 712.64 ;
     RECT  83.42 711.58 212.26 712.84 ;
     RECT  83.42 712.84 211.78 715.36 ;
     RECT  270.14 705.7 419.62 715.36 ;
     RECT  95.9 715.36 211.78 715.78 ;
     RECT  83.42 715.36 83.62 716.2 ;
     RECT  97.82 715.78 211.78 716.2 ;
     RECT  103.58 716.2 211.78 716.62 ;
     RECT  499.1 712.64 719.14 716.84 ;
     RECT  499.1 716.84 720.1 717.04 ;
     RECT  108.86 716.62 211.78 717.46 ;
     RECT  108.86 717.46 211.3 717.88 ;
     RECT  199.58 717.88 211.3 719.14 ;
     RECT  201.5 719.14 211.3 719.98 ;
     RECT  270.62 715.36 419.62 719.98 ;
     RECT  499.1 717.04 719.62 719.98 ;
     RECT  108.86 717.88 189.7 720.4 ;
     RECT  499.1 719.98 718.66 720.62 ;
     RECT  172.7 720.4 189.7 720.82 ;
     RECT  201.5 719.98 205.54 721.24 ;
     RECT  173.18 720.82 189.7 722.08 ;
     RECT  0.38 663.7 6.34 723.34 ;
     RECT  202.94 721.24 205.54 723.34 ;
     RECT  271.1 719.98 419.62 723.34 ;
     RECT  108.86 720.4 162.82 723.76 ;
     RECT  205.34 723.34 205.54 723.76 ;
     RECT  498.14 720.62 718.66 723.76 ;
     RECT  130.94 723.76 161.86 724.18 ;
     RECT  275.9 723.34 419.62 725.02 ;
     RECT  108.86 723.76 117.7 726.7 ;
     RECT  173.18 722.08 189.22 726.7 ;
     RECT  136.22 724.18 145.54 727.12 ;
     RECT  501.02 723.76 718.66 727.12 ;
     RECT  112.22 726.7 113.86 727.54 ;
     RECT  142.94 727.12 143.14 727.54 ;
     RECT  275.9 725.02 277.54 727.54 ;
     RECT  290.78 725.02 419.62 727.54 ;
     RECT  112.22 727.54 113.38 727.96 ;
     RECT  173.18 726.7 183.46 727.96 ;
     RECT  275.9 727.54 276.1 727.96 ;
     RECT  290.78 727.54 413.38 727.96 ;
     RECT  501.02 727.12 713.38 727.96 ;
     RECT  112.22 727.96 112.42 728.38 ;
     RECT  181.34 727.96 181.54 728.8 ;
     RECT  502.94 727.96 713.38 728.8 ;
     RECT  502.94 728.8 712.42 730.48 ;
     RECT  290.78 727.96 410.98 730.9 ;
     RECT  290.78 730.9 404.74 731.32 ;
     RECT  290.78 731.32 403.78 731.74 ;
     RECT  290.78 731.74 394.66 732.16 ;
     RECT  504.38 730.48 711.46 732.16 ;
     RECT  290.78 732.16 381.7 734.26 ;
     RECT  312.38 734.26 381.7 735.1 ;
     RECT  394.46 732.16 394.66 735.1 ;
     RECT  312.38 735.1 364.9 735.52 ;
     RECT  381.5 735.1 381.7 735.52 ;
     RECT  359.9 735.52 360.1 736.36 ;
     RECT  508.7 732.16 711.46 738.04 ;
     RECT  290.78 734.26 302.02 738.46 ;
     RECT  344.54 735.52 346.66 738.46 ;
     RECT  510.14 738.04 711.46 738.46 ;
     RECT  301.82 738.46 302.02 738.88 ;
     RECT  315.26 735.52 334.66 738.88 ;
     RECT  344.54 738.46 346.18 738.88 ;
     RECT  317.66 738.88 334.66 739.3 ;
     RECT  326.3 739.3 334.66 739.72 ;
     RECT  1.34 723.34 6.34 741.5 ;
     RECT  510.14 738.46 709.06 750.22 ;
     RECT  512.54 750.22 709.06 750.64 ;
     RECT  0.86 741.5 6.34 756.52 ;
     RECT  6.14 756.52 6.34 761.56 ;
     RECT  513.02 750.64 709.06 761.56 ;
     RECT  290.78 738.46 290.98 764.5 ;
     RECT  513.5 761.56 709.06 764.5 ;
     RECT  516.38 764.5 709.06 765.76 ;
     RECT  519.26 765.76 709.06 766.18 ;
     RECT  522.62 766.18 709.06 768.28 ;
     RECT  522.62 768.28 707.14 768.7 ;
     RECT  529.82 768.7 707.14 769.12 ;
     RECT  531.74 769.12 707.14 775.42 ;
     RECT  531.74 775.42 706.18 775.84 ;
     RECT  532.22 775.84 706.18 776.26 ;
     RECT  532.22 776.26 703.78 776.68 ;
     RECT  537.98 776.68 703.3 777.1 ;
     RECT  540.38 777.1 703.3 777.52 ;
     RECT  540.38 777.52 686.02 778.78 ;
     RECT  668.54 778.78 686.02 779.62 ;
     RECT  540.38 778.78 658.66 780.04 ;
     RECT  668.54 779.62 685.06 780.46 ;
     RECT  540.38 780.04 657.7 780.88 ;
     RECT  668.54 780.46 683.62 780.88 ;
     RECT  672.38 780.88 683.62 781.72 ;
     RECT  680.54 781.72 683.62 783.4 ;
     RECT  680.54 783.4 682.66 783.82 ;
     RECT  682.46 783.82 682.66 784.24 ;
     RECT  541.82 780.88 656.26 787.18 ;
     RECT  542.3 787.18 656.26 788.44 ;
     RECT  546.62 788.44 656.26 790.76 ;
     RECT  546.62 790.76 657.7 790.96 ;
     RECT  546.62 790.96 657.22 794.74 ;
     RECT  550.94 794.74 657.22 796 ;
     RECT  559.58 796 657.22 798.1 ;
     RECT  571.58 798.1 657.22 803.14 ;
     RECT  572.06 803.14 657.22 803.36 ;
     RECT  572.06 803.36 657.7 803.56 ;
     RECT  573.98 803.56 657.7 803.98 ;
     RECT  576.38 803.98 657.7 804.4 ;
     RECT  627.74 804.4 657.7 810.92 ;
     RECT  579.74 804.4 617.38 814.28 ;
     RECT  627.74 810.92 661.06 814.28 ;
     RECT  579.74 814.28 661.06 817.42 ;
     RECT  579.74 817.42 660.58 818.68 ;
     RECT  579.74 818.68 636.1 819.52 ;
     RECT  647.9 818.68 660.58 821.2 ;
     RECT  648.38 821.2 660.58 821.62 ;
     RECT  651.74 821.62 660.58 822.04 ;
     RECT  651.74 822.04 657.22 822.88 ;
     RECT  657.02 822.88 657.22 823.3 ;
     RECT  579.74 819.52 633.7 824.98 ;
     RECT  592.22 824.98 633.7 825.82 ;
     RECT  593.18 825.82 633.7 828.76 ;
     RECT  596.06 828.76 633.7 829.18 ;
     RECT  597.02 829.18 633.7 830.02 ;
     RECT  559.58 798.1 559.78 834.64 ;
     RECT  579.74 824.98 579.94 835.9 ;
     RECT  597.98 830.02 633.7 836.54 ;
     RECT  597.98 836.54 637.06 836.74 ;
     RECT  599.42 836.74 637.06 837.16 ;
     RECT  612.86 837.16 629.38 840.52 ;
     RECT  615.26 840.52 629.38 840.94 ;
     RECT  616.7 840.94 629.38 841.36 ;
     RECT  619.58 841.36 629.38 841.78 ;
     RECT  623.42 841.78 629.38 842.2 ;
     RECT  626.78 842.2 629.38 843.88 ;
     RECT  629.18 843.88 629.38 844.72 ;
    LAYER Metal4 ;
     RECT  0.38 273.74 0.86 273.94 ;
     RECT  0.38 763.88 1.06 764.08 ;
     RECT  0.38 549.26 1.34 549.46 ;
     RECT  0.38 619.4 1.34 619.6 ;
     RECT  0.38 690.38 1.34 698.56 ;
     RECT  1.34 548.84 1.54 549.88 ;
     RECT  0.86 269.12 1.82 273.94 ;
     RECT  0.86 288.86 1.82 289.06 ;
     RECT  0.38 594.2 1.82 595.24 ;
     RECT  1.82 592.1 2.02 595.24 ;
     RECT  1.34 619.4 2.02 628 ;
     RECT  1.82 642.92 2.02 644.8 ;
     RECT  1.34 299.36 2.3 299.56 ;
     RECT  1.34 321.62 2.3 321.82 ;
     RECT  1.54 549.68 2.5 549.88 ;
     RECT  2.02 627.8 2.98 628 ;
     RECT  1.82 269.12 3.26 289.06 ;
     RECT  2.3 299.36 3.26 305.02 ;
     RECT  1.34 689.54 3.26 698.56 ;
     RECT  0.38 400.58 3.46 400.78 ;
     RECT  3.26 678.2 3.46 701.08 ;
     RECT  3.26 269.12 3.74 305.02 ;
     RECT  2.3 321.62 4.22 322.24 ;
     RECT  1.82 231.32 4.7 231.52 ;
     RECT  3.74 495.5 5.38 495.7 ;
     RECT  3.74 514.82 5.38 515.02 ;
     RECT  2.02 594.2 7.1 595.24 ;
     RECT  3.26 183.02 10.46 183.22 ;
     RECT  2.78 254 11.42 254.2 ;
     RECT  11.42 248.12 12.38 254.2 ;
     RECT  4.22 321.62 12.86 326.86 ;
     RECT  9.5 356.06 13.34 356.26 ;
     RECT  7.1 441.32 13.82 446.56 ;
     RECT  7.1 393.44 17.66 393.64 ;
     RECT  4.7 223.76 18.14 231.52 ;
     RECT  10.46 183.02 18.62 184.06 ;
     RECT  9.98 367.82 19.58 368.02 ;
     RECT  19.1 377.9 19.58 378.1 ;
     RECT  17.66 392.18 20.06 393.64 ;
     RECT  20.06 390.5 20.54 393.64 ;
     RECT  12.38 246.44 24.86 254.2 ;
     RECT  13.34 352.28 25.82 356.26 ;
     RECT  19.58 367.82 26.78 378.1 ;
     RECT  20.54 388.4 26.78 393.64 ;
     RECT  29.18 523.64 29.66 527.2 ;
     RECT  3.26 552.2 31.1 552.4 ;
     RECT  11.9 337.58 32.06 337.78 ;
     RECT  7.1 632.42 32.06 635.56 ;
     RECT  25.82 352.28 32.54 356.68 ;
     RECT  25.34 480.8 33.02 481 ;
     RECT  3.26 504.32 33.02 504.52 ;
     RECT  18.62 464 34.46 464.2 ;
     RECT  33.02 474.08 34.46 481 ;
     RECT  33.02 504.32 34.46 512.08 ;
     RECT  34.46 497.6 34.94 512.08 ;
     RECT  29.66 522.8 34.94 527.2 ;
     RECT  3.74 269.12 35.9 311.74 ;
     RECT  34.94 497.6 35.9 527.2 ;
     RECT  34.46 464 36.86 481 ;
     RECT  35.9 493.82 36.86 527.2 ;
     RECT  31.1 552.2 38.3 554.08 ;
     RECT  38.3 546.32 38.98 554.08 ;
     RECT  37.34 537.5 39.26 537.7 ;
     RECT  38.98 546.32 39.26 552.4 ;
     RECT  35.9 266.18 39.94 311.74 ;
     RECT  36.86 493.4 40.42 527.2 ;
     RECT  40.42 516.08 40.7 527.2 ;
     RECT  39.26 537.5 40.7 552.4 ;
     RECT  40.42 493.4 45.22 504.94 ;
     RECT  45.22 493.4 45.5 494.86 ;
     RECT  40.7 516.08 45.7 552.4 ;
     RECT  39.26 205.7 48.58 205.9 ;
     RECT  45.7 516.5 49.54 552.4 ;
     RECT  32.06 336.74 50.3 337.78 ;
     RECT  32.54 349.34 50.3 356.68 ;
     RECT  36.86 464 50.3 481.84 ;
     RECT  49.54 552.2 50.3 552.4 ;
     RECT  39.94 269.12 50.78 311.74 ;
     RECT  12.86 321.62 50.78 327.7 ;
     RECT  50.3 463.58 52.7 483.94 ;
     RECT  52.7 463.16 54.14 483.94 ;
     RECT  45.5 492.98 54.14 494.86 ;
     RECT  13.82 441.32 56.06 449.92 ;
     RECT  50.78 269.12 56.54 327.7 ;
     RECT  50.3 336.74 56.54 356.68 ;
     RECT  50.78 429.98 56.54 430.18 ;
     RECT  56.54 269.12 57.22 356.68 ;
     RECT  54.14 463.16 57.22 494.86 ;
     RECT  45.22 504.32 57.98 504.94 ;
     RECT  49.54 516.5 57.98 539.38 ;
     RECT  18.14 220.82 58.46 231.52 ;
     RECT  57.98 504.32 59.14 539.38 ;
     RECT  50.3 198.14 59.42 198.34 ;
     RECT  58.46 220.82 59.42 235.72 ;
     RECT  7.1 594.2 59.42 602.38 ;
     RECT  32.06 628.22 59.9 635.56 ;
     RECT  59.42 198.14 60.1 198.76 ;
     RECT  57.22 463.16 60.38 493.18 ;
     RECT  59.42 218.72 60.58 235.72 ;
     RECT  7.1 612.68 61.34 617.5 ;
     RECT  59.9 628.22 61.34 637.66 ;
     RECT  7.1 648.38 61.34 668.32 ;
     RECT  57.22 321.62 62.3 356.68 ;
     RECT  26.78 367.82 62.3 393.64 ;
     RECT  7.1 584.96 62.3 585.16 ;
     RECT  7.1 406.04 64.22 408.76 ;
     RECT  50.3 552.2 64.42 553.66 ;
     RECT  61.34 612.68 64.7 617.92 ;
     RECT  61.34 628.22 64.7 668.32 ;
     RECT  62.3 321.62 64.9 393.64 ;
     RECT  59.14 504.32 64.9 538.54 ;
     RECT  59.42 594.2 65.18 602.8 ;
     RECT  64.7 612.68 65.18 668.32 ;
     RECT  60.38 462.74 65.38 493.18 ;
     RECT  57.22 269.12 65.66 311.74 ;
     RECT  64.9 321.62 65.66 356.68 ;
     RECT  64.22 402.26 65.86 408.76 ;
     RECT  65.38 479.96 65.86 493.18 ;
     RECT  65.18 594.2 65.86 668.32 ;
     RECT  62.3 579.5 66.14 585.16 ;
     RECT  65.86 594.2 66.14 617.5 ;
     RECT  3.46 700.88 66.14 701.08 ;
     RECT  65.66 269.12 66.82 356.68 ;
     RECT  66.14 579.5 66.82 617.5 ;
     RECT  66.82 269.12 67.1 311.74 ;
     RECT  7.1 569.84 67.1 570.04 ;
     RECT  66.82 579.5 67.1 602.8 ;
     RECT  60.58 218.72 67.58 231.52 ;
     RECT  56.06 440.9 68.54 449.92 ;
     RECT  65.38 462.74 68.54 470.5 ;
     RECT  60.1 198.56 69.22 198.76 ;
     RECT  67.1 569.84 69.22 602.8 ;
     RECT  69.22 569.84 69.98 602.38 ;
     RECT  69.98 564.8 70.18 602.38 ;
     RECT  64.9 504.32 70.46 534.76 ;
     RECT  70.18 564.8 71.14 585.16 ;
     RECT  68.54 440.9 71.62 470.5 ;
     RECT  68.54 553.88 71.9 554.08 ;
     RECT  71.14 564.8 71.9 570.04 ;
     RECT  66.14 700.46 72.38 701.08 ;
     RECT  64.9 367.82 72.86 393.64 ;
     RECT  70.46 500.96 73.54 534.76 ;
     RECT  56.54 429.56 73.82 430.18 ;
     RECT  71.62 459.8 73.82 470.5 ;
     RECT  65.86 479.96 73.82 489.82 ;
     RECT  65.86 628.22 74.3 668.32 ;
     RECT  3.46 678.2 74.3 691 ;
     RECT  72.86 367.82 74.5 395.74 ;
     RECT  67.1 266.6 75.26 311.74 ;
     RECT  66.82 321.62 75.26 356.68 ;
     RECT  73.82 459.8 75.26 489.82 ;
     RECT  73.54 500.96 75.26 529.3 ;
     RECT  71.9 553.88 77.18 570.04 ;
     RECT  75.26 459.8 77.86 529.3 ;
     RECT  74.3 628.22 77.86 691 ;
     RECT  75.74 538.76 78.82 538.96 ;
     RECT  72.38 700.46 78.82 701.5 ;
     RECT  74.78 417.38 79.1 417.58 ;
     RECT  70.18 594.2 79.1 602.38 ;
     RECT  67.58 216.62 80.54 231.52 ;
     RECT  24.86 244.76 80.54 254.2 ;
     RECT  77.86 628.22 80.74 637.66 ;
     RECT  18.62 179.66 81.02 184.06 ;
     RECT  78.82 700.88 81.02 701.5 ;
     RECT  80.54 216.62 82.18 254.2 ;
     RECT  77.86 529.1 82.18 529.3 ;
     RECT  65.86 406.04 82.46 408.76 ;
     RECT  79.1 417.38 82.46 418.42 ;
     RECT  73.82 429.14 82.94 430.18 ;
     RECT  71.62 440.9 82.94 449.92 ;
     RECT  57.02 164.12 83.9 164.32 ;
     RECT  75.26 266.6 84.58 356.68 ;
     RECT  82.46 406.04 85.34 418.42 ;
     RECT  82.94 429.14 85.34 449.92 ;
     RECT  77.86 459.8 85.34 518.8 ;
     RECT  79.1 594.2 86.02 602.8 ;
     RECT  74.5 367.82 88.22 393.64 ;
     RECT  85.34 402.26 88.22 418.42 ;
     RECT  88.22 367.82 88.42 418.42 ;
     RECT  77.86 648.38 88.7 691 ;
     RECT  81.02 700.88 89.38 708.64 ;
     RECT  88.42 367.82 89.86 396.16 ;
     RECT  85.82 198.56 90.62 198.76 ;
     RECT  84.58 269.12 90.62 356.68 ;
     RECT  89.86 367.82 90.62 393.64 ;
     RECT  77.18 549.68 91.3 570.04 ;
     RECT  91.3 549.68 92.54 558.28 ;
     RECT  90.62 269.12 92.74 393.64 ;
     RECT  66.82 612.68 93.5 617.5 ;
     RECT  80.74 628.22 93.5 635.56 ;
     RECT  85.34 429.14 93.7 518.8 ;
     RECT  93.7 429.14 93.98 430.18 ;
     RECT  88.42 406.04 96.1 417.58 ;
     RECT  93.7 440.9 96.1 518.8 ;
     RECT  93.5 612.68 96.86 635.56 ;
     RECT  88.7 645.02 96.86 691 ;
     RECT  92.74 269.12 97.06 356.68 ;
     RECT  90.62 198.56 97.34 202.12 ;
     RECT  83.9 163.7 97.54 164.32 ;
     RECT  93.98 426.62 97.54 430.18 ;
     RECT  92.54 542.54 97.54 558.28 ;
     RECT  97.34 195.62 98.02 202.12 ;
     RECT  97.54 542.54 98.98 554.08 ;
     RECT  97.54 163.7 99.46 163.9 ;
     RECT  98.02 195.62 100.42 201.7 ;
     RECT  81.02 179.66 100.7 184.9 ;
     RECT  89.38 700.88 100.7 701.08 ;
     RECT  100.42 199.4 100.9 201.7 ;
     RECT  97.06 269.12 100.9 337.78 ;
     RECT  96.1 406.04 100.9 415.06 ;
     RECT  86.02 594.2 101.18 602.38 ;
     RECT  96.86 612.68 101.18 691 ;
     RECT  82.18 218.72 101.66 254.2 ;
     RECT  92.74 367.82 103.58 393.64 ;
     RECT  97.54 429.14 103.58 430.18 ;
     RECT  96.1 440.9 103.58 508.3 ;
     RECT  100.9 199.4 105.7 201.28 ;
     RECT  103.58 429.14 105.98 508.3 ;
     RECT  71.14 584.96 105.98 585.16 ;
     RECT  101.18 594.2 105.98 691 ;
     RECT  100.7 700.88 105.98 702.34 ;
     RECT  105.98 425.36 106.94 508.3 ;
     RECT  96.1 518.6 106.94 518.8 ;
     RECT  101.66 217.04 107.42 254.2 ;
     RECT  106.94 419.06 107.42 518.8 ;
     RECT  105.98 584.96 109.82 691 ;
     RECT  100.9 269.12 111.26 311.74 ;
     RECT  100.9 321.62 111.26 327.7 ;
     RECT  109.82 584.96 111.94 691.42 ;
     RECT  100.7 179.66 112.22 190.78 ;
     RECT  91.3 569.84 113.18 570.04 ;
     RECT  111.74 153.62 113.38 153.82 ;
     RECT  111.26 269.12 114.14 327.7 ;
     RECT  114.14 265.76 114.34 327.7 ;
     RECT  112.22 179.66 115.1 196.24 ;
     RECT  113.18 569.84 115.3 571.72 ;
     RECT  107.42 213.26 116.26 254.2 ;
     RECT  103.58 365.3 116.54 393.64 ;
     RECT  100.9 406.04 116.54 408.76 ;
     RECT  116.26 213.26 117.22 233.2 ;
     RECT  116.54 365.3 117.22 408.76 ;
     RECT  97.06 349.34 117.5 356.68 ;
     RECT  105.98 700.88 118.94 708.64 ;
     RECT  117.5 349.34 121.54 357.1 ;
     RECT  98.98 547.58 121.82 554.08 ;
     RECT  111.94 584.96 121.82 617.5 ;
     RECT  115.1 172.94 122.5 198.34 ;
     RECT  111.94 628.22 125.38 691.42 ;
     RECT  117.22 213.26 126.82 231.52 ;
     RECT  126.82 216.2 127.1 231.52 ;
     RECT  116.26 244.76 127.1 254.2 ;
     RECT  117.22 367.82 129.7 408.76 ;
     RECT  121.82 583.7 129.7 617.5 ;
     RECT  121.54 349.34 129.98 356.68 ;
     RECT  129.7 367.82 129.98 395.32 ;
     RECT  107.42 419.06 130.46 519.64 ;
     RECT  127.1 216.2 130.66 254.2 ;
     RECT  129.7 584.12 131.14 617.5 ;
     RECT  129.98 349.34 132.58 395.32 ;
     RECT  118.94 700.88 132.58 716.2 ;
     RECT  122.5 178.82 132.86 198.34 ;
     RECT  121.82 547.58 132.86 557.86 ;
     RECT  127.1 169.16 133.34 169.36 ;
     RECT  132.86 178.82 133.34 198.76 ;
     RECT  133.34 169.16 133.54 198.76 ;
     RECT  132.86 547.58 133.82 561.64 ;
     RECT  115.3 571.1 133.82 571.72 ;
     RECT  130.46 419.06 134.5 523.42 ;
     RECT  132.58 700.88 134.5 715.78 ;
     RECT  133.54 171.68 136.42 198.76 ;
     RECT  136.42 196.04 136.9 198.76 ;
     RECT  129.7 404.78 138.34 408.76 ;
     RECT  138.34 405.62 139.58 408.76 ;
     RECT  134.5 419.06 139.58 519.64 ;
     RECT  132.58 367.82 139.78 395.32 ;
     RECT  133.82 547.58 139.78 571.72 ;
     RECT  131.14 584.96 140.54 617.5 ;
     RECT  125.38 628.22 140.54 691 ;
     RECT  139.78 549.26 141.22 571.72 ;
     RECT  130.66 217.46 141.7 254.2 ;
     RECT  139.78 367.82 142.46 393.64 ;
     RECT  139.58 405.62 143.9 519.64 ;
     RECT  141.7 220.82 144.1 254.2 ;
     RECT  100.9 336.74 145.34 337.78 ;
     RECT  132.58 349.34 145.34 356.68 ;
     RECT  140.54 584.96 146.02 691 ;
     RECT  134.5 700.88 146.98 708.64 ;
     RECT  141.22 549.68 147.46 571.72 ;
     RECT  144.1 243.5 149.38 254.2 ;
     RECT  145.34 336.74 149.86 356.68 ;
     RECT  142.94 209.48 150.34 209.68 ;
     RECT  144.1 220.82 151.1 231.52 ;
     RECT  114.34 269.12 151.1 327.7 ;
     RECT  149.86 336.74 151.1 338.2 ;
     RECT  143.9 405.62 151.1 523.84 ;
     RECT  147.26 538.76 151.1 538.96 ;
     RECT  147.46 570.68 151.3 571.72 ;
     RECT  146.02 612.68 151.3 691 ;
     RECT  142.46 366.56 152.54 393.64 ;
     RECT  151.1 405.62 152.54 538.96 ;
     RECT  147.46 549.68 152.54 561.64 ;
     RECT  151.1 215.78 152.74 231.52 ;
     RECT  151.1 269.12 153.02 338.2 ;
     RECT  136.42 171.68 153.5 184.06 ;
     RECT  136.9 198.56 153.5 198.76 ;
     RECT  151.1 709.7 154.46 709.9 ;
     RECT  149.86 349.34 154.94 356.68 ;
     RECT  152.54 366.56 154.94 538.96 ;
     RECT  154.94 349.34 155.62 538.96 ;
     RECT  155.62 402.68 156.86 538.96 ;
     RECT  154.46 709.7 157.06 710.32 ;
     RECT  155.62 349.34 158.02 393.64 ;
     RECT  156.86 402.68 158.02 539.38 ;
     RECT  158.02 539.18 158.3 539.38 ;
     RECT  152.54 549.26 158.3 561.64 ;
     RECT  153.5 171.68 158.78 198.76 ;
     RECT  158.3 539.18 158.98 561.64 ;
     RECT  153.02 265.76 160.22 338.2 ;
     RECT  160.22 264.92 160.9 338.2 ;
     RECT  157.06 710.12 161.86 710.32 ;
     RECT  158.3 719.78 161.86 719.98 ;
     RECT  152.74 220.82 162.14 231.52 ;
     RECT  162.14 220.4 163.1 231.52 ;
     RECT  158.78 171.68 163.78 202.96 ;
     RECT  146.02 584.96 164.06 602.38 ;
     RECT  151.3 612.68 164.06 668.32 ;
     RECT  163.78 179.66 164.26 202.96 ;
     RECT  151.3 677.78 165.02 691 ;
     RECT  146.98 700.88 165.02 701.08 ;
     RECT  163.1 216.2 165.5 231.52 ;
     RECT  149.38 244.76 165.5 254.2 ;
     RECT  151.3 571.1 165.5 571.72 ;
     RECT  164.06 584.96 165.5 668.32 ;
     RECT  158.98 539.18 165.7 553.66 ;
     RECT  165.5 216.2 166.94 254.2 ;
     RECT  158.02 367.82 166.94 393.64 ;
     RECT  165.02 165.38 167.14 165.58 ;
     RECT  166.94 366.98 167.14 393.64 ;
     RECT  167.14 367.4 167.62 393.64 ;
     RECT  160.9 268.28 168.86 338.2 ;
     RECT  158.02 349.34 168.86 356.68 ;
     RECT  167.62 367.82 168.86 393.64 ;
     RECT  158.02 402.68 168.86 529.72 ;
     RECT  168.86 367.82 169.06 529.72 ;
     RECT  164.26 198.56 170.02 202.96 ;
     RECT  168.86 268.28 170.98 356.68 ;
     RECT  165.7 549.26 171.26 553.66 ;
     RECT  165.7 539.18 172.22 539.38 ;
     RECT  170.98 268.28 172.42 337.78 ;
     RECT  165.5 569.84 174.34 668.32 ;
     RECT  174.34 569.84 175.78 576.34 ;
     RECT  166.94 213.68 177.7 254.2 ;
     RECT  169.06 367.82 177.7 408.76 ;
     RECT  177.7 214.52 177.98 254.2 ;
     RECT  164.26 179.66 178.46 184.06 ;
     RECT  177.98 214.52 178.66 260.5 ;
     RECT  178.66 240.14 179.62 260.5 ;
     RECT  179.62 240.14 180.1 254.2 ;
     RECT  170.98 349.34 180.38 356.68 ;
     RECT  172.42 269.12 181.34 337.78 ;
     RECT  180.38 349.34 181.34 357.1 ;
     RECT  178.46 179.66 182.3 187 ;
     RECT  170.02 198.56 182.3 200.86 ;
     RECT  172.22 538.76 182.3 539.38 ;
     RECT  171.26 549.26 182.3 557.44 ;
     RECT  181.34 269.12 182.5 357.1 ;
     RECT  182.3 538.76 182.98 557.44 ;
     RECT  182.5 349.34 183.94 357.1 ;
     RECT  182.98 545.48 183.94 557.44 ;
     RECT  183.94 545.48 184.42 554.08 ;
     RECT  182.5 269.12 185.38 338.2 ;
     RECT  177.7 405.62 186.34 408.76 ;
     RECT  182.3 198.56 187.1 201.7 ;
     RECT  174.34 584.96 187.58 668.32 ;
     RECT  180.1 244.76 188.54 254.2 ;
     RECT  175.78 569.84 189.02 573.4 ;
     RECT  169.34 138.08 189.5 138.28 ;
     RECT  189.5 138.08 189.7 139.96 ;
     RECT  185.38 269.12 189.7 337.78 ;
     RECT  189.02 569 189.98 573.4 ;
     RECT  188.54 242.24 191.14 254.2 ;
     RECT  187.58 584.96 191.14 669.16 ;
     RECT  184.42 549.26 191.62 554.08 ;
     RECT  189.98 563.54 192.1 573.4 ;
     RECT  189.7 321.62 192.58 337.78 ;
     RECT  187.1 198.14 192.86 201.7 ;
     RECT  191.62 549.68 193.82 554.08 ;
     RECT  192.1 563.54 193.82 570.46 ;
     RECT  194.3 152.78 195.26 152.98 ;
     RECT  191.14 244.34 195.26 254.2 ;
     RECT  189.7 269.12 195.26 311.74 ;
     RECT  194.3 169.16 195.46 169.36 ;
     RECT  195.26 244.34 196.42 311.74 ;
     RECT  169.06 419.06 196.42 529.72 ;
     RECT  195.26 152.78 197.38 155.08 ;
     RECT  193.82 549.68 197.38 570.46 ;
     RECT  191.14 584.96 197.66 668.32 ;
     RECT  197.38 152.78 197.86 152.98 ;
     RECT  197.38 549.68 197.86 570.04 ;
     RECT  196.42 422.42 198.34 529.72 ;
     RECT  197.66 580.34 198.34 668.32 ;
     RECT  192.58 336.74 199.58 337.78 ;
     RECT  198.34 422.42 199.78 523.84 ;
     RECT  200.06 534.56 201.02 534.76 ;
     RECT  196.42 266.6 201.22 311.74 ;
     RECT  201.02 534.56 201.22 538.12 ;
     RECT  196.42 244.34 201.5 254.2 ;
     RECT  189.7 139.76 201.7 139.96 ;
     RECT  192.86 198.14 201.7 202.54 ;
     RECT  198.34 584.96 201.7 668.32 ;
     RECT  201.7 198.14 202.18 200.86 ;
     RECT  165.02 677.78 202.46 701.08 ;
     RECT  201.7 647.54 203.14 668.32 ;
     RECT  201.22 268.28 203.42 311.74 ;
     RECT  202.46 677.78 204.38 704.86 ;
     RECT  183.94 349.34 204.86 356.68 ;
     RECT  177.7 367.82 204.86 393.64 ;
     RECT  197.86 549.68 204.86 559.96 ;
     RECT  202.18 198.56 205.06 200.86 ;
     RECT  203.42 268.28 205.34 312.58 ;
     RECT  192.58 321.62 205.34 327.7 ;
     RECT  204.86 547.58 206.5 559.96 ;
     RECT  205.34 268.28 206.98 327.7 ;
     RECT  204.86 349.34 207.74 393.64 ;
     RECT  206.5 549.68 208.7 559.96 ;
     RECT  197.86 569.84 208.7 570.04 ;
     RECT  199.58 336.74 209.18 338.2 ;
     RECT  207.74 348.5 209.18 393.64 ;
     RECT  201.5 243.08 209.38 254.2 ;
     RECT  206.98 268.28 209.66 311.74 ;
     RECT  209.18 336.74 209.66 393.64 ;
     RECT  178.66 214.52 209.86 231.52 ;
     RECT  209.38 244.34 210.14 254.2 ;
     RECT  201.7 584.96 210.62 602.38 ;
     RECT  204.38 677.78 210.82 709.06 ;
     RECT  210.82 700.88 211.3 709.06 ;
     RECT  205.06 200.66 211.78 200.86 ;
     RECT  209.66 336.74 212.06 394.06 ;
     RECT  199.78 424.94 212.06 523.84 ;
     RECT  203.14 648.38 212.06 668.32 ;
     RECT  208.7 549.68 212.26 570.04 ;
     RECT  209.66 265.76 212.74 311.74 ;
     RECT  210.62 584.96 212.74 603.22 ;
     RECT  211.3 700.88 212.74 704.86 ;
     RECT  212.06 336.74 213.22 395.32 ;
     RECT  210.14 244.34 213.7 255.04 ;
     RECT  212.26 558.5 214.18 570.04 ;
     RECT  213.22 336.74 214.66 338.2 ;
     RECT  206.98 321.2 216.38 327.7 ;
     RECT  214.66 336.74 216.38 337.78 ;
     RECT  213.22 348.5 216.86 395.32 ;
     RECT  216.86 348.5 217.82 397 ;
     RECT  186.34 406.04 217.82 408.76 ;
     RECT  215.9 146.48 218.5 146.68 ;
     RECT  212.06 418.64 218.5 523.84 ;
     RECT  213.7 244.76 218.78 255.04 ;
     RECT  212.74 269.12 219.26 311.74 ;
     RECT  216.38 321.2 219.26 337.78 ;
     RECT  212.06 644.18 219.46 668.32 ;
     RECT  209.86 220.82 220.22 231.52 ;
     RECT  217.82 348.5 222.34 408.76 ;
     RECT  182.3 179.66 223.1 187.42 ;
     RECT  201.7 612.68 224.54 635.56 ;
     RECT  214.18 569.84 225.02 570.04 ;
     RECT  214.18 558.5 225.22 559.96 ;
     RECT  212.74 584.96 225.5 602.38 ;
     RECT  218.78 244.76 225.98 257.98 ;
     RECT  219.26 269.12 225.98 337.78 ;
     RECT  220.22 220.82 227.42 233.62 ;
     RECT  225.98 244.76 228.38 337.78 ;
     RECT  222.34 348.5 228.38 356.68 ;
     RECT  223.1 175.46 228.86 187.42 ;
     RECT  228.86 171.68 229.54 187.42 ;
     RECT  201.22 537.92 229.82 538.12 ;
     RECT  229.82 537.92 230.02 541.48 ;
     RECT  221.18 209.48 230.3 209.68 ;
     RECT  218.5 421.16 230.98 523.84 ;
     RECT  229.54 171.68 232.22 184.06 ;
     RECT  225.5 584.96 232.9 602.8 ;
     RECT  232.22 164.96 233.38 184.06 ;
     RECT  225.02 569.84 233.38 572.56 ;
     RECT  222.34 367.82 233.66 408.76 ;
     RECT  227.42 220.82 234.82 236.14 ;
     RECT  233.66 366.14 234.82 408.76 ;
     RECT  230.3 205.7 235.58 209.68 ;
     RECT  234.82 220.82 235.58 234.88 ;
     RECT  232.9 584.96 235.58 602.38 ;
     RECT  219.46 648.38 236.54 668.32 ;
     RECT  230.78 112.04 237.02 112.24 ;
     RECT  230.3 145.64 237.5 145.84 ;
     RECT  224.54 612.68 237.7 637.66 ;
     RECT  235.58 205.7 238.18 234.88 ;
     RECT  238.18 205.7 238.66 205.9 ;
     RECT  237.02 112.04 239.14 115.18 ;
     RECT  239.14 112.04 239.42 112.24 ;
     RECT  230.98 421.58 239.42 523.84 ;
     RECT  239.42 110.36 239.62 112.24 ;
     RECT  233.38 171.68 239.62 184.06 ;
     RECT  239.62 112.04 240.1 112.24 ;
     RECT  237.5 144.8 240.86 146.68 ;
     RECT  240.86 144.8 242.5 150.88 ;
     RECT  234.82 367.82 242.78 408.76 ;
     RECT  239.42 421.16 242.78 523.84 ;
     RECT  236.54 647.12 242.98 668.32 ;
     RECT  225.22 559.76 243.26 559.96 ;
     RECT  237.5 160.76 244.9 160.96 ;
     RECT  238.18 216.2 246.14 234.88 ;
     RECT  228.38 244.76 246.14 356.68 ;
     RECT  230.02 541.28 247.1 541.48 ;
     RECT  243.26 553.46 247.1 559.96 ;
     RECT  246.14 216.2 247.58 356.68 ;
     RECT  242.78 367.82 247.58 523.84 ;
     RECT  247.1 541.28 248.74 559.96 ;
     RECT  247.58 367.82 249.02 530.98 ;
     RECT  248.74 541.28 249.02 541.48 ;
     RECT  247.58 212.42 249.7 356.68 ;
     RECT  233.38 569.84 249.98 570.04 ;
     RECT  249.7 212.42 250.18 259.24 ;
     RECT  249.02 367.82 250.18 541.48 ;
     RECT  250.18 541.28 251.14 541.48 ;
     RECT  249.98 569.84 251.14 575.5 ;
     RECT  250.18 212.42 251.62 255.04 ;
     RECT  250.18 367.82 251.62 532.66 ;
     RECT  248.74 553.46 251.62 559.96 ;
     RECT  242.5 145.64 251.9 150.88 ;
     RECT  235.58 584.54 251.9 602.38 ;
     RECT  210.82 677.78 251.9 691 ;
     RECT  212.74 700.88 251.9 701.08 ;
     RECT  251.62 559.76 252.1 559.96 ;
     RECT  242.98 648.38 252.86 668.32 ;
     RECT  251.9 677.78 252.86 701.08 ;
     RECT  251.9 580.34 254.02 602.8 ;
     RECT  249.7 269.12 256.42 356.68 ;
     RECT  256.42 348.5 258.14 356.68 ;
     RECT  256.42 269.12 259.1 337.78 ;
     RECT  251.62 212.42 259.58 254.2 ;
     RECT  258.14 348.5 259.58 359.2 ;
     RECT  251.62 367.82 259.58 530.98 ;
     RECT  259.58 348.5 259.78 530.98 ;
     RECT  239.62 179.66 260.06 184.06 ;
     RECT  259.78 348.5 261.22 523.42 ;
     RECT  259.58 209.48 262.94 254.2 ;
     RECT  259.1 262.82 262.94 337.78 ;
     RECT  251.9 165.38 263.14 165.58 ;
     RECT  251.9 145.64 263.62 156.76 ;
     RECT  252.86 648.38 264.38 701.08 ;
     RECT  264.38 647.96 264.58 701.08 ;
     RECT  258.14 197.72 264.86 197.92 ;
     RECT  262.94 209.48 264.86 337.78 ;
     RECT  263.62 145.64 265.82 151.72 ;
     RECT  251.14 569.84 265.82 570.04 ;
     RECT  265.82 561.86 266.78 570.04 ;
     RECT  265.82 143.96 266.98 151.72 ;
     RECT  260.06 179.66 267.26 186.58 ;
     RECT  264.86 197.72 267.46 337.78 ;
     RECT  264.58 647.96 268.9 668.32 ;
     RECT  254.02 584.12 269.18 602.8 ;
     RECT  237.7 612.68 269.66 635.56 ;
     RECT  268.9 647.96 269.66 656.14 ;
     RECT  267.46 209.9 270.14 337.78 ;
     RECT  261.22 348.5 270.14 522.58 ;
     RECT  270.14 209.9 270.34 522.58 ;
     RECT  260.54 130.1 272.06 130.3 ;
     RECT  266.98 143.96 272.06 149.2 ;
     RECT  272.06 130.1 272.74 149.2 ;
     RECT  270.34 367.4 272.74 522.58 ;
     RECT  272.74 136.4 273.7 149.2 ;
     RECT  264.58 678.2 273.98 701.08 ;
     RECT  271.58 716.42 273.98 716.62 ;
     RECT  270.34 209.9 274.18 357.94 ;
     RECT  268.9 668.12 274.18 668.32 ;
     RECT  273.7 143.96 274.66 149.2 ;
     RECT  267.46 197.72 274.94 197.92 ;
     RECT  266.78 561.02 274.94 570.04 ;
     RECT  269.18 582.44 274.94 602.8 ;
     RECT  274.18 209.9 276.58 356.68 ;
     RECT  274.94 561.02 276.58 602.8 ;
     RECT  276.58 561.02 278.5 561.22 ;
     RECT  274.94 195.2 279.26 197.92 ;
     RECT  269.66 612.68 279.26 656.14 ;
     RECT  269.66 92.3 281.38 92.5 ;
     RECT  267.26 176.72 281.66 186.58 ;
     RECT  279.26 195.2 281.66 202.96 ;
     RECT  276.58 212.42 282.34 356.68 ;
     RECT  279.26 612.68 282.34 662.44 ;
     RECT  273.02 107.84 283.3 108.04 ;
     RECT  276.58 569.84 283.58 602.8 ;
     RECT  282.34 612.68 283.58 656.14 ;
     RECT  281.66 176.72 283.78 202.96 ;
     RECT  273.98 678.2 284.06 716.62 ;
     RECT  284.06 671.06 284.74 716.62 ;
     RECT  283.1 164.54 285.22 164.74 ;
     RECT  283.78 179.66 286.46 202.96 ;
     RECT  282.34 212.42 286.46 257.14 ;
     RECT  284.74 671.06 286.46 716.2 ;
     RECT  286.46 179.66 286.66 257.14 ;
     RECT  286.46 666.86 286.66 716.2 ;
     RECT  283.58 569.84 288.1 656.14 ;
     RECT  288.1 569.84 288.38 602.38 ;
     RECT  286.66 666.86 290.02 712.42 ;
     RECT  286.66 197.72 290.5 257.14 ;
     RECT  288.38 569 292.42 602.38 ;
     RECT  290.02 670.22 292.42 712.42 ;
     RECT  274.66 145.22 292.9 149.2 ;
     RECT  292.42 670.22 292.9 708.64 ;
     RECT  272.74 367.4 293.18 408.76 ;
     RECT  282.34 266.18 293.38 356.68 ;
     RECT  290.5 202.76 294.34 257.14 ;
     RECT  293.18 365.72 294.34 408.76 ;
     RECT  292.42 569 296.54 585.16 ;
     RECT  292.9 145.22 297.22 145.42 ;
     RECT  296.54 563.54 298.66 585.16 ;
     RECT  286.94 101.12 299.14 101.32 ;
     RECT  293.38 266.18 302.02 337.78 ;
     RECT  272.74 418.22 302.02 522.58 ;
     RECT  292.9 670.22 302.02 701.08 ;
     RECT  294.34 207.8 302.3 257.14 ;
     RECT  302.02 266.18 302.3 311.74 ;
     RECT  302.02 420.74 302.3 522.58 ;
     RECT  283.58 548.84 302.3 549.04 ;
     RECT  302.02 670.22 302.3 690.16 ;
     RECT  302.3 207.8 302.5 311.74 ;
     RECT  302.02 321.62 302.5 337.78 ;
     RECT  302.3 548.84 302.5 554.5 ;
     RECT  288.1 612.68 302.5 656.14 ;
     RECT  302.02 699.2 302.5 701.08 ;
     RECT  302.3 420.74 302.98 524.26 ;
     RECT  302.5 548.84 302.98 554.08 ;
     RECT  302.5 336.74 304.7 337.78 ;
     RECT  293.38 348.5 304.7 356.68 ;
     RECT  302.3 539.18 305.18 539.38 ;
     RECT  302.98 548.84 305.18 549.04 ;
     RECT  302.5 648.38 306.14 656.14 ;
     RECT  302.3 668.54 306.14 690.16 ;
     RECT  298.66 569 307.1 585.16 ;
     RECT  292.42 594.2 307.1 602.38 ;
     RECT  304.7 336.74 308.54 356.68 ;
     RECT  294.34 367.4 308.54 408.76 ;
     RECT  305.18 539.18 308.54 549.04 ;
     RECT  302.5 321.62 312.38 327.7 ;
     RECT  308.54 336.74 312.38 408.76 ;
     RECT  306.14 648.38 313.54 690.16 ;
     RECT  312.38 107.42 313.82 107.62 ;
     RECT  313.82 99.44 314.3 107.62 ;
     RECT  308.54 537.08 314.78 549.04 ;
     RECT  312.38 321.62 314.98 408.76 ;
     RECT  314.98 336.74 315.26 408.76 ;
     RECT  302.98 420.74 315.26 522.58 ;
     RECT  314.3 99.44 315.74 108.04 ;
     RECT  304.7 198.56 315.74 198.76 ;
     RECT  302.5 207.8 315.74 208 ;
     RECT  315.26 336.74 316.42 522.58 ;
     RECT  311.42 133.88 316.7 134.08 ;
     RECT  315.26 156.56 316.7 156.76 ;
     RECT  286.66 179.66 316.7 184.06 ;
     RECT  307.1 569 316.7 602.38 ;
     RECT  316.7 156.56 317.38 160.96 ;
     RECT  315.74 93.14 318.14 108.04 ;
     RECT  316.7 130.52 319.1 134.08 ;
     RECT  316.7 178.82 319.1 184.9 ;
     RECT  317.38 159.08 319.3 160.96 ;
     RECT  318.14 88.1 320.54 108.04 ;
     RECT  319.1 171.26 320.54 184.9 ;
     RECT  319.3 159.5 321.22 160.96 ;
     RECT  320.54 88.1 321.7 111.4 ;
     RECT  316.42 336.74 321.7 408.76 ;
     RECT  321.7 99.44 321.98 111.4 ;
     RECT  321.98 99.44 322.46 112.24 ;
     RECT  322.46 99.44 322.94 116.02 ;
     RECT  320.54 171.26 322.94 188.68 ;
     RECT  315.74 198.56 322.94 208 ;
     RECT  321.7 88.1 323.14 88.3 ;
     RECT  302.5 220.82 323.42 311.74 ;
     RECT  321.22 159.92 323.9 160.96 ;
     RECT  322.94 171.26 323.9 208 ;
     RECT  311.9 712.64 325.34 712.84 ;
     RECT  319.1 130.52 325.82 140.8 ;
     RECT  318.62 149.42 325.82 149.62 ;
     RECT  313.54 667.28 326.3 690.16 ;
     RECT  302.5 700.88 326.3 701.08 ;
     RECT  323.9 159.92 326.98 208 ;
     RECT  325.34 712.64 326.98 718.72 ;
     RECT  326.98 160.34 327.94 208 ;
     RECT  316.42 417.38 328.22 522.58 ;
     RECT  326.3 667.28 328.9 701.08 ;
     RECT  325.82 130.52 330.34 149.62 ;
     RECT  328.22 417.38 330.34 526.36 ;
     RECT  328.9 688.28 330.34 701.08 ;
     RECT  314.78 537.08 331.1 554.08 ;
     RECT  316.7 568.58 331.1 602.38 ;
     RECT  331.1 537.08 331.3 602.38 ;
     RECT  328.9 667.28 331.3 678.4 ;
     RECT  327.94 160.76 331.58 208 ;
     RECT  323.42 217.04 331.58 311.74 ;
     RECT  314.98 321.62 332.06 327.7 ;
     RECT  331.3 561.44 332.26 602.38 ;
     RECT  302.5 612.68 332.54 635.56 ;
     RECT  313.54 648.38 332.54 656.14 ;
     RECT  321.7 336.74 332.74 356.68 ;
     RECT  332.06 321.2 333.02 327.7 ;
     RECT  332.74 336.74 333.02 337.78 ;
     RECT  330.34 130.52 333.22 139.96 ;
     RECT  331.58 160.76 334.46 311.74 ;
     RECT  333.02 321.2 334.46 337.78 ;
     RECT  332.26 568.58 335.14 602.38 ;
     RECT  334.46 160.76 336.1 337.78 ;
     RECT  322.94 99.44 337.34 119.8 ;
     RECT  336.1 194.78 338.02 337.78 ;
     RECT  332.06 73.4 339.26 73.6 ;
     RECT  337.34 92.72 339.26 119.8 ;
     RECT  330.34 420.74 339.74 526.36 ;
     RECT  331.3 537.08 339.74 549.04 ;
     RECT  336.1 160.76 339.94 184.9 ;
     RECT  339.74 420.74 339.94 549.04 ;
     RECT  339.26 73.4 340.22 77.8 ;
     RECT  339.26 88.94 340.22 119.8 ;
     RECT  339.94 420.74 340.42 538.96 ;
     RECT  340.22 73.4 341.38 119.8 ;
     RECT  340.42 420.74 341.38 530.98 ;
     RECT  341.38 73.4 342.34 100.06 ;
     RECT  342.34 88.94 342.82 100.06 ;
     RECT  335.14 569 342.82 602.38 ;
     RECT  341.38 111.62 343.1 119.8 ;
     RECT  333.22 130.52 343.1 134.08 ;
     RECT  342.34 73.4 343.3 77.8 ;
     RECT  342.82 88.94 343.78 92.92 ;
     RECT  330.34 688.28 343.78 690.16 ;
     RECT  343.1 111.62 344.26 134.08 ;
     RECT  338.02 194.78 344.74 197.08 ;
     RECT  332.54 612.68 344.74 656.14 ;
     RECT  344.26 114.56 345.02 134.08 ;
     RECT  321.7 367.82 345.7 408.76 ;
     RECT  341.38 420.74 345.7 526.36 ;
     RECT  330.34 149.42 345.98 149.62 ;
     RECT  332.74 348.5 346.46 356.68 ;
     RECT  345.7 367.82 346.46 406.24 ;
     RECT  339.94 164.12 346.66 184.9 ;
     RECT  331.3 669.8 346.66 678.4 ;
     RECT  344.74 612.68 347.14 651.1 ;
     RECT  344.74 195.2 347.42 197.08 ;
     RECT  338.02 207.8 347.42 337.78 ;
     RECT  346.46 348.5 347.62 406.24 ;
     RECT  347.14 612.68 348.58 640.6 ;
     RECT  346.66 164.96 348.86 184.9 ;
     RECT  343.78 92.72 349.06 92.92 ;
     RECT  345.7 517.34 349.06 526.36 ;
     RECT  345.98 726.92 349.54 727.12 ;
     RECT  349.06 518.6 350.02 526.36 ;
     RECT  345.02 114.56 352.7 134.5 ;
     RECT  343.3 73.4 352.9 74.02 ;
     RECT  345.98 149.42 353.66 154.24 ;
     RECT  352.7 113.72 354.34 139.96 ;
     RECT  347.14 650.9 354.62 651.1 ;
     RECT  346.46 659.72 354.62 659.92 ;
     RECT  339.94 548.84 355.58 549.04 ;
     RECT  343.58 557.66 355.58 557.86 ;
     RECT  353.66 149.42 356.26 155.92 ;
     RECT  354.62 650.9 356.26 659.92 ;
     RECT  348.86 164.96 356.54 186.58 ;
     RECT  347.42 195.2 356.54 337.78 ;
     RECT  346.66 669.8 357.5 670 ;
     RECT  356.54 164.96 357.7 337.78 ;
     RECT  330.34 700.88 358.46 701.08 ;
     RECT  343.78 688.28 360.86 688.48 ;
     RECT  357.7 165.8 361.06 337.78 ;
     RECT  356.26 149.42 362.02 149.62 ;
     RECT  354.34 114.98 362.3 139.96 ;
     RECT  360.86 688.28 362.5 690.16 ;
     RECT  358.46 700.88 362.78 706.12 ;
     RECT  362.3 114.98 364.7 147.52 ;
     RECT  362.5 689.96 364.7 690.16 ;
     RECT  362.78 699.2 364.7 706.12 ;
     RECT  342.82 594.2 364.9 602.38 ;
     RECT  357.5 77.6 366.14 77.8 ;
     RECT  356.26 650.9 366.62 656.14 ;
     RECT  361.06 167.9 367.3 337.78 ;
     RECT  366.14 77.6 367.58 81.16 ;
     RECT  357.5 666.86 367.58 670 ;
     RECT  367.58 77.18 368.06 81.16 ;
     RECT  364.7 114.56 368.26 147.52 ;
     RECT  367.58 99.86 369.02 100.06 ;
     RECT  366.62 650.9 369.22 656.56 ;
     RECT  364.7 689.96 369.7 706.12 ;
     RECT  369.02 99.86 370.18 106.78 ;
     RECT  369.22 650.9 370.18 656.14 ;
     RECT  370.18 99.86 371.42 100.06 ;
     RECT  369.7 699.2 371.62 706.12 ;
     RECT  368.06 77.18 371.9 81.58 ;
     RECT  371.42 92.3 371.9 100.06 ;
     RECT  355.58 548.84 373.34 557.86 ;
     RECT  342.82 569 373.34 584.74 ;
     RECT  367.3 168.32 375.26 337.78 ;
     RECT  347.62 348.5 375.26 356.68 ;
     RECT  375.26 168.32 376.22 356.68 ;
     RECT  368.54 157.4 377.18 157.6 ;
     RECT  371.9 77.18 379.78 100.06 ;
     RECT  368.26 121.7 380.54 147.52 ;
     RECT  377.18 156.98 380.54 157.6 ;
     RECT  367.58 666.44 380.74 670 ;
     RECT  371.62 700.88 381.7 706.12 ;
     RECT  380.54 121.7 381.98 157.6 ;
     RECT  376.22 167.06 381.98 356.68 ;
     RECT  373.34 548.84 382.94 584.74 ;
     RECT  364.9 594.2 382.94 601.96 ;
     RECT  370.18 650.9 383.62 651.94 ;
     RECT  369.7 689.96 384.58 690.16 ;
     RECT  379.58 66.26 386.02 66.46 ;
     RECT  379.78 77.6 386.98 100.06 ;
     RECT  381.98 121.7 387.94 356.68 ;
     RECT  386.98 80.96 388.22 100.06 ;
     RECT  350.02 518.6 388.7 522.58 ;
     RECT  387.94 121.7 389.38 337.78 ;
     RECT  380.74 666.86 391.58 670 ;
     RECT  389.38 121.7 392.26 201.7 ;
     RECT  388.22 80.96 394.18 100.9 ;
     RECT  394.18 92.3 394.66 100.9 ;
     RECT  392.26 121.7 394.94 147.52 ;
     RECT  394.94 115.82 395.14 147.52 ;
     RECT  392.26 156.14 395.14 201.7 ;
     RECT  382.94 548.84 395.14 601.96 ;
     RECT  383.62 650.9 395.9 651.1 ;
     RECT  394.66 92.3 396.1 100.48 ;
     RECT  395.14 115.82 396.1 126.1 ;
     RECT  391.58 666.86 396.58 678.4 ;
     RECT  396.1 92.3 397.06 100.06 ;
     RECT  396.58 666.86 397.06 670 ;
     RECT  381.7 700.88 397.54 701.08 ;
     RECT  347.62 367.82 399.26 406.24 ;
     RECT  394.18 81.38 401.38 81.58 ;
     RECT  395.14 569.84 401.66 601.96 ;
     RECT  348.58 612.68 401.66 635.56 ;
     RECT  395.14 137.66 402.14 147.52 ;
     RECT  395.14 156.14 402.14 157.6 ;
     RECT  389.38 213.26 402.14 337.78 ;
     RECT  387.94 348.5 402.14 356.68 ;
     RECT  397.06 92.3 402.62 99.64 ;
     RECT  395.9 645.44 402.82 651.1 ;
     RECT  401.66 569.84 403.1 635.56 ;
     RECT  395.14 168.32 404.06 201.7 ;
     RECT  399.26 367.82 404.54 410.02 ;
     RECT  388.22 51.98 404.74 52.18 ;
     RECT  402.14 137.66 405.02 157.6 ;
     RECT  404.06 166.64 405.02 201.7 ;
     RECT  388.7 518.6 405.02 523.42 ;
     RECT  405.02 137.66 405.5 201.7 ;
     RECT  395.14 548.84 405.5 561.22 ;
     RECT  403.1 569.84 405.5 637.24 ;
     RECT  397.06 669.8 405.5 670 ;
     RECT  396.1 121.7 406.46 126.1 ;
     RECT  402.82 648.8 406.94 651.1 ;
     RECT  405.5 548.84 408.1 637.24 ;
     RECT  405.5 137.66 408.86 202.96 ;
     RECT  402.14 213.26 408.86 356.68 ;
     RECT  402.62 88.52 410.78 99.64 ;
     RECT  406.46 118.76 410.78 126.1 ;
     RECT  404.54 367.82 410.78 411.28 ;
     RECT  345.7 420.74 410.78 508.3 ;
     RECT  408.1 569.84 411.26 637.24 ;
     RECT  406.94 648.8 411.26 652.78 ;
     RECT  411.26 569.84 411.74 652.78 ;
     RECT  405.5 661.82 411.74 670 ;
     RECT  410.78 86 412.7 99.64 ;
     RECT  411.74 569.84 412.9 670 ;
     RECT  392.54 539.6 413.66 539.8 ;
     RECT  413.66 538.76 413.86 539.8 ;
     RECT  408.86 137.66 414.34 356.68 ;
     RECT  405.02 518.6 414.34 528.46 ;
     RECT  414.34 137.66 415.58 337.78 ;
     RECT  410.78 118.76 417.02 126.94 ;
     RECT  410.78 46.94 417.22 47.14 ;
     RECT  417.02 114.98 417.5 126.94 ;
     RECT  417.5 114.56 417.7 126.94 ;
     RECT  415.58 136.4 417.7 337.78 ;
     RECT  410.78 367.82 417.7 508.3 ;
     RECT  408.1 548.84 417.7 561.22 ;
     RECT  413.86 538.76 421.34 538.96 ;
     RECT  417.7 121.7 421.54 126.94 ;
     RECT  414.34 518.6 421.54 523.42 ;
     RECT  421.34 538.34 421.54 538.96 ;
     RECT  412.7 83.48 422.78 99.64 ;
     RECT  421.54 538.76 423.46 538.96 ;
     RECT  412.9 576.56 424.22 670 ;
     RECT  422.78 83.48 426.14 100.06 ;
     RECT  424.22 571.52 428.06 670 ;
     RECT  417.7 549.68 431.42 561.22 ;
     RECT  428.06 570.68 431.42 670 ;
     RECT  426.14 83.48 431.62 108.04 ;
     RECT  421.54 519.86 431.9 523.42 ;
     RECT  417.7 137.66 432.38 337.78 ;
     RECT  421.54 125.9 433.54 126.94 ;
     RECT  417.7 367.82 433.82 507.88 ;
     RECT  431.9 519.86 433.82 527.62 ;
     RECT  431.42 549.68 434.02 670 ;
     RECT  433.82 367.82 436.9 527.62 ;
     RECT  431.62 83.48 437.38 100.48 ;
     RECT  434.02 570.68 437.86 670 ;
     RECT  414.34 348.5 440.06 356.68 ;
     RECT  436.9 367.82 440.06 523.42 ;
     RECT  437.86 571.94 441.02 670 ;
     RECT  432.38 137.66 441.5 338.2 ;
     RECT  441.5 136.82 441.98 338.2 ;
     RECT  440.06 348.5 441.98 523.42 ;
     RECT  437.38 86 442.46 100.48 ;
     RECT  433.54 125.9 445.34 126.1 ;
     RECT  441.98 136.82 445.34 523.42 ;
     RECT  445.34 125.9 448.42 523.42 ;
     RECT  441.02 571.94 448.42 670.42 ;
     RECT  427.1 50.72 448.9 50.92 ;
     RECT  448.42 367.82 449.86 523.42 ;
     RECT  448.42 576.14 450.82 670.42 ;
     RECT  448.42 125.9 451.58 356.68 ;
     RECT  442.46 86 453.5 107.62 ;
     RECT  451.58 118.76 453.5 356.68 ;
     RECT  450.82 576.14 453.7 670 ;
     RECT  453.7 669.38 455.62 670 ;
     RECT  434.02 549.68 455.9 561.22 ;
     RECT  453.5 86 456.86 356.68 ;
     RECT  449.86 522.38 456.86 523.42 ;
     RECT  455.9 545.9 458.5 561.22 ;
     RECT  449.86 367.82 460.22 507.88 ;
     RECT  458.5 549.68 460.22 561.22 ;
     RECT  453.7 576.14 460.42 655.72 ;
     RECT  456.86 85.16 460.9 356.68 ;
     RECT  460.9 85.16 461.38 169.78 ;
     RECT  460.42 576.14 461.38 642.28 ;
     RECT  461.38 576.14 461.86 635.56 ;
     RECT  456.86 522.38 463.58 528.04 ;
     RECT  460.22 549.68 465.02 562.06 ;
     RECT  460.22 367.82 467.42 509.14 ;
     RECT  461.86 576.14 467.9 601.96 ;
     RECT  460.9 178.82 468.38 356.68 ;
     RECT  467.42 367.82 468.38 509.98 ;
     RECT  461.38 114.98 468.58 169.78 ;
     RECT  463.58 520.28 468.86 528.04 ;
     RECT  466.94 539.6 468.86 539.8 ;
     RECT  455.42 54.5 469.54 54.7 ;
     RECT  468.38 178.82 469.82 509.98 ;
     RECT  468.86 520.28 469.82 539.8 ;
     RECT  468.58 124.64 470.3 169.78 ;
     RECT  469.82 178.82 470.3 539.8 ;
     RECT  467.9 574.04 471.46 601.96 ;
     RECT  461.38 85.16 471.74 105.1 ;
     RECT  468.58 114.98 471.74 115.18 ;
     RECT  470.3 124.64 473.38 539.8 ;
     RECT  473.38 178.4 473.86 539.8 ;
     RECT  471.46 574.04 473.86 584.74 ;
     RECT  473.86 419.9 475.1 539.8 ;
     RECT  465.02 549.68 475.1 565 ;
     RECT  475.1 419.9 475.3 565 ;
     RECT  471.74 85.16 477.7 115.18 ;
     RECT  477.7 85.16 479.62 111.82 ;
     RECT  473.38 124.64 482.3 169.78 ;
     RECT  473.86 178.4 482.3 411.28 ;
     RECT  479.62 85.16 482.5 109.3 ;
     RECT  482.5 85.16 484.22 105.1 ;
     RECT  482.3 124.64 484.22 411.28 ;
     RECT  484.22 122.96 484.42 411.28 ;
     RECT  475.3 419.9 484.7 561.22 ;
     RECT  461.86 613.1 484.7 635.56 ;
     RECT  484.42 178.82 485.66 411.28 ;
     RECT  484.7 419.9 485.66 561.64 ;
     RECT  473.86 576.14 485.66 584.74 ;
     RECT  484.22 80.96 489.02 105.1 ;
     RECT  484.7 613.1 489.22 640.6 ;
     RECT  489.02 80.54 489.5 105.1 ;
     RECT  484.42 122.96 489.5 169.36 ;
     RECT  455.62 669.8 489.5 670 ;
     RECT  471.46 594.62 489.98 601.96 ;
     RECT  489.5 115.4 490.66 169.36 ;
     RECT  490.66 122.96 492.1 169.36 ;
     RECT  489.5 669.8 492.86 671.26 ;
     RECT  492.1 124.64 494.02 169.36 ;
     RECT  489.98 594.62 494.98 602.8 ;
     RECT  492.86 669.8 495.46 678.4 ;
     RECT  460.42 650.9 498.14 651.1 ;
     RECT  489.5 72.98 498.82 105.1 ;
     RECT  498.14 650.9 499.1 652.36 ;
     RECT  496.7 705.08 499.1 705.28 ;
     RECT  495.46 669.8 499.78 670 ;
     RECT  499.1 650.9 500.06 655.72 ;
     RECT  494.98 594.62 500.54 601.96 ;
     RECT  498.82 84.74 503.14 105.1 ;
     RECT  499.58 728.18 503.14 728.38 ;
     RECT  500.06 650.9 503.62 656.56 ;
     RECT  499.1 705.08 503.62 708.64 ;
     RECT  498.82 72.98 504.1 75.28 ;
     RECT  503.14 88.52 504.1 105.1 ;
     RECT  489.22 613.1 504.38 637.66 ;
     RECT  503.62 650.9 504.58 655.72 ;
     RECT  494.02 125.9 504.86 169.36 ;
     RECT  485.66 178.82 504.86 584.74 ;
     RECT  503.9 114.98 505.34 115.18 ;
     RECT  504.86 125.9 505.34 584.74 ;
     RECT  500.54 593.78 505.34 601.96 ;
     RECT  503.62 708.02 506.3 708.64 ;
     RECT  505.34 125.9 506.5 601.96 ;
     RECT  505.82 674.84 507.26 675.04 ;
     RECT  504.38 613.1 507.46 640.6 ;
     RECT  506.3 708.02 507.74 716.2 ;
     RECT  506.78 738.68 509.18 738.88 ;
     RECT  506.5 532.46 510.34 601.96 ;
     RECT  510.34 534.56 511.58 601.96 ;
     RECT  507.46 613.1 511.58 635.56 ;
     RECT  509.18 738.68 512.26 743.08 ;
     RECT  504.1 88.52 512.54 100.06 ;
     RECT  507.26 674.84 512.74 683.44 ;
     RECT  507.74 708.02 512.74 720.4 ;
     RECT  513.02 758.42 514.46 758.62 ;
     RECT  505.82 67.94 514.94 68.14 ;
     RECT  512.74 708.02 515.14 715.78 ;
     RECT  512.74 683.24 516.1 683.44 ;
     RECT  512.54 88.52 516.38 100.48 ;
     RECT  515.14 708.02 516.38 715.36 ;
     RECT  512.26 742.88 516.38 743.08 ;
     RECT  504.58 650.9 516.86 651.1 ;
     RECT  511.58 534.56 517.54 635.56 ;
     RECT  516.38 85.16 518.02 100.48 ;
     RECT  512.06 692.48 518.02 692.68 ;
     RECT  516.38 742.88 518.02 746.44 ;
     RECT  516.38 701.3 518.3 715.36 ;
     RECT  517.54 534.56 518.5 601.96 ;
     RECT  514.46 758.42 518.78 761.56 ;
     RECT  506.5 125.9 518.98 523.84 ;
     RECT  518.5 534.56 518.98 601.54 ;
     RECT  514.94 67.94 519.26 74.02 ;
     RECT  516.86 650.9 520.9 656.56 ;
     RECT  518.78 758 521.38 761.56 ;
     RECT  518.02 88.52 521.66 100.48 ;
     RECT  505.34 112.46 521.66 115.18 ;
     RECT  520.9 650.9 522.34 656.14 ;
     RECT  518.02 745.4 522.34 746.44 ;
     RECT  521.66 88.52 523.58 115.18 ;
     RECT  518.98 125.9 523.58 523.42 ;
     RECT  518.3 700.88 523.78 715.36 ;
     RECT  521.38 758.42 523.78 761.56 ;
     RECT  522.34 652.58 524.26 656.14 ;
     RECT  523.78 700.88 524.26 704.86 ;
     RECT  524.26 700.88 525.22 704.44 ;
     RECT  519.26 64.58 525.7 74.02 ;
     RECT  523.78 760.52 525.7 761.56 ;
     RECT  523.1 678.2 527.14 678.4 ;
     RECT  525.22 702.56 527.62 704.44 ;
     RECT  518.98 542.96 529.34 601.54 ;
     RECT  523.58 88.52 530.3 523.42 ;
     RECT  529.34 542.96 531.46 602.8 ;
     RECT  524.26 655.94 531.74 656.14 ;
     RECT  531.74 655.94 533.86 663.28 ;
     RECT  525.7 67.94 534.14 74.02 ;
     RECT  530.3 88.52 534.14 527.2 ;
     RECT  531.46 542.96 534.14 561.64 ;
     RECT  533.86 663.08 534.14 663.28 ;
     RECT  525.7 761.36 534.62 761.56 ;
     RECT  534.14 663.08 535.3 670 ;
     RECT  522.34 745.4 536.54 745.6 ;
     RECT  535.3 669.8 536.74 670 ;
     RECT  534.14 67.94 537.5 527.2 ;
     RECT  534.14 536.24 537.5 561.64 ;
     RECT  523.78 715.16 538.66 715.36 ;
     RECT  534.62 760.94 539.14 761.56 ;
     RECT  539.14 760.94 539.62 761.14 ;
     RECT  536.54 744.98 540.38 745.6 ;
     RECT  531.26 693.32 541.06 693.52 ;
     RECT  537.5 67.94 541.34 561.64 ;
     RECT  527.62 702.56 541.34 702.76 ;
     RECT  541.34 67.94 541.54 562.06 ;
     RECT  517.54 613.1 542.3 635.56 ;
     RECT  541.54 114.56 542.5 562.06 ;
     RECT  539.9 727.34 542.5 727.54 ;
     RECT  540.38 738.68 543.26 745.6 ;
     RECT  541.54 67.94 543.74 104.26 ;
     RECT  541.34 694.58 544.42 702.76 ;
     RECT  543.74 59.54 546.34 104.26 ;
     RECT  546.34 59.54 546.82 100.48 ;
     RECT  542.5 114.56 546.82 561.64 ;
     RECT  542.3 613.1 547.1 636.82 ;
     RECT  542.78 718.94 547.1 721.24 ;
     RECT  547.1 712.22 547.3 721.24 ;
     RECT  547.1 613.1 547.58 643.54 ;
     RECT  544.42 697.52 549.7 702.76 ;
     RECT  546.82 67.94 551.62 100.48 ;
     RECT  546.82 122.54 552.38 561.64 ;
     RECT  552.38 122.54 553.82 562.06 ;
     RECT  531.46 571.94 553.82 602.8 ;
     RECT  553.82 122.54 554.3 602.8 ;
     RECT  547.58 613.1 554.3 643.96 ;
     RECT  549.7 697.94 554.3 702.76 ;
     RECT  547.3 712.22 554.3 712.42 ;
     RECT  553.82 786.98 554.3 787.18 ;
     RECT  554.3 677.36 554.78 677.56 ;
     RECT  554.3 785.72 554.78 787.18 ;
     RECT  543.26 734.06 555.26 745.6 ;
     RECT  554.3 122.54 555.46 643.96 ;
     RECT  554.78 784.04 555.74 787.18 ;
     RECT  551.62 67.94 556.22 99.64 ;
     RECT  554.78 677.36 556.22 682.6 ;
     RECT  556.22 677.36 557.38 683.44 ;
     RECT  557.38 677.78 558.14 683.44 ;
     RECT  556.22 64.58 558.34 99.64 ;
     RECT  554.3 722.3 558.62 722.5 ;
     RECT  555.26 731.12 558.62 745.6 ;
     RECT  554.3 756.32 558.62 756.52 ;
     RECT  558.62 756.32 559.1 760.3 ;
     RECT  558.62 722.3 560.54 745.6 ;
     RECT  559.1 756.32 560.54 761.56 ;
     RECT  555.46 123.38 560.74 643.96 ;
     RECT  558.14 677.78 560.74 689.32 ;
     RECT  560.74 689.12 561.98 689.32 ;
     RECT  554.3 697.94 561.98 712.42 ;
     RECT  558.34 69.2 562.66 99.64 ;
     RECT  559.1 659.72 562.94 659.92 ;
     RECT  555.74 784.04 565.06 788.44 ;
     RECT  561.02 113.3 565.34 113.5 ;
     RECT  560.74 123.38 565.34 141.64 ;
     RECT  561.98 689.12 565.34 712.42 ;
     RECT  560.54 722.3 565.34 761.56 ;
     RECT  562.66 96.08 565.54 99.64 ;
     RECT  560.74 152.36 565.82 643.96 ;
     RECT  560.74 677.78 566.02 677.98 ;
     RECT  565.34 689.12 566.02 761.56 ;
     RECT  561.5 772.28 566.02 772.48 ;
     RECT  565.34 113.3 566.3 141.64 ;
     RECT  562.66 69.2 566.98 86.2 ;
     RECT  565.06 784.04 567.74 785.92 ;
     RECT  566.98 70.04 568.9 86.2 ;
     RECT  562.94 659.72 568.9 663.28 ;
     RECT  567.74 783.62 568.9 785.92 ;
     RECT  568.9 659.72 569.38 662.86 ;
     RECT  566.3 103.64 569.66 141.64 ;
     RECT  565.82 152.36 569.66 647.74 ;
     RECT  569.66 103.64 569.86 647.74 ;
     RECT  568.9 76.76 570.82 86.2 ;
     RECT  568.9 783.62 570.82 784.24 ;
     RECT  569.66 678.62 571.3 678.82 ;
     RECT  570.82 784.04 571.3 784.24 ;
     RECT  571.58 802.52 572.54 802.72 ;
     RECT  569.86 124.22 572.74 647.74 ;
     RECT  572.54 802.52 573.5 803.56 ;
     RECT  570.82 76.76 574.18 81.16 ;
     RECT  572.74 152.36 575.42 647.74 ;
     RECT  566.02 689.12 575.9 689.32 ;
     RECT  566.02 697.94 575.9 761.56 ;
     RECT  572.74 124.22 576.1 141.64 ;
     RECT  569.38 662.66 576.1 662.86 ;
     RECT  573.5 799.16 578.98 803.56 ;
     RECT  575.42 152.36 579.46 651.94 ;
     RECT  578.98 799.16 579.46 803.14 ;
     RECT  579.46 802.52 580.42 803.14 ;
     RECT  576.1 124.22 580.7 138.7 ;
     RECT  579.46 152.36 580.9 644.8 ;
     RECT  574.46 674.84 581.18 675.04 ;
     RECT  574.18 78.02 581.38 81.16 ;
     RECT  580.42 802.52 581.38 802.72 ;
     RECT  575.9 689.12 581.86 761.56 ;
     RECT  581.18 780.68 582.14 780.88 ;
     RECT  580.7 123.8 582.82 138.7 ;
     RECT  580.9 152.36 582.82 643.96 ;
     RECT  581.86 689.96 583.78 761.56 ;
     RECT  569.86 103.64 584.06 115.18 ;
     RECT  581.18 674.84 584.54 676.72 ;
     RECT  571.1 92.3 584.74 92.5 ;
     RECT  582.82 124.22 584.74 138.7 ;
     RECT  584.06 103.22 585.02 115.18 ;
     RECT  585.02 103.22 585.7 115.6 ;
     RECT  582.14 780.68 586.94 781.3 ;
     RECT  584.54 669.8 587.9 676.72 ;
     RECT  584.74 138.5 588.38 138.7 ;
     RECT  585.7 103.64 589.54 115.6 ;
     RECT  587.9 669.38 589.82 676.72 ;
     RECT  586.94 780.68 589.82 788.44 ;
     RECT  588.38 138.5 590.02 143.74 ;
     RECT  584.74 124.22 590.98 129.88 ;
     RECT  582.82 152.36 591.26 186.58 ;
     RECT  582.82 195.2 591.26 643.96 ;
     RECT  585.5 658.88 591.26 659.08 ;
     RECT  590.02 138.5 591.94 138.7 ;
     RECT  591.26 658.88 592.22 659.5 ;
     RECT  591.26 152.36 592.7 643.96 ;
     RECT  592.22 655.52 592.7 659.5 ;
     RECT  592.7 152.36 593.18 659.5 ;
     RECT  589.82 669.38 593.18 678.4 ;
     RECT  589.82 780.26 593.38 788.44 ;
     RECT  593.38 783.62 593.66 788.44 ;
     RECT  593.18 152.36 593.86 678.4 ;
     RECT  583.78 689.96 593.86 760.72 ;
     RECT  581.38 80.96 594.82 81.16 ;
     RECT  593.86 689.96 594.82 712.42 ;
     RECT  593.86 152.36 595.3 274.36 ;
     RECT  593.86 722.3 595.3 760.72 ;
     RECT  593.66 783.62 596.06 795.58 ;
     RECT  593.86 284.24 596.74 678.4 ;
     RECT  596.06 783.62 598.18 796 ;
     RECT  596.74 655.52 599.62 678.4 ;
     RECT  598.18 783.62 599.62 788.44 ;
     RECT  595.3 748.76 600.86 760.72 ;
     RECT  589.54 115.4 601.54 115.6 ;
     RECT  590.98 124.22 601.54 124.42 ;
     RECT  593.18 136.82 602.3 137.02 ;
     RECT  602.3 133.88 602.78 137.02 ;
     RECT  595.3 152.36 603.26 270.16 ;
     RECT  603.26 149 603.46 270.16 ;
     RECT  600.86 748.76 603.46 761.56 ;
     RECT  595.3 722.3 603.94 738.88 ;
     RECT  603.46 748.76 603.94 760.72 ;
     RECT  602.78 133.88 604.7 139.96 ;
     RECT  603.46 195.2 604.7 270.16 ;
     RECT  596.74 284.24 604.7 643.96 ;
     RECT  603.94 732.8 604.7 738.88 ;
     RECT  603.94 748.76 604.7 759.04 ;
     RECT  603.26 821 604.7 821.2 ;
     RECT  589.54 103.64 604.9 105.94 ;
     RECT  603.46 149 604.9 186.58 ;
     RECT  594.82 691.22 605.18 712.42 ;
     RECT  604.7 128.84 605.86 139.96 ;
     RECT  599.62 783.62 605.86 783.82 ;
     RECT  604.7 195.2 606.34 643.96 ;
     RECT  604.7 821 607.58 826.24 ;
     RECT  606.34 195.2 607.78 637.24 ;
     RECT  605.86 128.84 608.74 129.04 ;
     RECT  599.62 655.94 609.02 669.16 ;
     RECT  607.58 818.06 609.02 826.24 ;
     RECT  605.86 139.76 609.7 139.96 ;
     RECT  607.58 807.56 609.98 807.76 ;
     RECT  605.18 684.92 610.94 712.84 ;
     RECT  607.78 195.2 612.58 614.98 ;
     RECT  610.94 682.82 612.86 712.84 ;
     RECT  604.9 153.2 613.06 184.06 ;
     RECT  609.98 806.72 613.06 807.76 ;
     RECT  607.78 624.44 613.54 637.24 ;
     RECT  609.02 654.68 613.82 669.16 ;
     RECT  612.86 678.62 613.82 712.84 ;
     RECT  613.82 654.68 614.3 712.84 ;
     RECT  603.94 723.14 614.3 724.18 ;
     RECT  613.06 806.72 614.78 807.34 ;
     RECT  614.78 805.46 614.98 807.34 ;
     RECT  614.98 805.46 615.94 806.92 ;
     RECT  609.5 99.86 616.22 100.06 ;
     RECT  612.86 111.2 616.22 111.4 ;
     RECT  609.02 818.06 616.42 833.8 ;
     RECT  614.3 654.68 616.7 724.18 ;
     RECT  604.7 732.8 616.7 759.04 ;
     RECT  612.58 284.24 617.18 614.98 ;
     RECT  613.54 624.44 617.18 635.56 ;
     RECT  615.94 805.46 617.38 805.66 ;
     RECT  613.34 788.24 617.86 788.44 ;
     RECT  616.22 99.86 618.34 111.4 ;
     RECT  616.7 126.74 618.62 126.94 ;
     RECT  618.34 111.2 619.78 111.4 ;
     RECT  618.62 126.32 619.78 126.94 ;
     RECT  617.18 284.24 619.78 635.56 ;
     RECT  616.7 654.68 619.78 759.04 ;
     RECT  612.58 195.2 620.06 270.16 ;
     RECT  613.06 153.2 622.18 181.12 ;
     RECT  622.18 155.3 622.46 181.12 ;
     RECT  620.06 189.74 622.46 270.16 ;
     RECT  618.34 99.86 623.14 100.48 ;
     RECT  616.42 826.04 623.42 833.8 ;
     RECT  622.46 155.3 623.62 270.16 ;
     RECT  623.14 100.28 624.1 100.48 ;
     RECT  619.78 655.94 624.58 759.04 ;
     RECT  619.78 284.24 624.86 614.98 ;
     RECT  619.78 624.44 625.54 635.56 ;
     RECT  624.38 803.36 626.3 803.56 ;
     RECT  624.58 656.78 627.46 759.04 ;
     RECT  625.54 633.68 627.74 635.56 ;
     RECT  606.14 776.48 627.94 776.68 ;
     RECT  627.46 661.82 629.86 759.04 ;
     RECT  626.3 802.94 630.34 803.56 ;
     RECT  619.78 126.32 631.3 126.52 ;
     RECT  630.34 802.94 631.3 803.14 ;
     RECT  623.42 826.04 631.3 837.16 ;
     RECT  631.3 826.04 632.26 826.24 ;
     RECT  625.54 624.44 633.22 624.64 ;
     RECT  629.86 667.7 633.7 759.04 ;
     RECT  633.7 667.7 636.1 675.88 ;
     RECT  631.3 836.54 636.1 837.16 ;
     RECT  636.1 836.54 637.06 836.74 ;
     RECT  624.86 282.98 637.34 614.98 ;
     RECT  623.62 191 638.78 270.16 ;
     RECT  623.62 155.3 638.98 181.12 ;
     RECT  636.1 667.7 639.26 675.04 ;
     RECT  638.78 191 639.46 273.94 ;
     RECT  633.7 684.92 639.46 759.04 ;
     RECT  639.26 663.08 639.74 675.04 ;
     RECT  639.46 690.8 639.94 759.04 ;
     RECT  638.98 177.98 640.22 181.12 ;
     RECT  639.46 191 640.22 270.16 ;
     RECT  638.3 145.64 640.9 145.84 ;
     RECT  637.34 282.98 641.18 615.82 ;
     RECT  639.94 721.88 641.18 759.04 ;
     RECT  641.18 282.98 641.66 617.5 ;
     RECT  639.74 655.94 644.26 675.04 ;
     RECT  627.74 633.68 646.18 639.76 ;
     RECT  644.26 655.94 646.18 670.84 ;
     RECT  639.94 691.22 646.18 712.84 ;
     RECT  641.66 282.98 646.46 617.92 ;
     RECT  641.18 721.88 646.66 762.4 ;
     RECT  646.46 282.98 647.14 624.64 ;
     RECT  646.18 655.94 648.38 667.9 ;
     RECT  624.86 815.54 648.38 815.74 ;
     RECT  646.18 700.88 648.58 712.84 ;
     RECT  646.66 744.98 649.06 762.4 ;
     RECT  648.38 653 649.34 667.9 ;
     RECT  648.58 700.88 649.54 701.5 ;
     RECT  646.18 633.68 650.5 638.5 ;
     RECT  648.38 813.86 650.78 815.74 ;
     RECT  649.34 652.16 651.46 667.9 ;
     RECT  647.14 282.98 651.94 617.5 ;
     RECT  651.94 296 652.42 617.5 ;
     RECT  650.78 813.02 652.7 815.74 ;
     RECT  649.06 745.82 652.9 762.4 ;
     RECT  651.46 652.16 653.38 657.4 ;
     RECT  640.22 177.98 653.66 270.16 ;
     RECT  650.5 633.68 653.86 636.4 ;
     RECT  652.9 747.5 653.86 762.4 ;
     RECT  653.66 177.98 655.3 271 ;
     RECT  651.46 667.7 655.3 667.9 ;
     RECT  653.86 750.44 655.3 762.4 ;
     RECT  648.58 712.22 655.58 712.84 ;
     RECT  646.66 721.88 655.58 736.36 ;
     RECT  652.7 813.02 655.78 818.68 ;
     RECT  651.94 282.98 656.54 283.18 ;
     RECT  655.3 186.8 657.02 271 ;
     RECT  656.54 282.56 657.02 283.18 ;
     RECT  652.42 296.42 657.5 617.5 ;
     RECT  655.78 813.44 658.66 818.68 ;
     RECT  655.58 712.22 659.14 736.36 ;
     RECT  658.66 818.48 659.62 818.68 ;
     RECT  655.3 750.86 660.58 751.06 ;
     RECT  657.02 186.8 661.34 283.18 ;
     RECT  657.5 296.42 662.5 620.44 ;
     RECT  638.98 156.14 662.98 169.36 ;
     RECT  662.5 296.42 662.98 615.82 ;
     RECT  659.14 727.76 662.98 736.36 ;
     RECT  661.34 186.8 663.74 285.7 ;
     RECT  662.98 296.42 663.74 614.56 ;
     RECT  653.38 654.68 665.66 657.4 ;
     RECT  653.86 633.68 667.1 635.56 ;
     RECT  659.14 712.22 667.3 718.3 ;
     RECT  662.98 727.76 667.78 727.96 ;
     RECT  665.66 652.16 668.06 657.4 ;
     RECT  661.34 773.12 668.54 773.32 ;
     RECT  667.1 625.7 668.74 635.56 ;
     RECT  668.06 652.16 669.5 659.5 ;
     RECT  667.3 712.22 669.5 712.84 ;
     RECT  649.54 700.88 670.46 701.08 ;
     RECT  668.54 773.12 670.66 776.26 ;
     RECT  662.98 161.18 671.9 169.36 ;
     RECT  663.74 179.66 671.9 614.56 ;
     RECT  669.5 645.86 671.9 662.44 ;
     RECT  670.66 773.12 672.1 773.32 ;
     RECT  671.9 161.18 673.06 614.56 ;
     RECT  670.46 697.52 674.3 701.08 ;
     RECT  669.5 710.54 674.3 712.84 ;
     RECT  673.06 161.18 675.94 613.3 ;
     RECT  671.9 645.86 675.94 667.9 ;
     RECT  668.74 633.68 676.22 635.56 ;
     RECT  675.94 645.86 676.22 663.7 ;
     RECT  674.3 697.52 676.42 712.84 ;
     RECT  676.42 705.08 678.34 712.84 ;
     RECT  678.34 710.54 679.58 712.84 ;
     RECT  675.94 161.18 680.26 294.52 ;
     RECT  679.58 710.54 680.26 720.4 ;
     RECT  676.22 633.68 681.5 663.7 ;
     RECT  680.26 161.18 682.18 271.84 ;
     RECT  682.46 694.16 683.42 694.36 ;
     RECT  680.26 720.2 683.42 720.4 ;
     RECT  682.46 760.94 683.9 761.14 ;
     RECT  680.26 282.56 684.1 294.52 ;
     RECT  681.5 632.42 684.58 663.7 ;
     RECT  675.94 303.14 684.86 613.3 ;
     RECT  683.9 758.42 684.86 761.14 ;
     RECT  682.18 186.8 685.06 271.84 ;
     RECT  684.1 285.5 685.34 294.52 ;
     RECT  684.86 303.14 685.34 618.34 ;
     RECT  680.54 677.36 685.34 677.56 ;
     RECT  683.42 689.96 685.34 694.36 ;
     RECT  684.58 645.86 685.54 663.7 ;
     RECT  685.34 677.36 685.54 694.36 ;
     RECT  682.18 161.18 686.02 176.08 ;
     RECT  685.54 658.88 686.3 663.7 ;
     RECT  686.3 658.88 686.5 671.26 ;
     RECT  686.5 660.14 686.98 671.26 ;
     RECT  685.54 681.98 687.46 694.36 ;
     RECT  683.42 720.2 687.46 724.6 ;
     RECT  680.26 710.54 688.22 710.74 ;
     RECT  684.86 758 688.22 761.14 ;
     RECT  686.98 660.56 688.42 671.26 ;
     RECT  688.22 705.08 688.42 710.74 ;
     RECT  688.42 660.56 688.9 660.76 ;
     RECT  685.54 648.38 689.38 648.58 ;
     RECT  685.34 285.5 690.82 618.34 ;
     RECT  685.06 186.8 691.78 269.74 ;
     RECT  688.22 758 691.78 761.56 ;
     RECT  691.78 186.8 692.26 267.22 ;
     RECT  690.82 285.5 692.74 614.56 ;
     RECT  687.46 689.96 693.7 694.36 ;
     RECT  687.46 723.56 693.98 724.6 ;
     RECT  688.42 705.08 694.18 705.28 ;
     RECT  692.74 285.5 694.66 613.3 ;
     RECT  692.26 186.8 696.58 220.18 ;
     RECT  694.66 320.36 697.06 613.3 ;
     RECT  693.7 689.96 697.54 690.58 ;
     RECT  691.78 758 698.02 758.62 ;
     RECT  692.26 228.8 698.98 267.22 ;
     RECT  693.98 723.56 699.46 727.96 ;
     RECT  688.42 670.22 699.74 671.26 ;
     RECT  698.3 768.92 699.74 769.12 ;
     RECT  697.54 689.96 700.42 690.16 ;
     RECT  699.74 669.38 700.9 671.26 ;
     RECT  696.58 186.8 701.38 218.5 ;
     RECT  697.34 747.08 701.38 747.28 ;
     RECT  698.98 228.8 701.86 252.94 ;
     RECT  697.06 447.62 702.34 613.3 ;
     RECT  700.9 671.06 702.34 671.26 ;
     RECT  698.02 758 702.82 758.2 ;
     RECT  699.74 768.92 702.82 773.74 ;
     RECT  698.98 267.02 703.78 267.22 ;
     RECT  701.86 228.8 704.26 230.26 ;
     RECT  702.82 773.54 704.74 773.74 ;
     RECT  694.66 285.5 705.22 305.44 ;
     RECT  705.22 293.9 705.7 305.44 ;
     RECT  705.5 654.68 705.7 655.3 ;
     RECT  697.06 320.36 706.18 439 ;
     RECT  705.7 654.68 706.18 654.88 ;
     RECT  702.34 454.76 707.14 613.3 ;
     RECT  705.5 775.22 707.14 775.42 ;
     RECT  707.14 557.66 707.62 613.3 ;
     RECT  684.58 632.42 707.9 635.56 ;
     RECT  705.98 269.12 708.38 269.32 ;
     RECT  705.02 705.08 708.38 705.28 ;
     RECT  699.46 727.34 708.38 727.54 ;
     RECT  707.14 454.76 709.06 546.94 ;
     RECT  707.62 557.66 709.06 560.8 ;
     RECT  707.9 632.42 709.34 638.5 ;
     RECT  709.06 454.76 710.02 546.1 ;
     RECT  705.7 303.14 710.3 305.44 ;
     RECT  706.18 320.36 710.3 429.76 ;
     RECT  710.02 454.76 710.5 542.32 ;
     RECT  708.38 727.34 710.5 727.96 ;
     RECT  710.5 727.34 711.46 727.54 ;
     RECT  709.06 559.34 711.94 560.8 ;
     RECT  708.38 704.66 712.22 705.28 ;
     RECT  710.5 521.12 712.42 542.32 ;
     RECT  707.62 571.1 712.42 613.3 ;
     RECT  712.22 697.52 712.42 709.06 ;
     RECT  712.42 708.86 712.7 709.06 ;
     RECT  712.42 538.34 713.38 542.32 ;
     RECT  710.3 303.14 713.86 429.76 ;
     RECT  709.34 629.9 713.86 638.5 ;
     RECT  713.86 629.9 714.14 637.66 ;
     RECT  710.5 454.76 714.62 510.82 ;
     RECT  713.38 538.76 714.82 542.32 ;
     RECT  714.14 629.06 715.58 637.66 ;
     RECT  712.42 697.52 715.58 697.72 ;
     RECT  715.58 693.32 715.78 697.72 ;
     RECT  714.62 448.04 716.26 510.82 ;
     RECT  714.82 542.12 716.26 542.32 ;
     RECT  704.26 229.64 716.74 230.26 ;
     RECT  712.42 521.12 716.74 527.62 ;
     RECT  712.7 708.86 716.74 712.84 ;
     RECT  708.38 269.12 717.22 270.16 ;
     RECT  712.42 571.1 717.7 599.86 ;
     RECT  716.74 708.86 717.7 709.06 ;
     RECT  713.86 308.18 718.18 429.76 ;
     RECT  716.74 521.12 718.66 526.78 ;
     RECT  716.26 491.3 718.94 510.82 ;
     RECT  718.66 521.12 718.94 526.36 ;
     RECT  718.18 316.58 719.14 429.76 ;
     RECT  715.78 693.32 719.14 693.52 ;
     RECT  701.86 240.14 719.9 252.94 ;
     RECT  715.58 624.86 719.9 637.66 ;
     RECT  719.14 316.58 720.1 422.2 ;
     RECT  706.18 438.8 720.38 439 ;
     RECT  716.26 448.04 720.38 481.84 ;
     RECT  718.46 545.9 720.38 546.1 ;
     RECT  701.38 186.8 720.58 216.82 ;
     RECT  719.9 622.76 721.06 637.66 ;
     RECT  709.82 647.96 721.06 648.16 ;
     RECT  705.7 293.9 722.02 294.1 ;
     RECT  721.06 622.76 722.02 634.3 ;
     RECT  720.38 545.9 722.3 549.88 ;
     RECT  711.94 560.18 722.3 560.8 ;
     RECT  722.3 545.9 722.5 560.8 ;
     RECT  722.02 622.76 723.46 633.88 ;
     RECT  717.7 571.1 724.42 599.02 ;
     RECT  720.1 319.52 725.38 422.2 ;
     RECT  722.5 549.68 725.38 560.8 ;
     RECT  723.46 624.86 725.38 633.88 ;
     RECT  717.22 269.96 725.66 270.16 ;
     RECT  720.38 438.8 726.14 481.84 ;
     RECT  725.38 319.52 726.34 421.78 ;
     RECT  725.38 553.04 726.34 560.8 ;
     RECT  725.38 632.84 726.34 633.88 ;
     RECT  726.34 319.52 726.82 420.52 ;
     RECT  726.34 553.46 726.82 560.8 ;
     RECT  726.14 438.8 728.06 482.26 ;
     RECT  718.94 491.3 728.06 526.36 ;
     RECT  726.82 319.52 728.54 394.06 ;
     RECT  724.42 571.1 729.7 594.82 ;
     RECT  728.54 316.58 730.18 394.06 ;
     RECT  728.06 438.8 730.18 526.36 ;
     RECT  730.18 438.8 730.66 512.5 ;
     RECT  729.7 571.1 730.66 586.84 ;
     RECT  730.66 438.8 730.94 481.42 ;
     RECT  730.66 490.04 731.14 512.5 ;
     RECT  730.66 571.1 731.62 576.76 ;
     RECT  725.66 267.44 731.9 270.16 ;
     RECT  726.82 554.3 732.58 560.8 ;
     RECT  686.02 161.18 734.5 169.36 ;
     RECT  732.58 560.18 734.78 560.8 ;
     RECT  734.3 309.44 734.98 309.64 ;
     RECT  730.18 322.88 735.74 394.06 ;
     RECT  731.9 267.44 736.7 275.2 ;
     RECT  730.94 431.66 737.38 481.42 ;
     RECT  737.38 448.04 739.78 481.42 ;
     RECT  731.62 571.1 740.26 576.34 ;
     RECT  712.42 608.9 740.54 613.3 ;
     RECT  737.66 541.28 740.74 541.48 ;
     RECT  734.78 560.18 741.5 561.64 ;
     RECT  740.26 571.1 741.5 575.92 ;
     RECT  717.02 228.8 741.98 229 ;
     RECT  719.9 239.72 741.98 252.94 ;
     RECT  741.5 560.18 741.98 575.92 ;
     RECT  731.14 491.3 742.18 512.5 ;
     RECT  734.5 162.02 742.66 169.36 ;
     RECT  736.7 265.76 743.42 275.2 ;
     RECT  726.82 407.72 743.42 420.52 ;
     RECT  737.38 431.66 743.42 439 ;
     RECT  735.74 322.88 743.9 395.32 ;
     RECT  741.98 228.8 744.1 252.94 ;
     RECT  742.94 537.08 744.1 537.28 ;
     RECT  741.98 557.24 744.58 575.92 ;
     RECT  743.42 262.82 745.06 275.2 ;
     RECT  743.9 322.88 745.06 396.16 ;
     RECT  744.58 557.24 746.02 571.3 ;
     RECT  743.42 407.72 746.78 439 ;
     RECT  720.58 186.8 746.98 214.3 ;
     RECT  746.02 557.24 749.86 561.64 ;
     RECT  749.86 557.24 750.14 560.8 ;
     RECT  745.06 326.24 750.34 396.16 ;
     RECT  750.14 556.82 750.34 560.8 ;
     RECT  745.82 315.32 751.58 315.52 ;
     RECT  750.34 393.86 751.58 396.16 ;
     RECT  746.78 407.72 751.58 443.62 ;
     RECT  742.18 491.3 752.54 507.46 ;
     RECT  730.18 521.12 752.54 526.36 ;
     RECT  737.66 296.84 753.02 297.04 ;
     RECT  751.58 307.76 753.02 315.52 ;
     RECT  750.34 556.82 753.02 557.02 ;
     RECT  745.06 262.82 753.22 271 ;
     RECT  753.02 296.84 753.22 315.52 ;
     RECT  750.34 326.24 753.22 383.56 ;
     RECT  751.58 393.86 753.22 443.62 ;
     RECT  753.22 311.96 753.7 315.52 ;
     RECT  740.54 608.9 753.7 613.72 ;
     RECT  753.02 553.88 755.14 557.02 ;
     RECT  744.1 239.72 756.1 252.94 ;
     RECT  753.22 270.8 756.1 271 ;
     RECT  753.22 326.24 756.1 344.08 ;
     RECT  752.54 491.3 756.1 526.36 ;
     RECT  756.1 239.72 756.38 241.18 ;
     RECT  753.22 296.84 757.82 302.92 ;
     RECT  756.38 541.7 758.3 541.9 ;
     RECT  746.98 205.7 758.98 214.3 ;
     RECT  758.3 538.34 758.98 541.9 ;
     RECT  756.1 252.32 759.26 252.94 ;
     RECT  755.14 554.3 759.26 557.02 ;
     RECT  759.26 554.3 759.46 557.44 ;
     RECT  756.1 494.24 760.22 526.36 ;
     RECT  759.26 252.32 760.9 255.88 ;
     RECT  756.38 236.78 761.18 241.18 ;
     RECT  753.22 353.54 761.18 383.56 ;
     RECT  761.18 353.54 761.66 384.82 ;
     RECT  753.22 393.86 761.66 442.78 ;
     RECT  759.46 556.4 761.86 557.44 ;
     RECT  757.82 296.42 762.14 302.92 ;
     RECT  753.7 311.96 762.14 313.84 ;
     RECT  761.86 556.4 762.82 556.6 ;
     RECT  762.14 296.42 763.3 315.94 ;
     RECT  761.66 353.54 764.06 442.78 ;
     RECT  760.22 494.24 764.74 532.66 ;
     RECT  761.18 236.36 765.5 241.18 ;
     RECT  763.3 296.42 765.5 312.16 ;
     RECT  760.7 275 766.46 275.2 ;
     RECT  756.1 326.24 767.14 343.24 ;
     RECT  764.74 494.24 767.62 526.36 ;
     RECT  766.46 274.16 768.38 275.2 ;
     RECT  768.38 274.16 768.58 277.72 ;
     RECT  764.06 353.54 768.58 444.04 ;
     RECT  765.5 235.94 769.82 241.18 ;
     RECT  760.9 252.74 769.82 255.88 ;
     RECT  768.58 275 770.02 277.72 ;
     RECT  768.86 571.52 770.02 571.72 ;
     RECT  768.58 353.54 771.46 443.62 ;
     RECT  739.78 454.76 772.42 481.42 ;
     RECT  772.22 598.82 772.9 599.02 ;
     RECT  767.14 337.16 773.38 343.24 ;
     RECT  767.62 507.26 773.38 526.36 ;
     RECT  771.46 355.64 773.86 443.62 ;
     RECT  773.86 402.68 774.34 443.2 ;
     RECT  774.34 402.68 774.82 425.98 ;
     RECT  767.14 326.24 775.3 326.44 ;
     RECT  774.82 402.68 775.3 422.62 ;
     RECT  773.86 355.64 775.78 384.82 ;
     RECT  775.3 402.68 775.78 421.36 ;
     RECT  773.38 511.46 775.78 526.36 ;
     RECT  765.5 289.28 776.26 312.16 ;
     RECT  767.62 494.24 776.26 497.8 ;
     RECT  776.26 289.28 776.74 307.96 ;
     RECT  775.78 407.3 776.74 421.36 ;
     RECT  776.26 494.24 776.74 494.44 ;
     RECT  774.34 435.86 778.18 443.2 ;
     RECT  772.42 454.76 778.18 479.32 ;
     RECT  776.74 289.28 778.66 304.18 ;
     RECT  775.78 512.3 778.66 526.36 ;
     RECT  776.74 418.64 779.14 421.36 ;
     RECT  778.18 438.8 779.14 443.2 ;
     RECT  779.14 438.8 779.62 440.68 ;
     RECT  726.34 633.68 780.1 633.88 ;
     RECT  778.66 516.5 780.58 526.36 ;
     RECT  773.86 393.86 781.54 394.06 ;
     RECT  769.82 235.94 782.02 255.88 ;
     RECT  730.66 586.22 782.5 586.84 ;
     RECT  780.58 518.18 782.98 525.94 ;
     RECT  753.7 608.9 783.46 609.52 ;
     RECT  782.98 521.12 783.94 525.94 ;
     RECT  778.18 457.28 784.42 479.32 ;
     RECT  784.42 457.28 784.9 472.6 ;
     RECT  782.5 586.22 784.9 586.42 ;
     RECT  776.74 408.98 785.38 409.6 ;
     RECT  784.9 458.12 785.38 472.6 ;
     RECT  783.46 609.32 785.38 609.52 ;
     RECT  773.38 338 785.86 343.24 ;
     RECT  782.02 235.94 787.3 252.94 ;
     RECT  778.66 289.28 787.3 296.62 ;
     RECT  787.3 235.94 788.74 241.18 ;
     RECT  770.02 277.52 788.74 277.72 ;
     RECT  787.3 296.42 788.74 296.62 ;
     RECT  775.78 355.64 788.74 383.56 ;
     RECT  785.38 408.98 790.18 409.18 ;
     RECT  785.38 458.12 792.58 465.88 ;
     RECT  792.58 458.12 793.54 459.58 ;
     RECT  788.74 355.64 795.46 381.04 ;
     RECT  758.98 205.7 802.66 213.88 ;
     RECT  793.54 458.12 802.66 458.32 ;
     RECT  783.94 521.12 802.66 521.32 ;
     RECT  742.66 169.16 806.5 169.36 ;
     RECT  787.3 252.74 806.5 252.94 ;
     RECT  785.86 343.04 806.5 343.24 ;
     RECT  795.46 355.64 806.5 365.92 ;
     RECT  795.46 380.84 806.5 381.04 ;
     RECT  779.14 418.64 806.5 420.52 ;
     RECT  779.62 438.8 806.5 439 ;
     RECT  806.5 356.9 807.46 357.1 ;
     RECT  746.98 186.8 808.42 194.56 ;
     RECT  808.42 194.36 809.86 194.56 ;
     RECT  802.66 205.7 810.82 213.46 ;
     RECT  810.82 205.7 811.3 205.9 ;
     RECT  788.74 240.98 811.78 241.18 ;
    LAYER Metal5 ;
     RECT  389.18 51.14 389.38 51.98 ;
     RECT  543.74 62.06 543.94 79.7 ;
     RECT  559.1 72.14 559.3 79.7 ;
     RECT  497.18 77.18 497.38 80.74 ;
     RECT  362.3 62.9 362.5 81.38 ;
     RECT  413.66 86 413.86 86.42 ;
     RECT  388.22 51.98 389.38 89.78 ;
     RECT  499.58 84.74 499.78 92.3 ;
     RECT  543.74 79.7 559.3 92.72 ;
     RECT  490.46 92.3 499.78 93.56 ;
     RECT  543.74 92.72 562.18 95.24 ;
     RECT  471.26 95.24 471.46 96.08 ;
     RECT  381.02 89.78 389.38 97.76 ;
     RECT  362.3 81.38 369.22 100.7 ;
     RECT  466.46 96.08 471.46 102.8 ;
     RECT  543.74 95.24 571.78 104.06 ;
     RECT  527.9 101.12 528.1 105.74 ;
     RECT  438.62 64.16 438.82 107.42 ;
     RECT  452.06 101.12 452.26 107.42 ;
     RECT  527.9 105.74 530.5 107.84 ;
     RECT  402.62 88.52 402.82 111.2 ;
     RECT  413.66 86.42 417.22 111.2 ;
     RECT  402.62 111.2 417.22 115.18 ;
     RECT  541.82 104.06 571.78 115.3 ;
     RECT  381.02 97.76 392.74 125.26 ;
     RECT  402.62 115.18 413.86 126.74 ;
     RECT  424.22 126.32 424.42 126.74 ;
     RECT  487.58 93.56 499.78 130.3 ;
     RECT  355.58 100.7 369.22 130.52 ;
     RECT  519.26 107.84 530.5 130.52 ;
     RECT  346.94 130.52 369.22 130.72 ;
     RECT  381.02 125.26 389.38 133.46 ;
     RECT  487.58 130.3 490.66 134.08 ;
     RECT  365.66 130.72 369.22 134.5 ;
     RECT  346.94 130.72 355.78 134.92 ;
     RECT  380.54 133.46 389.38 143.96 ;
     RECT  438.62 107.42 452.26 144.38 ;
     RECT  402.62 126.74 424.42 149 ;
     RECT  487.58 134.08 489.7 149 ;
     RECT  355.58 134.92 355.78 149.42 ;
     RECT  365.66 134.5 365.86 149.42 ;
     RECT  503.42 139.76 503.62 150.88 ;
     RECT  402.14 149 424.42 151.1 ;
     RECT  355.58 149.42 365.86 151.3 ;
     RECT  483.74 149 489.7 152.98 ;
     RECT  402.14 151.1 425.38 153.2 ;
     RECT  438.62 144.38 453.22 153.2 ;
     RECT  483.74 152.98 487.78 155.08 ;
     RECT  519.26 130.52 530.98 157.4 ;
     RECT  518.78 157.4 530.98 157.82 ;
     RECT  542.3 115.3 571.78 157.82 ;
     RECT  518.78 157.82 571.78 160.76 ;
     RECT  510.14 160.76 571.78 162.22 ;
     RECT  483.74 155.08 483.94 163.7 ;
     RECT  464.06 102.8 471.46 165.8 ;
     RECT  483.26 163.7 483.94 165.8 ;
     RECT  500.06 158.66 500.26 167.9 ;
     RECT  361.82 151.3 365.86 168.52 ;
     RECT  663.26 164.12 663.46 168.74 ;
     RECT  348.86 167.06 349.06 172.52 ;
     RECT  277.34 150.26 277.54 175.88 ;
     RECT  291.26 145.64 291.46 175.88 ;
     RECT  464.06 165.8 483.94 175.88 ;
     RECT  575.42 175.04 575.62 175.88 ;
     RECT  402.14 153.2 453.22 176.3 ;
     RECT  464.06 175.88 486.82 176.3 ;
     RECT  402.14 176.3 486.82 179.66 ;
     RECT  498.62 167.9 500.26 179.66 ;
     RECT  619.58 111.2 619.78 187.22 ;
     RECT  380.54 143.96 392.26 191.84 ;
     RECT  402.14 179.66 500.26 191.84 ;
     RECT  674.3 183.44 674.5 194.78 ;
     RECT  663.26 168.74 663.94 198.56 ;
     RECT  674.3 194.78 683.14 198.56 ;
     RECT  380.54 191.84 500.26 199.82 ;
     RECT  510.14 162.22 562.18 199.82 ;
     RECT  365.66 168.52 365.86 200.66 ;
     RECT  619.58 187.22 623.62 201.28 ;
     RECT  619.58 201.28 622.18 201.5 ;
     RECT  277.34 175.88 291.46 201.92 ;
     RECT  663.26 198.56 683.14 201.92 ;
     RECT  348.86 172.52 353.38 206.12 ;
     RECT  659.9 201.92 683.14 206.12 ;
     RECT  575.42 175.88 577.06 206.54 ;
     RECT  587.9 88.52 588.1 206.54 ;
     RECT  659.9 206.12 683.62 208.64 ;
     RECT  365.66 200.66 369.22 209.06 ;
     RECT  380.54 199.82 562.18 209.06 ;
     RECT  614.78 201.5 622.18 210.52 ;
     RECT  651.26 208.64 683.62 213.68 ;
     RECT  365.66 209.06 562.18 214.52 ;
     RECT  651.26 213.68 684.1 215.36 ;
     RECT  237.98 209.48 238.18 216.2 ;
     RECT  614.78 210.52 619.78 217.88 ;
     RECT  575.42 206.54 588.1 222.08 ;
     RECT  223.1 201.92 223.3 223.34 ;
     RECT  195.26 201.5 195.46 224.6 ;
     RECT  206.3 201.5 206.5 224.6 ;
     RECT  158.3 178.82 158.5 228.8 ;
     RECT  277.34 201.92 294.34 229.84 ;
     RECT  365.66 214.52 564.1 230.26 ;
     RECT  3.26 183.02 3.46 231.32 ;
     RECT  543.74 230.26 564.1 231.52 ;
     RECT  545.18 231.52 564.1 233.2 ;
     RECT  651.26 215.36 687.46 237.2 ;
     RECT  697.82 231.32 698.02 237.2 ;
     RECT  277.34 229.84 289.06 239.08 ;
     RECT  613.82 217.88 619.78 240.76 ;
     RECT  158.3 228.8 162.34 243.92 ;
     RECT  575.42 222.08 596.74 244.34 ;
     RECT  365.66 230.26 533.38 244.76 ;
     RECT  545.18 233.2 557.38 244.76 ;
     RECT  639.26 243.5 639.46 246.86 ;
     RECT  195.26 224.6 206.5 247.06 ;
     RECT  721.82 183.86 722.02 248.12 ;
     RECT  277.34 239.08 285.7 251.68 ;
     RECT  343.1 206.12 353.38 251.68 ;
     RECT  195.26 247.06 201.22 252.1 ;
     RECT  343.1 251.68 343.3 252.1 ;
     RECT  365.66 244.76 557.38 252.1 ;
     RECT  613.82 240.76 617.38 252.1 ;
     RECT  651.26 237.2 698.02 252.1 ;
     RECT  218.78 223.34 223.3 254.84 ;
     RECT  555.26 252.1 557.38 254.84 ;
     RECT  569.18 244.34 596.74 254.84 ;
     RECT  636.86 246.86 639.46 256.52 ;
     RECT  555.26 254.84 596.74 258.2 ;
     RECT  632.06 256.52 639.46 258.62 ;
     RECT  651.26 252.1 683.62 258.62 ;
     RECT  632.06 258.62 683.62 261.56 ;
     RECT  555.26 258.2 601.06 261.98 ;
     RECT  610.94 254.42 611.14 261.98 ;
     RECT  195.26 252.1 195.46 262.18 ;
     RECT  622.94 261.56 683.62 264.7 ;
     RECT  632.06 264.7 683.62 269.54 ;
     RECT  695.42 252.1 698.02 269.54 ;
     RECT  353.18 251.68 353.38 270.16 ;
     RECT  365.66 252.1 545.38 270.16 ;
     RECT  373.82 270.16 545.38 271.22 ;
     RECT  555.26 261.98 611.14 271.22 ;
     RECT  285.5 251.68 285.7 273.32 ;
     RECT  1.82 231.32 3.46 273.74 ;
     RECT  743.42 228.38 743.62 275 ;
     RECT  285.5 273.32 289.06 276.88 ;
     RECT  373.82 271.22 611.14 276.88 ;
     RECT  632.06 269.54 698.02 277.72 ;
     RECT  680.54 277.72 698.02 282.76 ;
     RECT  632.06 277.72 670.18 282.98 ;
     RECT  0.38 273.74 3.46 284.66 ;
     RECT  235.58 216.2 238.18 285.08 ;
     RECT  309.02 278.78 309.22 285.08 ;
     RECT  211.1 254.84 223.3 285.28 ;
     RECT  683.42 282.76 698.02 291.8 ;
     RECT  683.42 291.8 705.22 293.9 ;
     RECT  389.18 276.88 555.46 294.1 ;
     RECT  409.34 294.1 555.46 294.52 ;
     RECT  389.18 294.1 398.5 294.94 ;
     RECT  453.98 294.52 555.46 295.16 ;
     RECT  453.98 295.16 558.34 295.58 ;
     RECT  624.86 282.98 670.18 296.42 ;
     RECT  373.82 276.88 374.98 296.84 ;
     RECT  758.78 214.1 758.98 297.04 ;
     RECT  158.3 243.92 170.02 302.3 ;
     RECT  573.5 276.88 611.14 302.3 ;
     RECT  622.46 296.42 670.18 302.3 ;
     RECT  756.38 300.2 756.58 302.72 ;
     RECT  158.3 302.3 177.22 304.4 ;
     RECT  235.58 285.08 246.34 304.6 ;
     RECT  285.5 276.88 285.7 305.44 ;
     RECT  211.1 285.28 218.98 306.08 ;
     RECT  573.5 302.3 670.18 307.76 ;
     RECT  235.58 304.6 244.42 311.12 ;
     RECT  573.5 307.76 672.58 311.54 ;
     RECT  683.42 293.9 706.18 311.54 ;
     RECT  453.98 295.58 563.14 311.96 ;
     RECT  573.5 311.54 706.18 311.96 ;
     RECT  373.82 296.84 375.94 312.16 ;
     RECT  755.42 302.72 756.58 313.84 ;
     RECT  409.34 294.52 443.14 315.52 ;
     RECT  453.98 311.96 706.18 316.9 ;
     RECT  734.3 275 743.62 316.9 ;
     RECT  208.7 306.08 218.98 317.84 ;
     RECT  231.26 311.12 244.42 317.84 ;
     RECT  158.3 304.4 181.06 319.52 ;
     RECT  716.06 248.12 722.02 319.52 ;
     RECT  734.3 316.9 742.18 319.52 ;
     RECT  373.82 312.16 374.98 327.28 ;
     RECT  389.18 294.94 396.58 327.28 ;
     RECT  409.34 315.52 441.22 328.76 ;
     RECT  453.98 316.9 705.7 328.76 ;
     RECT  756.38 313.84 756.58 330.44 ;
     RECT  208.7 317.84 244.42 337.36 ;
     RECT  158.3 319.52 183.94 338 ;
     RECT  409.34 328.76 705.7 338.2 ;
     RECT  753.02 330.44 756.58 338.42 ;
     RECT  329.66 292.64 329.86 341.78 ;
     RECT  329.66 341.78 331.3 342.2 ;
     RECT  289.34 308.6 289.54 342.4 ;
     RECT  210.14 337.36 244.42 347.86 ;
     RECT  450.14 338.2 705.7 349.76 ;
     RECT  158.3 338 184.42 352.7 ;
     RECT  716.06 319.52 742.18 352.7 ;
     RECT  753.02 338.42 767.14 352.7 ;
     RECT  450.14 349.76 706.18 360.68 ;
     RECT  716.06 352.7 767.14 360.68 ;
     RECT  96.86 345.56 97.06 363.62 ;
     RECT  409.34 338.2 438.82 364.66 ;
     RECT  110.3 353.54 110.5 365.3 ;
     RECT  151.58 352.7 184.42 368.66 ;
     RECT  211.1 347.86 244.42 368.66 ;
     RECT  211.1 368.66 252.58 372.22 ;
     RECT  431.42 364.66 438.82 372.22 ;
     RECT  133.34 171.68 133.54 372.44 ;
     RECT  133.34 372.44 134.02 376.84 ;
     RECT  151.58 368.66 185.38 380.62 ;
     RECT  450.14 360.68 767.14 387.98 ;
     RECT  777.98 375.8 778.18 387.98 ;
     RECT  329.66 342.2 334.66 388.18 ;
     RECT  438.62 372.22 438.82 389.24 ;
     RECT  450.14 387.98 778.18 389.24 ;
     RECT  409.34 364.66 417.22 394.9 ;
     RECT  267.26 365.72 267.46 395.12 ;
     RECT  438.62 389.24 778.18 397.84 ;
     RECT  438.62 397.84 490.66 402.46 ;
     RECT  334.46 388.18 334.66 403.1 ;
     RECT  152.54 380.62 185.38 403.3 ;
     RECT  152.54 403.3 158.5 405.82 ;
     RECT  450.14 402.46 490.66 412.76 ;
     RECT  505.82 397.84 778.18 412.76 ;
     RECT  293.18 365.72 293.38 420.94 ;
     RECT  211.1 372.22 244.42 421.16 ;
     RECT  169.82 403.3 185.38 422.62 ;
     RECT  156.38 405.82 158.5 423.04 ;
     RECT  265.82 395.12 267.46 423.04 ;
     RECT  180.86 422.62 185.38 424.72 ;
     RECT  156.86 423.04 158.5 427.24 ;
     RECT  92.54 363.62 97.06 428.92 ;
     RECT  389.18 327.28 396.1 431.86 ;
     RECT  158.3 427.24 158.5 432.28 ;
     RECT  185.18 424.72 185.38 435.64 ;
     RECT  450.14 412.76 778.18 438.58 ;
     RECT  211.1 421.16 254.02 440.26 ;
     RECT  395.9 431.86 396.1 444.26 ;
     RECT  469.34 438.58 778.18 444.88 ;
     RECT  469.34 444.88 565.54 446.56 ;
     RECT  471.26 446.56 565.54 450.76 ;
     RECT  325.82 403.1 334.66 451.6 ;
     RECT  471.26 450.76 563.62 452.44 ;
     RECT  575.42 444.88 778.18 452.44 ;
     RECT  438.62 402.46 438.82 453.5 ;
     RECT  450.14 438.58 457.54 453.5 ;
     RECT  500.54 452.44 563.62 453.7 ;
     RECT  575.9 452.44 778.18 454.54 ;
     RECT  527.9 453.7 563.62 455.38 ;
     RECT  500.54 453.7 518.02 455.8 ;
     RECT  212.06 440.26 254.02 456.02 ;
     RECT  438.62 453.5 457.54 460.22 ;
     RECT  202.46 456.02 254.02 460.64 ;
     RECT  265.82 423.04 266.02 460.64 ;
     RECT  202.46 460.64 266.02 461.26 ;
     RECT  63.74 455.6 63.94 462.32 ;
     RECT  282.14 459.38 282.34 462.32 ;
     RECT  471.26 452.44 490.66 463.16 ;
     RECT  59.42 462.32 63.94 464 ;
     RECT  59.42 464 65.38 464.62 ;
     RECT  438.62 460.22 458.02 464.84 ;
     RECT  468.38 463.16 490.66 464.84 ;
     RECT  605.18 454.54 778.18 466.72 ;
     RECT  438.62 464.84 490.66 466.94 ;
     RECT  500.54 455.8 514.18 466.94 ;
     RECT  527.9 455.38 562.66 467.78 ;
     RECT  309.02 285.08 311.14 468.1 ;
     RECT  575.9 454.54 595.3 468.2 ;
     RECT  605.18 466.72 772.42 468.2 ;
     RECT  438.62 466.94 514.18 469.66 ;
     RECT  110.3 365.3 117.22 470.5 ;
     RECT  468.38 469.66 514.18 470.92 ;
     RECT  527.9 467.78 565.54 471.56 ;
     RECT  575.9 468.2 772.42 471.56 ;
     RECT  169.82 422.62 170.02 472.6 ;
     RECT  61.82 464.62 65.38 474.5 ;
     RECT  471.26 470.92 514.18 475.96 ;
     RECT  346.46 393.44 346.66 476.18 ;
     RECT  438.62 469.66 457.54 476.8 ;
     RECT  133.82 376.84 134.02 477.22 ;
     RECT  346.46 476.18 352.42 478.9 ;
     RECT  500.54 475.96 514.18 481.64 ;
     RECT  527.9 471.56 772.42 481.64 ;
     RECT  446.3 476.8 457.54 481.84 ;
     RECT  59.42 474.5 65.38 482.26 ;
     RECT  334.46 451.6 334.66 482.68 ;
     RECT  202.46 461.26 227.14 483.94 ;
     RECT  243.26 461.26 266.02 483.94 ;
     RECT  117.02 470.5 117.22 485.2 ;
     RECT  61.82 482.26 65.38 485.62 ;
     RECT  203.42 483.94 227.14 489.4 ;
     RECT  450.14 481.84 457.54 492.34 ;
     RECT  500.54 481.64 772.42 492.98 ;
     RECT  309.02 468.1 310.66 496.76 ;
     RECT  500.54 492.98 776.74 497.38 ;
     RECT  346.46 478.9 346.66 498.86 ;
     RECT  432.86 490.04 433.06 500.96 ;
     RECT  471.26 475.96 490.66 501.16 ;
     RECT  61.82 485.62 64.42 502 ;
     RECT  395.9 444.26 398.5 504.1 ;
     RECT  226.94 489.4 227.14 504.52 ;
     RECT  409.34 394.9 413.86 504.52 ;
     RECT  500.54 497.38 772.42 506.2 ;
     RECT  471.26 501.16 471.94 509.14 ;
     RECT  432.86 500.96 440.74 512.3 ;
     RECT  305.66 496.76 310.66 517.34 ;
     RECT  302.3 517.34 310.66 518.38 ;
     RECT  49.82 516.92 50.02 519.86 ;
     RECT  525.5 506.2 772.42 520.06 ;
     RECT  471.26 509.14 471.46 528.04 ;
     RECT  413.66 504.52 413.86 528.26 ;
     RECT  528.38 520.06 772.42 532.66 ;
     RECT  44.54 519.86 50.02 534.56 ;
     RECT  203.42 489.4 216.58 534.56 ;
     RECT  457.34 492.34 457.54 535.6 ;
     RECT  481.82 501.16 490.66 535.6 ;
     RECT  528.38 532.66 758.5 538.54 ;
     RECT  78.62 478.7 78.82 538.96 ;
     RECT  339.74 498.86 346.66 538.96 ;
     RECT  40.7 534.56 50.02 539.38 ;
     RECT  413.66 528.26 414.34 539.8 ;
     RECT  528.38 538.54 757.54 541.9 ;
     RECT  96.86 428.92 97.06 542.32 ;
     RECT  40.7 539.38 44.74 544.84 ;
     RECT  40.7 544.84 40.9 546.52 ;
     RECT  200.54 534.56 216.58 546.52 ;
     RECT  528.38 541.9 753.22 546.52 ;
     RECT  595.1 546.52 753.22 551.14 ;
     RECT  64.22 502 64.42 552.4 ;
     RECT  158.3 541.28 158.5 553.04 ;
     RECT  528.38 546.52 584.74 553.66 ;
     RECT  302.78 518.38 310.66 554.08 ;
     RECT  200.54 546.52 200.74 554.3 ;
     RECT  212.06 546.52 216.58 554.5 ;
     RECT  626.3 551.14 753.22 554.5 ;
     RECT  629.18 554.5 753.22 556.6 ;
     RECT  490.46 535.6 490.66 557.24 ;
     RECT  500.54 506.2 514.18 557.24 ;
     RECT  595.1 551.14 615.94 558.28 ;
     RECT  551.9 553.66 584.74 560.8 ;
     RECT  629.18 556.6 746.02 561.22 ;
     RECT  528.38 553.66 541.54 562.06 ;
     RECT  552.86 560.8 584.74 562.06 ;
     RECT  490.46 557.24 514.18 564.16 ;
     RECT  158.3 553.04 159.46 564.8 ;
     RECT  629.18 561.22 708.1 567.32 ;
     RECT  606.62 558.28 615.94 568.16 ;
     RECT  626.78 567.32 708.1 568.16 ;
     RECT  490.46 564.16 490.66 568.7 ;
     RECT  500.54 564.16 514.18 568.7 ;
     RECT  489.98 568.7 490.66 568.9 ;
     RECT  553.34 562.06 584.74 570.04 ;
     RECT  719.42 561.22 746.02 571.3 ;
     RECT  432.86 512.3 443.14 571.94 ;
     RECT  528.38 562.06 537.22 574.24 ;
     RECT  595.1 558.28 596.74 574.46 ;
     RECT  606.62 568.16 708.1 574.46 ;
     RECT  595.1 574.46 708.1 574.66 ;
     RECT  332.54 554.3 332.74 576.34 ;
     RECT  620.06 574.66 708.1 576.34 ;
     RECT  719.42 571.3 745.06 576.34 ;
     RECT  620.06 576.34 695.62 577.18 ;
     RECT  719.42 576.34 730.66 577.18 ;
     RECT  243.26 483.94 260.26 577.6 ;
     RECT  535.1 574.24 537.22 578.44 ;
     RECT  620.06 577.18 694.66 578.44 ;
     RECT  282.14 462.32 289.54 579.28 ;
     RECT  721.82 577.18 730.66 579.28 ;
     RECT  620.06 578.44 633.7 579.7 ;
     RECT  414.14 539.8 414.34 580.34 ;
     RECT  197.66 554.3 200.74 580.54 ;
     RECT  645.5 578.44 694.66 580.54 ;
     RECT  645.5 580.54 693.22 580.96 ;
     RECT  595.1 574.66 609.7 583.06 ;
     RECT  535.1 578.44 535.3 584.32 ;
     RECT  693.02 580.96 693.22 584.74 ;
     RECT  705.98 576.34 708.1 586 ;
     RECT  553.34 570.04 582.82 587.26 ;
     RECT  620.06 579.7 631.78 587.26 ;
     RECT  143.42 557.24 143.62 587.48 ;
     RECT  283.1 579.28 289.54 587.68 ;
     RECT  500.54 568.7 514.66 587.68 ;
     RECT  555.26 587.26 582.82 587.68 ;
     RECT  707.9 586 708.1 587.68 ;
     RECT  631.58 587.26 631.78 588.94 ;
     RECT  505.82 587.68 514.66 591.46 ;
     RECT  140.54 587.48 143.62 591.68 ;
     RECT  158.3 564.8 169.06 591.88 ;
     RECT  243.26 577.6 243.46 591.88 ;
     RECT  605.18 583.06 609.7 594.4 ;
     RECT  159.26 591.88 169.06 595.24 ;
     RECT  605.18 594.4 608.74 596.5 ;
     RECT  572.54 587.68 582.82 596.92 ;
     RECT  514.46 591.46 514.66 598.18 ;
     RECT  414.14 580.34 415.78 598.82 ;
     RECT  721.82 579.28 722.02 599.02 ;
     RECT  772.22 532.66 772.42 599.02 ;
     RECT  645.5 580.96 677.86 599.44 ;
     RECT  255.26 577.6 260.26 600.08 ;
     RECT  645.5 599.44 670.66 602.38 ;
     RECT  408.38 598.82 415.78 602.6 ;
     RECT  489.98 568.9 490.18 602.8 ;
     RECT  645.5 602.38 669.22 604.06 ;
     RECT  395.9 504.1 396.1 604.7 ;
     RECT  405.98 602.6 415.78 604.7 ;
     RECT  427.1 571.94 443.14 604.7 ;
     RECT  0.38 284.66 3.94 605.32 ;
     RECT  555.26 587.68 560.26 606.58 ;
     RECT  608.54 596.5 608.74 606.58 ;
     RECT  395.9 604.7 415.78 606.8 ;
     RECT  426.14 604.7 443.14 606.8 ;
     RECT  575.42 596.92 582.82 607 ;
     RECT  595.1 583.06 595.3 610.78 ;
     RECT  395.9 606.8 443.14 611.84 ;
     RECT  395.9 611.84 446.5 612.88 ;
     RECT  744.86 576.34 745.06 613.3 ;
     RECT  575.42 607 580.9 614.36 ;
     RECT  165.98 595.24 169.06 614.56 ;
     RECT  283.1 587.68 284.26 614.56 ;
     RECT  558.62 606.58 560.26 614.56 ;
     RECT  658.94 604.06 669.22 614.56 ;
     RECT  373.82 327.28 374.02 617.5 ;
     RECT  65.18 595.04 65.38 617.92 ;
     RECT  645.5 604.06 647.14 617.92 ;
     RECT  402.62 612.88 446.5 619.4 ;
     RECT  658.94 614.56 668.74 620.44 ;
     RECT  560.06 614.56 560.26 620.86 ;
     RECT  255.26 600.08 263.14 621.28 ;
     RECT  166.94 614.56 169.06 622.12 ;
     RECT  99.26 591.68 99.46 622.34 ;
     RECT  646.94 617.92 647.14 624.64 ;
     RECT  98.78 622.34 99.46 624.86 ;
     RECT  322.46 512.3 322.66 625.06 ;
     RECT  668.54 620.44 668.74 625.9 ;
     RECT  0.38 605.32 2.98 628 ;
     RECT  402.62 619.4 454.66 628.84 ;
     RECT  137.66 591.68 143.62 629.68 ;
     RECT  216.38 554.5 216.58 629.68 ;
     RECT  574.46 614.36 580.9 630.74 ;
     RECT  402.62 628.84 443.62 632.62 ;
     RECT  626.3 621.08 626.5 632.84 ;
     RECT  137.66 629.68 141.22 633.04 ;
     RECT  453.98 628.84 454.66 636.2 ;
     RECT  402.62 632.62 422.98 636.4 ;
     RECT  200.54 580.54 200.74 637.46 ;
     RECT  574.46 630.74 581.38 637.66 ;
     RECT  414.62 636.4 422.98 640.6 ;
     RECT  575.42 637.66 581.38 640.82 ;
     RECT  414.62 640.6 415.3 641.02 ;
     RECT  453.98 636.2 455.62 641.44 ;
     RECT  453.98 641.44 454.66 641.86 ;
     RECT  705.98 638.72 706.18 644.6 ;
     RECT  453.98 641.86 454.18 644.8 ;
     RECT  434.3 632.62 443.62 645.22 ;
     RECT  402.62 636.4 402.82 645.64 ;
     RECT  200.54 637.46 203.14 647.74 ;
     RECT  575.42 640.82 582.82 648.16 ;
     RECT  140.54 633.04 141.22 649.84 ;
     RECT  97.34 624.86 99.46 652.36 ;
     RECT  98.78 652.36 99.46 652.78 ;
     RECT  698.3 644.6 706.18 654.88 ;
     RECT  415.1 641.02 415.3 655.3 ;
     RECT  434.3 645.22 441.7 655.3 ;
     RECT  99.26 652.78 99.46 655.72 ;
     RECT  167.9 622.12 169.06 657.82 ;
     RECT  346.46 538.96 346.66 659.92 ;
     RECT  606.14 643.76 606.34 660.56 ;
     RECT  625.34 632.84 626.5 661.82 ;
     RECT  606.14 660.56 608.26 662.66 ;
     RECT  167.9 657.82 168.1 663.28 ;
     RECT  597.98 662.66 608.26 663.28 ;
     RECT  309.02 554.08 310.66 663.7 ;
     RECT  141.02 649.84 141.22 667.06 ;
     RECT  284.06 614.56 284.26 671.26 ;
     RECT  310.46 663.7 310.66 674.62 ;
     RECT  581.18 648.16 582.82 676.72 ;
     RECT  255.26 621.28 255.46 677.98 ;
     RECT  200.54 647.74 200.74 683.86 ;
     RECT  625.34 661.82 629.86 684.92 ;
     RECT  597.98 663.28 606.34 691.22 ;
     RECT  125.18 659.3 125.38 691.42 ;
     RECT  625.34 684.92 635.62 697.72 ;
     RECT  594.62 691.22 606.34 709.06 ;
     RECT  582.62 676.72 582.82 712.42 ;
     RECT  0.38 628 2.5 721.24 ;
     RECT  565.82 716.42 566.02 726.92 ;
     RECT  565.82 726.92 570.82 734.48 ;
     RECT  594.62 709.06 594.82 735.1 ;
     RECT  565.82 734.48 571.78 742.66 ;
     RECT  625.34 697.72 629.86 743.08 ;
     RECT  0.38 721.24 1.54 746.44 ;
     RECT  653.66 747.5 653.86 754 ;
     RECT  565.82 742.66 568.42 756.32 ;
     RECT  698.3 654.88 698.5 763.66 ;
     RECT  0.38 746.44 0.58 764.08 ;
     RECT  565.34 756.32 568.42 769.54 ;
     RECT  568.22 769.54 568.42 776.26 ;
     RECT  625.34 743.08 625.54 815.74 ;
     RECT  606.14 709.06 606.34 834.22 ;
  END
END cve2_core
END LIBRARY
