//Latest Update Date: 12th Nov, 2025
//Owner: B Nithin Reddy

//Interface
interface dff_if;
  
  logic clk;
  logic rst;
  logic din;
  logic dout;
  
endinterface
