module dm_top (clk_i,
    debug_req_o,
    dmactive_o,
    dmi_req_i_0_,
    dmi_req_i_10_,
    dmi_req_i_11_,
    dmi_req_i_12_,
    dmi_req_i_13_,
    dmi_req_i_14_,
    dmi_req_i_15_,
    dmi_req_i_16_,
    dmi_req_i_17_,
    dmi_req_i_18_,
    dmi_req_i_19_,
    dmi_req_i_1_,
    dmi_req_i_20_,
    dmi_req_i_21_,
    dmi_req_i_22_,
    dmi_req_i_23_,
    dmi_req_i_24_,
    dmi_req_i_25_,
    dmi_req_i_26_,
    dmi_req_i_27_,
    dmi_req_i_28_,
    dmi_req_i_29_,
    dmi_req_i_2_,
    dmi_req_i_30_,
    dmi_req_i_31_,
    dmi_req_i_32_,
    dmi_req_i_33_,
    dmi_req_i_34_,
    dmi_req_i_35_,
    dmi_req_i_36_,
    dmi_req_i_37_,
    dmi_req_i_38_,
    dmi_req_i_39_,
    dmi_req_i_3_,
    dmi_req_i_40_,
    dmi_req_i_4_,
    dmi_req_i_5_,
    dmi_req_i_6_,
    dmi_req_i_7_,
    dmi_req_i_8_,
    dmi_req_i_9_,
    dmi_req_ready_o,
    dmi_req_valid_i,
    dmi_resp_o_0_,
    dmi_resp_o_10_,
    dmi_resp_o_11_,
    dmi_resp_o_12_,
    dmi_resp_o_13_,
    dmi_resp_o_14_,
    dmi_resp_o_15_,
    dmi_resp_o_16_,
    dmi_resp_o_17_,
    dmi_resp_o_18_,
    dmi_resp_o_19_,
    dmi_resp_o_1_,
    dmi_resp_o_20_,
    dmi_resp_o_21_,
    dmi_resp_o_22_,
    dmi_resp_o_23_,
    dmi_resp_o_24_,
    dmi_resp_o_25_,
    dmi_resp_o_26_,
    dmi_resp_o_27_,
    dmi_resp_o_28_,
    dmi_resp_o_29_,
    dmi_resp_o_2_,
    dmi_resp_o_30_,
    dmi_resp_o_31_,
    dmi_resp_o_32_,
    dmi_resp_o_33_,
    dmi_resp_o_3_,
    dmi_resp_o_4_,
    dmi_resp_o_5_,
    dmi_resp_o_6_,
    dmi_resp_o_7_,
    dmi_resp_o_8_,
    dmi_resp_o_9_,
    dmi_resp_ready_i,
    dmi_resp_valid_o,
    dmi_rst_ni,
    hartinfo_i_0_,
    hartinfo_i_10_,
    hartinfo_i_11_,
    hartinfo_i_12_,
    hartinfo_i_13_,
    hartinfo_i_14_,
    hartinfo_i_15_,
    hartinfo_i_16_,
    hartinfo_i_17_,
    hartinfo_i_18_,
    hartinfo_i_19_,
    hartinfo_i_1_,
    hartinfo_i_20_,
    hartinfo_i_21_,
    hartinfo_i_22_,
    hartinfo_i_23_,
    hartinfo_i_24_,
    hartinfo_i_25_,
    hartinfo_i_26_,
    hartinfo_i_27_,
    hartinfo_i_28_,
    hartinfo_i_29_,
    hartinfo_i_2_,
    hartinfo_i_30_,
    hartinfo_i_31_,
    hartinfo_i_3_,
    hartinfo_i_4_,
    hartinfo_i_5_,
    hartinfo_i_6_,
    hartinfo_i_7_,
    hartinfo_i_8_,
    hartinfo_i_9_,
    master_add_o_0_,
    master_add_o_10_,
    master_add_o_11_,
    master_add_o_12_,
    master_add_o_13_,
    master_add_o_14_,
    master_add_o_15_,
    master_add_o_16_,
    master_add_o_17_,
    master_add_o_18_,
    master_add_o_19_,
    master_add_o_1_,
    master_add_o_20_,
    master_add_o_21_,
    master_add_o_22_,
    master_add_o_23_,
    master_add_o_24_,
    master_add_o_25_,
    master_add_o_26_,
    master_add_o_27_,
    master_add_o_28_,
    master_add_o_29_,
    master_add_o_2_,
    master_add_o_30_,
    master_add_o_31_,
    master_add_o_3_,
    master_add_o_4_,
    master_add_o_5_,
    master_add_o_6_,
    master_add_o_7_,
    master_add_o_8_,
    master_add_o_9_,
    master_be_o_0_,
    master_be_o_1_,
    master_be_o_2_,
    master_be_o_3_,
    master_gnt_i,
    master_r_err_i,
    master_r_other_err_i,
    master_r_rdata_i_0_,
    master_r_rdata_i_10_,
    master_r_rdata_i_11_,
    master_r_rdata_i_12_,
    master_r_rdata_i_13_,
    master_r_rdata_i_14_,
    master_r_rdata_i_15_,
    master_r_rdata_i_16_,
    master_r_rdata_i_17_,
    master_r_rdata_i_18_,
    master_r_rdata_i_19_,
    master_r_rdata_i_1_,
    master_r_rdata_i_20_,
    master_r_rdata_i_21_,
    master_r_rdata_i_22_,
    master_r_rdata_i_23_,
    master_r_rdata_i_24_,
    master_r_rdata_i_25_,
    master_r_rdata_i_26_,
    master_r_rdata_i_27_,
    master_r_rdata_i_28_,
    master_r_rdata_i_29_,
    master_r_rdata_i_2_,
    master_r_rdata_i_30_,
    master_r_rdata_i_31_,
    master_r_rdata_i_3_,
    master_r_rdata_i_4_,
    master_r_rdata_i_5_,
    master_r_rdata_i_6_,
    master_r_rdata_i_7_,
    master_r_rdata_i_8_,
    master_r_rdata_i_9_,
    master_r_valid_i,
    master_req_o,
    master_wdata_o_0_,
    master_wdata_o_10_,
    master_wdata_o_11_,
    master_wdata_o_12_,
    master_wdata_o_13_,
    master_wdata_o_14_,
    master_wdata_o_15_,
    master_wdata_o_16_,
    master_wdata_o_17_,
    master_wdata_o_18_,
    master_wdata_o_19_,
    master_wdata_o_1_,
    master_wdata_o_20_,
    master_wdata_o_21_,
    master_wdata_o_22_,
    master_wdata_o_23_,
    master_wdata_o_24_,
    master_wdata_o_25_,
    master_wdata_o_26_,
    master_wdata_o_27_,
    master_wdata_o_28_,
    master_wdata_o_29_,
    master_wdata_o_2_,
    master_wdata_o_30_,
    master_wdata_o_31_,
    master_wdata_o_3_,
    master_wdata_o_4_,
    master_wdata_o_5_,
    master_wdata_o_6_,
    master_wdata_o_7_,
    master_wdata_o_8_,
    master_wdata_o_9_,
    master_we_o,
    ndmreset_ack_i,
    ndmreset_o,
    next_dm_addr_i_0_,
    next_dm_addr_i_10_,
    next_dm_addr_i_11_,
    next_dm_addr_i_12_,
    next_dm_addr_i_13_,
    next_dm_addr_i_14_,
    next_dm_addr_i_15_,
    next_dm_addr_i_16_,
    next_dm_addr_i_17_,
    next_dm_addr_i_18_,
    next_dm_addr_i_19_,
    next_dm_addr_i_1_,
    next_dm_addr_i_20_,
    next_dm_addr_i_21_,
    next_dm_addr_i_22_,
    next_dm_addr_i_23_,
    next_dm_addr_i_24_,
    next_dm_addr_i_25_,
    next_dm_addr_i_26_,
    next_dm_addr_i_27_,
    next_dm_addr_i_28_,
    next_dm_addr_i_29_,
    next_dm_addr_i_2_,
    next_dm_addr_i_30_,
    next_dm_addr_i_31_,
    next_dm_addr_i_3_,
    next_dm_addr_i_4_,
    next_dm_addr_i_5_,
    next_dm_addr_i_6_,
    next_dm_addr_i_7_,
    next_dm_addr_i_8_,
    next_dm_addr_i_9_,
    rst_ni,
    slave_addr_i_0_,
    slave_addr_i_10_,
    slave_addr_i_11_,
    slave_addr_i_12_,
    slave_addr_i_13_,
    slave_addr_i_14_,
    slave_addr_i_15_,
    slave_addr_i_16_,
    slave_addr_i_17_,
    slave_addr_i_18_,
    slave_addr_i_19_,
    slave_addr_i_1_,
    slave_addr_i_20_,
    slave_addr_i_21_,
    slave_addr_i_22_,
    slave_addr_i_23_,
    slave_addr_i_24_,
    slave_addr_i_25_,
    slave_addr_i_26_,
    slave_addr_i_27_,
    slave_addr_i_28_,
    slave_addr_i_29_,
    slave_addr_i_2_,
    slave_addr_i_30_,
    slave_addr_i_31_,
    slave_addr_i_3_,
    slave_addr_i_4_,
    slave_addr_i_5_,
    slave_addr_i_6_,
    slave_addr_i_7_,
    slave_addr_i_8_,
    slave_addr_i_9_,
    slave_be_i_0_,
    slave_be_i_1_,
    slave_be_i_2_,
    slave_be_i_3_,
    slave_rdata_o_0_,
    slave_rdata_o_10_,
    slave_rdata_o_11_,
    slave_rdata_o_12_,
    slave_rdata_o_13_,
    slave_rdata_o_14_,
    slave_rdata_o_15_,
    slave_rdata_o_16_,
    slave_rdata_o_17_,
    slave_rdata_o_18_,
    slave_rdata_o_19_,
    slave_rdata_o_1_,
    slave_rdata_o_20_,
    slave_rdata_o_21_,
    slave_rdata_o_22_,
    slave_rdata_o_23_,
    slave_rdata_o_24_,
    slave_rdata_o_25_,
    slave_rdata_o_26_,
    slave_rdata_o_27_,
    slave_rdata_o_28_,
    slave_rdata_o_29_,
    slave_rdata_o_2_,
    slave_rdata_o_30_,
    slave_rdata_o_31_,
    slave_rdata_o_3_,
    slave_rdata_o_4_,
    slave_rdata_o_5_,
    slave_rdata_o_6_,
    slave_rdata_o_7_,
    slave_rdata_o_8_,
    slave_rdata_o_9_,
    slave_req_i,
    slave_wdata_i_0_,
    slave_wdata_i_10_,
    slave_wdata_i_11_,
    slave_wdata_i_12_,
    slave_wdata_i_13_,
    slave_wdata_i_14_,
    slave_wdata_i_15_,
    slave_wdata_i_16_,
    slave_wdata_i_17_,
    slave_wdata_i_18_,
    slave_wdata_i_19_,
    slave_wdata_i_1_,
    slave_wdata_i_20_,
    slave_wdata_i_21_,
    slave_wdata_i_22_,
    slave_wdata_i_23_,
    slave_wdata_i_24_,
    slave_wdata_i_25_,
    slave_wdata_i_26_,
    slave_wdata_i_27_,
    slave_wdata_i_28_,
    slave_wdata_i_29_,
    slave_wdata_i_2_,
    slave_wdata_i_30_,
    slave_wdata_i_31_,
    slave_wdata_i_3_,
    slave_wdata_i_4_,
    slave_wdata_i_5_,
    slave_wdata_i_6_,
    slave_wdata_i_7_,
    slave_wdata_i_8_,
    slave_wdata_i_9_,
    slave_we_i,
    testmode_i,
    unavailable_i);
 input clk_i;
 output debug_req_o;
 output dmactive_o;
 input dmi_req_i_0_;
 input dmi_req_i_10_;
 input dmi_req_i_11_;
 input dmi_req_i_12_;
 input dmi_req_i_13_;
 input dmi_req_i_14_;
 input dmi_req_i_15_;
 input dmi_req_i_16_;
 input dmi_req_i_17_;
 input dmi_req_i_18_;
 input dmi_req_i_19_;
 input dmi_req_i_1_;
 input dmi_req_i_20_;
 input dmi_req_i_21_;
 input dmi_req_i_22_;
 input dmi_req_i_23_;
 input dmi_req_i_24_;
 input dmi_req_i_25_;
 input dmi_req_i_26_;
 input dmi_req_i_27_;
 input dmi_req_i_28_;
 input dmi_req_i_29_;
 input dmi_req_i_2_;
 input dmi_req_i_30_;
 input dmi_req_i_31_;
 input dmi_req_i_32_;
 input dmi_req_i_33_;
 input dmi_req_i_34_;
 input dmi_req_i_35_;
 input dmi_req_i_36_;
 input dmi_req_i_37_;
 input dmi_req_i_38_;
 input dmi_req_i_39_;
 input dmi_req_i_3_;
 input dmi_req_i_40_;
 input dmi_req_i_4_;
 input dmi_req_i_5_;
 input dmi_req_i_6_;
 input dmi_req_i_7_;
 input dmi_req_i_8_;
 input dmi_req_i_9_;
 output dmi_req_ready_o;
 input dmi_req_valid_i;
 output dmi_resp_o_0_;
 output dmi_resp_o_10_;
 output dmi_resp_o_11_;
 output dmi_resp_o_12_;
 output dmi_resp_o_13_;
 output dmi_resp_o_14_;
 output dmi_resp_o_15_;
 output dmi_resp_o_16_;
 output dmi_resp_o_17_;
 output dmi_resp_o_18_;
 output dmi_resp_o_19_;
 output dmi_resp_o_1_;
 output dmi_resp_o_20_;
 output dmi_resp_o_21_;
 output dmi_resp_o_22_;
 output dmi_resp_o_23_;
 output dmi_resp_o_24_;
 output dmi_resp_o_25_;
 output dmi_resp_o_26_;
 output dmi_resp_o_27_;
 output dmi_resp_o_28_;
 output dmi_resp_o_29_;
 output dmi_resp_o_2_;
 output dmi_resp_o_30_;
 output dmi_resp_o_31_;
 output dmi_resp_o_32_;
 output dmi_resp_o_33_;
 output dmi_resp_o_3_;
 output dmi_resp_o_4_;
 output dmi_resp_o_5_;
 output dmi_resp_o_6_;
 output dmi_resp_o_7_;
 output dmi_resp_o_8_;
 output dmi_resp_o_9_;
 input dmi_resp_ready_i;
 output dmi_resp_valid_o;
 input dmi_rst_ni;
 input hartinfo_i_0_;
 input hartinfo_i_10_;
 input hartinfo_i_11_;
 input hartinfo_i_12_;
 input hartinfo_i_13_;
 input hartinfo_i_14_;
 input hartinfo_i_15_;
 input hartinfo_i_16_;
 input hartinfo_i_17_;
 input hartinfo_i_18_;
 input hartinfo_i_19_;
 input hartinfo_i_1_;
 input hartinfo_i_20_;
 input hartinfo_i_21_;
 input hartinfo_i_22_;
 input hartinfo_i_23_;
 input hartinfo_i_24_;
 input hartinfo_i_25_;
 input hartinfo_i_26_;
 input hartinfo_i_27_;
 input hartinfo_i_28_;
 input hartinfo_i_29_;
 input hartinfo_i_2_;
 input hartinfo_i_30_;
 input hartinfo_i_31_;
 input hartinfo_i_3_;
 input hartinfo_i_4_;
 input hartinfo_i_5_;
 input hartinfo_i_6_;
 input hartinfo_i_7_;
 input hartinfo_i_8_;
 input hartinfo_i_9_;
 output master_add_o_0_;
 output master_add_o_10_;
 output master_add_o_11_;
 output master_add_o_12_;
 output master_add_o_13_;
 output master_add_o_14_;
 output master_add_o_15_;
 output master_add_o_16_;
 output master_add_o_17_;
 output master_add_o_18_;
 output master_add_o_19_;
 output master_add_o_1_;
 output master_add_o_20_;
 output master_add_o_21_;
 output master_add_o_22_;
 output master_add_o_23_;
 output master_add_o_24_;
 output master_add_o_25_;
 output master_add_o_26_;
 output master_add_o_27_;
 output master_add_o_28_;
 output master_add_o_29_;
 output master_add_o_2_;
 output master_add_o_30_;
 output master_add_o_31_;
 output master_add_o_3_;
 output master_add_o_4_;
 output master_add_o_5_;
 output master_add_o_6_;
 output master_add_o_7_;
 output master_add_o_8_;
 output master_add_o_9_;
 output master_be_o_0_;
 output master_be_o_1_;
 output master_be_o_2_;
 output master_be_o_3_;
 input master_gnt_i;
 input master_r_err_i;
 input master_r_other_err_i;
 input master_r_rdata_i_0_;
 input master_r_rdata_i_10_;
 input master_r_rdata_i_11_;
 input master_r_rdata_i_12_;
 input master_r_rdata_i_13_;
 input master_r_rdata_i_14_;
 input master_r_rdata_i_15_;
 input master_r_rdata_i_16_;
 input master_r_rdata_i_17_;
 input master_r_rdata_i_18_;
 input master_r_rdata_i_19_;
 input master_r_rdata_i_1_;
 input master_r_rdata_i_20_;
 input master_r_rdata_i_21_;
 input master_r_rdata_i_22_;
 input master_r_rdata_i_23_;
 input master_r_rdata_i_24_;
 input master_r_rdata_i_25_;
 input master_r_rdata_i_26_;
 input master_r_rdata_i_27_;
 input master_r_rdata_i_28_;
 input master_r_rdata_i_29_;
 input master_r_rdata_i_2_;
 input master_r_rdata_i_30_;
 input master_r_rdata_i_31_;
 input master_r_rdata_i_3_;
 input master_r_rdata_i_4_;
 input master_r_rdata_i_5_;
 input master_r_rdata_i_6_;
 input master_r_rdata_i_7_;
 input master_r_rdata_i_8_;
 input master_r_rdata_i_9_;
 input master_r_valid_i;
 output master_req_o;
 output master_wdata_o_0_;
 output master_wdata_o_10_;
 output master_wdata_o_11_;
 output master_wdata_o_12_;
 output master_wdata_o_13_;
 output master_wdata_o_14_;
 output master_wdata_o_15_;
 output master_wdata_o_16_;
 output master_wdata_o_17_;
 output master_wdata_o_18_;
 output master_wdata_o_19_;
 output master_wdata_o_1_;
 output master_wdata_o_20_;
 output master_wdata_o_21_;
 output master_wdata_o_22_;
 output master_wdata_o_23_;
 output master_wdata_o_24_;
 output master_wdata_o_25_;
 output master_wdata_o_26_;
 output master_wdata_o_27_;
 output master_wdata_o_28_;
 output master_wdata_o_29_;
 output master_wdata_o_2_;
 output master_wdata_o_30_;
 output master_wdata_o_31_;
 output master_wdata_o_3_;
 output master_wdata_o_4_;
 output master_wdata_o_5_;
 output master_wdata_o_6_;
 output master_wdata_o_7_;
 output master_wdata_o_8_;
 output master_wdata_o_9_;
 output master_we_o;
 input ndmreset_ack_i;
 output ndmreset_o;
 input next_dm_addr_i_0_;
 input next_dm_addr_i_10_;
 input next_dm_addr_i_11_;
 input next_dm_addr_i_12_;
 input next_dm_addr_i_13_;
 input next_dm_addr_i_14_;
 input next_dm_addr_i_15_;
 input next_dm_addr_i_16_;
 input next_dm_addr_i_17_;
 input next_dm_addr_i_18_;
 input next_dm_addr_i_19_;
 input next_dm_addr_i_1_;
 input next_dm_addr_i_20_;
 input next_dm_addr_i_21_;
 input next_dm_addr_i_22_;
 input next_dm_addr_i_23_;
 input next_dm_addr_i_24_;
 input next_dm_addr_i_25_;
 input next_dm_addr_i_26_;
 input next_dm_addr_i_27_;
 input next_dm_addr_i_28_;
 input next_dm_addr_i_29_;
 input next_dm_addr_i_2_;
 input next_dm_addr_i_30_;
 input next_dm_addr_i_31_;
 input next_dm_addr_i_3_;
 input next_dm_addr_i_4_;
 input next_dm_addr_i_5_;
 input next_dm_addr_i_6_;
 input next_dm_addr_i_7_;
 input next_dm_addr_i_8_;
 input next_dm_addr_i_9_;
 input rst_ni;
 input slave_addr_i_0_;
 input slave_addr_i_10_;
 input slave_addr_i_11_;
 input slave_addr_i_12_;
 input slave_addr_i_13_;
 input slave_addr_i_14_;
 input slave_addr_i_15_;
 input slave_addr_i_16_;
 input slave_addr_i_17_;
 input slave_addr_i_18_;
 input slave_addr_i_19_;
 input slave_addr_i_1_;
 input slave_addr_i_20_;
 input slave_addr_i_21_;
 input slave_addr_i_22_;
 input slave_addr_i_23_;
 input slave_addr_i_24_;
 input slave_addr_i_25_;
 input slave_addr_i_26_;
 input slave_addr_i_27_;
 input slave_addr_i_28_;
 input slave_addr_i_29_;
 input slave_addr_i_2_;
 input slave_addr_i_30_;
 input slave_addr_i_31_;
 input slave_addr_i_3_;
 input slave_addr_i_4_;
 input slave_addr_i_5_;
 input slave_addr_i_6_;
 input slave_addr_i_7_;
 input slave_addr_i_8_;
 input slave_addr_i_9_;
 input slave_be_i_0_;
 input slave_be_i_1_;
 input slave_be_i_2_;
 input slave_be_i_3_;
 output slave_rdata_o_0_;
 output slave_rdata_o_10_;
 output slave_rdata_o_11_;
 output slave_rdata_o_12_;
 output slave_rdata_o_13_;
 output slave_rdata_o_14_;
 output slave_rdata_o_15_;
 output slave_rdata_o_16_;
 output slave_rdata_o_17_;
 output slave_rdata_o_18_;
 output slave_rdata_o_19_;
 output slave_rdata_o_1_;
 output slave_rdata_o_20_;
 output slave_rdata_o_21_;
 output slave_rdata_o_22_;
 output slave_rdata_o_23_;
 output slave_rdata_o_24_;
 output slave_rdata_o_25_;
 output slave_rdata_o_26_;
 output slave_rdata_o_27_;
 output slave_rdata_o_28_;
 output slave_rdata_o_29_;
 output slave_rdata_o_2_;
 output slave_rdata_o_30_;
 output slave_rdata_o_31_;
 output slave_rdata_o_3_;
 output slave_rdata_o_4_;
 output slave_rdata_o_5_;
 output slave_rdata_o_6_;
 output slave_rdata_o_7_;
 output slave_rdata_o_8_;
 output slave_rdata_o_9_;
 input slave_req_i;
 input slave_wdata_i_0_;
 input slave_wdata_i_10_;
 input slave_wdata_i_11_;
 input slave_wdata_i_12_;
 input slave_wdata_i_13_;
 input slave_wdata_i_14_;
 input slave_wdata_i_15_;
 input slave_wdata_i_16_;
 input slave_wdata_i_17_;
 input slave_wdata_i_18_;
 input slave_wdata_i_19_;
 input slave_wdata_i_1_;
 input slave_wdata_i_20_;
 input slave_wdata_i_21_;
 input slave_wdata_i_22_;
 input slave_wdata_i_23_;
 input slave_wdata_i_24_;
 input slave_wdata_i_25_;
 input slave_wdata_i_26_;
 input slave_wdata_i_27_;
 input slave_wdata_i_28_;
 input slave_wdata_i_29_;
 input slave_wdata_i_2_;
 input slave_wdata_i_30_;
 input slave_wdata_i_31_;
 input slave_wdata_i_3_;
 input slave_wdata_i_4_;
 input slave_wdata_i_5_;
 input slave_wdata_i_6_;
 input slave_wdata_i_7_;
 input slave_wdata_i_8_;
 input slave_wdata_i_9_;
 input slave_we_i;
 input testmode_i;
 input unavailable_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire net443;
 wire net442;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire net441;
 wire net440;
 wire _0602_;
 wire _0603_;
 wire net439;
 wire net438;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire net437;
 wire _0611_;
 wire _0612_;
 wire net436;
 wire _0614_;
 wire net435;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire net434;
 wire net433;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire net432;
 wire net431;
 wire _0626_;
 wire net430;
 wire net429;
 wire _0629_;
 wire net428;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire net427;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire net426;
 wire _0643_;
 wire net425;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire net424;
 wire net423;
 wire net422;
 wire _0655_;
 wire net421;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire net420;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire net419;
 wire net418;
 wire _0679_;
 wire net417;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire net416;
 wire _0687_;
 wire _0688_;
 wire net415;
 wire _0690_;
 wire _0691_;
 wire net414;
 wire _0693_;
 wire _0694_;
 wire net413;
 wire _0696_;
 wire _0697_;
 wire net412;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire net411;
 wire _0709_;
 wire _0710_;
 wire net410;
 wire _0712_;
 wire _0713_;
 wire net409;
 wire net408;
 wire net407;
 wire net406;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire net405;
 wire net404;
 wire net403;
 wire net402;
 wire net401;
 wire net400;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire net399;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire net398;
 wire _0741_;
 wire _0742_;
 wire net397;
 wire net396;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire net395;
 wire net394;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire net393;
 wire net392;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire net391;
 wire net390;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire net389;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire net388;
 wire _0802_;
 wire net387;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire net386;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire net385;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire net384;
 wire net383;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire net382;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire net381;
 wire _0860_;
 wire net380;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire net379;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire net378;
 wire net377;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire net376;
 wire net375;
 wire _0893_;
 wire net374;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire net373;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire net372;
 wire _0905_;
 wire _0906_;
 wire net371;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire net370;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire net369;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire net368;
 wire net367;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire net366;
 wire _0966_;
 wire _0967_;
 wire net365;
 wire _0969_;
 wire net364;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire net363;
 wire _0994_;
 wire net362;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire net361;
 wire net360;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire net359;
 wire _1029_;
 wire _1030_;
 wire net358;
 wire _1032_;
 wire net357;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire net356;
 wire net355;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire net354;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire net353;
 wire net352;
 wire net351;
 wire net350;
 wire net349;
 wire net348;
 wire net347;
 wire net346;
 wire net345;
 wire net344;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire net343;
 wire net342;
 wire net341;
 wire net340;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire net339;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire net338;
 wire net337;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire net336;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire net335;
 wire _1172_;
 wire net334;
 wire _1174_;
 wire net333;
 wire net332;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire net331;
 wire net330;
 wire net329;
 wire net328;
 wire _1184_;
 wire net327;
 wire _1186_;
 wire net326;
 wire net325;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire net324;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire net323;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire net322;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire net321;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire net320;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire net319;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire net318;
 wire net317;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire net316;
 wire net315;
 wire _1252_;
 wire net314;
 wire net313;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire net312;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire net311;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire net310;
 wire net309;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire net308;
 wire net307;
 wire net306;
 wire net305;
 wire net304;
 wire net303;
 wire _1299_;
 wire _1300_;
 wire net302;
 wire net301;
 wire _1303_;
 wire _1304_;
 wire net300;
 wire net299;
 wire _1307_;
 wire net298;
 wire net297;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire net296;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire net295;
 wire _1319_;
 wire net294;
 wire net293;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire net292;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire net291;
 wire net290;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire net289;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire net288;
 wire _1377_;
 wire net287;
 wire net286;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire net285;
 wire net284;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire net283;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire net282;
 wire _1396_;
 wire net281;
 wire net280;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire net279;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire net278;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire net277;
 wire net276;
 wire net275;
 wire _1435_;
 wire net274;
 wire net273;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire net272;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire net271;
 wire net270;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire net269;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire net268;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire net267;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire net266;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire net265;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire net264;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire net263;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire net262;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire net261;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire net260;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire net259;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire net258;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire net257;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire net256;
 wire net255;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire net254;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire net253;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire net252;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire net251;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire net250;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire net249;
 wire net248;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire net247;
 wire _1905_;
 wire _1906_;
 wire net246;
 wire net245;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire net244;
 wire net243;
 wire net242;
 wire _1920_;
 wire net241;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire net240;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire net239;
 wire _1936_;
 wire _1937_;
 wire net238;
 wire _1939_;
 wire net237;
 wire _1941_;
 wire net236;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire net235;
 wire net234;
 wire _1949_;
 wire _1950_;
 wire net233;
 wire net232;
 wire _1953_;
 wire _1954_;
 wire net231;
 wire _1956_;
 wire _1957_;
 wire net230;
 wire _1959_;
 wire _1960_;
 wire net229;
 wire _1962_;
 wire _1963_;
 wire net228;
 wire _1965_;
 wire _1966_;
 wire net227;
 wire _1968_;
 wire _1969_;
 wire net226;
 wire _1971_;
 wire _1972_;
 wire net225;
 wire _1974_;
 wire net224;
 wire _1976_;
 wire net223;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire net222;
 wire net221;
 wire _1984_;
 wire _1985_;
 wire net220;
 wire net219;
 wire _1988_;
 wire _1989_;
 wire net218;
 wire _1991_;
 wire _1992_;
 wire net217;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire net216;
 wire _1999_;
 wire _2000_;
 wire net215;
 wire _2002_;
 wire _2003_;
 wire net214;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire net213;
 wire _2012_;
 wire net212;
 wire net211;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire net210;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire net209;
 wire net208;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire net207;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire net206;
 wire net205;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire net204;
 wire net203;
 wire net202;
 wire _2098_;
 wire net201;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire net200;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire net199;
 wire _2122_;
 wire _2123_;
 wire net198;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire net197;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire net196;
 wire _2146_;
 wire net195;
 wire _2148_;
 wire _2149_;
 wire net194;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire net193;
 wire net192;
 wire net191;
 wire _2183_;
 wire net190;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire net189;
 wire net188;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire net187;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire net186;
 wire _2211_;
 wire _2212_;
 wire net185;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire net184;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire net183;
 wire _2236_;
 wire _2237_;
 wire net182;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire net181;
 wire _2266_;
 wire net180;
 wire net179;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire net178;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire net177;
 wire net176;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire net175;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire net174;
 wire net173;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire net172;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire net171;
 wire net170;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire net169;
 wire _2368_;
 wire net168;
 wire net167;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire net166;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire net165;
 wire net164;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire net163;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire net162;
 wire net161;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire net160;
 wire _2451_;
 wire net159;
 wire net158;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire net157;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire net156;
 wire net155;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire net154;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire net153;
 wire net152;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire net151;
 wire _2540_;
 wire _2541_;
 wire net150;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire net149;
 wire net148;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire net147;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire net146;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire net145;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire net144;
 wire _2613_;
 wire _2614_;
 wire net143;
 wire _2616_;
 wire _2617_;
 wire net142;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire net141;
 wire net140;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire net139;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire net138;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire net137;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire net136;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire net135;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire net134;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire net133;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire net132;
 wire net131;
 wire net130;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire net129;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire net128;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire net127;
 wire _2845_;
 wire _2846_;
 wire net126;
 wire _2848_;
 wire net125;
 wire net124;
 wire net123;
 wire _2852_;
 wire _2853_;
 wire net122;
 wire net121;
 wire _2856_;
 wire net120;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire net119;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire net118;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire net117;
 wire net116;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire net115;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire net114;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire net113;
 wire net112;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire net111;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire net110;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire net109;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire net108;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire net107;
 wire net106;
 wire net105;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire net104;
 wire _3034_;
 wire _3035_;
 wire net103;
 wire net102;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire net101;
 wire _3047_;
 wire _3048_;
 wire net100;
 wire net99;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire net98;
 wire _3066_;
 wire net97;
 wire net96;
 wire _3069_;
 wire _3070_;
 wire net95;
 wire _3072_;
 wire net94;
 wire _3074_;
 wire net93;
 wire net92;
 wire _3077_;
 wire _3078_;
 wire net91;
 wire net90;
 wire _3081_;
 wire _3082_;
 wire net89;
 wire net88;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire net87;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire net86;
 wire net85;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire net84;
 wire _3120_;
 wire net83;
 wire _3122_;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire net76;
 wire net75;
 wire net74;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire net73;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire net72;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire net71;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire net70;
 wire net69;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire net68;
 wire net67;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire net66;
 wire net65;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire net64;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire net63;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire net62;
 wire net61;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire net60;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire net59;
 wire net58;
 wire net57;
 wire _3229_;
 wire _3230_;
 wire net56;
 wire _3232_;
 wire net55;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire net54;
 wire net53;
 wire _3240_;
 wire _3241_;
 wire net52;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire net51;
 wire net50;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire net49;
 wire _3366_;
 wire net48;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire net47;
 wire net46;
 wire net45;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire net44;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire net43;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire net42;
 wire net41;
 wire _3707_;
 wire _3708_;
 wire net40;
 wire net39;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire net38;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire net37;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire net36;
 wire net35;
 wire _3770_;
 wire _3771_;
 wire net34;
 wire net33;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire net27;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire net26;
 wire _3792_;
 wire net25;
 wire net24;
 wire net23;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire net22;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire net21;
 wire net20;
 wire net19;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire net18;
 wire net17;
 wire _3815_;
 wire _3816_;
 wire net16;
 wire _3818_;
 wire _3819_;
 wire net15;
 wire _3821_;
 wire net14;
 wire _3823_;
 wire _3824_;
 wire net13;
 wire _3826_;
 wire _3827_;
 wire net12;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire net11;
 wire net10;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire net9;
 wire net8;
 wire net7;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire net6;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire net5;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire net4;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire net3;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire net2;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire net1;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire _4553_;
 wire _4554_;
 wire _4555_;
 wire _4556_;
 wire _4557_;
 wire _4558_;
 wire _4559_;
 wire _4560_;
 wire _4561_;
 wire _4562_;
 wire _4563_;
 wire _4564_;
 wire _4565_;
 wire _4566_;
 wire _4567_;
 wire _4568_;
 wire _4569_;
 wire _4570_;
 wire _4571_;
 wire _4572_;
 wire _4573_;
 wire _4574_;
 wire _4575_;
 wire _4576_;
 wire _4577_;
 wire _4578_;
 wire _4579_;
 wire _4580_;
 wire _4581_;
 wire _4582_;
 wire _4583_;
 wire _4584_;
 wire _4585_;
 wire _4586_;
 wire _4587_;
 wire _4588_;
 wire _4589_;
 wire _4590_;
 wire _4591_;
 wire _4592_;
 wire _4593_;
 wire _4594_;
 wire _4595_;
 wire _4596_;
 wire _4597_;
 wire _4598_;
 wire _4599_;
 wire _4600_;
 wire _4601_;
 wire _4602_;
 wire _4603_;
 wire _4604_;
 wire _4605_;
 wire _4606_;
 wire _4607_;
 wire _4608_;
 wire _4609_;
 wire _4610_;
 wire _4611_;
 wire _4612_;
 wire _4613_;
 wire _4614_;
 wire _4615_;
 wire _4616_;
 wire _4617_;
 wire _4618_;
 wire _4619_;
 wire _4620_;
 wire _4621_;
 wire _4622_;
 wire _4623_;
 wire _4624_;
 wire _4625_;
 wire _4626_;
 wire _4627_;
 wire _4628_;
 wire _4629_;
 wire _4630_;
 wire _4631_;
 wire _4632_;
 wire _4633_;
 wire _4634_;
 wire _4635_;
 wire _4636_;
 wire _4637_;
 wire _4638_;
 wire _4639_;
 wire _4640_;
 wire _4641_;
 wire _4642_;
 wire _4643_;
 wire _4644_;
 wire _4645_;
 wire _4646_;
 wire _4647_;
 wire _4648_;
 wire _4649_;
 wire _4650_;
 wire _4651_;
 wire _4652_;
 wire _4653_;
 wire _4654_;
 wire _4655_;
 wire _4656_;
 wire _4657_;
 wire _4658_;
 wire _4659_;
 wire _4660_;
 wire _4661_;
 wire _4662_;
 wire _4663_;
 wire _4664_;
 wire _4665_;
 wire _4666_;
 wire _4667_;
 wire _4668_;
 wire _4669_;
 wire _4670_;
 wire _4671_;
 wire _4672_;
 wire _4673_;
 wire _4674_;
 wire _4675_;
 wire _4676_;
 wire _4677_;
 wire _4678_;
 wire _4679_;
 wire _4680_;
 wire _4681_;
 wire _4682_;
 wire _4683_;
 wire _4684_;
 wire _4685_;
 wire _4686_;
 wire _4687_;
 wire _4688_;
 wire _4689_;
 wire _4690_;
 wire _4691_;
 wire _4692_;
 wire _4693_;
 wire _4694_;
 wire _4695_;
 wire _4696_;
 wire _4697_;
 wire _4698_;
 wire _4699_;
 wire _4700_;
 wire _4701_;
 wire _4702_;
 wire _4703_;
 wire _4704_;
 wire _4705_;
 wire _4706_;
 wire _4707_;
 wire _4708_;
 wire _4709_;
 wire _4710_;
 wire _4711_;
 wire _4712_;
 wire _4713_;
 wire _4714_;
 wire _4715_;
 wire _4716_;
 wire _4717_;
 wire _4718_;
 wire _4719_;
 wire _4720_;
 wire _4721_;
 wire _4722_;
 wire _4723_;
 wire _4724_;
 wire _4725_;
 wire _4726_;
 wire _4727_;
 wire _4728_;
 wire _4729_;
 wire _4730_;
 wire _4731_;
 wire _4732_;
 wire _4733_;
 wire _4734_;
 wire _4735_;
 wire _4736_;
 wire _4737_;
 wire _4738_;
 wire _4739_;
 wire _4740_;
 wire _4741_;
 wire _4742_;
 wire _4743_;
 wire _4744_;
 wire _4745_;
 wire _4746_;
 wire _4747_;
 wire _4748_;
 wire \clear_resumeack_$_AND__Y_A ;
 wire cmd_0_;
 wire \cmd_0__$_OR__A_B ;
 wire cmd_10_;
 wire cmd_11_;
 wire cmd_12_;
 wire cmd_14_;
 wire cmd_15_;
 wire cmd_16_;
 wire \cmd_16__$_NOT__A_Y ;
 wire cmd_17_;
 wire \cmd_17__$_NOT__A_Y ;
 wire cmd_18_;
 wire cmd_19_;
 wire \cmd_19__$_OR__B_A_$_OR__Y_B_$_AND__Y_A ;
 wire cmd_1_;
 wire cmd_20_;
 wire cmd_21_;
 wire cmd_22_;
 wire cmd_24_;
 wire cmd_25_;
 wire cmd_26_;
 wire cmd_27_;
 wire cmd_28_;
 wire cmd_29_;
 wire cmd_2_;
 wire cmd_30_;
 wire cmd_31_;
 wire cmd_3_;
 wire \cmd_3__$_NOT__A_Y ;
 wire cmd_4_;
 wire cmd_5_;
 wire \cmd_5__$_NOT__A_Y ;
 wire cmd_6_;
 wire cmd_7_;
 wire cmd_8_;
 wire cmd_9_;
 wire cmd_valid;
 wire cmd_valid_reg_D;
 wire data_csrs_mem_0_;
 wire data_csrs_mem_10_;
 wire data_csrs_mem_11_;
 wire data_csrs_mem_12_;
 wire data_csrs_mem_13_;
 wire data_csrs_mem_14_;
 wire data_csrs_mem_15_;
 wire data_csrs_mem_16_;
 wire data_csrs_mem_17_;
 wire data_csrs_mem_18_;
 wire data_csrs_mem_19_;
 wire data_csrs_mem_1_;
 wire data_csrs_mem_20_;
 wire data_csrs_mem_21_;
 wire data_csrs_mem_22_;
 wire data_csrs_mem_23_;
 wire data_csrs_mem_24_;
 wire data_csrs_mem_25_;
 wire data_csrs_mem_26_;
 wire data_csrs_mem_27_;
 wire data_csrs_mem_28_;
 wire data_csrs_mem_29_;
 wire data_csrs_mem_2_;
 wire data_csrs_mem_30_;
 wire data_csrs_mem_31_;
 wire data_csrs_mem_32_;
 wire data_csrs_mem_33_;
 wire data_csrs_mem_34_;
 wire data_csrs_mem_35_;
 wire data_csrs_mem_36_;
 wire data_csrs_mem_37_;
 wire data_csrs_mem_38_;
 wire data_csrs_mem_39_;
 wire data_csrs_mem_3_;
 wire data_csrs_mem_40_;
 wire data_csrs_mem_41_;
 wire data_csrs_mem_42_;
 wire data_csrs_mem_43_;
 wire data_csrs_mem_44_;
 wire data_csrs_mem_45_;
 wire data_csrs_mem_46_;
 wire data_csrs_mem_47_;
 wire data_csrs_mem_48_;
 wire data_csrs_mem_49_;
 wire data_csrs_mem_4_;
 wire data_csrs_mem_50_;
 wire data_csrs_mem_51_;
 wire data_csrs_mem_52_;
 wire data_csrs_mem_53_;
 wire data_csrs_mem_54_;
 wire data_csrs_mem_55_;
 wire data_csrs_mem_56_;
 wire data_csrs_mem_57_;
 wire data_csrs_mem_58_;
 wire data_csrs_mem_59_;
 wire data_csrs_mem_5_;
 wire data_csrs_mem_60_;
 wire data_csrs_mem_61_;
 wire data_csrs_mem_62_;
 wire data_csrs_mem_63_;
 wire data_csrs_mem_6_;
 wire data_csrs_mem_7_;
 wire data_csrs_mem_8_;
 wire data_csrs_mem_9_;
 wire halted;
 wire \i_dm_csrs.abstractauto_q_0_ ;
 wire \i_dm_csrs.abstractauto_q_16_ ;
 wire \i_dm_csrs.abstractauto_q_17_ ;
 wire \i_dm_csrs.abstractauto_q_18_ ;
 wire \i_dm_csrs.abstractauto_q_19_ ;
 wire \i_dm_csrs.abstractauto_q_1_ ;
 wire \i_dm_csrs.abstractauto_q_20_ ;
 wire \i_dm_csrs.abstractauto_q_21_ ;
 wire \i_dm_csrs.abstractauto_q_22_ ;
 wire \i_dm_csrs.abstractauto_q_23_ ;
 wire \i_dm_csrs.cmderr_q_0_ ;
 wire \i_dm_csrs.cmderr_q_0__reg_D ;
 wire \i_dm_csrs.cmderr_q_1_ ;
 wire \i_dm_csrs.cmderr_q_1__reg_D ;
 wire \i_dm_csrs.cmderr_q_2_ ;
 wire \i_dm_csrs.cmderr_q_2__reg_D ;
 wire \i_dm_csrs.dmstatus_11__$_AND__Y_A ;
 wire \i_dm_csrs.dmstatus_16_ ;
 wire \i_dm_csrs.dmstatus_18_ ;
 wire \i_dm_csrs.i_fifo.full_o_$_NOT__Y_A_$_OR__Y_B ;
 wire \i_dm_csrs.i_fifo.mem_q_0_ ;
 wire \i_dm_csrs.i_fifo.mem_q_10_ ;
 wire \i_dm_csrs.i_fifo.mem_q_11_ ;
 wire \i_dm_csrs.i_fifo.mem_q_12_ ;
 wire \i_dm_csrs.i_fifo.mem_q_13_ ;
 wire \i_dm_csrs.i_fifo.mem_q_14_ ;
 wire \i_dm_csrs.i_fifo.mem_q_15_ ;
 wire \i_dm_csrs.i_fifo.mem_q_16_ ;
 wire \i_dm_csrs.i_fifo.mem_q_17_ ;
 wire \i_dm_csrs.i_fifo.mem_q_18_ ;
 wire \i_dm_csrs.i_fifo.mem_q_19_ ;
 wire \i_dm_csrs.i_fifo.mem_q_1_ ;
 wire \i_dm_csrs.i_fifo.mem_q_20_ ;
 wire \i_dm_csrs.i_fifo.mem_q_21_ ;
 wire \i_dm_csrs.i_fifo.mem_q_22_ ;
 wire \i_dm_csrs.i_fifo.mem_q_23_ ;
 wire \i_dm_csrs.i_fifo.mem_q_24_ ;
 wire \i_dm_csrs.i_fifo.mem_q_25_ ;
 wire \i_dm_csrs.i_fifo.mem_q_26_ ;
 wire \i_dm_csrs.i_fifo.mem_q_27_ ;
 wire \i_dm_csrs.i_fifo.mem_q_28_ ;
 wire \i_dm_csrs.i_fifo.mem_q_29_ ;
 wire \i_dm_csrs.i_fifo.mem_q_2_ ;
 wire \i_dm_csrs.i_fifo.mem_q_30_ ;
 wire \i_dm_csrs.i_fifo.mem_q_31_ ;
 wire \i_dm_csrs.i_fifo.mem_q_32_ ;
 wire \i_dm_csrs.i_fifo.mem_q_33_ ;
 wire \i_dm_csrs.i_fifo.mem_q_34_ ;
 wire \i_dm_csrs.i_fifo.mem_q_35_ ;
 wire \i_dm_csrs.i_fifo.mem_q_36_ ;
 wire \i_dm_csrs.i_fifo.mem_q_37_ ;
 wire \i_dm_csrs.i_fifo.mem_q_38_ ;
 wire \i_dm_csrs.i_fifo.mem_q_39_ ;
 wire \i_dm_csrs.i_fifo.mem_q_3_ ;
 wire \i_dm_csrs.i_fifo.mem_q_40_ ;
 wire \i_dm_csrs.i_fifo.mem_q_41_ ;
 wire \i_dm_csrs.i_fifo.mem_q_42_ ;
 wire \i_dm_csrs.i_fifo.mem_q_43_ ;
 wire \i_dm_csrs.i_fifo.mem_q_44_ ;
 wire \i_dm_csrs.i_fifo.mem_q_45_ ;
 wire \i_dm_csrs.i_fifo.mem_q_46_ ;
 wire \i_dm_csrs.i_fifo.mem_q_47_ ;
 wire \i_dm_csrs.i_fifo.mem_q_48_ ;
 wire \i_dm_csrs.i_fifo.mem_q_49_ ;
 wire \i_dm_csrs.i_fifo.mem_q_4_ ;
 wire \i_dm_csrs.i_fifo.mem_q_50_ ;
 wire \i_dm_csrs.i_fifo.mem_q_51_ ;
 wire \i_dm_csrs.i_fifo.mem_q_52_ ;
 wire \i_dm_csrs.i_fifo.mem_q_53_ ;
 wire \i_dm_csrs.i_fifo.mem_q_54_ ;
 wire \i_dm_csrs.i_fifo.mem_q_55_ ;
 wire \i_dm_csrs.i_fifo.mem_q_56_ ;
 wire \i_dm_csrs.i_fifo.mem_q_57_ ;
 wire \i_dm_csrs.i_fifo.mem_q_58_ ;
 wire \i_dm_csrs.i_fifo.mem_q_59_ ;
 wire \i_dm_csrs.i_fifo.mem_q_5_ ;
 wire \i_dm_csrs.i_fifo.mem_q_60_ ;
 wire \i_dm_csrs.i_fifo.mem_q_61_ ;
 wire \i_dm_csrs.i_fifo.mem_q_62_ ;
 wire \i_dm_csrs.i_fifo.mem_q_63_ ;
 wire \i_dm_csrs.i_fifo.mem_q_64_ ;
 wire \i_dm_csrs.i_fifo.mem_q_65_ ;
 wire \i_dm_csrs.i_fifo.mem_q_66_ ;
 wire \i_dm_csrs.i_fifo.mem_q_67_ ;
 wire \i_dm_csrs.i_fifo.mem_q_6_ ;
 wire \i_dm_csrs.i_fifo.mem_q_7_ ;
 wire \i_dm_csrs.i_fifo.mem_q_8_ ;
 wire \i_dm_csrs.i_fifo.mem_q_9_ ;
 wire \i_dm_csrs.i_fifo.read_pointer_n ;
 wire \i_dm_csrs.i_fifo.read_pointer_q ;
 wire \i_dm_csrs.i_fifo.status_cnt_n_0_ ;
 wire \i_dm_csrs.i_fifo.status_cnt_q_0_ ;
 wire \i_dm_csrs.i_fifo.status_cnt_q_1_ ;
 wire \i_dm_csrs.i_fifo.write_pointer_n ;
 wire \i_dm_csrs.i_fifo.write_pointer_q ;
 wire \i_dm_csrs.progbuf_o_0_ ;
 wire \i_dm_csrs.progbuf_o_100_ ;
 wire \i_dm_csrs.progbuf_o_101_ ;
 wire \i_dm_csrs.progbuf_o_102_ ;
 wire \i_dm_csrs.progbuf_o_103_ ;
 wire \i_dm_csrs.progbuf_o_104_ ;
 wire \i_dm_csrs.progbuf_o_105_ ;
 wire \i_dm_csrs.progbuf_o_106_ ;
 wire \i_dm_csrs.progbuf_o_107_ ;
 wire \i_dm_csrs.progbuf_o_108_ ;
 wire \i_dm_csrs.progbuf_o_109_ ;
 wire \i_dm_csrs.progbuf_o_10_ ;
 wire \i_dm_csrs.progbuf_o_110_ ;
 wire \i_dm_csrs.progbuf_o_111_ ;
 wire \i_dm_csrs.progbuf_o_112_ ;
 wire \i_dm_csrs.progbuf_o_113_ ;
 wire \i_dm_csrs.progbuf_o_114_ ;
 wire \i_dm_csrs.progbuf_o_115_ ;
 wire \i_dm_csrs.progbuf_o_116_ ;
 wire \i_dm_csrs.progbuf_o_117_ ;
 wire \i_dm_csrs.progbuf_o_118_ ;
 wire \i_dm_csrs.progbuf_o_119_ ;
 wire \i_dm_csrs.progbuf_o_11_ ;
 wire \i_dm_csrs.progbuf_o_120_ ;
 wire \i_dm_csrs.progbuf_o_121_ ;
 wire \i_dm_csrs.progbuf_o_122_ ;
 wire \i_dm_csrs.progbuf_o_123_ ;
 wire \i_dm_csrs.progbuf_o_124_ ;
 wire \i_dm_csrs.progbuf_o_125_ ;
 wire \i_dm_csrs.progbuf_o_126_ ;
 wire \i_dm_csrs.progbuf_o_127_ ;
 wire \i_dm_csrs.progbuf_o_128_ ;
 wire \i_dm_csrs.progbuf_o_129_ ;
 wire \i_dm_csrs.progbuf_o_12_ ;
 wire \i_dm_csrs.progbuf_o_130_ ;
 wire \i_dm_csrs.progbuf_o_131_ ;
 wire \i_dm_csrs.progbuf_o_132_ ;
 wire \i_dm_csrs.progbuf_o_133_ ;
 wire \i_dm_csrs.progbuf_o_134_ ;
 wire \i_dm_csrs.progbuf_o_135_ ;
 wire \i_dm_csrs.progbuf_o_136_ ;
 wire \i_dm_csrs.progbuf_o_137_ ;
 wire \i_dm_csrs.progbuf_o_138_ ;
 wire \i_dm_csrs.progbuf_o_139_ ;
 wire \i_dm_csrs.progbuf_o_13_ ;
 wire \i_dm_csrs.progbuf_o_140_ ;
 wire \i_dm_csrs.progbuf_o_141_ ;
 wire \i_dm_csrs.progbuf_o_142_ ;
 wire \i_dm_csrs.progbuf_o_143_ ;
 wire \i_dm_csrs.progbuf_o_144_ ;
 wire \i_dm_csrs.progbuf_o_145_ ;
 wire \i_dm_csrs.progbuf_o_146_ ;
 wire \i_dm_csrs.progbuf_o_147_ ;
 wire \i_dm_csrs.progbuf_o_148_ ;
 wire \i_dm_csrs.progbuf_o_149_ ;
 wire \i_dm_csrs.progbuf_o_14_ ;
 wire \i_dm_csrs.progbuf_o_150_ ;
 wire \i_dm_csrs.progbuf_o_151_ ;
 wire \i_dm_csrs.progbuf_o_152_ ;
 wire \i_dm_csrs.progbuf_o_153_ ;
 wire \i_dm_csrs.progbuf_o_154_ ;
 wire \i_dm_csrs.progbuf_o_155_ ;
 wire \i_dm_csrs.progbuf_o_156_ ;
 wire \i_dm_csrs.progbuf_o_157_ ;
 wire \i_dm_csrs.progbuf_o_158_ ;
 wire \i_dm_csrs.progbuf_o_159_ ;
 wire \i_dm_csrs.progbuf_o_15_ ;
 wire \i_dm_csrs.progbuf_o_160_ ;
 wire \i_dm_csrs.progbuf_o_161_ ;
 wire \i_dm_csrs.progbuf_o_162_ ;
 wire \i_dm_csrs.progbuf_o_163_ ;
 wire \i_dm_csrs.progbuf_o_164_ ;
 wire \i_dm_csrs.progbuf_o_165_ ;
 wire \i_dm_csrs.progbuf_o_166_ ;
 wire \i_dm_csrs.progbuf_o_167_ ;
 wire \i_dm_csrs.progbuf_o_168_ ;
 wire \i_dm_csrs.progbuf_o_169_ ;
 wire \i_dm_csrs.progbuf_o_16_ ;
 wire \i_dm_csrs.progbuf_o_170_ ;
 wire \i_dm_csrs.progbuf_o_171_ ;
 wire \i_dm_csrs.progbuf_o_172_ ;
 wire \i_dm_csrs.progbuf_o_173_ ;
 wire \i_dm_csrs.progbuf_o_174_ ;
 wire \i_dm_csrs.progbuf_o_175_ ;
 wire \i_dm_csrs.progbuf_o_176_ ;
 wire \i_dm_csrs.progbuf_o_177_ ;
 wire \i_dm_csrs.progbuf_o_178_ ;
 wire \i_dm_csrs.progbuf_o_179_ ;
 wire \i_dm_csrs.progbuf_o_17_ ;
 wire \i_dm_csrs.progbuf_o_180_ ;
 wire \i_dm_csrs.progbuf_o_181_ ;
 wire \i_dm_csrs.progbuf_o_182_ ;
 wire \i_dm_csrs.progbuf_o_183_ ;
 wire \i_dm_csrs.progbuf_o_184_ ;
 wire \i_dm_csrs.progbuf_o_185_ ;
 wire \i_dm_csrs.progbuf_o_186_ ;
 wire \i_dm_csrs.progbuf_o_187_ ;
 wire \i_dm_csrs.progbuf_o_188_ ;
 wire \i_dm_csrs.progbuf_o_189_ ;
 wire \i_dm_csrs.progbuf_o_18_ ;
 wire \i_dm_csrs.progbuf_o_190_ ;
 wire \i_dm_csrs.progbuf_o_191_ ;
 wire \i_dm_csrs.progbuf_o_192_ ;
 wire \i_dm_csrs.progbuf_o_193_ ;
 wire \i_dm_csrs.progbuf_o_194_ ;
 wire \i_dm_csrs.progbuf_o_195_ ;
 wire \i_dm_csrs.progbuf_o_196_ ;
 wire \i_dm_csrs.progbuf_o_197_ ;
 wire \i_dm_csrs.progbuf_o_198_ ;
 wire \i_dm_csrs.progbuf_o_199_ ;
 wire \i_dm_csrs.progbuf_o_19_ ;
 wire \i_dm_csrs.progbuf_o_1_ ;
 wire \i_dm_csrs.progbuf_o_200_ ;
 wire \i_dm_csrs.progbuf_o_201_ ;
 wire \i_dm_csrs.progbuf_o_202_ ;
 wire \i_dm_csrs.progbuf_o_203_ ;
 wire \i_dm_csrs.progbuf_o_204_ ;
 wire \i_dm_csrs.progbuf_o_205_ ;
 wire \i_dm_csrs.progbuf_o_206_ ;
 wire \i_dm_csrs.progbuf_o_207_ ;
 wire \i_dm_csrs.progbuf_o_208_ ;
 wire \i_dm_csrs.progbuf_o_209_ ;
 wire \i_dm_csrs.progbuf_o_20_ ;
 wire \i_dm_csrs.progbuf_o_210_ ;
 wire \i_dm_csrs.progbuf_o_211_ ;
 wire \i_dm_csrs.progbuf_o_212_ ;
 wire \i_dm_csrs.progbuf_o_213_ ;
 wire \i_dm_csrs.progbuf_o_214_ ;
 wire \i_dm_csrs.progbuf_o_215_ ;
 wire \i_dm_csrs.progbuf_o_216_ ;
 wire \i_dm_csrs.progbuf_o_217_ ;
 wire \i_dm_csrs.progbuf_o_218_ ;
 wire \i_dm_csrs.progbuf_o_219_ ;
 wire \i_dm_csrs.progbuf_o_21_ ;
 wire \i_dm_csrs.progbuf_o_220_ ;
 wire \i_dm_csrs.progbuf_o_221_ ;
 wire \i_dm_csrs.progbuf_o_222_ ;
 wire \i_dm_csrs.progbuf_o_223_ ;
 wire \i_dm_csrs.progbuf_o_224_ ;
 wire \i_dm_csrs.progbuf_o_225_ ;
 wire \i_dm_csrs.progbuf_o_226_ ;
 wire \i_dm_csrs.progbuf_o_227_ ;
 wire \i_dm_csrs.progbuf_o_228_ ;
 wire \i_dm_csrs.progbuf_o_229_ ;
 wire \i_dm_csrs.progbuf_o_22_ ;
 wire \i_dm_csrs.progbuf_o_230_ ;
 wire \i_dm_csrs.progbuf_o_231_ ;
 wire \i_dm_csrs.progbuf_o_232_ ;
 wire \i_dm_csrs.progbuf_o_233_ ;
 wire \i_dm_csrs.progbuf_o_234_ ;
 wire \i_dm_csrs.progbuf_o_235_ ;
 wire \i_dm_csrs.progbuf_o_236_ ;
 wire \i_dm_csrs.progbuf_o_237_ ;
 wire \i_dm_csrs.progbuf_o_238_ ;
 wire \i_dm_csrs.progbuf_o_239_ ;
 wire \i_dm_csrs.progbuf_o_23_ ;
 wire \i_dm_csrs.progbuf_o_240_ ;
 wire \i_dm_csrs.progbuf_o_241_ ;
 wire \i_dm_csrs.progbuf_o_242_ ;
 wire \i_dm_csrs.progbuf_o_243_ ;
 wire \i_dm_csrs.progbuf_o_244_ ;
 wire \i_dm_csrs.progbuf_o_245_ ;
 wire \i_dm_csrs.progbuf_o_246_ ;
 wire \i_dm_csrs.progbuf_o_247_ ;
 wire \i_dm_csrs.progbuf_o_248_ ;
 wire \i_dm_csrs.progbuf_o_249_ ;
 wire \i_dm_csrs.progbuf_o_24_ ;
 wire \i_dm_csrs.progbuf_o_250_ ;
 wire \i_dm_csrs.progbuf_o_251_ ;
 wire \i_dm_csrs.progbuf_o_252_ ;
 wire \i_dm_csrs.progbuf_o_253_ ;
 wire \i_dm_csrs.progbuf_o_254_ ;
 wire \i_dm_csrs.progbuf_o_255_ ;
 wire \i_dm_csrs.progbuf_o_25_ ;
 wire \i_dm_csrs.progbuf_o_26_ ;
 wire \i_dm_csrs.progbuf_o_27_ ;
 wire \i_dm_csrs.progbuf_o_28_ ;
 wire \i_dm_csrs.progbuf_o_29_ ;
 wire \i_dm_csrs.progbuf_o_2_ ;
 wire \i_dm_csrs.progbuf_o_30_ ;
 wire \i_dm_csrs.progbuf_o_31_ ;
 wire \i_dm_csrs.progbuf_o_32_ ;
 wire \i_dm_csrs.progbuf_o_33_ ;
 wire \i_dm_csrs.progbuf_o_34_ ;
 wire \i_dm_csrs.progbuf_o_35_ ;
 wire \i_dm_csrs.progbuf_o_36_ ;
 wire \i_dm_csrs.progbuf_o_37_ ;
 wire \i_dm_csrs.progbuf_o_38_ ;
 wire \i_dm_csrs.progbuf_o_39_ ;
 wire \i_dm_csrs.progbuf_o_3_ ;
 wire \i_dm_csrs.progbuf_o_40_ ;
 wire \i_dm_csrs.progbuf_o_41_ ;
 wire \i_dm_csrs.progbuf_o_42_ ;
 wire \i_dm_csrs.progbuf_o_43_ ;
 wire \i_dm_csrs.progbuf_o_44_ ;
 wire \i_dm_csrs.progbuf_o_45_ ;
 wire \i_dm_csrs.progbuf_o_46_ ;
 wire \i_dm_csrs.progbuf_o_47_ ;
 wire \i_dm_csrs.progbuf_o_48_ ;
 wire \i_dm_csrs.progbuf_o_49_ ;
 wire \i_dm_csrs.progbuf_o_4_ ;
 wire \i_dm_csrs.progbuf_o_50_ ;
 wire \i_dm_csrs.progbuf_o_51_ ;
 wire \i_dm_csrs.progbuf_o_52_ ;
 wire \i_dm_csrs.progbuf_o_53_ ;
 wire \i_dm_csrs.progbuf_o_54_ ;
 wire \i_dm_csrs.progbuf_o_55_ ;
 wire \i_dm_csrs.progbuf_o_56_ ;
 wire \i_dm_csrs.progbuf_o_57_ ;
 wire \i_dm_csrs.progbuf_o_58_ ;
 wire \i_dm_csrs.progbuf_o_59_ ;
 wire \i_dm_csrs.progbuf_o_5_ ;
 wire \i_dm_csrs.progbuf_o_60_ ;
 wire \i_dm_csrs.progbuf_o_61_ ;
 wire \i_dm_csrs.progbuf_o_62_ ;
 wire \i_dm_csrs.progbuf_o_63_ ;
 wire \i_dm_csrs.progbuf_o_64_ ;
 wire \i_dm_csrs.progbuf_o_65_ ;
 wire \i_dm_csrs.progbuf_o_66_ ;
 wire \i_dm_csrs.progbuf_o_67_ ;
 wire \i_dm_csrs.progbuf_o_68_ ;
 wire \i_dm_csrs.progbuf_o_69_ ;
 wire \i_dm_csrs.progbuf_o_6_ ;
 wire \i_dm_csrs.progbuf_o_70_ ;
 wire \i_dm_csrs.progbuf_o_71_ ;
 wire \i_dm_csrs.progbuf_o_72_ ;
 wire \i_dm_csrs.progbuf_o_73_ ;
 wire \i_dm_csrs.progbuf_o_74_ ;
 wire \i_dm_csrs.progbuf_o_75_ ;
 wire \i_dm_csrs.progbuf_o_76_ ;
 wire \i_dm_csrs.progbuf_o_77_ ;
 wire \i_dm_csrs.progbuf_o_78_ ;
 wire \i_dm_csrs.progbuf_o_79_ ;
 wire \i_dm_csrs.progbuf_o_7_ ;
 wire \i_dm_csrs.progbuf_o_80_ ;
 wire \i_dm_csrs.progbuf_o_81_ ;
 wire \i_dm_csrs.progbuf_o_82_ ;
 wire \i_dm_csrs.progbuf_o_83_ ;
 wire \i_dm_csrs.progbuf_o_84_ ;
 wire \i_dm_csrs.progbuf_o_85_ ;
 wire \i_dm_csrs.progbuf_o_86_ ;
 wire \i_dm_csrs.progbuf_o_87_ ;
 wire \i_dm_csrs.progbuf_o_88_ ;
 wire \i_dm_csrs.progbuf_o_89_ ;
 wire \i_dm_csrs.progbuf_o_8_ ;
 wire \i_dm_csrs.progbuf_o_90_ ;
 wire \i_dm_csrs.progbuf_o_91_ ;
 wire \i_dm_csrs.progbuf_o_92_ ;
 wire \i_dm_csrs.progbuf_o_93_ ;
 wire \i_dm_csrs.progbuf_o_94_ ;
 wire \i_dm_csrs.progbuf_o_95_ ;
 wire \i_dm_csrs.progbuf_o_96_ ;
 wire \i_dm_csrs.progbuf_o_97_ ;
 wire \i_dm_csrs.progbuf_o_98_ ;
 wire \i_dm_csrs.progbuf_o_99_ ;
 wire \i_dm_csrs.progbuf_o_9_ ;
 wire \i_dm_csrs.resumereq_o ;
 wire \i_dm_csrs.resumereq_o_reg_D ;
 wire \i_dm_csrs.sbaccess_o_0_ ;
 wire \i_dm_csrs.sbaccess_o_1_ ;
 wire \i_dm_csrs.sbaccess_o_2_ ;
 wire \i_dm_csrs.sbaddr_q_32_ ;
 wire \i_dm_csrs.sbaddr_q_32__reg_D ;
 wire \i_dm_csrs.sbaddr_q_33_ ;
 wire \i_dm_csrs.sbaddr_q_33__reg_D ;
 wire \i_dm_csrs.sbaddr_q_34_ ;
 wire \i_dm_csrs.sbaddr_q_34__reg_D ;
 wire \i_dm_csrs.sbaddr_q_35_ ;
 wire \i_dm_csrs.sbaddr_q_35__reg_D ;
 wire \i_dm_csrs.sbaddr_q_36_ ;
 wire \i_dm_csrs.sbaddr_q_36__reg_D ;
 wire \i_dm_csrs.sbaddr_q_37_ ;
 wire \i_dm_csrs.sbaddr_q_37__reg_D ;
 wire \i_dm_csrs.sbaddr_q_38_ ;
 wire \i_dm_csrs.sbaddr_q_38__reg_D ;
 wire \i_dm_csrs.sbaddr_q_39_ ;
 wire \i_dm_csrs.sbaddr_q_39__reg_D ;
 wire \i_dm_csrs.sbaddr_q_40_ ;
 wire \i_dm_csrs.sbaddr_q_40__reg_D ;
 wire \i_dm_csrs.sbaddr_q_41_ ;
 wire \i_dm_csrs.sbaddr_q_41__reg_D ;
 wire \i_dm_csrs.sbaddr_q_42_ ;
 wire \i_dm_csrs.sbaddr_q_42__reg_D ;
 wire \i_dm_csrs.sbaddr_q_43_ ;
 wire \i_dm_csrs.sbaddr_q_43__reg_D ;
 wire \i_dm_csrs.sbaddr_q_44_ ;
 wire \i_dm_csrs.sbaddr_q_44__reg_D ;
 wire \i_dm_csrs.sbaddr_q_45_ ;
 wire \i_dm_csrs.sbaddr_q_45__reg_D ;
 wire \i_dm_csrs.sbaddr_q_46_ ;
 wire \i_dm_csrs.sbaddr_q_46__reg_D ;
 wire \i_dm_csrs.sbaddr_q_47_ ;
 wire \i_dm_csrs.sbaddr_q_47__reg_D ;
 wire \i_dm_csrs.sbaddr_q_48_ ;
 wire \i_dm_csrs.sbaddr_q_48__reg_D ;
 wire \i_dm_csrs.sbaddr_q_49_ ;
 wire \i_dm_csrs.sbaddr_q_49__reg_D ;
 wire \i_dm_csrs.sbaddr_q_50_ ;
 wire \i_dm_csrs.sbaddr_q_50__reg_D ;
 wire \i_dm_csrs.sbaddr_q_51_ ;
 wire \i_dm_csrs.sbaddr_q_51__reg_D ;
 wire \i_dm_csrs.sbaddr_q_52_ ;
 wire \i_dm_csrs.sbaddr_q_52__reg_D ;
 wire \i_dm_csrs.sbaddr_q_53_ ;
 wire \i_dm_csrs.sbaddr_q_53__reg_D ;
 wire \i_dm_csrs.sbaddr_q_54_ ;
 wire \i_dm_csrs.sbaddr_q_54__reg_D ;
 wire \i_dm_csrs.sbaddr_q_55_ ;
 wire \i_dm_csrs.sbaddr_q_55__reg_D ;
 wire \i_dm_csrs.sbaddr_q_56_ ;
 wire \i_dm_csrs.sbaddr_q_56__reg_D ;
 wire \i_dm_csrs.sbaddr_q_57_ ;
 wire \i_dm_csrs.sbaddr_q_57__reg_D ;
 wire \i_dm_csrs.sbaddr_q_58_ ;
 wire \i_dm_csrs.sbaddr_q_58__reg_D ;
 wire \i_dm_csrs.sbaddr_q_59_ ;
 wire \i_dm_csrs.sbaddr_q_59__reg_D ;
 wire \i_dm_csrs.sbaddr_q_60_ ;
 wire \i_dm_csrs.sbaddr_q_60__reg_D ;
 wire \i_dm_csrs.sbaddr_q_61_ ;
 wire \i_dm_csrs.sbaddr_q_61__reg_D ;
 wire \i_dm_csrs.sbaddr_q_62_ ;
 wire \i_dm_csrs.sbaddr_q_62__reg_D ;
 wire \i_dm_csrs.sbaddr_q_63_ ;
 wire \i_dm_csrs.sbaddr_q_63__reg_D ;
 wire \i_dm_csrs.sbautoincrement_o ;
 wire \i_dm_csrs.sbbusy_i_$_OR__Y_A_$_OR__A_B ;
 wire \i_dm_csrs.sbcs_q_0_ ;
 wire \i_dm_csrs.sbcs_q_12_ ;
 wire \i_dm_csrs.sbcs_q_13_ ;
 wire \i_dm_csrs.sbcs_q_14_ ;
 wire \i_dm_csrs.sbcs_q_15_ ;
 wire \i_dm_csrs.sbcs_q_20_ ;
 wire \i_dm_csrs.sbcs_q_21_ ;
 wire \i_dm_csrs.sbcs_q_21__reg_D ;
 wire \i_dm_csrs.sbcs_q_22_ ;
 wire \i_dm_csrs.sbcs_q_22__reg_D ;
 wire \i_dm_csrs.sbcs_q_23_ ;
 wire \i_dm_csrs.sbcs_q_24_ ;
 wire \i_dm_csrs.sbcs_q_25_ ;
 wire \i_dm_csrs.sbcs_q_26_ ;
 wire \i_dm_csrs.sbcs_q_27_ ;
 wire \i_dm_csrs.sbcs_q_28_ ;
 wire \i_dm_csrs.sbdata_o_0_ ;
 wire \i_dm_csrs.sbdata_o_10_ ;
 wire \i_dm_csrs.sbdata_o_11_ ;
 wire \i_dm_csrs.sbdata_o_12_ ;
 wire \i_dm_csrs.sbdata_o_13_ ;
 wire \i_dm_csrs.sbdata_o_14_ ;
 wire \i_dm_csrs.sbdata_o_15_ ;
 wire \i_dm_csrs.sbdata_o_16_ ;
 wire \i_dm_csrs.sbdata_o_17_ ;
 wire \i_dm_csrs.sbdata_o_18_ ;
 wire \i_dm_csrs.sbdata_o_19_ ;
 wire \i_dm_csrs.sbdata_o_1_ ;
 wire \i_dm_csrs.sbdata_o_20_ ;
 wire \i_dm_csrs.sbdata_o_21_ ;
 wire \i_dm_csrs.sbdata_o_22_ ;
 wire \i_dm_csrs.sbdata_o_23_ ;
 wire \i_dm_csrs.sbdata_o_24_ ;
 wire \i_dm_csrs.sbdata_o_25_ ;
 wire \i_dm_csrs.sbdata_o_26_ ;
 wire \i_dm_csrs.sbdata_o_27_ ;
 wire \i_dm_csrs.sbdata_o_28_ ;
 wire \i_dm_csrs.sbdata_o_29_ ;
 wire \i_dm_csrs.sbdata_o_2_ ;
 wire \i_dm_csrs.sbdata_o_30_ ;
 wire \i_dm_csrs.sbdata_o_31_ ;
 wire \i_dm_csrs.sbdata_o_3_ ;
 wire \i_dm_csrs.sbdata_o_4_ ;
 wire \i_dm_csrs.sbdata_o_5_ ;
 wire \i_dm_csrs.sbdata_o_6_ ;
 wire \i_dm_csrs.sbdata_o_7_ ;
 wire \i_dm_csrs.sbdata_o_8_ ;
 wire \i_dm_csrs.sbdata_o_9_ ;
 wire \i_dm_csrs.sbdata_q_32_ ;
 wire \i_dm_csrs.sbdata_q_33_ ;
 wire \i_dm_csrs.sbdata_q_34_ ;
 wire \i_dm_csrs.sbdata_q_35_ ;
 wire \i_dm_csrs.sbdata_q_36_ ;
 wire \i_dm_csrs.sbdata_q_37_ ;
 wire \i_dm_csrs.sbdata_q_38_ ;
 wire \i_dm_csrs.sbdata_q_39_ ;
 wire \i_dm_csrs.sbdata_q_40_ ;
 wire \i_dm_csrs.sbdata_q_41_ ;
 wire \i_dm_csrs.sbdata_q_42_ ;
 wire \i_dm_csrs.sbdata_q_43_ ;
 wire \i_dm_csrs.sbdata_q_44_ ;
 wire \i_dm_csrs.sbdata_q_45_ ;
 wire \i_dm_csrs.sbdata_q_46_ ;
 wire \i_dm_csrs.sbdata_q_47_ ;
 wire \i_dm_csrs.sbdata_q_48_ ;
 wire \i_dm_csrs.sbdata_q_49_ ;
 wire \i_dm_csrs.sbdata_q_50_ ;
 wire \i_dm_csrs.sbdata_q_51_ ;
 wire \i_dm_csrs.sbdata_q_52_ ;
 wire \i_dm_csrs.sbdata_q_53_ ;
 wire \i_dm_csrs.sbdata_q_54_ ;
 wire \i_dm_csrs.sbdata_q_55_ ;
 wire \i_dm_csrs.sbdata_q_56_ ;
 wire \i_dm_csrs.sbdata_q_57_ ;
 wire \i_dm_csrs.sbdata_q_58_ ;
 wire \i_dm_csrs.sbdata_q_59_ ;
 wire \i_dm_csrs.sbdata_q_60_ ;
 wire \i_dm_csrs.sbdata_q_61_ ;
 wire \i_dm_csrs.sbdata_q_62_ ;
 wire \i_dm_csrs.sbdata_q_63_ ;
 wire \i_dm_mem.abstract_cmd_132__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
 wire \i_dm_mem.fwd_rom_q ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_0_ ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_1_ ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2_ ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3_ ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__$_NOT__A_Y ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_2__$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
 wire \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_42__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
 wire \i_dm_mem.rdata_q_0_ ;
 wire \i_dm_mem.rdata_q_10_ ;
 wire \i_dm_mem.rdata_q_11_ ;
 wire \i_dm_mem.rdata_q_12_ ;
 wire \i_dm_mem.rdata_q_13_ ;
 wire \i_dm_mem.rdata_q_14_ ;
 wire \i_dm_mem.rdata_q_15_ ;
 wire \i_dm_mem.rdata_q_16_ ;
 wire \i_dm_mem.rdata_q_17_ ;
 wire \i_dm_mem.rdata_q_18_ ;
 wire \i_dm_mem.rdata_q_19_ ;
 wire \i_dm_mem.rdata_q_1_ ;
 wire \i_dm_mem.rdata_q_20_ ;
 wire \i_dm_mem.rdata_q_21_ ;
 wire \i_dm_mem.rdata_q_22_ ;
 wire \i_dm_mem.rdata_q_23_ ;
 wire \i_dm_mem.rdata_q_24_ ;
 wire \i_dm_mem.rdata_q_25_ ;
 wire \i_dm_mem.rdata_q_26_ ;
 wire \i_dm_mem.rdata_q_27_ ;
 wire \i_dm_mem.rdata_q_28_ ;
 wire \i_dm_mem.rdata_q_29_ ;
 wire \i_dm_mem.rdata_q_2_ ;
 wire \i_dm_mem.rdata_q_30_ ;
 wire \i_dm_mem.rdata_q_31_ ;
 wire \i_dm_mem.rdata_q_32_ ;
 wire \i_dm_mem.rdata_q_33_ ;
 wire \i_dm_mem.rdata_q_34_ ;
 wire \i_dm_mem.rdata_q_35_ ;
 wire \i_dm_mem.rdata_q_36_ ;
 wire \i_dm_mem.rdata_q_37_ ;
 wire \i_dm_mem.rdata_q_38_ ;
 wire \i_dm_mem.rdata_q_39_ ;
 wire \i_dm_mem.rdata_q_3_ ;
 wire \i_dm_mem.rdata_q_40_ ;
 wire \i_dm_mem.rdata_q_41_ ;
 wire \i_dm_mem.rdata_q_42_ ;
 wire \i_dm_mem.rdata_q_43_ ;
 wire \i_dm_mem.rdata_q_44_ ;
 wire \i_dm_mem.rdata_q_45_ ;
 wire \i_dm_mem.rdata_q_46_ ;
 wire \i_dm_mem.rdata_q_47_ ;
 wire \i_dm_mem.rdata_q_48_ ;
 wire \i_dm_mem.rdata_q_49_ ;
 wire \i_dm_mem.rdata_q_4_ ;
 wire \i_dm_mem.rdata_q_50_ ;
 wire \i_dm_mem.rdata_q_51_ ;
 wire \i_dm_mem.rdata_q_52_ ;
 wire \i_dm_mem.rdata_q_53_ ;
 wire \i_dm_mem.rdata_q_54_ ;
 wire \i_dm_mem.rdata_q_55_ ;
 wire \i_dm_mem.rdata_q_56_ ;
 wire \i_dm_mem.rdata_q_57_ ;
 wire \i_dm_mem.rdata_q_58_ ;
 wire \i_dm_mem.rdata_q_59_ ;
 wire \i_dm_mem.rdata_q_5_ ;
 wire \i_dm_mem.rdata_q_60_ ;
 wire \i_dm_mem.rdata_q_61_ ;
 wire \i_dm_mem.rdata_q_62_ ;
 wire \i_dm_mem.rdata_q_63_ ;
 wire \i_dm_mem.rdata_q_6_ ;
 wire \i_dm_mem.rdata_q_7_ ;
 wire \i_dm_mem.rdata_q_8_ ;
 wire \i_dm_mem.rdata_q_9_ ;
 wire \i_dm_mem.resuming_d ;
 wire \i_dm_mem.state_q_0_ ;
 wire \i_dm_mem.state_q_0__$_NOT__A_Y ;
 wire \i_dm_mem.state_q_1_ ;
 wire \i_dm_mem.state_q_1__$_NOT__A_Y ;
 wire \i_dm_mem.word_enable32_q ;
 wire \i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_A ;
 wire \i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_B ;
 wire \i_dm_sba.sbaccess_mask_3_ ;
 wire \i_dm_sba.sbaccess_mask_3__$_AND__B_A_$_AND__Y_A ;
 wire \i_dm_sba.state_q_0_ ;
 wire \i_dm_sba.state_q_0__$_NOT__A_Y ;
 wire \i_dm_sba.state_q_1_ ;
 wire \i_dm_sba.state_q_1__$_NOT__A_Y ;
 wire \i_dm_sba.state_q_2_ ;
 wire \master_add_o[0]_reg_D ;
 wire \master_add_o[10]_reg_D ;
 wire \master_add_o[11]_reg_D ;
 wire \master_add_o[12]_reg_D ;
 wire \master_add_o[13]_reg_D ;
 wire \master_add_o[14]_reg_D ;
 wire \master_add_o[15]_reg_D ;
 wire \master_add_o[16]_reg_D ;
 wire \master_add_o[17]_reg_D ;
 wire \master_add_o[18]_reg_D ;
 wire \master_add_o[19]_reg_D ;
 wire \master_add_o[1]_reg_D ;
 wire \master_add_o[20]_reg_D ;
 wire \master_add_o[21]_reg_D ;
 wire \master_add_o[22]_reg_D ;
 wire \master_add_o[23]_reg_D ;
 wire \master_add_o[24]_reg_D ;
 wire \master_add_o[25]_reg_D ;
 wire \master_add_o[26]_reg_D ;
 wire \master_add_o[27]_reg_D ;
 wire \master_add_o[28]_reg_D ;
 wire \master_add_o[29]_reg_D ;
 wire \master_add_o[2]_reg_D ;
 wire \master_add_o[30]_reg_D ;
 wire \master_add_o[31]_reg_D ;
 wire \master_add_o[3]_reg_D ;
 wire \master_add_o[4]_reg_D ;
 wire \master_add_o[5]_reg_D ;
 wire \master_add_o[6]_reg_D ;
 wire \master_add_o[7]_reg_D ;
 wire \master_add_o[8]_reg_D ;
 wire \master_add_o[9]_reg_D ;
 wire \ndmreset_o_reg_E_$_AND__Y_B_$_OR__Y_A ;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire clknet_leaf_0_clk_i;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_leaf_35_clk_i;
 wire clknet_leaf_36_clk_i;
 wire clknet_leaf_37_clk_i;
 wire clknet_leaf_39_clk_i;
 wire clknet_leaf_40_clk_i;
 wire clknet_leaf_41_clk_i;
 wire clknet_leaf_42_clk_i;
 wire clknet_leaf_43_clk_i;
 wire clknet_leaf_44_clk_i;
 wire clknet_leaf_45_clk_i;
 wire clknet_leaf_46_clk_i;
 wire clknet_leaf_47_clk_i;
 wire clknet_leaf_48_clk_i;
 wire clknet_leaf_49_clk_i;
 wire clknet_leaf_50_clk_i;
 wire clknet_leaf_51_clk_i;
 wire clknet_leaf_52_clk_i;
 wire clknet_leaf_53_clk_i;
 wire clknet_leaf_54_clk_i;
 wire clknet_leaf_56_clk_i;
 wire clknet_leaf_57_clk_i;
 wire clknet_leaf_58_clk_i;
 wire clknet_leaf_59_clk_i;
 wire clknet_leaf_60_clk_i;
 wire clknet_leaf_61_clk_i;
 wire clknet_leaf_62_clk_i;
 wire clknet_leaf_63_clk_i;
 wire clknet_leaf_64_clk_i;
 wire clknet_leaf_65_clk_i;
 wire clknet_leaf_66_clk_i;
 wire clknet_leaf_67_clk_i;
 wire clknet_leaf_68_clk_i;
 wire clknet_leaf_69_clk_i;
 wire clknet_leaf_70_clk_i;
 wire clknet_leaf_71_clk_i;
 wire clknet_leaf_72_clk_i;
 wire clknet_leaf_73_clk_i;
 wire clknet_leaf_74_clk_i;
 wire clknet_leaf_75_clk_i;
 wire clknet_leaf_76_clk_i;
 wire clknet_leaf_77_clk_i;
 wire clknet_leaf_78_clk_i;
 wire clknet_leaf_79_clk_i;
 wire clknet_leaf_81_clk_i;
 wire clknet_leaf_82_clk_i;
 wire clknet_leaf_83_clk_i;
 wire clknet_leaf_84_clk_i;
 wire clknet_leaf_85_clk_i;
 wire clknet_leaf_86_clk_i;
 wire clknet_leaf_87_clk_i;
 wire clknet_leaf_88_clk_i;
 wire clknet_leaf_89_clk_i;
 wire clknet_leaf_90_clk_i;
 wire clknet_leaf_91_clk_i;
 wire clknet_leaf_92_clk_i;
 wire clknet_leaf_93_clk_i;
 wire clknet_leaf_94_clk_i;
 wire clknet_leaf_95_clk_i;
 wire clknet_leaf_96_clk_i;
 wire clknet_leaf_97_clk_i;
 wire clknet_leaf_98_clk_i;
 wire clknet_leaf_99_clk_i;
 wire clknet_leaf_100_clk_i;
 wire clknet_leaf_101_clk_i;
 wire clknet_leaf_102_clk_i;
 wire clknet_leaf_103_clk_i;
 wire clknet_leaf_104_clk_i;
 wire clknet_0_clk_i;
 wire clknet_4_0_0_clk_i;
 wire clknet_4_1_0_clk_i;
 wire clknet_4_2_0_clk_i;
 wire clknet_4_3_0_clk_i;
 wire clknet_4_4_0_clk_i;
 wire clknet_4_5_0_clk_i;
 wire clknet_4_6_0_clk_i;
 wire clknet_4_7_0_clk_i;
 wire clknet_4_8_0_clk_i;
 wire clknet_4_9_0_clk_i;
 wire clknet_4_10_0_clk_i;
 wire clknet_4_11_0_clk_i;
 wire clknet_4_12_0_clk_i;
 wire clknet_4_13_0_clk_i;
 wire clknet_4_14_0_clk_i;
 wire clknet_4_15_0_clk_i;

 sg13g2_buf_16 fanout443 (.X(net443),
    .A(net450));
 sg13g2_buf_16 fanout442 (.X(net442),
    .A(net443));
 sg13g2_nor2b_1 _4751_ (.A(dmi_req_i_40_),
    .B_N(dmi_req_i_38_),
    .Y(_0594_));
 sg13g2_nand2b_2 _4752_ (.Y(_0595_),
    .B(_0594_),
    .A_N(net130));
 sg13g2_nor3_2 _4753_ (.A(net134),
    .B(net133),
    .C(_0595_),
    .Y(_0596_));
 sg13g2_nand2b_1 _4754_ (.Y(_0597_),
    .B(dmi_req_i_33_),
    .A_N(dmi_req_i_32_));
 sg13g2_or2_2 _4755_ (.X(dmi_req_ready_o),
    .B(\i_dm_csrs.i_fifo.full_o_$_NOT__Y_A_$_OR__Y_B ),
    .A(\i_dm_csrs.i_fifo.status_cnt_q_0_ ));
 sg13g2_nand2_2 _4756_ (.Y(_0598_),
    .A(dmi_req_valid_i),
    .B(dmi_req_ready_o));
 sg13g2_nor2_2 _4757_ (.A(_0597_),
    .B(_0598_),
    .Y(_0599_));
 sg13g2_buf_2 fanout441 (.A(_3116_),
    .X(net441));
 sg13g2_buf_2 fanout440 (.A(_0713_),
    .X(net440));
 sg13g2_nor2_2 _4760_ (.A(net162),
    .B(net155),
    .Y(_0602_));
 sg13g2_nand4_1 _4761_ (.B(_0596_),
    .C(_0599_),
    .A(net210),
    .Y(_0603_),
    .D(_0602_));
 sg13g2_a21oi_1 _4762_ (.A1(\i_dm_csrs.dmstatus_18_ ),
    .A2(_0603_),
    .Y(_0002_),
    .B1(ndmreset_ack_i));
 sg13g2_buf_4 fanout439 (.X(net439),
    .A(_1912_));
 sg13g2_buf_4 fanout438 (.X(net438),
    .A(net439));
 sg13g2_nand2_2 _4765_ (.Y(_0606_),
    .A(net245),
    .B(net84));
 sg13g2_nor2_1 _4766_ (.A(\i_dm_mem.state_q_0_ ),
    .B(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .Y(_0607_));
 sg13g2_a21oi_1 _4767_ (.A1(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .A2(\i_dm_mem.state_q_1_ ),
    .Y(_0608_),
    .B1(\i_dm_mem.state_q_0__$_NOT__A_Y ));
 sg13g2_nor2_2 _4768_ (.A(_0607_),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_buf_4 fanout437 (.X(net437),
    .A(_1912_));
 sg13g2_nor2b_2 _4770_ (.A(dmi_req_i_32_),
    .B_N(dmi_req_i_33_),
    .Y(_0611_));
 sg13g2_and2_2 _4771_ (.A(dmi_req_valid_i),
    .B(dmi_req_ready_o),
    .X(_0612_));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(net437));
 sg13g2_nand2_2 _4773_ (.Y(_0614_),
    .A(_0611_),
    .B(net44));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(net437));
 sg13g2_nor2_1 _4775_ (.A(net133),
    .B(dmi_req_i_40_),
    .Y(_0616_));
 sg13g2_nor2b_1 _4776_ (.A(net131),
    .B_N(dmi_req_i_38_),
    .Y(_0617_));
 sg13g2_nand2_1 _4777_ (.Y(_0618_),
    .A(_0616_),
    .B(_0617_));
 sg13g2_buf_4 fanout434 (.X(net434),
    .A(_2451_));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(net434));
 sg13g2_nand3_1 _4780_ (.B(net145),
    .C(net135),
    .A(net177),
    .Y(_0621_));
 sg13g2_or2_1 _4781_ (.X(_0622_),
    .B(_0621_),
    .A(_0618_));
 sg13g2_nor2_2 _4782_ (.A(_0614_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_buf_4 fanout432 (.X(net432),
    .A(_2451_));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(net432));
 sg13g2_a21oi_2 _4785_ (.B1(net641),
    .Y(_0626_),
    .A2(_0623_),
    .A1(_0609_));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(net432));
 sg13g2_buf_8 fanout429 (.A(_2541_),
    .X(net429));
 sg13g2_nand2_2 _4788_ (.Y(_0629_),
    .A(cmd_0_),
    .B(net417));
 sg13g2_o21ai_1 _4789_ (.B1(_0629_),
    .Y(_0003_),
    .A1(_0606_),
    .A2(net417));
 sg13g2_buf_16 fanout428 (.X(net428),
    .A(net429));
 sg13g2_nand2_1 _4791_ (.Y(_0631_),
    .A(net85),
    .B(net243));
 sg13g2_nand2_1 _4792_ (.Y(_0632_),
    .A(cmd_10_),
    .B(net419));
 sg13g2_o21ai_1 _4793_ (.B1(_0632_),
    .Y(_0004_),
    .A1(net419),
    .A2(_0631_));
 sg13g2_nand2_1 _4794_ (.Y(_0633_),
    .A(net85),
    .B(net241));
 sg13g2_nand2_2 _4795_ (.Y(_0634_),
    .A(cmd_11_),
    .B(net416));
 sg13g2_o21ai_1 _4796_ (.B1(_0634_),
    .Y(_0005_),
    .A1(net416),
    .A2(_0633_));
 sg13g2_nand2_2 _4797_ (.Y(_0635_),
    .A(net85),
    .B(net239));
 sg13g2_buf_2 fanout427 (.A(_2564_),
    .X(net427));
 sg13g2_nand2_2 _4799_ (.Y(_0637_),
    .A(cmd_12_),
    .B(net418));
 sg13g2_o21ai_1 _4800_ (.B1(_0637_),
    .Y(_0006_),
    .A1(net415),
    .A2(_0635_));
 sg13g2_nand2_1 _4801_ (.Y(_0638_),
    .A(net85),
    .B(net237));
 sg13g2_nand2_2 _4802_ (.Y(_0639_),
    .A(cmd_14_),
    .B(net415));
 sg13g2_o21ai_1 _4803_ (.B1(_0639_),
    .Y(_0007_),
    .A1(net415),
    .A2(_0638_));
 sg13g2_nand2_2 _4804_ (.Y(_0640_),
    .A(net85),
    .B(net235));
 sg13g2_nand2_2 _4805_ (.Y(_0641_),
    .A(cmd_15_),
    .B(net416));
 sg13g2_o21ai_1 _4806_ (.B1(_0641_),
    .Y(_0008_),
    .A1(net416),
    .A2(_0640_));
 sg13g2_buf_2 fanout426 (.A(_2944_),
    .X(net426));
 sg13g2_nand2_2 _4808_ (.Y(_0643_),
    .A(net86),
    .B(net233));
 sg13g2_buf_8 fanout425 (.A(_2944_),
    .X(net425));
 sg13g2_nand2_2 _4810_ (.Y(_0645_),
    .A(cmd_16_),
    .B(net415));
 sg13g2_o21ai_1 _4811_ (.B1(_0645_),
    .Y(_0009_),
    .A1(net415),
    .A2(_0643_));
 sg13g2_nand2_2 _4812_ (.Y(_0646_),
    .A(net86),
    .B(net231));
 sg13g2_nand2_2 _4813_ (.Y(_0647_),
    .A(cmd_17_),
    .B(net414));
 sg13g2_o21ai_1 _4814_ (.B1(_0647_),
    .Y(_0010_),
    .A1(net414),
    .A2(_0646_));
 sg13g2_nand2_2 _4815_ (.Y(_0648_),
    .A(net86),
    .B(net229));
 sg13g2_nand2_1 _4816_ (.Y(_0649_),
    .A(cmd_18_),
    .B(net414));
 sg13g2_o21ai_1 _4817_ (.B1(_0649_),
    .Y(_0011_),
    .A1(net414),
    .A2(_0648_));
 sg13g2_nand2_2 _4818_ (.Y(_0650_),
    .A(net86),
    .B(net227));
 sg13g2_nand2_2 _4819_ (.Y(_0651_),
    .A(cmd_19_),
    .B(net414));
 sg13g2_o21ai_1 _4820_ (.B1(_0651_),
    .Y(_0012_),
    .A1(net414),
    .A2(_0650_));
 sg13g2_buf_2 fanout424 (.A(_3451_),
    .X(net424));
 sg13g2_buf_8 fanout423 (.A(_0626_),
    .X(net423));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_nand2_2 _4824_ (.Y(_0655_),
    .A(net88),
    .B(net225));
 sg13g2_buf_16 fanout421 (.X(net421),
    .A(net423));
 sg13g2_nand2_1 _4826_ (.Y(_0657_),
    .A(cmd_1_),
    .B(net418));
 sg13g2_o21ai_1 _4827_ (.B1(_0657_),
    .Y(_0013_),
    .A1(net418),
    .A2(_0655_));
 sg13g2_nand2_2 _4828_ (.Y(_0658_),
    .A(net84),
    .B(net223));
 sg13g2_nand2_1 _4829_ (.Y(_0659_),
    .A(cmd_20_),
    .B(net416));
 sg13g2_o21ai_1 _4830_ (.B1(_0659_),
    .Y(_0014_),
    .A1(net415),
    .A2(_0658_));
 sg13g2_nand2_2 _4831_ (.Y(_0660_),
    .A(net84),
    .B(net221));
 sg13g2_nand2_1 _4832_ (.Y(_0661_),
    .A(cmd_21_),
    .B(net415));
 sg13g2_o21ai_1 _4833_ (.B1(_0661_),
    .Y(_0015_),
    .A1(net415),
    .A2(_0660_));
 sg13g2_nand2_2 _4834_ (.Y(_0662_),
    .A(net84),
    .B(net219));
 sg13g2_nand2_1 _4835_ (.Y(_0663_),
    .A(cmd_22_),
    .B(net420));
 sg13g2_o21ai_1 _4836_ (.B1(_0663_),
    .Y(_0016_),
    .A1(net420),
    .A2(_0662_));
 sg13g2_buf_8 fanout420 (.A(_0626_),
    .X(net420));
 sg13g2_nand2_1 _4838_ (.Y(_0665_),
    .A(net89),
    .B(net217));
 sg13g2_nand2_2 _4839_ (.Y(_0666_),
    .A(cmd_24_),
    .B(net421));
 sg13g2_o21ai_1 _4840_ (.B1(_0666_),
    .Y(_0017_),
    .A1(net421),
    .A2(_0665_));
 sg13g2_nand2_1 _4841_ (.Y(_0667_),
    .A(net89),
    .B(net215));
 sg13g2_nand2_2 _4842_ (.Y(_0668_),
    .A(cmd_25_),
    .B(net421));
 sg13g2_o21ai_1 _4843_ (.B1(_0668_),
    .Y(_0018_),
    .A1(net421),
    .A2(_0667_));
 sg13g2_nand2_1 _4844_ (.Y(_0669_),
    .A(net89),
    .B(net213));
 sg13g2_nand2_2 _4845_ (.Y(_0670_),
    .A(cmd_26_),
    .B(net421));
 sg13g2_o21ai_1 _4846_ (.B1(_0670_),
    .Y(_0019_),
    .A1(net421),
    .A2(_0669_));
 sg13g2_nand2_1 _4847_ (.Y(_0671_),
    .A(net89),
    .B(net211));
 sg13g2_nand2_2 _4848_ (.Y(_0672_),
    .A(cmd_27_),
    .B(net421));
 sg13g2_o21ai_1 _4849_ (.B1(_0672_),
    .Y(_0020_),
    .A1(net421),
    .A2(_0671_));
 sg13g2_nand2_1 _4850_ (.Y(_0673_),
    .A(net88),
    .B(net209));
 sg13g2_nand2_2 _4851_ (.Y(_0674_),
    .A(cmd_28_),
    .B(net423));
 sg13g2_o21ai_1 _4852_ (.B1(_0674_),
    .Y(_0021_),
    .A1(net423),
    .A2(_0673_));
 sg13g2_nand2_1 _4853_ (.Y(_0675_),
    .A(net88),
    .B(net207));
 sg13g2_nand2_1 _4854_ (.Y(_0676_),
    .A(cmd_29_),
    .B(net423));
 sg13g2_o21ai_1 _4855_ (.B1(_0676_),
    .Y(_0022_),
    .A1(net423),
    .A2(_0675_));
 sg13g2_buf_16 fanout419 (.X(net419),
    .A(net420));
 sg13g2_buf_16 fanout418 (.X(net418),
    .A(net419));
 sg13g2_nand2_2 _4858_ (.Y(_0679_),
    .A(net88),
    .B(net205));
 sg13g2_buf_16 fanout417 (.X(net417),
    .A(net418));
 sg13g2_nand2_1 _4860_ (.Y(_0681_),
    .A(cmd_2_),
    .B(net418));
 sg13g2_o21ai_1 _4861_ (.B1(_0681_),
    .Y(_0023_),
    .A1(net417),
    .A2(_0679_));
 sg13g2_nand2_2 _4862_ (.Y(_0682_),
    .A(net203),
    .B(net86));
 sg13g2_nand2_2 _4863_ (.Y(_0683_),
    .A(cmd_30_),
    .B(net422));
 sg13g2_o21ai_1 _4864_ (.B1(_0683_),
    .Y(_0024_),
    .A1(net422),
    .A2(_0682_));
 sg13g2_nand2_2 _4865_ (.Y(_0684_),
    .A(net84),
    .B(net201));
 sg13g2_nand2_2 _4866_ (.Y(_0685_),
    .A(cmd_31_),
    .B(net422));
 sg13g2_o21ai_1 _4867_ (.B1(_0685_),
    .Y(_0025_),
    .A1(net422),
    .A2(_0684_));
 sg13g2_buf_16 fanout416 (.X(net416),
    .A(net420));
 sg13g2_nand2_2 _4869_ (.Y(_0687_),
    .A(net88),
    .B(net128));
 sg13g2_nand2_2 _4870_ (.Y(_0688_),
    .A(cmd_3_),
    .B(net417));
 sg13g2_o21ai_1 _4871_ (.B1(_0688_),
    .Y(_0026_),
    .A1(net417),
    .A2(_0687_));
 sg13g2_buf_16 fanout415 (.X(net415),
    .A(net416));
 sg13g2_nand2_2 _4873_ (.Y(_0690_),
    .A(net88),
    .B(net126));
 sg13g2_nand2_1 _4874_ (.Y(_0691_),
    .A(cmd_4_),
    .B(net418));
 sg13g2_o21ai_1 _4875_ (.B1(_0691_),
    .Y(_0027_),
    .A1(net417),
    .A2(_0690_));
 sg13g2_buf_16 fanout414 (.X(net414),
    .A(net420));
 sg13g2_nand2_2 _4877_ (.Y(_0693_),
    .A(net88),
    .B(net124));
 sg13g2_nand2_2 _4878_ (.Y(_0694_),
    .A(cmd_5_),
    .B(net417));
 sg13g2_o21ai_1 _4879_ (.B1(_0694_),
    .Y(_0028_),
    .A1(net417),
    .A2(_0693_));
 sg13g2_buf_8 fanout413 (.A(_1151_),
    .X(net413));
 sg13g2_nand2_1 _4881_ (.Y(_0696_),
    .A(net86),
    .B(net122));
 sg13g2_nand2_2 _4882_ (.Y(_0697_),
    .A(cmd_6_),
    .B(net416));
 sg13g2_o21ai_1 _4883_ (.B1(_0697_),
    .Y(_0029_),
    .A1(net416),
    .A2(_0696_));
 sg13g2_buf_16 fanout412 (.X(net412),
    .A(net413));
 sg13g2_nand2_1 _4885_ (.Y(_0699_),
    .A(net86),
    .B(net120));
 sg13g2_nand2_2 _4886_ (.Y(_0700_),
    .A(cmd_7_),
    .B(net414));
 sg13g2_o21ai_1 _4887_ (.B1(_0700_),
    .Y(_0030_),
    .A1(net414),
    .A2(_0699_));
 sg13g2_nand2_2 _4888_ (.Y(_0701_),
    .A(net86),
    .B(net118));
 sg13g2_nand2_2 _4889_ (.Y(_0702_),
    .A(cmd_8_),
    .B(net419));
 sg13g2_o21ai_1 _4890_ (.B1(_0702_),
    .Y(_0031_),
    .A1(net419),
    .A2(_0701_));
 sg13g2_nand2_1 _4891_ (.Y(_0703_),
    .A(net85),
    .B(net116));
 sg13g2_nand2_2 _4892_ (.Y(_0704_),
    .A(cmd_9_),
    .B(net419));
 sg13g2_o21ai_1 _4893_ (.B1(_0704_),
    .Y(_0032_),
    .A1(net420),
    .A2(_0703_));
 sg13g2_nand2_1 _4894_ (.Y(_0705_),
    .A(net642),
    .B(slave_we_i));
 sg13g2_nor2_1 _4895_ (.A(slave_addr_i_10_),
    .B(slave_addr_i_11_),
    .Y(_0706_));
 sg13g2_and2_2 _4896_ (.A(slave_addr_i_9_),
    .B(_0706_),
    .X(_0707_));
 sg13g2_buf_16 fanout411 (.X(net411),
    .A(net413));
 sg13g2_nor4_1 _4898_ (.A(net102),
    .B(net654),
    .C(slave_addr_i_5_),
    .D(net644),
    .Y(_0709_));
 sg13g2_and3_1 _4899_ (.X(_0710_),
    .A(slave_addr_i_7_),
    .B(slave_addr_i_8_),
    .C(_0709_));
 sg13g2_buf_8 fanout410 (.A(_1277_),
    .X(net410));
 sg13g2_and2_1 _4901_ (.A(_0707_),
    .B(net555),
    .X(_0712_));
 sg13g2_nor2b_1 _4902_ (.A(_0705_),
    .B_N(net38),
    .Y(_0713_));
 sg13g2_buf_16 fanout409 (.X(net409),
    .A(net410));
 sg13g2_buf_16 fanout408 (.X(net408),
    .A(net409));
 sg13g2_buf_16 fanout407 (.X(net407),
    .A(net408));
 sg13g2_buf_16 fanout406 (.X(net406),
    .A(net409));
 sg13g2_nor2b_1 _4907_ (.A(net178),
    .B_N(net245),
    .Y(_0718_));
 sg13g2_o21ai_1 _4908_ (.B1(net88),
    .Y(_0719_),
    .A1(net26),
    .A2(_0718_));
 sg13g2_nor2b_1 _4909_ (.A(slave_addr_i_2_),
    .B_N(net25),
    .Y(_0720_));
 sg13g2_and2_1 _4910_ (.A(slave_be_i_0_),
    .B(_0720_),
    .X(_0721_));
 sg13g2_buf_16 fanout405 (.X(net405),
    .A(net410));
 sg13g2_buf_8 fanout404 (.A(_2554_),
    .X(net404));
 sg13g2_buf_2 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_1 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_2 fanout401 (.A(net402),
    .X(net401));
 sg13g2_buf_1 fanout400 (.A(net402),
    .X(net400));
 sg13g2_inv_1 _4917_ (.Y(_0728_),
    .A(net134));
 sg13g2_nor2_2 _4918_ (.A(net144),
    .B(net46),
    .Y(_0729_));
 sg13g2_nor3_2 _4919_ (.A(net132),
    .B(dmi_req_i_40_),
    .C(dmi_req_i_38_),
    .Y(_0730_));
 sg13g2_nand3b_1 _4920_ (.B(_0729_),
    .C(_0730_),
    .Y(_0731_),
    .A_N(net130));
 sg13g2_nand2_2 _4921_ (.Y(_0732_),
    .A(_0599_),
    .B(net556));
 sg13g2_nor3_2 _4922_ (.A(net163),
    .B(_0731_),
    .C(_0732_),
    .Y(_0733_));
 sg13g2_nor2_2 _4923_ (.A(net641),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nor2_2 _4924_ (.A(net27),
    .B(_0734_),
    .Y(_0735_));
 sg13g2_buf_2 fanout399 (.A(net400),
    .X(net399));
 sg13g2_a21oi_2 _4926_ (.B1(net384),
    .Y(_0737_),
    .A2(_0721_),
    .A1(slave_wdata_i_0_));
 sg13g2_nor2_1 _4927_ (.A(net641),
    .B(net33),
    .Y(_0738_));
 sg13g2_nand2b_2 _4928_ (.Y(_0739_),
    .B(_0738_),
    .A_N(_0733_));
 sg13g2_buf_8 fanout398 (.A(_2554_),
    .X(net398));
 sg13g2_o21ai_1 _4930_ (.B1(net380),
    .Y(_0741_),
    .A1(_0719_),
    .A2(net387));
 sg13g2_nand2_1 _4931_ (.Y(_0742_),
    .A(data_csrs_mem_0_),
    .B(_0741_));
 sg13g2_o21ai_1 _4932_ (.B1(_0742_),
    .Y(_0033_),
    .A1(_0719_),
    .A2(_0737_));
 sg13g2_buf_1 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_2 fanout396 (.A(net398),
    .X(net396));
 sg13g2_nor2b_1 _4935_ (.A(net179),
    .B_N(net243),
    .Y(_0745_));
 sg13g2_o21ai_1 _4936_ (.B1(net87),
    .Y(_0746_),
    .A1(net26),
    .A2(_0745_));
 sg13g2_and2_1 _4937_ (.A(slave_be_i_1_),
    .B(_0720_),
    .X(_0747_));
 sg13g2_buf_1 fanout395 (.A(_2554_),
    .X(net395));
 sg13g2_buf_2 fanout394 (.A(net395),
    .X(net394));
 sg13g2_a21oi_2 _4940_ (.B1(net385),
    .Y(_0750_),
    .A2(net375),
    .A1(slave_wdata_i_10_));
 sg13g2_o21ai_1 _4941_ (.B1(net380),
    .Y(_0751_),
    .A1(_0746_),
    .A2(_0747_));
 sg13g2_nand2_1 _4942_ (.Y(_0752_),
    .A(data_csrs_mem_10_),
    .B(_0751_));
 sg13g2_o21ai_1 _4943_ (.B1(_0752_),
    .Y(_0034_),
    .A1(_0746_),
    .A2(_0750_));
 sg13g2_buf_8 fanout393 (.A(_2732_),
    .X(net393));
 sg13g2_buf_16 fanout392 (.X(net392),
    .A(net393));
 sg13g2_nor2b_1 _4946_ (.A(net180),
    .B_N(net241),
    .Y(_0755_));
 sg13g2_o21ai_1 _4947_ (.B1(net84),
    .Y(_0756_),
    .A1(net28),
    .A2(_0755_));
 sg13g2_a21oi_2 _4948_ (.B1(net382),
    .Y(_0757_),
    .A2(net375),
    .A1(slave_wdata_i_11_));
 sg13g2_o21ai_1 _4949_ (.B1(net377),
    .Y(_0758_),
    .A1(net375),
    .A2(_0756_));
 sg13g2_nand2_1 _4950_ (.Y(_0759_),
    .A(data_csrs_mem_11_),
    .B(_0758_));
 sg13g2_o21ai_1 _4951_ (.B1(_0759_),
    .Y(_0035_),
    .A1(_0756_),
    .A2(_0757_));
 sg13g2_nor2b_1 _4952_ (.A(net180),
    .B_N(net239),
    .Y(_0760_));
 sg13g2_o21ai_1 _4953_ (.B1(net84),
    .Y(_0761_),
    .A1(net28),
    .A2(_0760_));
 sg13g2_a21oi_2 _4954_ (.B1(net381),
    .Y(_0762_),
    .A2(net375),
    .A1(slave_wdata_i_12_));
 sg13g2_o21ai_1 _4955_ (.B1(net376),
    .Y(_0763_),
    .A1(net375),
    .A2(_0761_));
 sg13g2_nand2_1 _4956_ (.Y(_0764_),
    .A(data_csrs_mem_12_),
    .B(_0763_));
 sg13g2_o21ai_1 _4957_ (.B1(_0764_),
    .Y(_0036_),
    .A1(_0761_),
    .A2(_0762_));
 sg13g2_nor2b_1 _4958_ (.A(net180),
    .B_N(net801),
    .Y(_0765_));
 sg13g2_o21ai_1 _4959_ (.B1(net84),
    .Y(_0766_),
    .A1(net28),
    .A2(_0765_));
 sg13g2_a21oi_2 _4960_ (.B1(net381),
    .Y(_0767_),
    .A2(net375),
    .A1(slave_wdata_i_13_));
 sg13g2_o21ai_1 _4961_ (.B1(net376),
    .Y(_0768_),
    .A1(net375),
    .A2(_0766_));
 sg13g2_nand2_1 _4962_ (.Y(_0769_),
    .A(data_csrs_mem_13_),
    .B(_0768_));
 sg13g2_o21ai_1 _4963_ (.B1(_0769_),
    .Y(_0037_),
    .A1(_0766_),
    .A2(_0767_));
 sg13g2_nor2b_1 _4964_ (.A(net180),
    .B_N(net237),
    .Y(_0770_));
 sg13g2_o21ai_1 _4965_ (.B1(net83),
    .Y(_0771_),
    .A1(net27),
    .A2(_0770_));
 sg13g2_a21oi_2 _4966_ (.B1(net385),
    .Y(_0772_),
    .A2(net374),
    .A1(slave_wdata_i_14_));
 sg13g2_o21ai_1 _4967_ (.B1(net380),
    .Y(_0773_),
    .A1(net374),
    .A2(_0771_));
 sg13g2_nand2_1 _4968_ (.Y(_0774_),
    .A(data_csrs_mem_14_),
    .B(_0773_));
 sg13g2_o21ai_1 _4969_ (.B1(_0774_),
    .Y(_0038_),
    .A1(_0771_),
    .A2(_0772_));
 sg13g2_nor2b_1 _4970_ (.A(net180),
    .B_N(net235),
    .Y(_0775_));
 sg13g2_o21ai_1 _4971_ (.B1(net83),
    .Y(_0776_),
    .A1(net27),
    .A2(_0775_));
 sg13g2_a21oi_2 _4972_ (.B1(net385),
    .Y(_0777_),
    .A2(net374),
    .A1(slave_wdata_i_15_));
 sg13g2_o21ai_1 _4973_ (.B1(net380),
    .Y(_0778_),
    .A1(net374),
    .A2(_0776_));
 sg13g2_nand2_1 _4974_ (.Y(_0779_),
    .A(data_csrs_mem_15_),
    .B(_0778_));
 sg13g2_o21ai_1 _4975_ (.B1(_0779_),
    .Y(_0039_),
    .A1(_0776_),
    .A2(_0777_));
 sg13g2_nor2b_1 _4976_ (.A(net179),
    .B_N(net233),
    .Y(_0780_));
 sg13g2_o21ai_1 _4977_ (.B1(net87),
    .Y(_0781_),
    .A1(net26),
    .A2(_0780_));
 sg13g2_and2_1 _4978_ (.A(slave_be_i_2_),
    .B(_0720_),
    .X(_0782_));
 sg13g2_buf_16 fanout391 (.X(net391),
    .A(net393));
 sg13g2_buf_16 fanout390 (.X(net390),
    .A(net391));
 sg13g2_a21oi_2 _4981_ (.B1(net382),
    .Y(_0785_),
    .A2(net373),
    .A1(slave_wdata_i_16_));
 sg13g2_o21ai_1 _4982_ (.B1(net377),
    .Y(_0786_),
    .A1(_0781_),
    .A2(net373));
 sg13g2_nand2_1 _4983_ (.Y(_0787_),
    .A(data_csrs_mem_16_),
    .B(_0786_));
 sg13g2_o21ai_1 _4984_ (.B1(_0787_),
    .Y(_0040_),
    .A1(_0781_),
    .A2(_0785_));
 sg13g2_nor2b_1 _4985_ (.A(net180),
    .B_N(net231),
    .Y(_0788_));
 sg13g2_buf_16 fanout389 (.X(net389),
    .A(net393));
 sg13g2_o21ai_1 _4987_ (.B1(net90),
    .Y(_0790_),
    .A1(net27),
    .A2(_0788_));
 sg13g2_a21oi_2 _4988_ (.B1(net382),
    .Y(_0791_),
    .A2(net372),
    .A1(slave_wdata_i_17_));
 sg13g2_o21ai_1 _4989_ (.B1(net377),
    .Y(_0792_),
    .A1(net372),
    .A2(_0790_));
 sg13g2_nand2_1 _4990_ (.Y(_0793_),
    .A(data_csrs_mem_17_),
    .B(_0792_));
 sg13g2_o21ai_1 _4991_ (.B1(_0793_),
    .Y(_0041_),
    .A1(_0790_),
    .A2(_0791_));
 sg13g2_nor2b_1 _4992_ (.A(net179),
    .B_N(net229),
    .Y(_0794_));
 sg13g2_o21ai_1 _4993_ (.B1(net90),
    .Y(_0795_),
    .A1(net27),
    .A2(_0794_));
 sg13g2_a21oi_2 _4994_ (.B1(net382),
    .Y(_0796_),
    .A2(net372),
    .A1(slave_wdata_i_18_));
 sg13g2_o21ai_1 _4995_ (.B1(net377),
    .Y(_0797_),
    .A1(net371),
    .A2(_0795_));
 sg13g2_nand2_1 _4996_ (.Y(_0798_),
    .A(data_csrs_mem_18_),
    .B(_0797_));
 sg13g2_o21ai_1 _4997_ (.B1(_0798_),
    .Y(_0042_),
    .A1(_0795_),
    .A2(_0796_));
 sg13g2_nor2b_1 _4998_ (.A(net179),
    .B_N(net227),
    .Y(_0799_));
 sg13g2_o21ai_1 _4999_ (.B1(net90),
    .Y(_0800_),
    .A1(net27),
    .A2(_0799_));
 sg13g2_buf_2 fanout388 (.A(_3097_),
    .X(net388));
 sg13g2_a21oi_2 _5001_ (.B1(net383),
    .Y(_0802_),
    .A2(net372),
    .A1(slave_wdata_i_19_));
 sg13g2_buf_2 fanout387 (.A(_0721_),
    .X(net387));
 sg13g2_o21ai_1 _5003_ (.B1(net378),
    .Y(_0804_),
    .A1(net371),
    .A2(_0800_));
 sg13g2_nand2_1 _5004_ (.Y(_0805_),
    .A(data_csrs_mem_19_),
    .B(_0804_));
 sg13g2_o21ai_1 _5005_ (.B1(_0805_),
    .Y(_0043_),
    .A1(_0800_),
    .A2(_0802_));
 sg13g2_nor2b_1 _5006_ (.A(net179),
    .B_N(net225),
    .Y(_0806_));
 sg13g2_o21ai_1 _5007_ (.B1(net90),
    .Y(_0807_),
    .A1(net27),
    .A2(_0806_));
 sg13g2_a21oi_2 _5008_ (.B1(net384),
    .Y(_0808_),
    .A2(net387),
    .A1(slave_wdata_i_1_));
 sg13g2_o21ai_1 _5009_ (.B1(net379),
    .Y(_0809_),
    .A1(net387),
    .A2(_0807_));
 sg13g2_nand2_1 _5010_ (.Y(_0810_),
    .A(data_csrs_mem_1_),
    .B(_0809_));
 sg13g2_o21ai_1 _5011_ (.B1(_0810_),
    .Y(_0044_),
    .A1(_0807_),
    .A2(_0808_));
 sg13g2_buf_2 fanout386 (.A(net387),
    .X(net386));
 sg13g2_nor2b_1 _5013_ (.A(net181),
    .B_N(net223),
    .Y(_0812_));
 sg13g2_o21ai_1 _5014_ (.B1(net90),
    .Y(_0813_),
    .A1(net27),
    .A2(_0812_));
 sg13g2_a21oi_2 _5015_ (.B1(net382),
    .Y(_0814_),
    .A2(net371),
    .A1(slave_wdata_i_20_));
 sg13g2_o21ai_1 _5016_ (.B1(net377),
    .Y(_0815_),
    .A1(net371),
    .A2(_0813_));
 sg13g2_nand2_1 _5017_ (.Y(_0816_),
    .A(data_csrs_mem_20_),
    .B(_0815_));
 sg13g2_o21ai_1 _5018_ (.B1(_0816_),
    .Y(_0045_),
    .A1(_0813_),
    .A2(_0814_));
 sg13g2_buf_8 fanout385 (.A(_0735_),
    .X(net385));
 sg13g2_nor2b_1 _5020_ (.A(net181),
    .B_N(net221),
    .Y(_0818_));
 sg13g2_o21ai_1 _5021_ (.B1(net90),
    .Y(_0819_),
    .A1(net29),
    .A2(_0818_));
 sg13g2_a21oi_2 _5022_ (.B1(net382),
    .Y(_0820_),
    .A2(net371),
    .A1(slave_wdata_i_21_));
 sg13g2_o21ai_1 _5023_ (.B1(net377),
    .Y(_0821_),
    .A1(net371),
    .A2(_0819_));
 sg13g2_nand2_1 _5024_ (.Y(_0822_),
    .A(data_csrs_mem_21_),
    .B(_0821_));
 sg13g2_o21ai_1 _5025_ (.B1(_0822_),
    .Y(_0046_),
    .A1(_0819_),
    .A2(_0820_));
 sg13g2_nor2b_1 _5026_ (.A(net181),
    .B_N(net219),
    .Y(_0823_));
 sg13g2_o21ai_1 _5027_ (.B1(net89),
    .Y(_0824_),
    .A1(net29),
    .A2(_0823_));
 sg13g2_a21oi_2 _5028_ (.B1(net382),
    .Y(_0825_),
    .A2(net371),
    .A1(slave_wdata_i_22_));
 sg13g2_o21ai_1 _5029_ (.B1(net377),
    .Y(_0826_),
    .A1(net371),
    .A2(_0824_));
 sg13g2_nand2_1 _5030_ (.Y(_0827_),
    .A(data_csrs_mem_22_),
    .B(_0826_));
 sg13g2_o21ai_1 _5031_ (.B1(_0827_),
    .Y(_0047_),
    .A1(_0824_),
    .A2(_0825_));
 sg13g2_nor2b_1 _5032_ (.A(net181),
    .B_N(net798),
    .Y(_0828_));
 sg13g2_o21ai_1 _5033_ (.B1(net89),
    .Y(_0829_),
    .A1(net29),
    .A2(_0828_));
 sg13g2_a21oi_2 _5034_ (.B1(net381),
    .Y(_0830_),
    .A2(net373),
    .A1(slave_wdata_i_23_));
 sg13g2_o21ai_1 _5035_ (.B1(net376),
    .Y(_0831_),
    .A1(net373),
    .A2(_0829_));
 sg13g2_nand2_1 _5036_ (.Y(_0832_),
    .A(data_csrs_mem_23_),
    .B(_0831_));
 sg13g2_o21ai_1 _5037_ (.B1(_0832_),
    .Y(_0048_),
    .A1(_0829_),
    .A2(_0830_));
 sg13g2_nor2b_1 _5038_ (.A(net179),
    .B_N(net217),
    .Y(_0833_));
 sg13g2_o21ai_1 _5039_ (.B1(net87),
    .Y(_0834_),
    .A1(net25),
    .A2(_0833_));
 sg13g2_and2_1 _5040_ (.A(slave_be_i_3_),
    .B(_0720_),
    .X(_0835_));
 sg13g2_buf_16 fanout384 (.X(net384),
    .A(net385));
 sg13g2_buf_8 fanout383 (.A(_0735_),
    .X(net383));
 sg13g2_a21oi_2 _5043_ (.B1(net381),
    .Y(_0838_),
    .A2(net369),
    .A1(slave_wdata_i_24_));
 sg13g2_o21ai_1 _5044_ (.B1(net376),
    .Y(_0839_),
    .A1(_0834_),
    .A2(_0835_));
 sg13g2_nand2_1 _5045_ (.Y(_0840_),
    .A(data_csrs_mem_24_),
    .B(_0839_));
 sg13g2_o21ai_1 _5046_ (.B1(_0840_),
    .Y(_0049_),
    .A1(_0834_),
    .A2(_0838_));
 sg13g2_nor2b_1 _5047_ (.A(net181),
    .B_N(net215),
    .Y(_0841_));
 sg13g2_o21ai_1 _5048_ (.B1(net89),
    .Y(_0842_),
    .A1(net29),
    .A2(_0841_));
 sg13g2_a21oi_2 _5049_ (.B1(net381),
    .Y(_0843_),
    .A2(net370),
    .A1(slave_wdata_i_25_));
 sg13g2_o21ai_1 _5050_ (.B1(net376),
    .Y(_0844_),
    .A1(net370),
    .A2(_0842_));
 sg13g2_nand2_1 _5051_ (.Y(_0845_),
    .A(data_csrs_mem_25_),
    .B(_0844_));
 sg13g2_o21ai_1 _5052_ (.B1(_0845_),
    .Y(_0050_),
    .A1(_0842_),
    .A2(_0843_));
 sg13g2_nor2b_1 _5053_ (.A(net181),
    .B_N(net213),
    .Y(_0846_));
 sg13g2_o21ai_1 _5054_ (.B1(net89),
    .Y(_0847_),
    .A1(net29),
    .A2(_0846_));
 sg13g2_a21oi_2 _5055_ (.B1(net381),
    .Y(_0848_),
    .A2(net369),
    .A1(slave_wdata_i_26_));
 sg13g2_o21ai_1 _5056_ (.B1(net376),
    .Y(_0849_),
    .A1(net369),
    .A2(_0847_));
 sg13g2_nand2_1 _5057_ (.Y(_0850_),
    .A(data_csrs_mem_26_),
    .B(_0849_));
 sg13g2_o21ai_1 _5058_ (.B1(_0850_),
    .Y(_0051_),
    .A1(_0847_),
    .A2(_0848_));
 sg13g2_nor2b_1 _5059_ (.A(net181),
    .B_N(net211),
    .Y(_0851_));
 sg13g2_buf_16 fanout382 (.X(net382),
    .A(net383));
 sg13g2_o21ai_1 _5061_ (.B1(net91),
    .Y(_0853_),
    .A1(net28),
    .A2(_0851_));
 sg13g2_a21oi_2 _5062_ (.B1(net381),
    .Y(_0854_),
    .A2(net370),
    .A1(slave_wdata_i_27_));
 sg13g2_o21ai_1 _5063_ (.B1(net376),
    .Y(_0855_),
    .A1(net370),
    .A2(_0853_));
 sg13g2_nand2_1 _5064_ (.Y(_0856_),
    .A(data_csrs_mem_27_),
    .B(_0855_));
 sg13g2_o21ai_1 _5065_ (.B1(_0856_),
    .Y(_0052_),
    .A1(_0853_),
    .A2(_0854_));
 sg13g2_nor2b_1 _5066_ (.A(net181),
    .B_N(net209),
    .Y(_0857_));
 sg13g2_o21ai_1 _5067_ (.B1(net91),
    .Y(_0858_),
    .A1(net28),
    .A2(_0857_));
 sg13g2_buf_16 fanout381 (.X(net381),
    .A(net383));
 sg13g2_a21oi_2 _5069_ (.B1(net382),
    .Y(_0860_),
    .A2(net370),
    .A1(slave_wdata_i_28_));
 sg13g2_buf_8 fanout380 (.A(_0739_),
    .X(net380));
 sg13g2_o21ai_1 _5071_ (.B1(net377),
    .Y(_0862_),
    .A1(net370),
    .A2(_0858_));
 sg13g2_nand2_1 _5072_ (.Y(_0863_),
    .A(data_csrs_mem_28_),
    .B(_0862_));
 sg13g2_o21ai_1 _5073_ (.B1(_0863_),
    .Y(_0053_),
    .A1(_0858_),
    .A2(_0860_));
 sg13g2_nor2b_1 _5074_ (.A(net180),
    .B_N(net207),
    .Y(_0864_));
 sg13g2_o21ai_1 _5075_ (.B1(net91),
    .Y(_0865_),
    .A1(net28),
    .A2(_0864_));
 sg13g2_a21oi_2 _5076_ (.B1(net381),
    .Y(_0866_),
    .A2(net369),
    .A1(slave_wdata_i_29_));
 sg13g2_o21ai_1 _5077_ (.B1(net376),
    .Y(_0867_),
    .A1(net369),
    .A2(_0865_));
 sg13g2_nand2_1 _5078_ (.Y(_0868_),
    .A(data_csrs_mem_29_),
    .B(_0867_));
 sg13g2_o21ai_1 _5079_ (.B1(_0868_),
    .Y(_0054_),
    .A1(_0865_),
    .A2(_0866_));
 sg13g2_nor2b_1 _5080_ (.A(net180),
    .B_N(net205),
    .Y(_0869_));
 sg13g2_o21ai_1 _5081_ (.B1(net91),
    .Y(_0870_),
    .A1(net28),
    .A2(_0869_));
 sg13g2_a21oi_2 _5082_ (.B1(net384),
    .Y(_0871_),
    .A2(net386),
    .A1(slave_wdata_i_2_));
 sg13g2_o21ai_1 _5083_ (.B1(net379),
    .Y(_0872_),
    .A1(net386),
    .A2(_0870_));
 sg13g2_nand2_1 _5084_ (.Y(_0873_),
    .A(data_csrs_mem_2_),
    .B(_0872_));
 sg13g2_o21ai_1 _5085_ (.B1(_0873_),
    .Y(_0055_),
    .A1(_0870_),
    .A2(_0871_));
 sg13g2_nor2b_1 _5086_ (.A(net178),
    .B_N(net203),
    .Y(_0874_));
 sg13g2_o21ai_1 _5087_ (.B1(net91),
    .Y(_0875_),
    .A1(net28),
    .A2(_0874_));
 sg13g2_a21oi_2 _5088_ (.B1(net383),
    .Y(_0876_),
    .A2(net370),
    .A1(slave_wdata_i_30_));
 sg13g2_o21ai_1 _5089_ (.B1(net378),
    .Y(_0877_),
    .A1(net369),
    .A2(_0875_));
 sg13g2_nand2_1 _5090_ (.Y(_0878_),
    .A(data_csrs_mem_30_),
    .B(_0877_));
 sg13g2_o21ai_1 _5091_ (.B1(_0878_),
    .Y(_0056_),
    .A1(_0875_),
    .A2(_0876_));
 sg13g2_buf_8 fanout379 (.A(_0739_),
    .X(net379));
 sg13g2_nor2b_1 _5093_ (.A(net178),
    .B_N(net201),
    .Y(_0880_));
 sg13g2_o21ai_1 _5094_ (.B1(net91),
    .Y(_0881_),
    .A1(net30),
    .A2(_0880_));
 sg13g2_a21oi_2 _5095_ (.B1(net383),
    .Y(_0882_),
    .A2(net369),
    .A1(slave_wdata_i_31_));
 sg13g2_o21ai_1 _5096_ (.B1(net378),
    .Y(_0883_),
    .A1(net369),
    .A2(_0881_));
 sg13g2_nand2_1 _5097_ (.Y(_0884_),
    .A(data_csrs_mem_31_),
    .B(_0883_));
 sg13g2_o21ai_1 _5098_ (.B1(_0884_),
    .Y(_0057_),
    .A1(_0881_),
    .A2(_0882_));
 sg13g2_buf_8 fanout378 (.A(_0739_),
    .X(net378));
 sg13g2_buf_16 fanout377 (.X(net377),
    .A(net378));
 sg13g2_and2_1 _5101_ (.A(net245),
    .B(net165),
    .X(_0887_));
 sg13g2_o21ai_1 _5102_ (.B1(net87),
    .Y(_0888_),
    .A1(net26),
    .A2(_0887_));
 sg13g2_and2_1 _5103_ (.A(slave_addr_i_2_),
    .B(net33),
    .X(_0889_));
 sg13g2_and2_1 _5104_ (.A(slave_be_i_0_),
    .B(_0889_),
    .X(_0890_));
 sg13g2_buf_16 fanout376 (.X(net376),
    .A(net378));
 sg13g2_buf_2 fanout375 (.A(_0747_),
    .X(net375));
 sg13g2_inv_2 _5107_ (.Y(_0893_),
    .A(net641));
 sg13g2_buf_2 fanout374 (.A(net375),
    .X(net374));
 sg13g2_inv_1 _5109_ (.Y(_0895_),
    .A(net144));
 sg13g2_nand2_2 _5110_ (.Y(_0896_),
    .A(net600),
    .B(net134));
 sg13g2_inv_1 _5111_ (.Y(_0897_),
    .A(_0730_));
 sg13g2_nor3_1 _5112_ (.A(net130),
    .B(_0896_),
    .C(_0897_),
    .Y(_0898_));
 sg13g2_buf_2 fanout373 (.A(_0782_),
    .X(net373));
 sg13g2_or2_2 _5114_ (.X(_0900_),
    .B(_0608_),
    .A(_0607_));
 sg13g2_nor2_2 _5115_ (.A(_0614_),
    .B(_0900_),
    .Y(_0901_));
 sg13g2_nand3_1 _5116_ (.B(net538),
    .C(_0901_),
    .A(net183),
    .Y(_0902_));
 sg13g2_a21oi_2 _5117_ (.B1(net26),
    .Y(_0903_),
    .A2(_0902_),
    .A1(_0893_));
 sg13g2_buf_1 fanout372 (.A(net373),
    .X(net372));
 sg13g2_a21oi_2 _5119_ (.B1(net365),
    .Y(_0905_),
    .A2(net368),
    .A1(slave_wdata_i_0_));
 sg13g2_nand2_1 _5120_ (.Y(_0906_),
    .A(_0738_),
    .B(_0902_));
 sg13g2_buf_2 fanout371 (.A(net373),
    .X(net371));
 sg13g2_o21ai_1 _5122_ (.B1(net360),
    .Y(_0908_),
    .A1(_0888_),
    .A2(net368));
 sg13g2_nand2_1 _5123_ (.Y(_0909_),
    .A(data_csrs_mem_32_),
    .B(_0908_));
 sg13g2_o21ai_1 _5124_ (.B1(_0909_),
    .Y(_0058_),
    .A1(_0888_),
    .A2(_0905_));
 sg13g2_and2_1 _5125_ (.A(net225),
    .B(net164),
    .X(_0910_));
 sg13g2_o21ai_1 _5126_ (.B1(net91),
    .Y(_0911_),
    .A1(net30),
    .A2(_0910_));
 sg13g2_a21oi_2 _5127_ (.B1(net365),
    .Y(_0912_),
    .A2(net368),
    .A1(slave_wdata_i_1_));
 sg13g2_o21ai_1 _5128_ (.B1(net360),
    .Y(_0913_),
    .A1(net368),
    .A2(_0911_));
 sg13g2_nand2_1 _5129_ (.Y(_0914_),
    .A(data_csrs_mem_33_),
    .B(_0913_));
 sg13g2_o21ai_1 _5130_ (.B1(_0914_),
    .Y(_0059_),
    .A1(_0911_),
    .A2(_0912_));
 sg13g2_and2_1 _5131_ (.A(net205),
    .B(net164),
    .X(_0915_));
 sg13g2_o21ai_1 _5132_ (.B1(net91),
    .Y(_0916_),
    .A1(net30),
    .A2(_0915_));
 sg13g2_a21oi_2 _5133_ (.B1(net364),
    .Y(_0917_),
    .A2(net367),
    .A1(slave_wdata_i_2_));
 sg13g2_o21ai_1 _5134_ (.B1(net359),
    .Y(_0918_),
    .A1(net367),
    .A2(_0916_));
 sg13g2_nand2_1 _5135_ (.Y(_0919_),
    .A(data_csrs_mem_34_),
    .B(_0918_));
 sg13g2_o21ai_1 _5136_ (.B1(_0919_),
    .Y(_0060_),
    .A1(_0916_),
    .A2(_0917_));
 sg13g2_buf_2 fanout370 (.A(_0835_),
    .X(net370));
 sg13g2_and2_1 _5138_ (.A(net128),
    .B(net167),
    .X(_0921_));
 sg13g2_o21ai_1 _5139_ (.B1(net90),
    .Y(_0922_),
    .A1(net30),
    .A2(_0921_));
 sg13g2_a21oi_2 _5140_ (.B1(net364),
    .Y(_0923_),
    .A2(net367),
    .A1(slave_wdata_i_3_));
 sg13g2_o21ai_1 _5141_ (.B1(net359),
    .Y(_0924_),
    .A1(net367),
    .A2(_0922_));
 sg13g2_nand2_1 _5142_ (.Y(_0925_),
    .A(data_csrs_mem_35_),
    .B(_0924_));
 sg13g2_o21ai_1 _5143_ (.B1(_0925_),
    .Y(_0061_),
    .A1(_0922_),
    .A2(_0923_));
 sg13g2_and2_1 _5144_ (.A(net126),
    .B(net167),
    .X(_0926_));
 sg13g2_o21ai_1 _5145_ (.B1(net90),
    .Y(_0927_),
    .A1(net30),
    .A2(_0926_));
 sg13g2_a21oi_2 _5146_ (.B1(net364),
    .Y(_0928_),
    .A2(net367),
    .A1(slave_wdata_i_4_));
 sg13g2_o21ai_1 _5147_ (.B1(net359),
    .Y(_0929_),
    .A1(net367),
    .A2(_0927_));
 sg13g2_nand2_1 _5148_ (.Y(_0930_),
    .A(data_csrs_mem_36_),
    .B(_0929_));
 sg13g2_o21ai_1 _5149_ (.B1(_0930_),
    .Y(_0062_),
    .A1(_0927_),
    .A2(_0928_));
 sg13g2_and2_1 _5150_ (.A(net124),
    .B(net167),
    .X(_0931_));
 sg13g2_buf_2 fanout369 (.A(net370),
    .X(net369));
 sg13g2_o21ai_1 _5152_ (.B1(net93),
    .Y(_0933_),
    .A1(net30),
    .A2(_0931_));
 sg13g2_a21oi_2 _5153_ (.B1(net364),
    .Y(_0934_),
    .A2(net368),
    .A1(slave_wdata_i_5_));
 sg13g2_o21ai_1 _5154_ (.B1(net359),
    .Y(_0935_),
    .A1(net368),
    .A2(_0933_));
 sg13g2_nand2_1 _5155_ (.Y(_0936_),
    .A(data_csrs_mem_37_),
    .B(_0935_));
 sg13g2_o21ai_1 _5156_ (.B1(_0936_),
    .Y(_0063_),
    .A1(_0933_),
    .A2(_0934_));
 sg13g2_and2_1 _5157_ (.A(net122),
    .B(net167),
    .X(_0937_));
 sg13g2_o21ai_1 _5158_ (.B1(net93),
    .Y(_0938_),
    .A1(net30),
    .A2(_0937_));
 sg13g2_a21oi_2 _5159_ (.B1(net364),
    .Y(_0939_),
    .A2(net368),
    .A1(slave_wdata_i_6_));
 sg13g2_o21ai_1 _5160_ (.B1(net359),
    .Y(_0940_),
    .A1(net368),
    .A2(_0938_));
 sg13g2_nand2_1 _5161_ (.Y(_0941_),
    .A(data_csrs_mem_38_),
    .B(_0940_));
 sg13g2_o21ai_1 _5162_ (.B1(_0941_),
    .Y(_0064_),
    .A1(_0938_),
    .A2(_0939_));
 sg13g2_and2_1 _5163_ (.A(net120),
    .B(net167),
    .X(_0942_));
 sg13g2_o21ai_1 _5164_ (.B1(net92),
    .Y(_0943_),
    .A1(net29),
    .A2(_0942_));
 sg13g2_a21oi_2 _5165_ (.B1(net364),
    .Y(_0944_),
    .A2(net367),
    .A1(slave_wdata_i_7_));
 sg13g2_o21ai_1 _5166_ (.B1(net359),
    .Y(_0945_),
    .A1(net367),
    .A2(_0943_));
 sg13g2_nand2_1 _5167_ (.Y(_0946_),
    .A(data_csrs_mem_39_),
    .B(_0945_));
 sg13g2_o21ai_1 _5168_ (.B1(_0946_),
    .Y(_0065_),
    .A1(_0943_),
    .A2(_0944_));
 sg13g2_nor2b_1 _5169_ (.A(net178),
    .B_N(net128),
    .Y(_0947_));
 sg13g2_o21ai_1 _5170_ (.B1(net92),
    .Y(_0948_),
    .A1(net29),
    .A2(_0947_));
 sg13g2_a21oi_2 _5171_ (.B1(net385),
    .Y(_0949_),
    .A2(net387),
    .A1(slave_wdata_i_3_));
 sg13g2_o21ai_1 _5172_ (.B1(net379),
    .Y(_0950_),
    .A1(net386),
    .A2(_0948_));
 sg13g2_nand2_1 _5173_ (.Y(_0951_),
    .A(data_csrs_mem_3_),
    .B(_0950_));
 sg13g2_o21ai_1 _5174_ (.B1(_0951_),
    .Y(_0066_),
    .A1(_0948_),
    .A2(_0949_));
 sg13g2_and2_1 _5175_ (.A(net118),
    .B(net165),
    .X(_0952_));
 sg13g2_o21ai_1 _5176_ (.B1(net87),
    .Y(_0953_),
    .A1(net26),
    .A2(_0952_));
 sg13g2_and2_1 _5177_ (.A(slave_be_i_1_),
    .B(_0889_),
    .X(_0954_));
 sg13g2_buf_2 fanout368 (.A(_0890_),
    .X(net368));
 sg13g2_buf_2 fanout367 (.A(_0890_),
    .X(net367));
 sg13g2_a21oi_2 _5180_ (.B1(net364),
    .Y(_0957_),
    .A2(net355),
    .A1(slave_wdata_i_8_));
 sg13g2_o21ai_1 _5181_ (.B1(net359),
    .Y(_0958_),
    .A1(_0953_),
    .A2(net355));
 sg13g2_nand2_1 _5182_ (.Y(_0959_),
    .A(data_csrs_mem_40_),
    .B(_0958_));
 sg13g2_o21ai_1 _5183_ (.B1(_0959_),
    .Y(_0067_),
    .A1(_0953_),
    .A2(_0957_));
 sg13g2_and2_1 _5184_ (.A(net116),
    .B(net167),
    .X(_0960_));
 sg13g2_o21ai_1 _5185_ (.B1(net92),
    .Y(_0961_),
    .A1(net29),
    .A2(_0960_));
 sg13g2_a21oi_2 _5186_ (.B1(net364),
    .Y(_0962_),
    .A2(net355),
    .A1(slave_wdata_i_9_));
 sg13g2_o21ai_1 _5187_ (.B1(net360),
    .Y(_0963_),
    .A1(net356),
    .A2(_0961_));
 sg13g2_nand2_1 _5188_ (.Y(_0964_),
    .A(data_csrs_mem_41_),
    .B(_0963_));
 sg13g2_o21ai_1 _5189_ (.B1(_0964_),
    .Y(_0068_),
    .A1(_0961_),
    .A2(_0962_));
 sg13g2_buf_8 fanout366 (.A(_0903_),
    .X(net366));
 sg13g2_and2_1 _5191_ (.A(net243),
    .B(net167),
    .X(_0966_));
 sg13g2_o21ai_1 _5192_ (.B1(net92),
    .Y(_0967_),
    .A1(net32),
    .A2(_0966_));
 sg13g2_buf_16 fanout365 (.X(net365),
    .A(net366));
 sg13g2_a21oi_2 _5194_ (.B1(net365),
    .Y(_0969_),
    .A2(net356),
    .A1(slave_wdata_i_10_));
 sg13g2_buf_16 fanout364 (.X(net364),
    .A(net365));
 sg13g2_o21ai_1 _5196_ (.B1(net360),
    .Y(_0971_),
    .A1(net355),
    .A2(_0967_));
 sg13g2_nand2_1 _5197_ (.Y(_0972_),
    .A(data_csrs_mem_42_),
    .B(_0971_));
 sg13g2_o21ai_1 _5198_ (.B1(_0972_),
    .Y(_0069_),
    .A1(_0967_),
    .A2(_0969_));
 sg13g2_and2_1 _5199_ (.A(net241),
    .B(net166),
    .X(_0973_));
 sg13g2_o21ai_1 _5200_ (.B1(net92),
    .Y(_0974_),
    .A1(net31),
    .A2(_0973_));
 sg13g2_a21oi_2 _5201_ (.B1(net365),
    .Y(_0975_),
    .A2(net356),
    .A1(slave_wdata_i_11_));
 sg13g2_o21ai_1 _5202_ (.B1(net360),
    .Y(_0976_),
    .A1(net355),
    .A2(_0974_));
 sg13g2_nand2_1 _5203_ (.Y(_0977_),
    .A(data_csrs_mem_43_),
    .B(_0976_));
 sg13g2_o21ai_1 _5204_ (.B1(_0977_),
    .Y(_0070_),
    .A1(_0974_),
    .A2(_0975_));
 sg13g2_and2_1 _5205_ (.A(net239),
    .B(net166),
    .X(_0978_));
 sg13g2_o21ai_1 _5206_ (.B1(net92),
    .Y(_0979_),
    .A1(net31),
    .A2(_0978_));
 sg13g2_a21oi_2 _5207_ (.B1(net362),
    .Y(_0980_),
    .A2(net356),
    .A1(slave_wdata_i_12_));
 sg13g2_o21ai_1 _5208_ (.B1(net357),
    .Y(_0981_),
    .A1(net356),
    .A2(_0979_));
 sg13g2_nand2_1 _5209_ (.Y(_0982_),
    .A(data_csrs_mem_44_),
    .B(_0981_));
 sg13g2_o21ai_1 _5210_ (.B1(_0982_),
    .Y(_0071_),
    .A1(_0979_),
    .A2(_0980_));
 sg13g2_and2_1 _5211_ (.A(net161),
    .B(net801),
    .X(_0983_));
 sg13g2_o21ai_1 _5212_ (.B1(net92),
    .Y(_0984_),
    .A1(net31),
    .A2(_0983_));
 sg13g2_a21oi_2 _5213_ (.B1(net362),
    .Y(_0985_),
    .A2(net356),
    .A1(slave_wdata_i_13_));
 sg13g2_o21ai_1 _5214_ (.B1(net359),
    .Y(_0986_),
    .A1(net356),
    .A2(_0984_));
 sg13g2_nand2_1 _5215_ (.Y(_0987_),
    .A(data_csrs_mem_45_),
    .B(_0986_));
 sg13g2_o21ai_1 _5216_ (.B1(_0987_),
    .Y(_0072_),
    .A1(_0984_),
    .A2(_0985_));
 sg13g2_and2_1 _5217_ (.A(net237),
    .B(net166),
    .X(_0988_));
 sg13g2_o21ai_1 _5218_ (.B1(net92),
    .Y(_0989_),
    .A1(net31),
    .A2(_0988_));
 sg13g2_a21oi_2 _5219_ (.B1(net365),
    .Y(_0990_),
    .A2(_0954_),
    .A1(slave_wdata_i_14_));
 sg13g2_o21ai_1 _5220_ (.B1(net360),
    .Y(_0991_),
    .A1(net355),
    .A2(_0989_));
 sg13g2_nand2_1 _5221_ (.Y(_0992_),
    .A(data_csrs_mem_46_),
    .B(_0991_));
 sg13g2_o21ai_1 _5222_ (.B1(_0992_),
    .Y(_0073_),
    .A1(_0989_),
    .A2(_0990_));
 sg13g2_buf_16 fanout363 (.X(net363),
    .A(net366));
 sg13g2_and2_1 _5224_ (.A(net235),
    .B(net169),
    .X(_0994_));
 sg13g2_buf_16 fanout362 (.X(net362),
    .A(net363));
 sg13g2_o21ai_1 _5226_ (.B1(net94),
    .Y(_0996_),
    .A1(net31),
    .A2(_0994_));
 sg13g2_a21oi_2 _5227_ (.B1(net365),
    .Y(_0997_),
    .A2(net355),
    .A1(slave_wdata_i_15_));
 sg13g2_o21ai_1 _5228_ (.B1(net360),
    .Y(_0998_),
    .A1(net355),
    .A2(_0996_));
 sg13g2_nand2_1 _5229_ (.Y(_0999_),
    .A(data_csrs_mem_47_),
    .B(_0998_));
 sg13g2_o21ai_1 _5230_ (.B1(_0999_),
    .Y(_0074_),
    .A1(_0996_),
    .A2(_0997_));
 sg13g2_and2_1 _5231_ (.A(net233),
    .B(net165),
    .X(_1000_));
 sg13g2_o21ai_1 _5232_ (.B1(net87),
    .Y(_1001_),
    .A1(net26),
    .A2(_1000_));
 sg13g2_and2_1 _5233_ (.A(slave_be_i_2_),
    .B(_0889_),
    .X(_1002_));
 sg13g2_buf_8 fanout361 (.A(_0906_),
    .X(net361));
 sg13g2_buf_16 fanout360 (.X(net360),
    .A(net361));
 sg13g2_a21oi_2 _5236_ (.B1(net363),
    .Y(_1005_),
    .A2(net354),
    .A1(slave_wdata_i_16_));
 sg13g2_o21ai_1 _5237_ (.B1(net358),
    .Y(_1006_),
    .A1(_1001_),
    .A2(net354));
 sg13g2_nand2_1 _5238_ (.Y(_1007_),
    .A(data_csrs_mem_48_),
    .B(_1006_));
 sg13g2_o21ai_1 _5239_ (.B1(_1007_),
    .Y(_0075_),
    .A1(_1001_),
    .A2(_1005_));
 sg13g2_and2_1 _5240_ (.A(net231),
    .B(net168),
    .X(_1008_));
 sg13g2_o21ai_1 _5241_ (.B1(net94),
    .Y(_1009_),
    .A1(net31),
    .A2(_1008_));
 sg13g2_a21oi_2 _5242_ (.B1(net363),
    .Y(_1010_),
    .A2(net353),
    .A1(slave_wdata_i_17_));
 sg13g2_o21ai_1 _5243_ (.B1(net358),
    .Y(_1011_),
    .A1(net353),
    .A2(_1009_));
 sg13g2_nand2_1 _5244_ (.Y(_1012_),
    .A(data_csrs_mem_49_),
    .B(_1011_));
 sg13g2_o21ai_1 _5245_ (.B1(_1012_),
    .Y(_0076_),
    .A1(_1009_),
    .A2(_1010_));
 sg13g2_nor2b_1 _5246_ (.A(net177),
    .B_N(net126),
    .Y(_1013_));
 sg13g2_o21ai_1 _5247_ (.B1(net94),
    .Y(_1014_),
    .A1(net31),
    .A2(_1013_));
 sg13g2_a21oi_1 _5248_ (.A1(slave_wdata_i_4_),
    .A2(net387),
    .Y(_1015_),
    .B1(net385));
 sg13g2_o21ai_1 _5249_ (.B1(net379),
    .Y(_1016_),
    .A1(net386),
    .A2(_1014_));
 sg13g2_nand2_1 _5250_ (.Y(_1017_),
    .A(data_csrs_mem_4_),
    .B(_1016_));
 sg13g2_o21ai_1 _5251_ (.B1(_1017_),
    .Y(_0077_),
    .A1(_1014_),
    .A2(_1015_));
 sg13g2_and2_1 _5252_ (.A(net229),
    .B(net168),
    .X(_1018_));
 sg13g2_o21ai_1 _5253_ (.B1(net94),
    .Y(_1019_),
    .A1(net31),
    .A2(_1018_));
 sg13g2_a21oi_2 _5254_ (.B1(net363),
    .Y(_1020_),
    .A2(net353),
    .A1(slave_wdata_i_18_));
 sg13g2_o21ai_1 _5255_ (.B1(net358),
    .Y(_1021_),
    .A1(net352),
    .A2(_1019_));
 sg13g2_nand2_1 _5256_ (.Y(_1022_),
    .A(data_csrs_mem_50_),
    .B(_1021_));
 sg13g2_o21ai_1 _5257_ (.B1(_1022_),
    .Y(_0078_),
    .A1(_1019_),
    .A2(_1020_));
 sg13g2_and2_1 _5258_ (.A(net227),
    .B(net168),
    .X(_1023_));
 sg13g2_o21ai_1 _5259_ (.B1(net93),
    .Y(_1024_),
    .A1(net30),
    .A2(_1023_));
 sg13g2_a21oi_2 _5260_ (.B1(net363),
    .Y(_1025_),
    .A2(net353),
    .A1(slave_wdata_i_19_));
 sg13g2_o21ai_1 _5261_ (.B1(net358),
    .Y(_1026_),
    .A1(net352),
    .A2(_1024_));
 sg13g2_nand2_1 _5262_ (.Y(_1027_),
    .A(data_csrs_mem_51_),
    .B(_1026_));
 sg13g2_o21ai_1 _5263_ (.B1(_1027_),
    .Y(_0079_),
    .A1(_1024_),
    .A2(_1025_));
 sg13g2_buf_16 fanout359 (.X(net359),
    .A(net360));
 sg13g2_and2_1 _5265_ (.A(net223),
    .B(net168),
    .X(_1029_));
 sg13g2_o21ai_1 _5266_ (.B1(net93),
    .Y(_1030_),
    .A1(net33),
    .A2(_1029_));
 sg13g2_buf_16 fanout358 (.X(net358),
    .A(net361));
 sg13g2_a21oi_2 _5268_ (.B1(net366),
    .Y(_1032_),
    .A2(net352),
    .A1(slave_wdata_i_20_));
 sg13g2_buf_16 fanout357 (.X(net357),
    .A(net358));
 sg13g2_o21ai_1 _5270_ (.B1(net361),
    .Y(_1034_),
    .A1(net352),
    .A2(_1030_));
 sg13g2_nand2_1 _5271_ (.Y(_1035_),
    .A(data_csrs_mem_52_),
    .B(_1034_));
 sg13g2_o21ai_1 _5272_ (.B1(_1035_),
    .Y(_0080_),
    .A1(_1030_),
    .A2(_1032_));
 sg13g2_and2_1 _5273_ (.A(net221),
    .B(net168),
    .X(_1036_));
 sg13g2_o21ai_1 _5274_ (.B1(net93),
    .Y(_1037_),
    .A1(net33),
    .A2(_1036_));
 sg13g2_a21oi_2 _5275_ (.B1(net366),
    .Y(_1038_),
    .A2(net352),
    .A1(slave_wdata_i_21_));
 sg13g2_o21ai_1 _5276_ (.B1(net361),
    .Y(_1039_),
    .A1(net352),
    .A2(_1037_));
 sg13g2_nand2_1 _5277_ (.Y(_1040_),
    .A(data_csrs_mem_53_),
    .B(_1039_));
 sg13g2_o21ai_1 _5278_ (.B1(_1040_),
    .Y(_0081_),
    .A1(_1037_),
    .A2(_1038_));
 sg13g2_and2_1 _5279_ (.A(net219),
    .B(net168),
    .X(_1041_));
 sg13g2_o21ai_1 _5280_ (.B1(net93),
    .Y(_1042_),
    .A1(net33),
    .A2(_1041_));
 sg13g2_a21oi_1 _5281_ (.A1(slave_wdata_i_22_),
    .A2(net352),
    .Y(_1043_),
    .B1(net366));
 sg13g2_o21ai_1 _5282_ (.B1(net358),
    .Y(_1044_),
    .A1(net352),
    .A2(_1042_));
 sg13g2_nand2_1 _5283_ (.Y(_1045_),
    .A(data_csrs_mem_54_),
    .B(_1044_));
 sg13g2_o21ai_1 _5284_ (.B1(_1045_),
    .Y(_0082_),
    .A1(_1042_),
    .A2(_1043_));
 sg13g2_and2_1 _5285_ (.A(net161),
    .B(net798),
    .X(_1046_));
 sg13g2_o21ai_1 _5286_ (.B1(net93),
    .Y(_1047_),
    .A1(net32),
    .A2(_1046_));
 sg13g2_a21oi_2 _5287_ (.B1(net363),
    .Y(_1048_),
    .A2(net354),
    .A1(slave_wdata_i_23_));
 sg13g2_o21ai_1 _5288_ (.B1(net358),
    .Y(_1049_),
    .A1(net354),
    .A2(_1047_));
 sg13g2_nand2_1 _5289_ (.Y(_1050_),
    .A(data_csrs_mem_55_),
    .B(_1049_));
 sg13g2_o21ai_1 _5290_ (.B1(_1050_),
    .Y(_0083_),
    .A1(_1047_),
    .A2(_1048_));
 sg13g2_and2_1 _5291_ (.A(net217),
    .B(net165),
    .X(_1051_));
 sg13g2_o21ai_1 _5292_ (.B1(net87),
    .Y(_1052_),
    .A1(net26),
    .A2(_1051_));
 sg13g2_and2_1 _5293_ (.A(slave_be_i_3_),
    .B(_0889_),
    .X(_1053_));
 sg13g2_buf_2 fanout356 (.A(_0954_),
    .X(net356));
 sg13g2_buf_2 fanout355 (.A(net356),
    .X(net355));
 sg13g2_a21oi_2 _5296_ (.B1(net362),
    .Y(_1056_),
    .A2(net350),
    .A1(slave_wdata_i_24_));
 sg13g2_o21ai_1 _5297_ (.B1(net357),
    .Y(_1057_),
    .A1(_1052_),
    .A2(_1053_));
 sg13g2_nand2_1 _5298_ (.Y(_1058_),
    .A(data_csrs_mem_56_),
    .B(_1057_));
 sg13g2_o21ai_1 _5299_ (.B1(_1058_),
    .Y(_0084_),
    .A1(_1052_),
    .A2(_1056_));
 sg13g2_and2_1 _5300_ (.A(net215),
    .B(net168),
    .X(_1059_));
 sg13g2_o21ai_1 _5301_ (.B1(net93),
    .Y(_1060_),
    .A1(net32),
    .A2(_1059_));
 sg13g2_a21oi_2 _5302_ (.B1(net362),
    .Y(_1061_),
    .A2(net351),
    .A1(slave_wdata_i_25_));
 sg13g2_o21ai_1 _5303_ (.B1(net357),
    .Y(_1062_),
    .A1(net351),
    .A2(_1060_));
 sg13g2_nand2_1 _5304_ (.Y(_1063_),
    .A(data_csrs_mem_57_),
    .B(_1062_));
 sg13g2_o21ai_1 _5305_ (.B1(_1063_),
    .Y(_0085_),
    .A1(_1060_),
    .A2(_1061_));
 sg13g2_and2_1 _5306_ (.A(net213),
    .B(net168),
    .X(_1064_));
 sg13g2_buf_2 fanout354 (.A(_1002_),
    .X(net354));
 sg13g2_o21ai_1 _5308_ (.B1(net95),
    .Y(_1066_),
    .A1(net32),
    .A2(_1064_));
 sg13g2_a21oi_2 _5309_ (.B1(net362),
    .Y(_1067_),
    .A2(net350),
    .A1(slave_wdata_i_26_));
 sg13g2_o21ai_1 _5310_ (.B1(net357),
    .Y(_1068_),
    .A1(net350),
    .A2(_1066_));
 sg13g2_nand2_1 _5311_ (.Y(_1069_),
    .A(data_csrs_mem_58_),
    .B(_1068_));
 sg13g2_o21ai_1 _5312_ (.B1(_1069_),
    .Y(_0086_),
    .A1(_1066_),
    .A2(_1067_));
 sg13g2_and2_1 _5313_ (.A(net211),
    .B(net167),
    .X(_1070_));
 sg13g2_o21ai_1 _5314_ (.B1(net95),
    .Y(_1071_),
    .A1(net32),
    .A2(_1070_));
 sg13g2_a21oi_2 _5315_ (.B1(net363),
    .Y(_1072_),
    .A2(net351),
    .A1(slave_wdata_i_27_));
 sg13g2_o21ai_1 _5316_ (.B1(net357),
    .Y(_1073_),
    .A1(net351),
    .A2(_1071_));
 sg13g2_nand2_1 _5317_ (.Y(_1074_),
    .A(data_csrs_mem_59_),
    .B(_1073_));
 sg13g2_o21ai_1 _5318_ (.B1(_1074_),
    .Y(_0087_),
    .A1(_1071_),
    .A2(_1072_));
 sg13g2_nor2b_1 _5319_ (.A(net177),
    .B_N(net124),
    .Y(_1075_));
 sg13g2_o21ai_1 _5320_ (.B1(net95),
    .Y(_1076_),
    .A1(net32),
    .A2(_1075_));
 sg13g2_a21oi_2 _5321_ (.B1(net384),
    .Y(_1077_),
    .A2(net387),
    .A1(slave_wdata_i_5_));
 sg13g2_o21ai_1 _5322_ (.B1(net380),
    .Y(_1078_),
    .A1(net387),
    .A2(_1076_));
 sg13g2_nand2_1 _5323_ (.Y(_1079_),
    .A(data_csrs_mem_5_),
    .B(_1078_));
 sg13g2_o21ai_1 _5324_ (.B1(_1079_),
    .Y(_0088_),
    .A1(_1076_),
    .A2(_1077_));
 sg13g2_and2_1 _5325_ (.A(net209),
    .B(net165),
    .X(_1080_));
 sg13g2_o21ai_1 _5326_ (.B1(net95),
    .Y(_1081_),
    .A1(net32),
    .A2(_1080_));
 sg13g2_a21oi_2 _5327_ (.B1(net363),
    .Y(_1082_),
    .A2(net351),
    .A1(slave_wdata_i_28_));
 sg13g2_o21ai_1 _5328_ (.B1(net358),
    .Y(_1083_),
    .A1(net351),
    .A2(_1081_));
 sg13g2_nand2_1 _5329_ (.Y(_1084_),
    .A(data_csrs_mem_60_),
    .B(_1083_));
 sg13g2_o21ai_1 _5330_ (.B1(_1084_),
    .Y(_0089_),
    .A1(_1081_),
    .A2(_1082_));
 sg13g2_and2_1 _5331_ (.A(net207),
    .B(net165),
    .X(_1085_));
 sg13g2_o21ai_1 _5332_ (.B1(net95),
    .Y(_1086_),
    .A1(net32),
    .A2(_1085_));
 sg13g2_a21oi_2 _5333_ (.B1(net362),
    .Y(_1087_),
    .A2(net350),
    .A1(slave_wdata_i_29_));
 sg13g2_o21ai_1 _5334_ (.B1(net357),
    .Y(_1088_),
    .A1(net350),
    .A2(_1086_));
 sg13g2_nand2_1 _5335_ (.Y(_1089_),
    .A(data_csrs_mem_61_),
    .B(_1088_));
 sg13g2_o21ai_1 _5336_ (.B1(_1089_),
    .Y(_0090_),
    .A1(_1086_),
    .A2(_1087_));
 sg13g2_and2_1 _5337_ (.A(net203),
    .B(net165),
    .X(_1090_));
 sg13g2_o21ai_1 _5338_ (.B1(net95),
    .Y(_1091_),
    .A1(net25),
    .A2(_1090_));
 sg13g2_a21oi_2 _5339_ (.B1(net362),
    .Y(_1092_),
    .A2(net351),
    .A1(slave_wdata_i_30_));
 sg13g2_o21ai_1 _5340_ (.B1(net357),
    .Y(_1093_),
    .A1(net350),
    .A2(_1091_));
 sg13g2_nand2_1 _5341_ (.Y(_1094_),
    .A(data_csrs_mem_62_),
    .B(_1093_));
 sg13g2_o21ai_1 _5342_ (.B1(_1094_),
    .Y(_0091_),
    .A1(_1091_),
    .A2(_1092_));
 sg13g2_and2_1 _5343_ (.A(net201),
    .B(net165),
    .X(_1095_));
 sg13g2_o21ai_1 _5344_ (.B1(net94),
    .Y(_1096_),
    .A1(net25),
    .A2(_1095_));
 sg13g2_a21oi_2 _5345_ (.B1(net362),
    .Y(_1097_),
    .A2(net350),
    .A1(slave_wdata_i_31_));
 sg13g2_o21ai_1 _5346_ (.B1(net357),
    .Y(_1098_),
    .A1(net350),
    .A2(_1096_));
 sg13g2_nand2_1 _5347_ (.Y(_1099_),
    .A(data_csrs_mem_63_),
    .B(_1098_));
 sg13g2_o21ai_1 _5348_ (.B1(_1099_),
    .Y(_0092_),
    .A1(_1096_),
    .A2(_1097_));
 sg13g2_nor2b_1 _5349_ (.A(net177),
    .B_N(net122),
    .Y(_1100_));
 sg13g2_o21ai_1 _5350_ (.B1(net94),
    .Y(_1101_),
    .A1(net25),
    .A2(_1100_));
 sg13g2_a21oi_2 _5351_ (.B1(net384),
    .Y(_1102_),
    .A2(net386),
    .A1(slave_wdata_i_6_));
 sg13g2_o21ai_1 _5352_ (.B1(net379),
    .Y(_1103_),
    .A1(net386),
    .A2(_1101_));
 sg13g2_nand2_1 _5353_ (.Y(_1104_),
    .A(data_csrs_mem_6_),
    .B(_1103_));
 sg13g2_o21ai_1 _5354_ (.B1(_1104_),
    .Y(_0093_),
    .A1(_1101_),
    .A2(_1102_));
 sg13g2_nor2b_1 _5355_ (.A(net177),
    .B_N(net120),
    .Y(_1105_));
 sg13g2_o21ai_1 _5356_ (.B1(net94),
    .Y(_1106_),
    .A1(net25),
    .A2(_1105_));
 sg13g2_a21oi_2 _5357_ (.B1(net384),
    .Y(_1107_),
    .A2(net386),
    .A1(slave_wdata_i_7_));
 sg13g2_o21ai_1 _5358_ (.B1(net379),
    .Y(_1108_),
    .A1(net386),
    .A2(_1106_));
 sg13g2_nand2_1 _5359_ (.Y(_1109_),
    .A(data_csrs_mem_7_),
    .B(_1108_));
 sg13g2_o21ai_1 _5360_ (.B1(_1109_),
    .Y(_0094_),
    .A1(_1106_),
    .A2(_1107_));
 sg13g2_nor2b_1 _5361_ (.A(net177),
    .B_N(net118),
    .Y(_1110_));
 sg13g2_o21ai_1 _5362_ (.B1(net94),
    .Y(_1111_),
    .A1(net25),
    .A2(_1110_));
 sg13g2_a21oi_2 _5363_ (.B1(net384),
    .Y(_1112_),
    .A2(net374),
    .A1(slave_wdata_i_8_));
 sg13g2_o21ai_1 _5364_ (.B1(net379),
    .Y(_1113_),
    .A1(net374),
    .A2(_1111_));
 sg13g2_nand2_1 _5365_ (.Y(_1114_),
    .A(data_csrs_mem_8_),
    .B(_1113_));
 sg13g2_o21ai_1 _5366_ (.B1(_1114_),
    .Y(_0095_),
    .A1(_1111_),
    .A2(_1112_));
 sg13g2_nor2b_1 _5367_ (.A(net177),
    .B_N(net116),
    .Y(_1115_));
 sg13g2_o21ai_1 _5368_ (.B1(net87),
    .Y(_1116_),
    .A1(net25),
    .A2(_1115_));
 sg13g2_a21oi_2 _5369_ (.B1(net384),
    .Y(_1117_),
    .A2(net374),
    .A1(slave_wdata_i_9_));
 sg13g2_o21ai_1 _5370_ (.B1(net379),
    .Y(_1118_),
    .A1(net374),
    .A2(_1116_));
 sg13g2_nand2_1 _5371_ (.Y(_1119_),
    .A(data_csrs_mem_9_),
    .B(_1118_));
 sg13g2_o21ai_1 _5372_ (.B1(_1119_),
    .Y(_0096_),
    .A1(_1116_),
    .A2(_1117_));
 sg13g2_nand3_1 _5373_ (.B(_0599_),
    .C(_0602_),
    .A(_0596_),
    .Y(_1120_));
 sg13g2_nand3_1 _5374_ (.B(_0893_),
    .C(_1120_),
    .A(debug_req_o),
    .Y(_1121_));
 sg13g2_o21ai_1 _5375_ (.B1(_1121_),
    .Y(_0097_),
    .A1(_1120_),
    .A2(_0684_));
 sg13g2_buf_1 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_2 fanout352 (.A(net354),
    .X(net352));
 sg13g2_mux2_1 _5378_ (.A0(net246),
    .A1(net98),
    .S(_1120_),
    .X(_0098_));
 sg13g2_buf_2 fanout351 (.A(_1053_),
    .X(net351));
 sg13g2_buf_2 fanout350 (.A(net351),
    .X(net350));
 sg13g2_mux2_2 _5381_ (.A0(\i_dm_csrs.i_fifo.mem_q_33_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_67_ ),
    .S(net635),
    .X(dmi_resp_o_33_));
 sg13g2_mux2_2 _5382_ (.A0(\i_dm_csrs.i_fifo.mem_q_32_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_66_ ),
    .S(net634),
    .X(dmi_resp_o_32_));
 sg13g2_mux2_2 _5383_ (.A0(\i_dm_csrs.i_fifo.mem_q_23_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_57_ ),
    .S(net637),
    .X(dmi_resp_o_23_));
 sg13g2_mux2_2 _5384_ (.A0(\i_dm_csrs.i_fifo.mem_q_22_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_56_ ),
    .S(net638),
    .X(dmi_resp_o_22_));
 sg13g2_mux2_2 _5385_ (.A0(\i_dm_csrs.i_fifo.mem_q_21_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_55_ ),
    .S(net637),
    .X(dmi_resp_o_21_));
 sg13g2_mux2_2 _5386_ (.A0(\i_dm_csrs.i_fifo.mem_q_20_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_54_ ),
    .S(net635),
    .X(dmi_resp_o_20_));
 sg13g2_mux2_2 _5387_ (.A0(\i_dm_csrs.i_fifo.mem_q_19_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_53_ ),
    .S(net637),
    .X(dmi_resp_o_19_));
 sg13g2_mux2_2 _5388_ (.A0(\i_dm_csrs.i_fifo.mem_q_18_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_52_ ),
    .S(net635),
    .X(dmi_resp_o_18_));
 sg13g2_mux2_2 _5389_ (.A0(\i_dm_csrs.i_fifo.mem_q_17_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_51_ ),
    .S(net638),
    .X(dmi_resp_o_17_));
 sg13g2_mux2_2 _5390_ (.A0(\i_dm_csrs.i_fifo.mem_q_16_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_50_ ),
    .S(net634),
    .X(dmi_resp_o_16_));
 sg13g2_buf_8 fanout349 (.A(_1903_),
    .X(net349));
 sg13g2_mux2_2 _5392_ (.A0(\i_dm_csrs.i_fifo.mem_q_15_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_49_ ),
    .S(net635),
    .X(dmi_resp_o_15_));
 sg13g2_mux2_2 _5393_ (.A0(\i_dm_csrs.i_fifo.mem_q_14_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_48_ ),
    .S(net638),
    .X(dmi_resp_o_14_));
 sg13g2_mux2_2 _5394_ (.A0(\i_dm_csrs.i_fifo.mem_q_31_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_65_ ),
    .S(net634),
    .X(dmi_resp_o_31_));
 sg13g2_mux2_2 _5395_ (.A0(\i_dm_csrs.i_fifo.mem_q_13_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_47_ ),
    .S(net634),
    .X(dmi_resp_o_13_));
 sg13g2_mux2_2 _5396_ (.A0(\i_dm_csrs.i_fifo.mem_q_12_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_46_ ),
    .S(net637),
    .X(dmi_resp_o_12_));
 sg13g2_mux2_2 _5397_ (.A0(\i_dm_csrs.i_fifo.mem_q_11_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_45_ ),
    .S(net635),
    .X(dmi_resp_o_11_));
 sg13g2_mux2_2 _5398_ (.A0(\i_dm_csrs.i_fifo.mem_q_10_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_44_ ),
    .S(net635),
    .X(dmi_resp_o_10_));
 sg13g2_mux2_2 _5399_ (.A0(\i_dm_csrs.i_fifo.mem_q_9_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_43_ ),
    .S(net637),
    .X(dmi_resp_o_9_));
 sg13g2_mux2_2 _5400_ (.A0(\i_dm_csrs.i_fifo.mem_q_8_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_42_ ),
    .S(net634),
    .X(dmi_resp_o_8_));
 sg13g2_mux2_2 _5401_ (.A0(\i_dm_csrs.i_fifo.mem_q_7_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_41_ ),
    .S(net634),
    .X(dmi_resp_o_7_));
 sg13g2_buf_16 fanout348 (.X(net348),
    .A(net349));
 sg13g2_mux2_2 _5403_ (.A0(\i_dm_csrs.i_fifo.mem_q_6_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_40_ ),
    .S(net635),
    .X(dmi_resp_o_6_));
 sg13g2_mux2_2 _5404_ (.A0(\i_dm_csrs.i_fifo.mem_q_5_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_39_ ),
    .S(net634),
    .X(dmi_resp_o_5_));
 sg13g2_mux2_2 _5405_ (.A0(\i_dm_csrs.i_fifo.mem_q_4_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_38_ ),
    .S(\i_dm_csrs.i_fifo.read_pointer_q ),
    .X(dmi_resp_o_4_));
 sg13g2_mux2_2 _5406_ (.A0(\i_dm_csrs.i_fifo.mem_q_30_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_64_ ),
    .S(net637),
    .X(dmi_resp_o_30_));
 sg13g2_mux2_2 _5407_ (.A0(\i_dm_csrs.i_fifo.mem_q_3_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_37_ ),
    .S(net638),
    .X(dmi_resp_o_3_));
 sg13g2_mux2_2 _5408_ (.A0(\i_dm_csrs.i_fifo.mem_q_2_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_36_ ),
    .S(net638),
    .X(dmi_resp_o_2_));
 sg13g2_mux2_2 _5409_ (.A0(\i_dm_csrs.i_fifo.mem_q_1_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_35_ ),
    .S(net636),
    .X(dmi_resp_o_1_));
 sg13g2_mux2_2 _5410_ (.A0(\i_dm_csrs.i_fifo.mem_q_0_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_34_ ),
    .S(net635),
    .X(dmi_resp_o_0_));
 sg13g2_mux2_2 _5411_ (.A0(\i_dm_csrs.i_fifo.mem_q_29_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_63_ ),
    .S(net636),
    .X(dmi_resp_o_29_));
 sg13g2_mux2_2 _5412_ (.A0(\i_dm_csrs.i_fifo.mem_q_28_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_62_ ),
    .S(net636),
    .X(dmi_resp_o_28_));
 sg13g2_mux2_2 _5413_ (.A0(\i_dm_csrs.i_fifo.mem_q_27_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_61_ ),
    .S(net637),
    .X(dmi_resp_o_27_));
 sg13g2_mux2_2 _5414_ (.A0(\i_dm_csrs.i_fifo.mem_q_26_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_60_ ),
    .S(net637),
    .X(dmi_resp_o_26_));
 sg13g2_mux2_2 _5415_ (.A0(\i_dm_csrs.i_fifo.mem_q_25_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_59_ ),
    .S(net638),
    .X(dmi_resp_o_25_));
 sg13g2_mux2_2 _5416_ (.A0(\i_dm_csrs.i_fifo.mem_q_24_ ),
    .A1(\i_dm_csrs.i_fifo.mem_q_58_ ),
    .S(net634),
    .X(dmi_resp_o_24_));
 sg13g2_or2_2 _5417_ (.X(dmi_resp_valid_o),
    .B(\i_dm_csrs.i_fifo.status_cnt_q_1_ ),
    .A(\i_dm_csrs.i_fifo.status_cnt_q_0_ ));
 sg13g2_buf_16 fanout347 (.X(net347),
    .A(net348));
 sg13g2_buf_16 fanout346 (.X(net346),
    .A(net348));
 sg13g2_buf_8 fanout345 (.A(_1903_),
    .X(net345));
 sg13g2_buf_16 fanout344 (.X(net344),
    .A(net345));
 sg13g2_or2_1 _5422_ (.X(_1132_),
    .B(slave_addr_i_11_),
    .A(slave_addr_i_9_));
 sg13g2_nor2_1 _5423_ (.A(net100),
    .B(net644),
    .Y(_1133_));
 sg13g2_nor3_2 _5424_ (.A(slave_addr_i_0_),
    .B(slave_addr_i_1_),
    .C(slave_addr_i_2_),
    .Y(_1134_));
 sg13g2_nor2b_2 _5425_ (.A(slave_addr_i_7_),
    .B_N(slave_addr_i_8_),
    .Y(_1135_));
 sg13g2_nand3_1 _5426_ (.B(_1134_),
    .C(_1135_),
    .A(_1133_),
    .Y(_1136_));
 sg13g2_or4_2 _5427_ (.A(slave_addr_i_10_),
    .B(_0705_),
    .C(_1132_),
    .D(_1136_),
    .X(_1137_));
 sg13g2_nor3_2 _5428_ (.A(slave_wdata_i_0_),
    .B(net103),
    .C(_1137_),
    .Y(_1138_));
 sg13g2_buf_16 fanout343 (.X(net343),
    .A(net344));
 sg13g2_buf_16 fanout342 (.X(net342),
    .A(net343));
 sg13g2_buf_16 fanout341 (.X(net341),
    .A(net345));
 sg13g2_buf_16 fanout340 (.X(net340),
    .A(net341));
 sg13g2_nand2_1 _5433_ (.Y(_1143_),
    .A(net662),
    .B(_1138_));
 sg13g2_o21ai_1 _5434_ (.B1(_1143_),
    .Y(_1144_),
    .A1(halted),
    .A2(_1138_));
 sg13g2_nor2_2 _5435_ (.A(ndmreset_o),
    .B(_1144_),
    .Y(_0099_));
 sg13g2_inv_1 _5436_ (.Y(_1145_),
    .A(dmi_req_i_40_));
 sg13g2_nand3_1 _5437_ (.B(_1145_),
    .C(_0617_),
    .A(net133),
    .Y(_1146_));
 sg13g2_buf_16 fanout339 (.X(net339),
    .A(net341));
 sg13g2_nor3_2 _5439_ (.A(net162),
    .B(net146),
    .C(net140),
    .Y(_1148_));
 sg13g2_nand2b_1 _5440_ (.Y(_1149_),
    .B(_1148_),
    .A_N(_1146_));
 sg13g2_inv_1 _5441_ (.Y(_1150_),
    .A(_1149_));
 sg13g2_a21oi_2 _5442_ (.B1(net639),
    .Y(_1151_),
    .A2(_1150_),
    .A1(_0901_));
 sg13g2_buf_8 fanout338 (.A(_2010_),
    .X(net338));
 sg13g2_buf_16 fanout337 (.X(net337),
    .A(net338));
 sg13g2_nand2_2 _5445_ (.Y(_1154_),
    .A(\i_dm_csrs.abstractauto_q_0_ ),
    .B(net413));
 sg13g2_o21ai_1 _5446_ (.B1(_1154_),
    .Y(_0100_),
    .A1(_0606_),
    .A2(net413));
 sg13g2_nand2_2 _5447_ (.Y(_1155_),
    .A(\i_dm_csrs.abstractauto_q_16_ ),
    .B(net411));
 sg13g2_o21ai_1 _5448_ (.B1(_1155_),
    .Y(_0101_),
    .A1(_0643_),
    .A2(net411));
 sg13g2_nand2_2 _5449_ (.Y(_1156_),
    .A(\i_dm_csrs.abstractauto_q_17_ ),
    .B(net411));
 sg13g2_o21ai_1 _5450_ (.B1(_1156_),
    .Y(_0102_),
    .A1(_0646_),
    .A2(net411));
 sg13g2_nand2_2 _5451_ (.Y(_1157_),
    .A(\i_dm_csrs.abstractauto_q_18_ ),
    .B(net412));
 sg13g2_o21ai_1 _5452_ (.B1(_1157_),
    .Y(_0103_),
    .A1(_0648_),
    .A2(net412));
 sg13g2_nand2_2 _5453_ (.Y(_1158_),
    .A(\i_dm_csrs.abstractauto_q_19_ ),
    .B(net411));
 sg13g2_o21ai_1 _5454_ (.B1(_1158_),
    .Y(_0104_),
    .A1(_0650_),
    .A2(net411));
 sg13g2_nand2_2 _5455_ (.Y(_1159_),
    .A(\i_dm_csrs.abstractauto_q_1_ ),
    .B(net413));
 sg13g2_o21ai_1 _5456_ (.B1(_1159_),
    .Y(_0105_),
    .A1(_0655_),
    .A2(net413));
 sg13g2_nand2_2 _5457_ (.Y(_1160_),
    .A(\i_dm_csrs.abstractauto_q_20_ ),
    .B(net412));
 sg13g2_o21ai_1 _5458_ (.B1(_1160_),
    .Y(_0106_),
    .A1(_0658_),
    .A2(net412));
 sg13g2_nand2_2 _5459_ (.Y(_1161_),
    .A(\i_dm_csrs.abstractauto_q_21_ ),
    .B(net411));
 sg13g2_o21ai_1 _5460_ (.B1(_1161_),
    .Y(_0107_),
    .A1(_0660_),
    .A2(net411));
 sg13g2_nand2_2 _5461_ (.Y(_1162_),
    .A(\i_dm_csrs.abstractauto_q_22_ ),
    .B(net412));
 sg13g2_o21ai_1 _5462_ (.B1(_1162_),
    .Y(_0108_),
    .A1(_0662_),
    .A2(net412));
 sg13g2_nand2_2 _5463_ (.Y(_1163_),
    .A(net85),
    .B(net799));
 sg13g2_nand2_1 _5464_ (.Y(_1164_),
    .A(\i_dm_csrs.abstractauto_q_23_ ),
    .B(net413));
 sg13g2_o21ai_1 _5465_ (.B1(_1164_),
    .Y(_0109_),
    .A1(net413),
    .A2(_1163_));
 sg13g2_inv_8 _5466_ (.Y(_1165_),
    .A(net83));
 sg13g2_buf_8 fanout336 (.A(net338),
    .X(net336));
 sg13g2_o21ai_1 _5468_ (.B1(_0730_),
    .Y(_1167_),
    .A1(net130),
    .A2(_0729_));
 sg13g2_nor2_1 _5469_ (.A(_0597_),
    .B(_1167_),
    .Y(_1168_));
 sg13g2_nor2b_2 _5470_ (.A(dmi_req_i_33_),
    .B_N(dmi_req_i_32_),
    .Y(_1169_));
 sg13g2_nor2_1 _5471_ (.A(_1168_),
    .B(_1169_),
    .Y(_1170_));
 sg13g2_buf_16 fanout335 (.X(net335),
    .A(net338));
 sg13g2_inv_1 _5473_ (.Y(_1172_),
    .A(net161));
 sg13g2_buf_8 fanout334 (.A(_2010_),
    .X(net334));
 sg13g2_nand2_1 _5475_ (.Y(_1174_),
    .A(net590),
    .B(\i_dm_csrs.abstractauto_q_0_ ));
 sg13g2_buf_16 fanout333 (.X(net333),
    .A(net334));
 sg13g2_buf_16 fanout332 (.X(net332),
    .A(net333));
 sg13g2_nand2_1 _5478_ (.Y(_1177_),
    .A(net183),
    .B(\i_dm_csrs.abstractauto_q_1_ ));
 sg13g2_a21oi_1 _5479_ (.A1(_1174_),
    .A2(_1177_),
    .Y(_1178_),
    .B1(_0896_));
 sg13g2_and2_1 _5480_ (.A(net130),
    .B(_0730_),
    .X(_1179_));
 sg13g2_buf_16 fanout331 (.X(net331),
    .A(net333));
 sg13g2_buf_8 fanout330 (.A(_2010_),
    .X(net330));
 sg13g2_buf_16 fanout329 (.X(net329),
    .A(net330));
 sg13g2_buf_16 fanout328 (.X(net328),
    .A(net330));
 sg13g2_mux4_1 _5485_ (.S0(net169),
    .A0(\i_dm_csrs.abstractauto_q_16_ ),
    .A1(\i_dm_csrs.abstractauto_q_17_ ),
    .A2(\i_dm_csrs.abstractauto_q_18_ ),
    .A3(\i_dm_csrs.abstractauto_q_19_ ),
    .S1(dmi_req_i_35_),
    .X(_1184_));
 sg13g2_buf_8 fanout327 (.A(_2179_),
    .X(net327));
 sg13g2_mux4_1 _5487_ (.S0(net171),
    .A0(\i_dm_csrs.abstractauto_q_20_ ),
    .A1(\i_dm_csrs.abstractauto_q_21_ ),
    .A2(\i_dm_csrs.abstractauto_q_22_ ),
    .A3(\i_dm_csrs.abstractauto_q_23_ ),
    .S1(dmi_req_i_35_),
    .X(_1186_));
 sg13g2_buf_16 fanout326 (.X(net326),
    .A(net327));
 sg13g2_buf_8 fanout325 (.A(net327),
    .X(net325));
 sg13g2_mux2_1 _5490_ (.A0(_1184_),
    .A1(_1186_),
    .S(net136),
    .X(_1189_));
 sg13g2_a22oi_1 _5491_ (.Y(_1190_),
    .B1(net583),
    .B2(_1189_),
    .A2(_1178_),
    .A1(net539));
 sg13g2_nor4_1 _5492_ (.A(net132),
    .B(_0598_),
    .C(_1170_),
    .D(_1190_),
    .Y(_1191_));
 sg13g2_nor2_1 _5493_ (.A(_0623_),
    .B(_1191_),
    .Y(_1192_));
 sg13g2_nor3_1 _5494_ (.A(net597),
    .B(_0900_),
    .C(_1192_),
    .Y(cmd_valid_reg_D));
 sg13g2_nand2_1 _5495_ (.Y(_1193_),
    .A(net109),
    .B(net656));
 sg13g2_nor2_1 _5496_ (.A(_1137_),
    .B(_1193_),
    .Y(_1194_));
 sg13g2_or2_1 _5497_ (.X(_1195_),
    .B(cmd_15_),
    .A(cmd_14_));
 sg13g2_nor2_2 _5498_ (.A(cmd_16_),
    .B(\cmd_16__$_NOT__A_Y ),
    .Y(_1196_));
 sg13g2_nor2b_1 _5499_ (.A(_1196_),
    .B_N(cmd_17_),
    .Y(_1197_));
 sg13g2_mux2_1 _5500_ (.A0(cmd_19_),
    .A1(_1195_),
    .S(_1197_),
    .X(_1198_));
 sg13g2_inv_1 _5501_ (.Y(_1199_),
    .A(cmd_22_));
 sg13g2_nor4_2 _5502_ (.A(cmd_24_),
    .B(cmd_25_),
    .C(cmd_26_),
    .Y(_1200_),
    .D(cmd_27_));
 sg13g2_nor4_2 _5503_ (.A(cmd_28_),
    .B(cmd_29_),
    .C(cmd_30_),
    .Y(_1201_),
    .D(cmd_31_));
 sg13g2_and2_1 _5504_ (.A(_1200_),
    .B(_1201_),
    .X(_1202_));
 sg13g2_buf_16 fanout324 (.X(net324),
    .A(net327));
 sg13g2_nand3_1 _5506_ (.B(cmd_21_),
    .C(cmd_20_),
    .A(\cmd_19__$_OR__B_A_$_OR__Y_B_$_AND__Y_A ),
    .Y(_1204_));
 sg13g2_nand3_1 _5507_ (.B(_1202_),
    .C(_1204_),
    .A(_1199_),
    .Y(_1205_));
 sg13g2_nor2_2 _5508_ (.A(_1198_),
    .B(_1205_),
    .Y(_1206_));
 sg13g2_o21ai_1 _5509_ (.B1(_1206_),
    .Y(_1207_),
    .A1(halted),
    .A2(_0900_));
 sg13g2_nand3_1 _5510_ (.B(_1149_),
    .C(_1167_),
    .A(_0622_),
    .Y(_1208_));
 sg13g2_buf_8 fanout323 (.A(_2179_),
    .X(net323));
 sg13g2_nor2_1 _5512_ (.A(net161),
    .B(net600),
    .Y(_1210_));
 sg13g2_nor2b_2 _5513_ (.A(_0618_),
    .B_N(net548),
    .Y(_1211_));
 sg13g2_nand2_1 _5514_ (.Y(_1212_),
    .A(net141),
    .B(_1211_));
 sg13g2_a21oi_1 _5515_ (.A1(net118),
    .A2(_0609_),
    .Y(_1213_),
    .B1(_1212_));
 sg13g2_nor4_2 _5516_ (.A(\i_dm_csrs.cmderr_q_1_ ),
    .B(\i_dm_csrs.cmderr_q_2_ ),
    .C(_0614_),
    .Y(_1214_),
    .D(_0609_));
 sg13g2_or2_1 _5517_ (.X(_1215_),
    .B(_1214_),
    .A(\i_dm_csrs.cmderr_q_0_ ));
 sg13g2_o21ai_1 _5518_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1208_),
    .A2(_1213_));
 sg13g2_nor2_1 _5519_ (.A(net556),
    .B(_1167_),
    .Y(_1217_));
 sg13g2_nand2_2 _5520_ (.Y(_1218_),
    .A(net44),
    .B(_1169_));
 sg13g2_nor3_1 _5521_ (.A(\i_dm_csrs.cmderr_q_1_ ),
    .B(\i_dm_csrs.cmderr_q_2_ ),
    .C(_1218_),
    .Y(_1219_));
 sg13g2_a21oi_1 _5522_ (.A1(_1217_),
    .A2(_1219_),
    .Y(_1220_),
    .B1(\i_dm_csrs.cmderr_q_0_ ));
 sg13g2_inv_1 _5523_ (.Y(_1221_),
    .A(dmi_req_i_38_));
 sg13g2_buf_16 fanout322 (.X(net322),
    .A(net323));
 sg13g2_nand2_1 _5525_ (.Y(_1223_),
    .A(net155),
    .B(_0617_));
 sg13g2_o21ai_1 _5526_ (.B1(_1223_),
    .Y(_1224_),
    .A1(net147),
    .A2(dmi_req_i_38_));
 sg13g2_a22oi_1 _5527_ (.Y(_1225_),
    .B1(_1224_),
    .B2(net141),
    .A2(_1221_),
    .A1(net131));
 sg13g2_nand2b_1 _5528_ (.Y(_1226_),
    .B(_0616_),
    .A_N(_1225_));
 sg13g2_a21oi_1 _5529_ (.A1(_1149_),
    .A2(_1226_),
    .Y(_1227_),
    .B1(_0614_));
 sg13g2_or2_1 _5530_ (.X(_1228_),
    .B(_1227_),
    .A(_1220_));
 sg13g2_a22oi_1 _5531_ (.Y(_1229_),
    .B1(_1216_),
    .B2(_1228_),
    .A2(_1207_),
    .A1(cmd_valid));
 sg13g2_buf_16 fanout321 (.X(net321),
    .A(net322));
 sg13g2_o21ai_1 _5533_ (.B1(net98),
    .Y(_1231_),
    .A1(_1194_),
    .A2(_1229_));
 sg13g2_inv_1 _5534_ (.Y(\i_dm_csrs.cmderr_q_0__reg_D ),
    .A(_1231_));
 sg13g2_inv_1 _5535_ (.Y(_1232_),
    .A(_1206_));
 sg13g2_a21oi_1 _5536_ (.A1(cmd_valid),
    .A2(_1232_),
    .Y(_1233_),
    .B1(_1194_));
 sg13g2_nand2_1 _5537_ (.Y(_1234_),
    .A(halted),
    .B(_1206_));
 sg13g2_nand3_1 _5538_ (.B(net556),
    .C(_1234_),
    .A(cmd_valid),
    .Y(_1235_));
 sg13g2_buf_16 fanout320 (.X(net320),
    .A(net322));
 sg13g2_nor3_2 _5540_ (.A(_0732_),
    .B(_1208_),
    .C(_1212_),
    .Y(_1237_));
 sg13g2_nand2_1 _5541_ (.Y(_1238_),
    .A(net117),
    .B(_1237_));
 sg13g2_nand3_1 _5542_ (.B(_1235_),
    .C(_1238_),
    .A(\i_dm_csrs.cmderr_q_1_ ),
    .Y(_1239_));
 sg13g2_a21oi_1 _5543_ (.A1(_1233_),
    .A2(_1239_),
    .Y(\i_dm_csrs.cmderr_q_1__reg_D ),
    .B1(net597));
 sg13g2_buf_8 fanout319 (.A(_2179_),
    .X(net319));
 sg13g2_nand2_1 _5545_ (.Y(_1241_),
    .A(net244),
    .B(_1237_));
 sg13g2_nand2_1 _5546_ (.Y(_1242_),
    .A(\i_dm_csrs.cmderr_q_2_ ),
    .B(_1241_));
 sg13g2_nand2_1 _5547_ (.Y(_1243_),
    .A(net95),
    .B(_1233_));
 sg13g2_a21oi_1 _5548_ (.A1(_1235_),
    .A2(_1242_),
    .Y(\i_dm_csrs.cmderr_q_2__reg_D ),
    .B1(_1243_));
 sg13g2_mux2_1 _5549_ (.A0(net203),
    .A1(\i_dm_csrs.resumereq_o ),
    .S(_1120_),
    .X(_1244_));
 sg13g2_buf_16 fanout318 (.X(net318),
    .A(net319));
 sg13g2_buf_16 fanout317 (.X(net317),
    .A(net319));
 sg13g2_a21oi_1 _5552_ (.A1(\i_dm_csrs.resumereq_o ),
    .A2(\i_dm_csrs.dmstatus_16_ ),
    .Y(_1247_),
    .B1(net598));
 sg13g2_and2_1 _5553_ (.A(_1244_),
    .B(_1247_),
    .X(\i_dm_csrs.resumereq_o_reg_D ));
 sg13g2_and2_2 _5554_ (.A(net130),
    .B(_0594_),
    .X(_1248_));
 sg13g2_and2_1 _5555_ (.A(net132),
    .B(_1248_),
    .X(_1249_));
 sg13g2_buf_8 fanout316 (.A(_2264_),
    .X(net316));
 sg13g2_buf_16 fanout315 (.X(net315),
    .A(net316));
 sg13g2_inv_1 _5558_ (.Y(_1252_),
    .A(\i_dm_csrs.sbcs_q_22_ ));
 sg13g2_buf_16 fanout314 (.X(net314),
    .A(net315));
 sg13g2_buf_16 fanout313 (.X(net313),
    .A(net315));
 sg13g2_nor3_2 _5561_ (.A(\i_dm_sba.state_q_2_ ),
    .B(\i_dm_sba.state_q_0_ ),
    .C(\i_dm_sba.state_q_1_ ),
    .Y(_1255_));
 sg13g2_a21oi_1 _5562_ (.A1(_1252_),
    .A2(net41),
    .Y(_1256_),
    .B1(_0896_));
 sg13g2_a21oi_1 _5563_ (.A1(net42),
    .A2(_1256_),
    .Y(_1257_),
    .B1(_1217_));
 sg13g2_inv_1 _5564_ (.Y(_1258_),
    .A(net132));
 sg13g2_nor2_1 _5565_ (.A(net134),
    .B(_1258_),
    .Y(_1259_));
 sg13g2_buf_8 fanout312 (.A(_2264_),
    .X(net312));
 sg13g2_nor2_1 _5567_ (.A(net600),
    .B(net46),
    .Y(_1261_));
 sg13g2_o21ai_1 _5568_ (.B1(net178),
    .Y(_1262_),
    .A1(_1259_),
    .A2(_1261_));
 sg13g2_nand3_1 _5569_ (.B(net134),
    .C(net132),
    .A(net589),
    .Y(_1263_));
 sg13g2_a21o_1 _5570_ (.A2(_1263_),
    .A1(_1262_),
    .B1(net131),
    .X(_1264_));
 sg13g2_o21ai_1 _5571_ (.B1(dmi_req_i_38_),
    .Y(_1265_),
    .A1(net130),
    .A2(_0729_));
 sg13g2_nand2_1 _5572_ (.Y(_1266_),
    .A(net156),
    .B(net132));
 sg13g2_o21ai_1 _5573_ (.B1(_1266_),
    .Y(_1267_),
    .A1(net132),
    .A2(_1265_));
 sg13g2_o21ai_1 _5574_ (.B1(_1258_),
    .Y(_1268_),
    .A1(net130),
    .A2(_0729_));
 sg13g2_and2_1 _5575_ (.A(_1221_),
    .B(_1268_),
    .X(_1269_));
 sg13g2_nor4_2 _5576_ (.A(dmi_req_i_40_),
    .B(_1218_),
    .C(_1267_),
    .Y(_1270_),
    .D(_1269_));
 sg13g2_nor2_2 _5577_ (.A(net161),
    .B(net140),
    .Y(_1271_));
 sg13g2_nor3_1 _5578_ (.A(_1145_),
    .B(net131),
    .C(dmi_req_i_38_),
    .Y(_1272_));
 sg13g2_a22oi_1 _5579_ (.Y(_1273_),
    .B1(_1272_),
    .B2(_1271_),
    .A2(_1248_),
    .A1(net134));
 sg13g2_nor3_1 _5580_ (.A(net147),
    .B(net133),
    .C(_1273_),
    .Y(_1274_));
 sg13g2_a21oi_1 _5581_ (.A1(_1271_),
    .A2(net42),
    .Y(_1275_),
    .B1(_1274_));
 sg13g2_nor2_1 _5582_ (.A(_1218_),
    .B(_1275_),
    .Y(_1276_));
 sg13g2_a21oi_2 _5583_ (.B1(_1276_),
    .Y(_1277_),
    .A2(_1270_),
    .A1(_1264_));
 sg13g2_buf_16 fanout311 (.X(net311),
    .A(net312));
 sg13g2_nand2_2 _5585_ (.Y(_1279_),
    .A(net133),
    .B(_1248_));
 sg13g2_o21ai_1 _5586_ (.B1(_1279_),
    .Y(_1280_),
    .A1(net146),
    .A2(_1146_));
 sg13g2_a22oi_1 _5587_ (.Y(_1281_),
    .B1(_1280_),
    .B2(_1271_),
    .A2(net43),
    .A1(net600));
 sg13g2_nand2_1 _5588_ (.Y(_1282_),
    .A(_1226_),
    .B(_1281_));
 sg13g2_nor2_1 _5589_ (.A(net600),
    .B(_1271_),
    .Y(_1283_));
 sg13g2_o21ai_1 _5590_ (.B1(net556),
    .Y(_1284_),
    .A1(_1279_),
    .A2(_1283_));
 sg13g2_buf_16 fanout310 (.X(net310),
    .A(net311));
 sg13g2_buf_16 fanout309 (.X(net309),
    .A(net310));
 sg13g2_o21ai_1 _5593_ (.B1(_1271_),
    .Y(_1287_),
    .A1(net600),
    .A2(_1252_));
 sg13g2_o21ai_1 _5594_ (.B1(_1287_),
    .Y(_1288_),
    .A1(net148),
    .A2(\i_dm_csrs.sbcs_q_22_ ));
 sg13g2_nand3_1 _5595_ (.B(_1288_),
    .C(net41),
    .A(net43),
    .Y(_1289_));
 sg13g2_nand4_1 _5596_ (.B(_1282_),
    .C(_1284_),
    .A(_0599_),
    .Y(_1290_),
    .D(_1289_));
 sg13g2_o21ai_1 _5597_ (.B1(_1290_),
    .Y(_1291_),
    .A1(_1257_),
    .A2(net405));
 sg13g2_and2_1 _5598_ (.A(\i_dm_csrs.i_fifo.write_pointer_n ),
    .B(net44),
    .X(_1292_));
 sg13g2_buf_16 fanout308 (.X(net308),
    .A(net310));
 sg13g2_buf_16 fanout307 (.X(net307),
    .A(net312));
 sg13g2_mux2_1 _5601_ (.A0(\i_dm_csrs.i_fifo.mem_q_0_ ),
    .A1(_1291_),
    .S(net489),
    .X(_0110_));
 sg13g2_buf_16 fanout306 (.X(net306),
    .A(net307));
 sg13g2_buf_16 fanout305 (.X(net305),
    .A(net307));
 sg13g2_buf_8 fanout304 (.A(_2366_),
    .X(net304));
 sg13g2_buf_16 fanout303 (.X(net303),
    .A(net304));
 sg13g2_mux4_1 _5606_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_8_ ),
    .A1(\i_dm_csrs.progbuf_o_72_ ),
    .A2(\i_dm_csrs.progbuf_o_40_ ),
    .A3(\i_dm_csrs.progbuf_o_104_ ),
    .S1(net194),
    .X(_1299_));
 sg13g2_mux4_1 _5607_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_136_ ),
    .A1(\i_dm_csrs.progbuf_o_200_ ),
    .A2(\i_dm_csrs.progbuf_o_168_ ),
    .A3(\i_dm_csrs.progbuf_o_232_ ),
    .S1(net194),
    .X(_1300_));
 sg13g2_buf_16 fanout302 (.X(net302),
    .A(net303));
 sg13g2_buf_16 fanout301 (.X(net301),
    .A(net302));
 sg13g2_mux2_2 _5610_ (.A0(_1299_),
    .A1(_1300_),
    .S(net139),
    .X(_1303_));
 sg13g2_nand3_1 _5611_ (.B(\i_dm_csrs.cmderr_q_0_ ),
    .C(_1211_),
    .A(net142),
    .Y(_1304_));
 sg13g2_buf_8 fanout300 (.A(_2366_),
    .X(net300));
 sg13g2_buf_16 fanout299 (.X(net299),
    .A(net300));
 sg13g2_nand2_1 _5614_ (.Y(_1307_),
    .A(net155),
    .B(\i_dm_csrs.sbaddr_q_40_ ));
 sg13g2_buf_16 fanout298 (.X(net298),
    .A(net299));
 sg13g2_buf_16 fanout297 (.X(net297),
    .A(net299));
 sg13g2_nand3_1 _5617_ (.B(net601),
    .C(master_add_o_8_),
    .A(net184),
    .Y(_1310_));
 sg13g2_o21ai_1 _5618_ (.B1(_1310_),
    .Y(_1311_),
    .A1(net162),
    .A2(_1307_));
 sg13g2_nand3_1 _5619_ (.B(net42),
    .C(_1311_),
    .A(net47),
    .Y(_1312_));
 sg13g2_buf_16 fanout296 (.X(net296),
    .A(net300));
 sg13g2_mux2_1 _5621_ (.A0(\i_dm_csrs.sbdata_o_8_ ),
    .A1(\i_dm_csrs.sbdata_q_40_ ),
    .S(net172),
    .X(_1314_));
 sg13g2_or3_2 _5622_ (.A(\i_dm_sba.state_q_2_ ),
    .B(\i_dm_sba.state_q_0_ ),
    .C(\i_dm_sba.state_q_1_ ),
    .X(_1315_));
 sg13g2_nor3_2 _5623_ (.A(\i_dm_csrs.sbcs_q_22_ ),
    .B(_0896_),
    .C(_1315_),
    .Y(_1316_));
 sg13g2_and2_1 _5624_ (.A(net42),
    .B(_1316_),
    .X(_1317_));
 sg13g2_buf_16 fanout295 (.X(net295),
    .A(net296));
 sg13g2_nand3b_1 _5626_ (.B(_1258_),
    .C(net47),
    .Y(_1319_),
    .A_N(_0595_));
 sg13g2_buf_8 fanout294 (.A(net300),
    .X(net294));
 sg13g2_buf_16 fanout293 (.X(net293),
    .A(net300));
 sg13g2_nor2b_1 _5629_ (.A(net155),
    .B_N(net161),
    .Y(_1322_));
 sg13g2_nor2b_2 _5630_ (.A(unavailable_i),
    .B_N(net580),
    .Y(_1323_));
 sg13g2_a22oi_1 _5631_ (.Y(_1324_),
    .B1(_1323_),
    .B2(halted),
    .A2(net547),
    .A1(hartinfo_i_8_));
 sg13g2_mux2_1 _5632_ (.A0(data_csrs_mem_8_),
    .A1(data_csrs_mem_40_),
    .S(net161),
    .X(_1325_));
 sg13g2_and2_1 _5633_ (.A(net134),
    .B(net581),
    .X(_1326_));
 sg13g2_nor2b_1 _5634_ (.A(_1146_),
    .B_N(_1326_),
    .Y(_1327_));
 sg13g2_buf_8 fanout292 (.A(_2449_),
    .X(net292));
 sg13g2_a22oi_1 _5636_ (.Y(_1329_),
    .B1(net535),
    .B2(next_dm_addr_i_8_),
    .A2(_1325_),
    .A1(net538));
 sg13g2_o21ai_1 _5637_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1319_),
    .A2(_1324_));
 sg13g2_a21oi_1 _5638_ (.A1(_1314_),
    .A2(net485),
    .Y(_1331_),
    .B1(_1330_));
 sg13g2_nand3_1 _5639_ (.B(_1312_),
    .C(_1331_),
    .A(_1304_),
    .Y(_1332_));
 sg13g2_a21oi_2 _5640_ (.B1(_1332_),
    .Y(_1333_),
    .A2(_1303_),
    .A1(net584));
 sg13g2_nor2_2 _5641_ (.A(net409),
    .B(_1333_),
    .Y(_1334_));
 sg13g2_mux2_1 _5642_ (.A0(\i_dm_csrs.i_fifo.mem_q_10_ ),
    .A1(_1334_),
    .S(net489),
    .X(_0111_));
 sg13g2_mux4_1 _5643_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_9_ ),
    .A1(\i_dm_csrs.progbuf_o_73_ ),
    .A2(\i_dm_csrs.progbuf_o_41_ ),
    .A3(\i_dm_csrs.progbuf_o_105_ ),
    .S1(net194),
    .X(_1335_));
 sg13g2_mux4_1 _5644_ (.S0(net148),
    .A0(\i_dm_csrs.progbuf_o_137_ ),
    .A1(\i_dm_csrs.progbuf_o_201_ ),
    .A2(\i_dm_csrs.progbuf_o_169_ ),
    .A3(\i_dm_csrs.progbuf_o_233_ ),
    .S1(net194),
    .X(_1336_));
 sg13g2_mux2_1 _5645_ (.A0(_1335_),
    .A1(_1336_),
    .S(net136),
    .X(_1337_));
 sg13g2_nand3_1 _5646_ (.B(\i_dm_csrs.cmderr_q_1_ ),
    .C(_1211_),
    .A(net142),
    .Y(_1338_));
 sg13g2_nand2_1 _5647_ (.Y(_1339_),
    .A(net155),
    .B(\i_dm_csrs.sbaddr_q_41_ ));
 sg13g2_nand3_1 _5648_ (.B(net602),
    .C(master_add_o_9_),
    .A(net184),
    .Y(_1340_));
 sg13g2_o21ai_1 _5649_ (.B1(_1340_),
    .Y(_1341_),
    .A1(net162),
    .A2(_1339_));
 sg13g2_nand3_1 _5650_ (.B(net42),
    .C(_1341_),
    .A(net47),
    .Y(_1342_));
 sg13g2_mux2_1 _5651_ (.A0(\i_dm_csrs.sbdata_o_9_ ),
    .A1(\i_dm_csrs.sbdata_q_41_ ),
    .S(net164),
    .X(_1343_));
 sg13g2_a22oi_1 _5652_ (.Y(_1344_),
    .B1(_1323_),
    .B2(halted),
    .A2(net547),
    .A1(hartinfo_i_9_));
 sg13g2_mux2_1 _5653_ (.A0(data_csrs_mem_9_),
    .A1(data_csrs_mem_41_),
    .S(net161),
    .X(_1345_));
 sg13g2_a22oi_1 _5654_ (.Y(_1346_),
    .B1(_1345_),
    .B2(net538),
    .A2(net533),
    .A1(next_dm_addr_i_9_));
 sg13g2_o21ai_1 _5655_ (.B1(_1346_),
    .Y(_1347_),
    .A1(_1319_),
    .A2(_1344_));
 sg13g2_a21oi_1 _5656_ (.A1(net485),
    .A2(_1343_),
    .Y(_1348_),
    .B1(_1347_));
 sg13g2_nand3_1 _5657_ (.B(_1342_),
    .C(_1348_),
    .A(_1338_),
    .Y(_1349_));
 sg13g2_a21oi_2 _5658_ (.B1(_1349_),
    .Y(_1350_),
    .A2(_1337_),
    .A1(net584));
 sg13g2_nor2_2 _5659_ (.A(net406),
    .B(_1350_),
    .Y(_1351_));
 sg13g2_mux2_1 _5660_ (.A0(\i_dm_csrs.i_fifo.mem_q_11_ ),
    .A1(_1351_),
    .S(net489),
    .X(_0112_));
 sg13g2_mux4_1 _5661_ (.S0(net148),
    .A0(\i_dm_csrs.progbuf_o_10_ ),
    .A1(\i_dm_csrs.progbuf_o_74_ ),
    .A2(\i_dm_csrs.progbuf_o_42_ ),
    .A3(\i_dm_csrs.progbuf_o_106_ ),
    .S1(net194),
    .X(_1352_));
 sg13g2_mux4_1 _5662_ (.S0(net148),
    .A0(\i_dm_csrs.progbuf_o_138_ ),
    .A1(\i_dm_csrs.progbuf_o_202_ ),
    .A2(\i_dm_csrs.progbuf_o_170_ ),
    .A3(\i_dm_csrs.progbuf_o_234_ ),
    .S1(net193),
    .X(_1353_));
 sg13g2_mux2_1 _5663_ (.A0(_1352_),
    .A1(_1353_),
    .S(net136),
    .X(_1354_));
 sg13g2_and2_2 _5664_ (.A(_1248_),
    .B(_1259_),
    .X(_1355_));
 sg13g2_buf_16 fanout291 (.X(net291),
    .A(net292));
 sg13g2_buf_16 fanout290 (.X(net290),
    .A(net291));
 sg13g2_nor2b_2 _5667_ (.A(net155),
    .B_N(\i_dm_csrs.sbcs_q_0_ ),
    .Y(_1358_));
 sg13g2_a21oi_1 _5668_ (.A1(net155),
    .A2(\i_dm_csrs.sbaddr_q_42_ ),
    .Y(_1359_),
    .B1(_1358_));
 sg13g2_nand3_1 _5669_ (.B(net601),
    .C(master_add_o_10_),
    .A(net183),
    .Y(_1360_));
 sg13g2_o21ai_1 _5670_ (.B1(_1360_),
    .Y(_1361_),
    .A1(net173),
    .A2(_1359_));
 sg13g2_nand2_1 _5671_ (.Y(_1362_),
    .A(net531),
    .B(_1361_));
 sg13g2_and2_1 _5672_ (.A(net135),
    .B(_1211_),
    .X(_1363_));
 sg13g2_and2_1 _5673_ (.A(_0596_),
    .B(net548),
    .X(_1364_));
 sg13g2_buf_16 fanout289 (.X(net289),
    .A(net291));
 sg13g2_a22oi_1 _5675_ (.Y(_1366_),
    .B1(net528),
    .B2(hartinfo_i_10_),
    .A2(_1363_),
    .A1(\i_dm_csrs.cmderr_q_2_ ));
 sg13g2_mux2_1 _5676_ (.A0(\i_dm_csrs.sbdata_o_10_ ),
    .A1(\i_dm_csrs.sbdata_q_42_ ),
    .S(net169),
    .X(_1367_));
 sg13g2_nor2b_1 _5677_ (.A(net177),
    .B_N(data_csrs_mem_10_),
    .Y(_1368_));
 sg13g2_a21oi_1 _5678_ (.A1(data_csrs_mem_42_),
    .A2(net183),
    .Y(_1369_),
    .B1(_1368_));
 sg13g2_nand3_1 _5679_ (.B(_0596_),
    .C(_1323_),
    .A(\i_dm_csrs.dmstatus_11__$_AND__Y_A ),
    .Y(_1370_));
 sg13g2_o21ai_1 _5680_ (.B1(_1370_),
    .Y(_1371_),
    .A1(_0731_),
    .A2(_1369_));
 sg13g2_a221oi_1 _5681_ (.B2(net483),
    .C1(_1371_),
    .B1(_1367_),
    .A1(next_dm_addr_i_10_),
    .Y(_1372_),
    .A2(net533));
 sg13g2_nand3_1 _5682_ (.B(_1366_),
    .C(_1372_),
    .A(_1362_),
    .Y(_1373_));
 sg13g2_a21oi_2 _5683_ (.B1(_1373_),
    .Y(_1374_),
    .A2(_1354_),
    .A1(net585));
 sg13g2_nor2_2 _5684_ (.A(net407),
    .B(_1374_),
    .Y(_1375_));
 sg13g2_mux2_1 _5685_ (.A0(\i_dm_csrs.i_fifo.mem_q_12_ ),
    .A1(_1375_),
    .S(net491),
    .X(_0113_));
 sg13g2_buf_8 fanout288 (.A(_2449_),
    .X(net288));
 sg13g2_mux4_1 _5687_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_11_ ),
    .A1(\i_dm_csrs.progbuf_o_75_ ),
    .A2(\i_dm_csrs.progbuf_o_43_ ),
    .A3(\i_dm_csrs.progbuf_o_107_ ),
    .S1(net192),
    .X(_1377_));
 sg13g2_buf_16 fanout287 (.X(net287),
    .A(net288));
 sg13g2_buf_16 fanout286 (.X(net286),
    .A(net287));
 sg13g2_mux4_1 _5690_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_139_ ),
    .A1(\i_dm_csrs.progbuf_o_203_ ),
    .A2(\i_dm_csrs.progbuf_o_171_ ),
    .A3(\i_dm_csrs.progbuf_o_235_ ),
    .S1(net196),
    .X(_1380_));
 sg13g2_mux2_1 _5691_ (.A0(_1377_),
    .A1(_1380_),
    .S(net139),
    .X(_1381_));
 sg13g2_nand2_1 _5692_ (.Y(_1382_),
    .A(net582),
    .B(_1381_));
 sg13g2_mux2_1 _5693_ (.A0(\i_dm_csrs.sbdata_o_11_ ),
    .A1(\i_dm_csrs.sbdata_q_43_ ),
    .S(net170),
    .X(_1383_));
 sg13g2_buf_8 fanout285 (.A(_2449_),
    .X(net285));
 sg13g2_buf_16 fanout284 (.X(net284),
    .A(net285));
 sg13g2_nand2_1 _5696_ (.Y(_1386_),
    .A(next_dm_addr_i_11_),
    .B(net533));
 sg13g2_nand2_1 _5697_ (.Y(_1387_),
    .A(net156),
    .B(\i_dm_csrs.sbaddr_q_43_ ));
 sg13g2_nand3_1 _5698_ (.B(net601),
    .C(master_add_o_11_),
    .A(net184),
    .Y(_1388_));
 sg13g2_o21ai_1 _5699_ (.B1(_1388_),
    .Y(_1389_),
    .A1(net163),
    .A2(_1387_));
 sg13g2_mux2_1 _5700_ (.A0(data_csrs_mem_11_),
    .A1(data_csrs_mem_43_),
    .S(net171),
    .X(_1390_));
 sg13g2_buf_16 fanout283 (.X(net283),
    .A(net285));
 sg13g2_a22oi_1 _5702_ (.Y(_1392_),
    .B1(_1390_),
    .B2(net537),
    .A2(_1389_),
    .A1(net530));
 sg13g2_nand3_1 _5703_ (.B(_1386_),
    .C(_1392_),
    .A(_1370_),
    .Y(_1393_));
 sg13g2_a221oi_1 _5704_ (.B2(net483),
    .C1(_1393_),
    .B1(_1383_),
    .A1(hartinfo_i_11_),
    .Y(_1394_),
    .A2(net527));
 sg13g2_buf_2 fanout282 (.A(_2611_),
    .X(net282));
 sg13g2_a21oi_2 _5706_ (.B1(net405),
    .Y(_1396_),
    .A2(_1394_),
    .A1(_1382_));
 sg13g2_mux2_1 _5707_ (.A0(\i_dm_csrs.i_fifo.mem_q_13_ ),
    .A1(_1396_),
    .S(net488),
    .X(_0114_));
 sg13g2_buf_8 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_16 fanout280 (.X(net280),
    .A(net281));
 sg13g2_and2_1 _5710_ (.A(net144),
    .B(\i_dm_csrs.sbaddr_q_44_ ),
    .X(_1399_));
 sg13g2_a21oi_1 _5711_ (.A1(net605),
    .A2(\i_dm_csrs.sbcs_q_12_ ),
    .Y(_1400_),
    .B1(_1399_));
 sg13g2_nand3_1 _5712_ (.B(net605),
    .C(master_add_o_12_),
    .A(net184),
    .Y(_1401_));
 sg13g2_o21ai_1 _5713_ (.B1(_1401_),
    .Y(_1402_),
    .A1(net174),
    .A2(_1400_));
 sg13g2_buf_8 fanout279 (.A(net282),
    .X(net279));
 sg13g2_mux2_1 _5715_ (.A0(\i_dm_csrs.sbdata_o_12_ ),
    .A1(\i_dm_csrs.sbdata_q_44_ ),
    .S(net174),
    .X(_1404_));
 sg13g2_a22oi_1 _5716_ (.Y(_1405_),
    .B1(_1404_),
    .B2(_1316_),
    .A2(_1402_),
    .A1(net47));
 sg13g2_mux4_1 _5717_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_12_ ),
    .A1(\i_dm_csrs.progbuf_o_76_ ),
    .A2(\i_dm_csrs.progbuf_o_44_ ),
    .A3(\i_dm_csrs.progbuf_o_108_ ),
    .S1(net192),
    .X(_1406_));
 sg13g2_mux4_1 _5718_ (.S0(net144),
    .A0(\i_dm_csrs.progbuf_o_140_ ),
    .A1(\i_dm_csrs.progbuf_o_204_ ),
    .A2(\i_dm_csrs.progbuf_o_172_ ),
    .A3(\i_dm_csrs.progbuf_o_236_ ),
    .S1(net192),
    .X(_1407_));
 sg13g2_mux2_2 _5719_ (.A0(_1406_),
    .A1(_1407_),
    .S(net135),
    .X(_1408_));
 sg13g2_buf_2 fanout278 (.A(_3135_),
    .X(net278));
 sg13g2_a22oi_1 _5721_ (.Y(_1410_),
    .B1(net580),
    .B2(unavailable_i),
    .A2(net547),
    .A1(hartinfo_i_12_));
 sg13g2_mux2_1 _5722_ (.A0(data_csrs_mem_12_),
    .A1(data_csrs_mem_44_),
    .S(net162),
    .X(_1411_));
 sg13g2_a22oi_1 _5723_ (.Y(_1412_),
    .B1(_1411_),
    .B2(net536),
    .A2(net534),
    .A1(next_dm_addr_i_12_));
 sg13g2_o21ai_1 _5724_ (.B1(_1412_),
    .Y(_1413_),
    .A1(_1319_),
    .A2(_1410_));
 sg13g2_a221oi_1 _5725_ (.B2(net582),
    .C1(_1413_),
    .B1(_1408_),
    .A1(_0900_),
    .Y(_1414_),
    .A2(_1363_));
 sg13g2_o21ai_1 _5726_ (.B1(_1414_),
    .Y(_1415_),
    .A1(_1279_),
    .A2(_1405_));
 sg13g2_nor2b_2 _5727_ (.A(net408),
    .B_N(_1415_),
    .Y(_1416_));
 sg13g2_mux2_1 _5728_ (.A0(\i_dm_csrs.i_fifo.mem_q_14_ ),
    .A1(_1416_),
    .S(net492),
    .X(_0115_));
 sg13g2_mux4_1 _5729_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_13_ ),
    .A1(\i_dm_csrs.progbuf_o_77_ ),
    .A2(\i_dm_csrs.progbuf_o_45_ ),
    .A3(\i_dm_csrs.progbuf_o_109_ ),
    .S1(net192),
    .X(_1417_));
 sg13g2_mux4_1 _5730_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_141_ ),
    .A1(\i_dm_csrs.progbuf_o_205_ ),
    .A2(\i_dm_csrs.progbuf_o_173_ ),
    .A3(\i_dm_csrs.progbuf_o_237_ ),
    .S1(net196),
    .X(_1418_));
 sg13g2_mux2_2 _5731_ (.A0(_1417_),
    .A1(_1418_),
    .S(net139),
    .X(_1419_));
 sg13g2_nand2_1 _5732_ (.Y(_1420_),
    .A(net584),
    .B(_1419_));
 sg13g2_mux2_1 _5733_ (.A0(\i_dm_csrs.sbdata_o_13_ ),
    .A1(\i_dm_csrs.sbdata_q_45_ ),
    .S(net173),
    .X(_1421_));
 sg13g2_and2_1 _5734_ (.A(net144),
    .B(\i_dm_csrs.sbaddr_q_45_ ),
    .X(_1422_));
 sg13g2_a21oi_1 _5735_ (.A1(net605),
    .A2(\i_dm_csrs.sbcs_q_13_ ),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_nand3_1 _5736_ (.B(net601),
    .C(master_add_o_13_),
    .A(net183),
    .Y(_1424_));
 sg13g2_o21ai_1 _5737_ (.B1(_1424_),
    .Y(_1425_),
    .A1(net164),
    .A2(_1423_));
 sg13g2_a22oi_1 _5738_ (.Y(_1426_),
    .B1(net580),
    .B2(unavailable_i),
    .A2(net547),
    .A1(hartinfo_i_13_));
 sg13g2_mux2_1 _5739_ (.A0(data_csrs_mem_13_),
    .A1(data_csrs_mem_45_),
    .S(net169),
    .X(_1427_));
 sg13g2_a22oi_1 _5740_ (.Y(_1428_),
    .B1(_1427_),
    .B2(net537),
    .A2(net535),
    .A1(next_dm_addr_i_13_));
 sg13g2_o21ai_1 _5741_ (.B1(_1428_),
    .Y(_1429_),
    .A1(_1319_),
    .A2(_1426_));
 sg13g2_a221oi_1 _5742_ (.B2(net531),
    .C1(_1429_),
    .B1(_1425_),
    .A1(net485),
    .Y(_1430_),
    .A2(_1421_));
 sg13g2_a21oi_2 _5743_ (.B1(net410),
    .Y(_1431_),
    .A2(_1430_),
    .A1(_1420_));
 sg13g2_mux2_1 _5744_ (.A0(\i_dm_csrs.i_fifo.mem_q_15_ ),
    .A1(_1431_),
    .S(net489),
    .X(_0116_));
 sg13g2_buf_1 fanout277 (.A(net278),
    .X(net277));
 sg13g2_buf_1 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_mux4_1 _5748_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_14_ ),
    .A1(\i_dm_csrs.progbuf_o_78_ ),
    .A2(\i_dm_csrs.progbuf_o_46_ ),
    .A3(\i_dm_csrs.progbuf_o_110_ ),
    .S1(net197),
    .X(_1435_));
 sg13g2_buf_2 fanout274 (.A(net276),
    .X(net274));
 sg13g2_buf_2 fanout273 (.A(net274),
    .X(net273));
 sg13g2_mux4_1 _5751_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_142_ ),
    .A1(\i_dm_csrs.progbuf_o_206_ ),
    .A2(\i_dm_csrs.progbuf_o_174_ ),
    .A3(\i_dm_csrs.progbuf_o_238_ ),
    .S1(net198),
    .X(_1438_));
 sg13g2_mux2_2 _5752_ (.A0(_1435_),
    .A1(_1438_),
    .S(net137),
    .X(_1439_));
 sg13g2_mux2_1 _5753_ (.A0(\i_dm_csrs.sbdata_o_14_ ),
    .A1(\i_dm_csrs.sbdata_q_46_ ),
    .S(net164),
    .X(_1440_));
 sg13g2_buf_8 fanout272 (.A(_1916_),
    .X(net272));
 sg13g2_and2_1 _5755_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_46_ ),
    .X(_1442_));
 sg13g2_a21oi_1 _5756_ (.A1(net602),
    .A2(\i_dm_csrs.sbcs_q_14_ ),
    .Y(_1443_),
    .B1(_1442_));
 sg13g2_nand3_1 _5757_ (.B(net601),
    .C(master_add_o_14_),
    .A(net183),
    .Y(_1444_));
 sg13g2_o21ai_1 _5758_ (.B1(_1444_),
    .Y(_1445_),
    .A1(net172),
    .A2(_1443_));
 sg13g2_nand2_1 _5759_ (.Y(_1446_),
    .A(net531),
    .B(_1445_));
 sg13g2_nand2_1 _5760_ (.Y(_1447_),
    .A(hartinfo_i_14_),
    .B(net527));
 sg13g2_mux2_1 _5761_ (.A0(data_csrs_mem_14_),
    .A1(data_csrs_mem_46_),
    .S(net164),
    .X(_1448_));
 sg13g2_a22oi_1 _5762_ (.Y(_1449_),
    .B1(_1448_),
    .B2(net538),
    .A2(net535),
    .A1(next_dm_addr_i_14_));
 sg13g2_nand3_1 _5763_ (.B(_1447_),
    .C(_1449_),
    .A(_1446_),
    .Y(_1450_));
 sg13g2_a221oi_1 _5764_ (.B2(net484),
    .C1(_1450_),
    .B1(_1440_),
    .A1(net583),
    .Y(_1451_),
    .A2(_1439_));
 sg13g2_nor2_2 _5765_ (.A(net406),
    .B(_1451_),
    .Y(_1452_));
 sg13g2_mux2_1 _5766_ (.A0(\i_dm_csrs.i_fifo.mem_q_16_ ),
    .A1(_1452_),
    .S(net488),
    .X(_0117_));
 sg13g2_mux4_1 _5767_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_15_ ),
    .A1(\i_dm_csrs.progbuf_o_79_ ),
    .A2(\i_dm_csrs.progbuf_o_47_ ),
    .A3(\i_dm_csrs.progbuf_o_111_ ),
    .S1(net197),
    .X(_1453_));
 sg13g2_mux4_1 _5768_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_143_ ),
    .A1(\i_dm_csrs.progbuf_o_207_ ),
    .A2(\i_dm_csrs.progbuf_o_175_ ),
    .A3(\i_dm_csrs.progbuf_o_239_ ),
    .S1(net198),
    .X(_1454_));
 sg13g2_mux2_2 _5769_ (.A0(_1453_),
    .A1(_1454_),
    .S(net137),
    .X(_1455_));
 sg13g2_mux2_1 _5770_ (.A0(\i_dm_csrs.sbdata_o_15_ ),
    .A1(\i_dm_csrs.sbdata_q_47_ ),
    .S(net164),
    .X(_1456_));
 sg13g2_and2_1 _5771_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_47_ ),
    .X(_1457_));
 sg13g2_a21oi_1 _5772_ (.A1(net603),
    .A2(\i_dm_csrs.sbcs_q_15_ ),
    .Y(_1458_),
    .B1(_1457_));
 sg13g2_nand3_1 _5773_ (.B(net602),
    .C(master_add_o_15_),
    .A(net182),
    .Y(_1459_));
 sg13g2_o21ai_1 _5774_ (.B1(_1459_),
    .Y(_1460_),
    .A1(net172),
    .A2(_1458_));
 sg13g2_nand2_1 _5775_ (.Y(_1461_),
    .A(net531),
    .B(_1460_));
 sg13g2_nand2_1 _5776_ (.Y(_1462_),
    .A(hartinfo_i_15_),
    .B(net528));
 sg13g2_mux2_1 _5777_ (.A0(data_csrs_mem_15_),
    .A1(data_csrs_mem_47_),
    .S(net164),
    .X(_1463_));
 sg13g2_a22oi_1 _5778_ (.Y(_1464_),
    .B1(_1463_),
    .B2(net539),
    .A2(net534),
    .A1(next_dm_addr_i_15_));
 sg13g2_nand3_1 _5779_ (.B(_1462_),
    .C(_1464_),
    .A(_1461_),
    .Y(_1465_));
 sg13g2_a221oi_1 _5780_ (.B2(net484),
    .C1(_1465_),
    .B1(_1456_),
    .A1(net586),
    .Y(_1466_),
    .A2(_1455_));
 sg13g2_nor2_2 _5781_ (.A(net407),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_mux2_1 _5782_ (.A0(\i_dm_csrs.i_fifo.mem_q_17_ ),
    .A1(_1467_),
    .S(net492),
    .X(_0118_));
 sg13g2_mux2_1 _5783_ (.A0(\i_dm_csrs.sbdata_o_16_ ),
    .A1(\i_dm_csrs.sbdata_q_48_ ),
    .S(net169),
    .X(_1468_));
 sg13g2_mux2_1 _5784_ (.A0(\i_dm_csrs.sbautoincrement_o ),
    .A1(\i_dm_csrs.sbaddr_q_48_ ),
    .S(net144),
    .X(_1469_));
 sg13g2_nand2_1 _5785_ (.Y(_1470_),
    .A(net590),
    .B(_1469_));
 sg13g2_nand3_1 _5786_ (.B(net605),
    .C(master_add_o_16_),
    .A(net182),
    .Y(_1471_));
 sg13g2_a21oi_1 _5787_ (.A1(_1470_),
    .A2(_1471_),
    .Y(_1472_),
    .B1(net138));
 sg13g2_a21o_1 _5788_ (.A2(_1468_),
    .A1(_1316_),
    .B1(_1472_),
    .X(_1473_));
 sg13g2_mux4_1 _5789_ (.S0(net148),
    .A0(\i_dm_csrs.progbuf_o_16_ ),
    .A1(\i_dm_csrs.progbuf_o_80_ ),
    .A2(\i_dm_csrs.progbuf_o_48_ ),
    .A3(\i_dm_csrs.progbuf_o_112_ ),
    .S1(net196),
    .X(_1474_));
 sg13g2_buf_16 fanout271 (.X(net271),
    .A(net272));
 sg13g2_buf_8 fanout270 (.A(net272),
    .X(net270));
 sg13g2_mux4_1 _5792_ (.S0(net159),
    .A0(\i_dm_csrs.progbuf_o_144_ ),
    .A1(\i_dm_csrs.progbuf_o_208_ ),
    .A2(\i_dm_csrs.progbuf_o_176_ ),
    .A3(\i_dm_csrs.progbuf_o_240_ ),
    .S1(net199),
    .X(_1477_));
 sg13g2_mux2_1 _5793_ (.A0(_1474_),
    .A1(_1477_),
    .S(net136),
    .X(_1478_));
 sg13g2_a22oi_1 _5794_ (.Y(_1479_),
    .B1(net580),
    .B2(\i_dm_csrs.dmstatus_16_ ),
    .A2(net547),
    .A1(hartinfo_i_16_));
 sg13g2_nor3_2 _5795_ (.A(net148),
    .B(_1258_),
    .C(_0595_),
    .Y(_1480_));
 sg13g2_nand3_1 _5796_ (.B(net135),
    .C(next_dm_addr_i_16_),
    .A(net184),
    .Y(_1481_));
 sg13g2_buf_16 fanout269 (.X(net269),
    .A(net272));
 sg13g2_nand3_1 _5798_ (.B(\i_dm_csrs.abstractauto_q_16_ ),
    .C(net46),
    .A(net588),
    .Y(_1483_));
 sg13g2_nand2_1 _5799_ (.Y(_1484_),
    .A(_1481_),
    .B(_1483_));
 sg13g2_mux2_1 _5800_ (.A0(data_csrs_mem_16_),
    .A1(data_csrs_mem_48_),
    .S(net163),
    .X(_1485_));
 sg13g2_a22oi_1 _5801_ (.Y(_1486_),
    .B1(_1485_),
    .B2(net537),
    .A2(_1484_),
    .A1(net526));
 sg13g2_o21ai_1 _5802_ (.B1(_1486_),
    .Y(_1487_),
    .A1(_1319_),
    .A2(_1479_));
 sg13g2_a221oi_1 _5803_ (.B2(net583),
    .C1(_1487_),
    .B1(_1478_),
    .A1(net43),
    .Y(_1488_),
    .A2(_1473_));
 sg13g2_nor2_2 _5804_ (.A(net406),
    .B(_1488_),
    .Y(_1489_));
 sg13g2_buf_4 fanout268 (.X(net268),
    .A(_1916_));
 sg13g2_mux2_1 _5806_ (.A0(\i_dm_csrs.i_fifo.mem_q_18_ ),
    .A1(_1489_),
    .S(net490),
    .X(_0119_));
 sg13g2_mux2_1 _5807_ (.A0(\i_dm_csrs.sbdata_o_17_ ),
    .A1(\i_dm_csrs.sbdata_q_49_ ),
    .S(net170),
    .X(_1491_));
 sg13g2_mux4_1 _5808_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_17_ ),
    .A1(\i_dm_csrs.progbuf_o_81_ ),
    .A2(\i_dm_csrs.progbuf_o_49_ ),
    .A3(\i_dm_csrs.progbuf_o_113_ ),
    .S1(net199),
    .X(_1492_));
 sg13g2_mux4_1 _5809_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_145_ ),
    .A1(\i_dm_csrs.progbuf_o_209_ ),
    .A2(\i_dm_csrs.progbuf_o_177_ ),
    .A3(\i_dm_csrs.progbuf_o_241_ ),
    .S1(net199),
    .X(_1493_));
 sg13g2_mux2_2 _5810_ (.A0(_1492_),
    .A1(_1493_),
    .S(net136),
    .X(_1494_));
 sg13g2_nand2_2 _5811_ (.Y(_1495_),
    .A(_1248_),
    .B(_1259_));
 sg13g2_inv_2 _5812_ (.Y(_1496_),
    .A(net632));
 sg13g2_buf_16 fanout267 (.X(net267),
    .A(net268));
 sg13g2_nand2_1 _5814_ (.Y(_1498_),
    .A(net160),
    .B(\i_dm_csrs.sbaddr_q_49_ ));
 sg13g2_o21ai_1 _5815_ (.B1(_1498_),
    .Y(_1499_),
    .A1(net148),
    .A2(_1496_));
 sg13g2_a22oi_1 _5816_ (.Y(_1500_),
    .B1(_1499_),
    .B2(net590),
    .A2(_1322_),
    .A1(master_add_o_17_));
 sg13g2_mux2_1 _5817_ (.A0(data_csrs_mem_17_),
    .A1(data_csrs_mem_49_),
    .S(net171),
    .X(_1501_));
 sg13g2_buf_16 fanout266 (.X(net266),
    .A(net267));
 sg13g2_nand3_1 _5819_ (.B(net140),
    .C(next_dm_addr_i_17_),
    .A(net185),
    .Y(_1503_));
 sg13g2_nand3_1 _5820_ (.B(\i_dm_csrs.abstractauto_q_17_ ),
    .C(net45),
    .A(net588),
    .Y(_1504_));
 sg13g2_nand2_1 _5821_ (.Y(_1505_),
    .A(_1503_),
    .B(_1504_));
 sg13g2_a22oi_1 _5822_ (.Y(_1506_),
    .B1(net580),
    .B2(\i_dm_csrs.dmstatus_16_ ),
    .A2(net547),
    .A1(hartinfo_i_17_));
 sg13g2_nor2_1 _5823_ (.A(_1319_),
    .B(_1506_),
    .Y(_1507_));
 sg13g2_a221oi_1 _5824_ (.B2(net526),
    .C1(_1507_),
    .B1(_1505_),
    .A1(net536),
    .Y(_1508_),
    .A2(_1501_));
 sg13g2_o21ai_1 _5825_ (.B1(_1508_),
    .Y(_1509_),
    .A1(_1495_),
    .A2(_1500_));
 sg13g2_a221oi_1 _5826_ (.B2(net587),
    .C1(_1509_),
    .B1(_1494_),
    .A1(net486),
    .Y(_1510_),
    .A2(_1491_));
 sg13g2_nor2_2 _5827_ (.A(net407),
    .B(_1510_),
    .Y(_1511_));
 sg13g2_mux2_1 _5828_ (.A0(\i_dm_csrs.i_fifo.mem_q_19_ ),
    .A1(_1511_),
    .S(net491),
    .X(_0120_));
 sg13g2_mux2_1 _5829_ (.A0(\i_dm_csrs.i_fifo.mem_q_1_ ),
    .A1(_1291_),
    .S(net489),
    .X(_0121_));
 sg13g2_mux2_1 _5830_ (.A0(\i_dm_csrs.sbdata_o_18_ ),
    .A1(\i_dm_csrs.sbdata_q_50_ ),
    .S(net170),
    .X(_1512_));
 sg13g2_mux4_1 _5831_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_18_ ),
    .A1(\i_dm_csrs.progbuf_o_82_ ),
    .A2(\i_dm_csrs.progbuf_o_50_ ),
    .A3(\i_dm_csrs.progbuf_o_114_ ),
    .S1(net199),
    .X(_1513_));
 sg13g2_mux4_1 _5832_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_146_ ),
    .A1(\i_dm_csrs.progbuf_o_210_ ),
    .A2(\i_dm_csrs.progbuf_o_178_ ),
    .A3(\i_dm_csrs.progbuf_o_242_ ),
    .S1(net199),
    .X(_1514_));
 sg13g2_mux2_2 _5833_ (.A0(_1513_),
    .A1(_1514_),
    .S(net136),
    .X(_1515_));
 sg13g2_buf_16 fanout265 (.X(net265),
    .A(net267));
 sg13g2_inv_2 _5835_ (.Y(_1517_),
    .A(net630));
 sg13g2_nand2_1 _5836_ (.Y(_1518_),
    .A(net160),
    .B(\i_dm_csrs.sbaddr_q_50_ ));
 sg13g2_o21ai_1 _5837_ (.B1(_1518_),
    .Y(_1519_),
    .A1(net147),
    .A2(_1517_));
 sg13g2_a22oi_1 _5838_ (.Y(_1520_),
    .B1(_1519_),
    .B2(net590),
    .A2(net581),
    .A1(master_add_o_18_));
 sg13g2_mux2_1 _5839_ (.A0(data_csrs_mem_18_),
    .A1(data_csrs_mem_50_),
    .S(net171),
    .X(_1521_));
 sg13g2_nand3_1 _5840_ (.B(net140),
    .C(next_dm_addr_i_18_),
    .A(net185),
    .Y(_1522_));
 sg13g2_nand3_1 _5841_ (.B(net47),
    .C(\i_dm_csrs.abstractauto_q_18_ ),
    .A(net588),
    .Y(_1523_));
 sg13g2_nand2_1 _5842_ (.Y(_1524_),
    .A(_1522_),
    .B(_1523_));
 sg13g2_a22oi_1 _5843_ (.Y(_1525_),
    .B1(net580),
    .B2(\i_dm_csrs.dmstatus_18_ ),
    .A2(net547),
    .A1(hartinfo_i_18_));
 sg13g2_nor2_1 _5844_ (.A(_1319_),
    .B(_1525_),
    .Y(_1526_));
 sg13g2_a221oi_1 _5845_ (.B2(net526),
    .C1(_1526_),
    .B1(_1524_),
    .A1(net536),
    .Y(_1527_),
    .A2(_1521_));
 sg13g2_o21ai_1 _5846_ (.B1(_1527_),
    .Y(_1528_),
    .A1(_1495_),
    .A2(_1520_));
 sg13g2_a221oi_1 _5847_ (.B2(net587),
    .C1(_1528_),
    .B1(_1515_),
    .A1(net487),
    .Y(_1529_),
    .A2(_1512_));
 sg13g2_nor2_2 _5848_ (.A(net406),
    .B(_1529_),
    .Y(_1530_));
 sg13g2_mux2_1 _5849_ (.A0(\i_dm_csrs.i_fifo.mem_q_20_ ),
    .A1(_1530_),
    .S(net489),
    .X(_0122_));
 sg13g2_mux2_1 _5850_ (.A0(\i_dm_csrs.sbdata_o_19_ ),
    .A1(\i_dm_csrs.sbdata_q_51_ ),
    .S(net170),
    .X(_1531_));
 sg13g2_mux4_1 _5851_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_19_ ),
    .A1(\i_dm_csrs.progbuf_o_83_ ),
    .A2(\i_dm_csrs.progbuf_o_51_ ),
    .A3(\i_dm_csrs.progbuf_o_115_ ),
    .S1(net199),
    .X(_1532_));
 sg13g2_mux4_1 _5852_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_147_ ),
    .A1(\i_dm_csrs.progbuf_o_211_ ),
    .A2(\i_dm_csrs.progbuf_o_179_ ),
    .A3(\i_dm_csrs.progbuf_o_243_ ),
    .S1(net199),
    .X(_1533_));
 sg13g2_mux2_1 _5853_ (.A0(_1532_),
    .A1(_1533_),
    .S(net135),
    .X(_1534_));
 sg13g2_buf_16 fanout264 (.X(net264),
    .A(net268));
 sg13g2_inv_2 _5855_ (.Y(_1536_),
    .A(net628));
 sg13g2_nand2_1 _5856_ (.Y(_1537_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_51_ ));
 sg13g2_o21ai_1 _5857_ (.B1(_1537_),
    .Y(_1538_),
    .A1(net147),
    .A2(_1536_));
 sg13g2_a22oi_1 _5858_ (.Y(_1539_),
    .B1(_1538_),
    .B2(net590),
    .A2(net581),
    .A1(master_add_o_19_));
 sg13g2_mux2_1 _5859_ (.A0(data_csrs_mem_19_),
    .A1(data_csrs_mem_51_),
    .S(net171),
    .X(_1540_));
 sg13g2_nand3_1 _5860_ (.B(net140),
    .C(next_dm_addr_i_19_),
    .A(net185),
    .Y(_1541_));
 sg13g2_nand3_1 _5861_ (.B(net46),
    .C(\i_dm_csrs.abstractauto_q_19_ ),
    .A(net588),
    .Y(_1542_));
 sg13g2_nand2_1 _5862_ (.Y(_1543_),
    .A(_1541_),
    .B(_1542_));
 sg13g2_a22oi_1 _5863_ (.Y(_1544_),
    .B1(net580),
    .B2(\i_dm_csrs.dmstatus_18_ ),
    .A2(net547),
    .A1(hartinfo_i_19_));
 sg13g2_nor2_1 _5864_ (.A(_1319_),
    .B(_1544_),
    .Y(_1545_));
 sg13g2_a221oi_1 _5865_ (.B2(net526),
    .C1(_1545_),
    .B1(_1543_),
    .A1(net536),
    .Y(_1546_),
    .A2(_1540_));
 sg13g2_o21ai_1 _5866_ (.B1(_1546_),
    .Y(_1547_),
    .A1(_1495_),
    .A2(_1539_));
 sg13g2_a221oi_1 _5867_ (.B2(net587),
    .C1(_1547_),
    .B1(_1534_),
    .A1(net486),
    .Y(_1548_),
    .A2(_1531_));
 sg13g2_nor2_2 _5868_ (.A(net407),
    .B(_1548_),
    .Y(_1549_));
 sg13g2_mux2_1 _5869_ (.A0(\i_dm_csrs.i_fifo.mem_q_21_ ),
    .A1(_1549_),
    .S(net491),
    .X(_0123_));
 sg13g2_buf_16 fanout263 (.X(net263),
    .A(net264));
 sg13g2_mux4_1 _5871_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_20_ ),
    .A1(\i_dm_csrs.progbuf_o_84_ ),
    .A2(\i_dm_csrs.progbuf_o_52_ ),
    .A3(\i_dm_csrs.progbuf_o_116_ ),
    .S1(net197),
    .X(_1551_));
 sg13g2_mux4_1 _5872_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_148_ ),
    .A1(\i_dm_csrs.progbuf_o_212_ ),
    .A2(\i_dm_csrs.progbuf_o_180_ ),
    .A3(\i_dm_csrs.progbuf_o_244_ ),
    .S1(net198),
    .X(_1552_));
 sg13g2_mux2_2 _5873_ (.A0(_1551_),
    .A1(_1552_),
    .S(net137),
    .X(_1553_));
 sg13g2_buf_16 fanout262 (.X(net262),
    .A(net264));
 sg13g2_mux2_1 _5875_ (.A0(\i_dm_csrs.sbdata_o_20_ ),
    .A1(\i_dm_csrs.sbdata_q_52_ ),
    .S(net176),
    .X(_1555_));
 sg13g2_and2_1 _5876_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_52_ ),
    .X(_1556_));
 sg13g2_a21oi_1 _5877_ (.A1(net605),
    .A2(\i_dm_csrs.sbcs_q_20_ ),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_nand3_1 _5878_ (.B(net605),
    .C(master_add_o_20_),
    .A(net182),
    .Y(_1558_));
 sg13g2_o21ai_1 _5879_ (.B1(_1558_),
    .Y(_1559_),
    .A1(net174),
    .A2(_1557_));
 sg13g2_nand2_1 _5880_ (.Y(_1560_),
    .A(net532),
    .B(_1559_));
 sg13g2_nand2_1 _5881_ (.Y(_1561_),
    .A(hartinfo_i_20_),
    .B(net529));
 sg13g2_nand3_1 _5882_ (.B(net140),
    .C(next_dm_addr_i_20_),
    .A(net185),
    .Y(_1562_));
 sg13g2_nand3_1 _5883_ (.B(net46),
    .C(\i_dm_csrs.abstractauto_q_20_ ),
    .A(net588),
    .Y(_1563_));
 sg13g2_nand2_1 _5884_ (.Y(_1564_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_buf_8 fanout261 (.A(_2094_),
    .X(net261));
 sg13g2_mux2_1 _5886_ (.A0(data_csrs_mem_20_),
    .A1(data_csrs_mem_52_),
    .S(net189),
    .X(_1566_));
 sg13g2_a22oi_1 _5887_ (.Y(_1567_),
    .B1(_1566_),
    .B2(net540),
    .A2(_1564_),
    .A1(net526));
 sg13g2_nand3_1 _5888_ (.B(_1561_),
    .C(_1567_),
    .A(_1560_),
    .Y(_1568_));
 sg13g2_a221oi_1 _5889_ (.B2(net486),
    .C1(_1568_),
    .B1(_1555_),
    .A1(net586),
    .Y(_1569_),
    .A2(_1553_));
 sg13g2_nor2_2 _5890_ (.A(net408),
    .B(_1569_),
    .Y(_1570_));
 sg13g2_mux2_1 _5891_ (.A0(\i_dm_csrs.i_fifo.mem_q_22_ ),
    .A1(_1570_),
    .S(net492),
    .X(_0124_));
 sg13g2_mux4_1 _5892_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_21_ ),
    .A1(\i_dm_csrs.progbuf_o_85_ ),
    .A2(\i_dm_csrs.progbuf_o_53_ ),
    .A3(\i_dm_csrs.progbuf_o_117_ ),
    .S1(net197),
    .X(_1571_));
 sg13g2_mux4_1 _5893_ (.S0(net146),
    .A0(\i_dm_csrs.progbuf_o_149_ ),
    .A1(\i_dm_csrs.progbuf_o_213_ ),
    .A2(\i_dm_csrs.progbuf_o_181_ ),
    .A3(\i_dm_csrs.progbuf_o_245_ ),
    .S1(net198),
    .X(_1572_));
 sg13g2_mux2_2 _5894_ (.A0(_1571_),
    .A1(_1572_),
    .S(net137),
    .X(_1573_));
 sg13g2_mux2_1 _5895_ (.A0(\i_dm_csrs.sbdata_o_21_ ),
    .A1(\i_dm_csrs.sbdata_q_53_ ),
    .S(net175),
    .X(_1574_));
 sg13g2_and2_1 _5896_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_53_ ),
    .X(_1575_));
 sg13g2_a21oi_1 _5897_ (.A1(net605),
    .A2(\i_dm_csrs.sbcs_q_21_ ),
    .Y(_1576_),
    .B1(_1575_));
 sg13g2_nand3_1 _5898_ (.B(net604),
    .C(master_add_o_21_),
    .A(net186),
    .Y(_1577_));
 sg13g2_o21ai_1 _5899_ (.B1(_1577_),
    .Y(_1578_),
    .A1(net174),
    .A2(_1576_));
 sg13g2_nand2_1 _5900_ (.Y(_1579_),
    .A(net532),
    .B(_1578_));
 sg13g2_buf_16 fanout260 (.X(net260),
    .A(net261));
 sg13g2_nand2_1 _5902_ (.Y(_1581_),
    .A(hartinfo_i_21_),
    .B(net529));
 sg13g2_nand3_1 _5903_ (.B(net140),
    .C(next_dm_addr_i_21_),
    .A(net185),
    .Y(_1582_));
 sg13g2_nand3_1 _5904_ (.B(net46),
    .C(\i_dm_csrs.abstractauto_q_21_ ),
    .A(net588),
    .Y(_1583_));
 sg13g2_nand2_1 _5905_ (.Y(_1584_),
    .A(_1582_),
    .B(_1583_));
 sg13g2_mux2_1 _5906_ (.A0(data_csrs_mem_21_),
    .A1(data_csrs_mem_53_),
    .S(net189),
    .X(_1585_));
 sg13g2_a22oi_1 _5907_ (.Y(_1586_),
    .B1(_1585_),
    .B2(net536),
    .A2(_1584_),
    .A1(net526));
 sg13g2_nand3_1 _5908_ (.B(_1581_),
    .C(_1586_),
    .A(_1579_),
    .Y(_1587_));
 sg13g2_a221oi_1 _5909_ (.B2(net486),
    .C1(_1587_),
    .B1(_1574_),
    .A1(net586),
    .Y(_1588_),
    .A2(_1573_));
 sg13g2_nor2_2 _5910_ (.A(net408),
    .B(_1588_),
    .Y(_1589_));
 sg13g2_mux2_1 _5911_ (.A0(\i_dm_csrs.i_fifo.mem_q_23_ ),
    .A1(_1589_),
    .S(net491),
    .X(_0125_));
 sg13g2_mux4_1 _5912_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_22_ ),
    .A1(\i_dm_csrs.progbuf_o_86_ ),
    .A2(\i_dm_csrs.progbuf_o_54_ ),
    .A3(\i_dm_csrs.progbuf_o_118_ ),
    .S1(net197),
    .X(_1590_));
 sg13g2_mux4_1 _5913_ (.S0(net146),
    .A0(\i_dm_csrs.progbuf_o_150_ ),
    .A1(\i_dm_csrs.progbuf_o_214_ ),
    .A2(\i_dm_csrs.progbuf_o_182_ ),
    .A3(\i_dm_csrs.progbuf_o_246_ ),
    .S1(net198),
    .X(_1591_));
 sg13g2_mux2_1 _5914_ (.A0(_1590_),
    .A1(_1591_),
    .S(net137),
    .X(_1592_));
 sg13g2_mux2_1 _5915_ (.A0(\i_dm_csrs.sbdata_o_22_ ),
    .A1(\i_dm_csrs.sbdata_q_54_ ),
    .S(net175),
    .X(_1593_));
 sg13g2_nand2_1 _5916_ (.Y(_1594_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_54_ ));
 sg13g2_o21ai_1 _5917_ (.B1(_1594_),
    .Y(_1595_),
    .A1(net146),
    .A2(_1252_));
 sg13g2_a22oi_1 _5918_ (.Y(_1596_),
    .B1(_1595_),
    .B2(net590),
    .A2(net581),
    .A1(master_add_o_22_));
 sg13g2_nand3_1 _5919_ (.B(net139),
    .C(next_dm_addr_i_22_),
    .A(net182),
    .Y(_1597_));
 sg13g2_nand3_1 _5920_ (.B(net46),
    .C(\i_dm_csrs.abstractauto_q_22_ ),
    .A(net588),
    .Y(_1598_));
 sg13g2_nand2_1 _5921_ (.Y(_1599_),
    .A(_1597_),
    .B(_1598_));
 sg13g2_nor2b_1 _5922_ (.A(net183),
    .B_N(data_csrs_mem_22_),
    .Y(_1600_));
 sg13g2_a21oi_1 _5923_ (.A1(data_csrs_mem_54_),
    .A2(net179),
    .Y(_1601_),
    .B1(_1600_));
 sg13g2_nor2_1 _5924_ (.A(_0731_),
    .B(_1601_),
    .Y(_1602_));
 sg13g2_a221oi_1 _5925_ (.B2(_1599_),
    .C1(_1602_),
    .B1(net526),
    .A1(hartinfo_i_22_),
    .Y(_1603_),
    .A2(net528));
 sg13g2_o21ai_1 _5926_ (.B1(_1603_),
    .Y(_1604_),
    .A1(_1495_),
    .A2(_1596_));
 sg13g2_a221oi_1 _5927_ (.B2(net485),
    .C1(_1604_),
    .B1(_1593_),
    .A1(net583),
    .Y(_1605_),
    .A2(_1592_));
 sg13g2_nor2_2 _5928_ (.A(net406),
    .B(_1605_),
    .Y(_1606_));
 sg13g2_mux2_1 _5929_ (.A0(\i_dm_csrs.i_fifo.mem_q_24_ ),
    .A1(_1606_),
    .S(net488),
    .X(_0126_));
 sg13g2_mux4_1 _5930_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_23_ ),
    .A1(\i_dm_csrs.progbuf_o_87_ ),
    .A2(\i_dm_csrs.progbuf_o_55_ ),
    .A3(\i_dm_csrs.progbuf_o_119_ ),
    .S1(net196),
    .X(_1607_));
 sg13g2_mux4_1 _5931_ (.S0(net146),
    .A0(\i_dm_csrs.progbuf_o_151_ ),
    .A1(\i_dm_csrs.progbuf_o_215_ ),
    .A2(\i_dm_csrs.progbuf_o_183_ ),
    .A3(\i_dm_csrs.progbuf_o_247_ ),
    .S1(net198),
    .X(_1608_));
 sg13g2_mux2_2 _5932_ (.A0(_1607_),
    .A1(_1608_),
    .S(net137),
    .X(_1609_));
 sg13g2_mux2_1 _5933_ (.A0(\i_dm_csrs.sbdata_o_23_ ),
    .A1(\i_dm_csrs.sbdata_q_55_ ),
    .S(net175),
    .X(_1610_));
 sg13g2_and2_1 _5934_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_55_ ),
    .X(_1611_));
 sg13g2_a21oi_1 _5935_ (.A1(net604),
    .A2(\i_dm_csrs.sbcs_q_23_ ),
    .Y(_1612_),
    .B1(_1611_));
 sg13g2_nand3_1 _5936_ (.B(net604),
    .C(master_add_o_23_),
    .A(net186),
    .Y(_1613_));
 sg13g2_o21ai_1 _5937_ (.B1(_1613_),
    .Y(_1614_),
    .A1(net174),
    .A2(_1612_));
 sg13g2_nand2_1 _5938_ (.Y(_1615_),
    .A(net532),
    .B(_1614_));
 sg13g2_nand2_1 _5939_ (.Y(_1616_),
    .A(hartinfo_i_23_),
    .B(net529));
 sg13g2_nand3_1 _5940_ (.B(net139),
    .C(next_dm_addr_i_23_),
    .A(net184),
    .Y(_1617_));
 sg13g2_nand3_1 _5941_ (.B(net46),
    .C(\i_dm_csrs.abstractauto_q_23_ ),
    .A(net588),
    .Y(_1618_));
 sg13g2_nand2_1 _5942_ (.Y(_1619_),
    .A(_1617_),
    .B(_1618_));
 sg13g2_mux2_1 _5943_ (.A0(data_csrs_mem_23_),
    .A1(data_csrs_mem_55_),
    .S(net189),
    .X(_1620_));
 sg13g2_a22oi_1 _5944_ (.Y(_1621_),
    .B1(_1620_),
    .B2(net539),
    .A2(_1619_),
    .A1(net526));
 sg13g2_nand3_1 _5945_ (.B(_1616_),
    .C(_1621_),
    .A(_1615_),
    .Y(_1622_));
 sg13g2_a221oi_1 _5946_ (.B2(net487),
    .C1(_1622_),
    .B1(_1610_),
    .A1(net587),
    .Y(_1623_),
    .A2(_1609_));
 sg13g2_nor2_2 _5947_ (.A(net407),
    .B(_1623_),
    .Y(_1624_));
 sg13g2_mux2_1 _5948_ (.A0(\i_dm_csrs.i_fifo.mem_q_25_ ),
    .A1(_1624_),
    .S(net492),
    .X(_0127_));
 sg13g2_mux4_1 _5949_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_24_ ),
    .A1(\i_dm_csrs.progbuf_o_88_ ),
    .A2(\i_dm_csrs.progbuf_o_56_ ),
    .A3(\i_dm_csrs.progbuf_o_120_ ),
    .S1(net196),
    .X(_1625_));
 sg13g2_mux4_1 _5950_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_152_ ),
    .A1(\i_dm_csrs.progbuf_o_216_ ),
    .A2(\i_dm_csrs.progbuf_o_184_ ),
    .A3(\i_dm_csrs.progbuf_o_248_ ),
    .S1(net197),
    .X(_1626_));
 sg13g2_mux2_2 _5951_ (.A0(_1625_),
    .A1(_1626_),
    .S(net137),
    .X(_1627_));
 sg13g2_mux2_1 _5952_ (.A0(\i_dm_csrs.sbdata_o_24_ ),
    .A1(\i_dm_csrs.sbdata_q_56_ ),
    .S(net175),
    .X(_1628_));
 sg13g2_buf_8 fanout259 (.A(net261),
    .X(net259));
 sg13g2_and2_1 _5954_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_56_ ),
    .X(_1630_));
 sg13g2_a21oi_1 _5955_ (.A1(net606),
    .A2(\i_dm_csrs.sbcs_q_24_ ),
    .Y(_1631_),
    .B1(_1630_));
 sg13g2_nand3_1 _5956_ (.B(net604),
    .C(master_add_o_24_),
    .A(net186),
    .Y(_1632_));
 sg13g2_o21ai_1 _5957_ (.B1(_1632_),
    .Y(_1633_),
    .A1(net174),
    .A2(_1631_));
 sg13g2_nand2_1 _5958_ (.Y(_1634_),
    .A(_1355_),
    .B(_1633_));
 sg13g2_nand2_1 _5959_ (.Y(_1635_),
    .A(hartinfo_i_24_),
    .B(net529));
 sg13g2_mux2_1 _5960_ (.A0(data_csrs_mem_24_),
    .A1(data_csrs_mem_56_),
    .S(net176),
    .X(_1636_));
 sg13g2_a22oi_1 _5961_ (.Y(_1637_),
    .B1(_1636_),
    .B2(net537),
    .A2(net535),
    .A1(next_dm_addr_i_24_));
 sg13g2_nand3_1 _5962_ (.B(_1635_),
    .C(_1637_),
    .A(_1634_),
    .Y(_1638_));
 sg13g2_a221oi_1 _5963_ (.B2(net486),
    .C1(_1638_),
    .B1(_1628_),
    .A1(net586),
    .Y(_1639_),
    .A2(_1627_));
 sg13g2_nor2_2 _5964_ (.A(net408),
    .B(_1639_),
    .Y(_1640_));
 sg13g2_mux2_1 _5965_ (.A0(\i_dm_csrs.i_fifo.mem_q_26_ ),
    .A1(_1640_),
    .S(net491),
    .X(_0128_));
 sg13g2_mux4_1 _5966_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_25_ ),
    .A1(\i_dm_csrs.progbuf_o_89_ ),
    .A2(\i_dm_csrs.progbuf_o_57_ ),
    .A3(\i_dm_csrs.progbuf_o_121_ ),
    .S1(net196),
    .X(_1641_));
 sg13g2_mux4_1 _5967_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_153_ ),
    .A1(\i_dm_csrs.progbuf_o_217_ ),
    .A2(\i_dm_csrs.progbuf_o_185_ ),
    .A3(\i_dm_csrs.progbuf_o_249_ ),
    .S1(net193),
    .X(_1642_));
 sg13g2_mux2_2 _5968_ (.A0(_1641_),
    .A1(_1642_),
    .S(net138),
    .X(_1643_));
 sg13g2_mux2_1 _5969_ (.A0(\i_dm_csrs.sbdata_o_25_ ),
    .A1(\i_dm_csrs.sbdata_q_57_ ),
    .S(net175),
    .X(_1644_));
 sg13g2_and2_1 _5970_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_57_ ),
    .X(_1645_));
 sg13g2_a21oi_1 _5971_ (.A1(net606),
    .A2(\i_dm_csrs.sbcs_q_25_ ),
    .Y(_1646_),
    .B1(_1645_));
 sg13g2_nand3_1 _5972_ (.B(net604),
    .C(master_add_o_25_),
    .A(net186),
    .Y(_1647_));
 sg13g2_o21ai_1 _5973_ (.B1(_1647_),
    .Y(_1648_),
    .A1(net174),
    .A2(_1646_));
 sg13g2_nand2_1 _5974_ (.Y(_1649_),
    .A(_1355_),
    .B(_1648_));
 sg13g2_nand2_1 _5975_ (.Y(_1650_),
    .A(hartinfo_i_25_),
    .B(net529));
 sg13g2_mux2_1 _5976_ (.A0(data_csrs_mem_25_),
    .A1(data_csrs_mem_57_),
    .S(net176),
    .X(_1651_));
 sg13g2_a22oi_1 _5977_ (.Y(_1652_),
    .B1(_1651_),
    .B2(net537),
    .A2(net535),
    .A1(next_dm_addr_i_25_));
 sg13g2_nand3_1 _5978_ (.B(_1650_),
    .C(_1652_),
    .A(_1649_),
    .Y(_1653_));
 sg13g2_a221oi_1 _5979_ (.B2(net486),
    .C1(_1653_),
    .B1(_1644_),
    .A1(net586),
    .Y(_1654_),
    .A2(_1643_));
 sg13g2_nor2_2 _5980_ (.A(net407),
    .B(_1654_),
    .Y(_1655_));
 sg13g2_buf_16 fanout258 (.X(net258),
    .A(net261));
 sg13g2_mux2_1 _5982_ (.A0(\i_dm_csrs.i_fifo.mem_q_27_ ),
    .A1(_1655_),
    .S(net491),
    .X(_0129_));
 sg13g2_mux4_1 _5983_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_26_ ),
    .A1(\i_dm_csrs.progbuf_o_90_ ),
    .A2(\i_dm_csrs.progbuf_o_58_ ),
    .A3(\i_dm_csrs.progbuf_o_122_ ),
    .S1(net196),
    .X(_1657_));
 sg13g2_mux4_1 _5984_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_154_ ),
    .A1(\i_dm_csrs.progbuf_o_218_ ),
    .A2(\i_dm_csrs.progbuf_o_186_ ),
    .A3(\i_dm_csrs.progbuf_o_250_ ),
    .S1(net193),
    .X(_1658_));
 sg13g2_mux2_2 _5985_ (.A0(_1657_),
    .A1(_1658_),
    .S(net138),
    .X(_1659_));
 sg13g2_mux2_1 _5986_ (.A0(\i_dm_csrs.sbdata_o_26_ ),
    .A1(\i_dm_csrs.sbdata_q_58_ ),
    .S(net175),
    .X(_1660_));
 sg13g2_and2_1 _5987_ (.A(net143),
    .B(\i_dm_csrs.sbaddr_q_58_ ),
    .X(_1661_));
 sg13g2_a21oi_1 _5988_ (.A1(net606),
    .A2(\i_dm_csrs.sbcs_q_26_ ),
    .Y(_1662_),
    .B1(_1661_));
 sg13g2_nand3_1 _5989_ (.B(net604),
    .C(master_add_o_26_),
    .A(net186),
    .Y(_1663_));
 sg13g2_o21ai_1 _5990_ (.B1(_1663_),
    .Y(_1664_),
    .A1(net173),
    .A2(_1662_));
 sg13g2_nand2_2 _5991_ (.Y(_1665_),
    .A(net532),
    .B(_1664_));
 sg13g2_nand2_1 _5992_ (.Y(_1666_),
    .A(hartinfo_i_26_),
    .B(net528));
 sg13g2_mux2_1 _5993_ (.A0(data_csrs_mem_26_),
    .A1(data_csrs_mem_58_),
    .S(net176),
    .X(_1667_));
 sg13g2_a22oi_1 _5994_ (.Y(_1668_),
    .B1(_1667_),
    .B2(net536),
    .A2(net534),
    .A1(next_dm_addr_i_26_));
 sg13g2_nand3_1 _5995_ (.B(_1666_),
    .C(_1668_),
    .A(_1665_),
    .Y(_1669_));
 sg13g2_a221oi_1 _5996_ (.B2(net484),
    .C1(_1669_),
    .B1(_1660_),
    .A1(net583),
    .Y(_1670_),
    .A2(_1659_));
 sg13g2_nor2_2 _5997_ (.A(net406),
    .B(_1670_),
    .Y(_1671_));
 sg13g2_mux2_1 _5998_ (.A0(\i_dm_csrs.i_fifo.mem_q_28_ ),
    .A1(_1671_),
    .S(net490),
    .X(_0130_));
 sg13g2_mux2_1 _5999_ (.A0(\i_dm_csrs.sbdata_o_27_ ),
    .A1(\i_dm_csrs.sbdata_q_59_ ),
    .S(net169),
    .X(_1672_));
 sg13g2_mux2_1 _6000_ (.A0(\i_dm_csrs.sbcs_q_27_ ),
    .A1(\i_dm_csrs.sbaddr_q_59_ ),
    .S(net144),
    .X(_1673_));
 sg13g2_nand2_1 _6001_ (.Y(_1674_),
    .A(net591),
    .B(_1673_));
 sg13g2_nand3_1 _6002_ (.B(net605),
    .C(master_add_o_27_),
    .A(net182),
    .Y(_1675_));
 sg13g2_a21oi_1 _6003_ (.A1(_1674_),
    .A2(_1675_),
    .Y(_1676_),
    .B1(net138));
 sg13g2_a21o_1 _6004_ (.A2(_1672_),
    .A1(_1316_),
    .B1(_1676_),
    .X(_1677_));
 sg13g2_mux4_1 _6005_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_27_ ),
    .A1(\i_dm_csrs.progbuf_o_91_ ),
    .A2(\i_dm_csrs.progbuf_o_59_ ),
    .A3(\i_dm_csrs.progbuf_o_123_ ),
    .S1(net199),
    .X(_1678_));
 sg13g2_mux4_1 _6006_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_155_ ),
    .A1(\i_dm_csrs.progbuf_o_219_ ),
    .A2(\i_dm_csrs.progbuf_o_187_ ),
    .A3(\i_dm_csrs.progbuf_o_251_ ),
    .S1(net195),
    .X(_1679_));
 sg13g2_mux2_1 _6007_ (.A0(_1678_),
    .A1(_1679_),
    .S(net135),
    .X(_1680_));
 sg13g2_nand2_1 _6008_ (.Y(_1681_),
    .A(next_dm_addr_i_27_),
    .B(net580));
 sg13g2_nor2_1 _6009_ (.A(_1146_),
    .B(_1681_),
    .Y(_1682_));
 sg13g2_o21ai_1 _6010_ (.B1(net142),
    .Y(_1683_),
    .A1(_1211_),
    .A2(_1682_));
 sg13g2_mux2_1 _6011_ (.A0(data_csrs_mem_27_),
    .A1(data_csrs_mem_59_),
    .S(net162),
    .X(_1684_));
 sg13g2_a22oi_1 _6012_ (.Y(_1685_),
    .B1(_1684_),
    .B2(net536),
    .A2(net528),
    .A1(hartinfo_i_27_));
 sg13g2_nand2_1 _6013_ (.Y(_1686_),
    .A(_1683_),
    .B(_1685_));
 sg13g2_a221oi_1 _6014_ (.B2(net583),
    .C1(_1686_),
    .B1(_1680_),
    .A1(net43),
    .Y(_1687_),
    .A2(_1677_));
 sg13g2_nor2_1 _6015_ (.A(net409),
    .B(_1687_),
    .Y(_1688_));
 sg13g2_mux2_1 _6016_ (.A0(\i_dm_csrs.i_fifo.mem_q_29_ ),
    .A1(_1688_),
    .S(net490),
    .X(_0131_));
 sg13g2_mux2_1 _6017_ (.A0(\i_dm_csrs.sbdata_o_0_ ),
    .A1(\i_dm_csrs.sbdata_q_32_ ),
    .S(net172),
    .X(_1689_));
 sg13g2_nand2_1 _6018_ (.Y(_1690_),
    .A(\i_dm_csrs.abstractauto_q_0_ ),
    .B(_1271_));
 sg13g2_nand3_1 _6019_ (.B(net135),
    .C(next_dm_addr_i_0_),
    .A(net178),
    .Y(_1691_));
 sg13g2_nand2_1 _6020_ (.Y(_1692_),
    .A(_1690_),
    .B(_1691_));
 sg13g2_a21oi_1 _6021_ (.A1(net156),
    .A2(\i_dm_csrs.sbaddr_q_32_ ),
    .Y(_1693_),
    .B1(_1358_));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_2094_));
 sg13g2_nand3_1 _6023_ (.B(net602),
    .C(net51),
    .A(net184),
    .Y(_1695_));
 sg13g2_o21ai_1 _6024_ (.B1(_1695_),
    .Y(_1696_),
    .A1(net162),
    .A2(_1693_));
 sg13g2_a22oi_1 _6025_ (.Y(_1697_),
    .B1(_1696_),
    .B2(net531),
    .A2(_1692_),
    .A1(_1480_));
 sg13g2_inv_1 _6026_ (.Y(_1698_),
    .A(_1697_));
 sg13g2_a221oi_1 _6027_ (.B2(_1689_),
    .C1(_1698_),
    .B1(net485),
    .A1(halted),
    .Y(_1699_),
    .A2(_1274_));
 sg13g2_mux4_1 _6028_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_0_ ),
    .A1(\i_dm_csrs.progbuf_o_64_ ),
    .A2(\i_dm_csrs.progbuf_o_32_ ),
    .A3(\i_dm_csrs.progbuf_o_96_ ),
    .S1(net195),
    .X(_1700_));
 sg13g2_mux4_1 _6029_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_128_ ),
    .A1(\i_dm_csrs.progbuf_o_192_ ),
    .A2(\i_dm_csrs.progbuf_o_160_ ),
    .A3(\i_dm_csrs.progbuf_o_224_ ),
    .S1(net194),
    .X(_1701_));
 sg13g2_mux2_1 _6030_ (.A0(_1700_),
    .A1(_1701_),
    .S(net136),
    .X(_1702_));
 sg13g2_inv_1 _6031_ (.Y(_1703_),
    .A(halted));
 sg13g2_nor2_1 _6032_ (.A(_1703_),
    .B(net600),
    .Y(_1704_));
 sg13g2_a22oi_1 _6033_ (.Y(_1705_),
    .B1(_1704_),
    .B2(_0596_),
    .A2(net538),
    .A1(data_csrs_mem_32_));
 sg13g2_nand2_2 _6034_ (.Y(_1706_),
    .A(hartinfo_i_0_),
    .B(net149));
 sg13g2_o21ai_1 _6035_ (.B1(_1706_),
    .Y(_1707_),
    .A1(net597),
    .A2(net146));
 sg13g2_a221oi_1 _6036_ (.B2(_0596_),
    .C1(net163),
    .B1(_1707_),
    .A1(data_csrs_mem_0_),
    .Y(_1708_),
    .A2(net538));
 sg13g2_a21oi_1 _6037_ (.A1(net179),
    .A2(_1705_),
    .Y(_1709_),
    .B1(_1708_));
 sg13g2_a21oi_1 _6038_ (.A1(net583),
    .A2(_1702_),
    .Y(_1710_),
    .B1(_1709_));
 sg13g2_a21oi_2 _6039_ (.B1(net405),
    .Y(_1711_),
    .A2(_1710_),
    .A1(_1699_));
 sg13g2_mux2_1 _6040_ (.A0(\i_dm_csrs.i_fifo.mem_q_2_ ),
    .A1(_1711_),
    .S(net492),
    .X(_0132_));
 sg13g2_mux4_1 _6041_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_28_ ),
    .A1(\i_dm_csrs.progbuf_o_92_ ),
    .A2(\i_dm_csrs.progbuf_o_60_ ),
    .A3(\i_dm_csrs.progbuf_o_124_ ),
    .S1(net196),
    .X(_1712_));
 sg13g2_mux4_1 _6042_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_156_ ),
    .A1(\i_dm_csrs.progbuf_o_220_ ),
    .A2(\i_dm_csrs.progbuf_o_188_ ),
    .A3(\i_dm_csrs.progbuf_o_252_ ),
    .S1(net193),
    .X(_1713_));
 sg13g2_mux2_2 _6043_ (.A0(_1712_),
    .A1(_1713_),
    .S(net138),
    .X(_1714_));
 sg13g2_mux2_1 _6044_ (.A0(\i_dm_csrs.sbdata_o_28_ ),
    .A1(\i_dm_csrs.sbdata_q_60_ ),
    .S(net175),
    .X(_1715_));
 sg13g2_and2_1 _6045_ (.A(net144),
    .B(\i_dm_csrs.sbaddr_q_60_ ),
    .X(_1716_));
 sg13g2_a21oi_1 _6046_ (.A1(net604),
    .A2(\i_dm_csrs.sbcs_q_28_ ),
    .Y(_1717_),
    .B1(_1716_));
 sg13g2_nand3_1 _6047_ (.B(net604),
    .C(master_add_o_28_),
    .A(net186),
    .Y(_1718_));
 sg13g2_o21ai_1 _6048_ (.B1(_1718_),
    .Y(_1719_),
    .A1(net173),
    .A2(_1717_));
 sg13g2_nand2_1 _6049_ (.Y(_1720_),
    .A(net532),
    .B(_1719_));
 sg13g2_nand2_1 _6050_ (.Y(_1721_),
    .A(hartinfo_i_28_),
    .B(net529));
 sg13g2_mux2_1 _6051_ (.A0(data_csrs_mem_28_),
    .A1(data_csrs_mem_60_),
    .S(net176),
    .X(_1722_));
 sg13g2_a22oi_1 _6052_ (.Y(_1723_),
    .B1(_1722_),
    .B2(net536),
    .A2(net534),
    .A1(next_dm_addr_i_28_));
 sg13g2_nand3_1 _6053_ (.B(_1721_),
    .C(_1723_),
    .A(_1720_),
    .Y(_1724_));
 sg13g2_a221oi_1 _6054_ (.B2(net486),
    .C1(_1724_),
    .B1(_1715_),
    .A1(net587),
    .Y(_1725_),
    .A2(_1714_));
 sg13g2_nor2_2 _6055_ (.A(net407),
    .B(_1725_),
    .Y(_1726_));
 sg13g2_mux2_1 _6056_ (.A0(\i_dm_csrs.i_fifo.mem_q_30_ ),
    .A1(_1726_),
    .S(net492),
    .X(_0133_));
 sg13g2_mux4_1 _6057_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_29_ ),
    .A1(\i_dm_csrs.progbuf_o_93_ ),
    .A2(\i_dm_csrs.progbuf_o_61_ ),
    .A3(\i_dm_csrs.progbuf_o_125_ ),
    .S1(net197),
    .X(_1727_));
 sg13g2_mux4_1 _6058_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_157_ ),
    .A1(\i_dm_csrs.progbuf_o_221_ ),
    .A2(\i_dm_csrs.progbuf_o_189_ ),
    .A3(\i_dm_csrs.progbuf_o_253_ ),
    .S1(net192),
    .X(_1728_));
 sg13g2_mux2_2 _6059_ (.A0(_1727_),
    .A1(_1728_),
    .S(net138),
    .X(_1729_));
 sg13g2_mux2_1 _6060_ (.A0(\i_dm_csrs.sbdata_o_29_ ),
    .A1(\i_dm_csrs.sbdata_q_61_ ),
    .S(net175),
    .X(_1730_));
 sg13g2_a21oi_1 _6061_ (.A1(net157),
    .A2(\i_dm_csrs.sbaddr_q_61_ ),
    .Y(_1731_),
    .B1(_1358_));
 sg13g2_nand3_1 _6062_ (.B(net602),
    .C(master_add_o_29_),
    .A(net185),
    .Y(_1732_));
 sg13g2_o21ai_1 _6063_ (.B1(_1732_),
    .Y(_1733_),
    .A1(net173),
    .A2(_1731_));
 sg13g2_nand2_2 _6064_ (.Y(_1734_),
    .A(net532),
    .B(_1733_));
 sg13g2_nand2_1 _6065_ (.Y(_1735_),
    .A(hartinfo_i_29_),
    .B(net529));
 sg13g2_mux2_1 _6066_ (.A0(data_csrs_mem_29_),
    .A1(data_csrs_mem_61_),
    .S(net176),
    .X(_1736_));
 sg13g2_a22oi_1 _6067_ (.Y(_1737_),
    .B1(_1736_),
    .B2(net537),
    .A2(net535),
    .A1(next_dm_addr_i_29_));
 sg13g2_nand3_1 _6068_ (.B(_1735_),
    .C(_1737_),
    .A(_1734_),
    .Y(_1738_));
 sg13g2_a221oi_1 _6069_ (.B2(net483),
    .C1(_1738_),
    .B1(_1730_),
    .A1(net582),
    .Y(_1739_),
    .A2(_1729_));
 sg13g2_nor2_2 _6070_ (.A(net406),
    .B(_1739_),
    .Y(_1740_));
 sg13g2_mux2_1 _6071_ (.A0(\i_dm_csrs.i_fifo.mem_q_31_ ),
    .A1(_1740_),
    .S(net488),
    .X(_0134_));
 sg13g2_mux2_1 _6072_ (.A0(\i_dm_csrs.sbdata_o_30_ ),
    .A1(\i_dm_csrs.sbdata_q_62_ ),
    .S(net170),
    .X(_1741_));
 sg13g2_mux4_1 _6073_ (.S0(net154),
    .A0(\i_dm_csrs.progbuf_o_30_ ),
    .A1(\i_dm_csrs.progbuf_o_94_ ),
    .A2(\i_dm_csrs.progbuf_o_62_ ),
    .A3(\i_dm_csrs.progbuf_o_126_ ),
    .S1(net198),
    .X(_1742_));
 sg13g2_mux4_1 _6074_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_158_ ),
    .A1(\i_dm_csrs.progbuf_o_222_ ),
    .A2(\i_dm_csrs.progbuf_o_190_ ),
    .A3(\i_dm_csrs.progbuf_o_254_ ),
    .S1(net194),
    .X(_1743_));
 sg13g2_mux2_2 _6075_ (.A0(_1742_),
    .A1(_1743_),
    .S(net135),
    .X(_1744_));
 sg13g2_inv_2 _6076_ (.Y(_1745_),
    .A(\i_dm_csrs.resumereq_o ));
 sg13g2_nand2_1 _6077_ (.Y(_1746_),
    .A(net155),
    .B(hartinfo_i_30_));
 sg13g2_o21ai_1 _6078_ (.B1(_1746_),
    .Y(_1747_),
    .A1(_1745_),
    .A2(net147));
 sg13g2_nor2b_1 _6079_ (.A(_0618_),
    .B_N(_1271_),
    .Y(_1748_));
 sg13g2_a22oi_1 _6080_ (.Y(_1749_),
    .B1(_1747_),
    .B2(_1748_),
    .A2(net533),
    .A1(next_dm_addr_i_30_));
 sg13g2_nand2_1 _6081_ (.Y(_1750_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_62_ ));
 sg13g2_nand3_1 _6082_ (.B(net606),
    .C(master_add_o_30_),
    .A(net178),
    .Y(_1751_));
 sg13g2_o21ai_1 _6083_ (.B1(_1751_),
    .Y(_1752_),
    .A1(net173),
    .A2(_1750_));
 sg13g2_mux2_2 _6084_ (.A0(data_csrs_mem_30_),
    .A1(data_csrs_mem_62_),
    .S(net162),
    .X(_1753_));
 sg13g2_a22oi_1 _6085_ (.Y(_1754_),
    .B1(_1753_),
    .B2(net539),
    .A2(_1752_),
    .A1(net530));
 sg13g2_nand2_1 _6086_ (.Y(_1755_),
    .A(_1749_),
    .B(_1754_));
 sg13g2_a221oi_1 _6087_ (.B2(net583),
    .C1(_1755_),
    .B1(_1744_),
    .A1(net485),
    .Y(_1756_),
    .A2(_1741_));
 sg13g2_nor2_2 _6088_ (.A(net406),
    .B(_1756_),
    .Y(_1757_));
 sg13g2_mux2_1 _6089_ (.A0(\i_dm_csrs.i_fifo.mem_q_32_ ),
    .A1(_1757_),
    .S(net488),
    .X(_0135_));
 sg13g2_mux2_1 _6090_ (.A0(\i_dm_csrs.sbdata_o_31_ ),
    .A1(\i_dm_csrs.sbdata_q_63_ ),
    .S(net170),
    .X(_1758_));
 sg13g2_mux4_1 _6091_ (.S0(net153),
    .A0(\i_dm_csrs.progbuf_o_31_ ),
    .A1(\i_dm_csrs.progbuf_o_95_ ),
    .A2(\i_dm_csrs.progbuf_o_63_ ),
    .A3(\i_dm_csrs.progbuf_o_127_ ),
    .S1(net198),
    .X(_1759_));
 sg13g2_mux4_1 _6092_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_159_ ),
    .A1(\i_dm_csrs.progbuf_o_223_ ),
    .A2(\i_dm_csrs.progbuf_o_191_ ),
    .A3(\i_dm_csrs.progbuf_o_255_ ),
    .S1(net194),
    .X(_1760_));
 sg13g2_mux2_2 _6093_ (.A0(_1759_),
    .A1(_1760_),
    .S(net136),
    .X(_1761_));
 sg13g2_mux2_1 _6094_ (.A0(debug_req_o),
    .A1(hartinfo_i_31_),
    .S(net146),
    .X(_1762_));
 sg13g2_a22oi_1 _6095_ (.Y(_1763_),
    .B1(_1748_),
    .B2(_1762_),
    .A2(net534),
    .A1(next_dm_addr_i_31_));
 sg13g2_nand2_1 _6096_ (.Y(_1764_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_63_ ));
 sg13g2_nand3_1 _6097_ (.B(net603),
    .C(master_add_o_31_),
    .A(net178),
    .Y(_1765_));
 sg13g2_o21ai_1 _6098_ (.B1(_1765_),
    .Y(_1766_),
    .A1(net173),
    .A2(_1764_));
 sg13g2_mux2_1 _6099_ (.A0(data_csrs_mem_31_),
    .A1(data_csrs_mem_63_),
    .S(net163),
    .X(_1767_));
 sg13g2_a22oi_1 _6100_ (.Y(_1768_),
    .B1(_1767_),
    .B2(net538),
    .A2(_1766_),
    .A1(net531));
 sg13g2_nand2_1 _6101_ (.Y(_1769_),
    .A(_1763_),
    .B(_1768_));
 sg13g2_a221oi_1 _6102_ (.B2(net586),
    .C1(_1769_),
    .B1(_1761_),
    .A1(net485),
    .Y(_1770_),
    .A2(_1758_));
 sg13g2_nor2_2 _6103_ (.A(net408),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_mux2_1 _6104_ (.A0(\i_dm_csrs.i_fifo.mem_q_33_ ),
    .A1(_1771_),
    .S(net490),
    .X(_0136_));
 sg13g2_and2_1 _6105_ (.A(\i_dm_csrs.i_fifo.write_pointer_q ),
    .B(net44),
    .X(_1772_));
 sg13g2_buf_16 fanout256 (.X(net256),
    .A(net257));
 sg13g2_buf_16 fanout255 (.X(net255),
    .A(net256));
 sg13g2_mux2_1 _6108_ (.A0(\i_dm_csrs.i_fifo.mem_q_34_ ),
    .A1(_1291_),
    .S(net479),
    .X(_0137_));
 sg13g2_mux2_1 _6109_ (.A0(\i_dm_csrs.i_fifo.mem_q_35_ ),
    .A1(_1291_),
    .S(net479),
    .X(_0138_));
 sg13g2_mux2_1 _6110_ (.A0(\i_dm_csrs.i_fifo.mem_q_36_ ),
    .A1(_1711_),
    .S(net482),
    .X(_0139_));
 sg13g2_mux4_1 _6111_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_1_ ),
    .A1(\i_dm_csrs.progbuf_o_65_ ),
    .A2(\i_dm_csrs.progbuf_o_33_ ),
    .A3(\i_dm_csrs.progbuf_o_97_ ),
    .S1(net192),
    .X(_1775_));
 sg13g2_mux4_1 _6112_ (.S0(net151),
    .A0(\i_dm_csrs.progbuf_o_129_ ),
    .A1(\i_dm_csrs.progbuf_o_193_ ),
    .A2(\i_dm_csrs.progbuf_o_161_ ),
    .A3(\i_dm_csrs.progbuf_o_225_ ),
    .S1(net195),
    .X(_1776_));
 sg13g2_mux2_2 _6113_ (.A0(_1775_),
    .A1(_1776_),
    .S(net139),
    .X(_1777_));
 sg13g2_nand2_1 _6114_ (.Y(_1778_),
    .A(net584),
    .B(_1777_));
 sg13g2_a21oi_1 _6115_ (.A1(net156),
    .A2(\i_dm_csrs.sbaddr_q_33_ ),
    .Y(_1779_),
    .B1(_1358_));
 sg13g2_buf_4 fanout254 (.X(net254),
    .A(_2094_));
 sg13g2_nand3_1 _6117_ (.B(net602),
    .C(master_add_o_1_),
    .A(net185),
    .Y(_1781_));
 sg13g2_o21ai_1 _6118_ (.B1(_1781_),
    .Y(_1782_),
    .A1(net163),
    .A2(_1779_));
 sg13g2_mux2_1 _6119_ (.A0(\i_dm_csrs.sbdata_o_1_ ),
    .A1(\i_dm_csrs.sbdata_q_33_ ),
    .S(net170),
    .X(_1783_));
 sg13g2_mux2_1 _6120_ (.A0(data_csrs_mem_1_),
    .A1(data_csrs_mem_33_),
    .S(net169),
    .X(_1784_));
 sg13g2_nand2_1 _6121_ (.Y(_1785_),
    .A(net538),
    .B(_1784_));
 sg13g2_nand3_1 _6122_ (.B(net139),
    .C(next_dm_addr_i_1_),
    .A(net183),
    .Y(_1786_));
 sg13g2_nand3_1 _6123_ (.B(\i_dm_csrs.abstractauto_q_1_ ),
    .C(net45),
    .A(net590),
    .Y(_1787_));
 sg13g2_nand2_1 _6124_ (.Y(_1788_),
    .A(_1786_),
    .B(_1787_));
 sg13g2_o21ai_1 _6125_ (.B1(net600),
    .Y(_1789_),
    .A1(ndmreset_o),
    .A2(net169));
 sg13g2_nand2_1 _6126_ (.Y(_1790_),
    .A(hartinfo_i_1_),
    .B(net548));
 sg13g2_nand2_1 _6127_ (.Y(_1791_),
    .A(_1789_),
    .B(_1790_));
 sg13g2_a22oi_1 _6128_ (.Y(_1792_),
    .B1(_1791_),
    .B2(_0596_),
    .A2(_1788_),
    .A1(_1480_));
 sg13g2_nand3_1 _6129_ (.B(_1785_),
    .C(_1792_),
    .A(_1212_),
    .Y(_1793_));
 sg13g2_a221oi_1 _6130_ (.B2(net485),
    .C1(_1793_),
    .B1(_1783_),
    .A1(net531),
    .Y(_1794_),
    .A2(_1782_));
 sg13g2_a21oi_2 _6131_ (.B1(net410),
    .Y(_1795_),
    .A2(_1794_),
    .A1(_1778_));
 sg13g2_mux2_1 _6132_ (.A0(\i_dm_csrs.i_fifo.mem_q_37_ ),
    .A1(_1795_),
    .S(net482),
    .X(_0140_));
 sg13g2_mux4_1 _6133_ (.S0(net152),
    .A0(\i_dm_csrs.progbuf_o_2_ ),
    .A1(\i_dm_csrs.progbuf_o_66_ ),
    .A2(\i_dm_csrs.progbuf_o_34_ ),
    .A3(\i_dm_csrs.progbuf_o_98_ ),
    .S1(net197),
    .X(_1796_));
 sg13g2_mux4_1 _6134_ (.S0(net145),
    .A0(\i_dm_csrs.progbuf_o_130_ ),
    .A1(\i_dm_csrs.progbuf_o_194_ ),
    .A2(\i_dm_csrs.progbuf_o_162_ ),
    .A3(\i_dm_csrs.progbuf_o_226_ ),
    .S1(net192),
    .X(_1797_));
 sg13g2_mux2_2 _6135_ (.A0(_1796_),
    .A1(_1797_),
    .S(net138),
    .X(_1798_));
 sg13g2_mux2_1 _6136_ (.A0(\i_dm_csrs.sbdata_o_2_ ),
    .A1(\i_dm_csrs.sbdata_q_34_ ),
    .S(net174),
    .X(_1799_));
 sg13g2_a21oi_1 _6137_ (.A1(net157),
    .A2(\i_dm_csrs.sbaddr_q_34_ ),
    .Y(_1800_),
    .B1(_1358_));
 sg13g2_buf_8 fanout253 (.A(net254),
    .X(net253));
 sg13g2_nand3_1 _6139_ (.B(net602),
    .C(net50),
    .A(net185),
    .Y(_1802_));
 sg13g2_o21ai_1 _6140_ (.B1(_1802_),
    .Y(_1803_),
    .A1(net173),
    .A2(_1800_));
 sg13g2_nand2_1 _6141_ (.Y(_1804_),
    .A(net530),
    .B(_1803_));
 sg13g2_nand2_1 _6142_ (.Y(_1805_),
    .A(hartinfo_i_2_),
    .B(net527));
 sg13g2_mux2_1 _6143_ (.A0(data_csrs_mem_2_),
    .A1(data_csrs_mem_34_),
    .S(net176),
    .X(_1806_));
 sg13g2_a22oi_1 _6144_ (.Y(_1807_),
    .B1(_1806_),
    .B2(net537),
    .A2(net535),
    .A1(next_dm_addr_i_2_));
 sg13g2_nand3_1 _6145_ (.B(_1805_),
    .C(_1807_),
    .A(_1804_),
    .Y(_1808_));
 sg13g2_a221oi_1 _6146_ (.B2(net486),
    .C1(_1808_),
    .B1(_1799_),
    .A1(net586),
    .Y(_1809_),
    .A2(_1798_));
 sg13g2_nor2_2 _6147_ (.A(net407),
    .B(_1809_),
    .Y(_1810_));
 sg13g2_mux2_1 _6148_ (.A0(\i_dm_csrs.i_fifo.mem_q_38_ ),
    .A1(_1810_),
    .S(net481),
    .X(_0141_));
 sg13g2_mux4_1 _6149_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_131_ ),
    .A1(\i_dm_csrs.progbuf_o_195_ ),
    .A2(\i_dm_csrs.progbuf_o_163_ ),
    .A3(\i_dm_csrs.progbuf_o_227_ ),
    .S1(net192),
    .X(_1811_));
 sg13g2_mux4_1 _6150_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_3_ ),
    .A1(\i_dm_csrs.progbuf_o_67_ ),
    .A2(\i_dm_csrs.progbuf_o_35_ ),
    .A3(\i_dm_csrs.progbuf_o_99_ ),
    .S1(net195),
    .X(_1812_));
 sg13g2_mux2_1 _6151_ (.A0(_1811_),
    .A1(_1812_),
    .S(net45),
    .X(_1813_));
 sg13g2_nand2_1 _6152_ (.Y(_1814_),
    .A(net582),
    .B(_1813_));
 sg13g2_mux2_1 _6153_ (.A0(\i_dm_csrs.sbdata_o_3_ ),
    .A1(\i_dm_csrs.sbdata_q_35_ ),
    .S(net170),
    .X(_1815_));
 sg13g2_and2_1 _6154_ (.A(data_csrs_mem_35_),
    .B(net163),
    .X(_1816_));
 sg13g2_a21oi_1 _6155_ (.A1(data_csrs_mem_3_),
    .A2(net591),
    .Y(_1817_),
    .B1(_1816_));
 sg13g2_nand2_1 _6156_ (.Y(_1818_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_35_ ));
 sg13g2_buf_16 fanout252 (.X(net252),
    .A(net254));
 sg13g2_nand3_1 _6158_ (.B(net602),
    .C(master_add_o_3_),
    .A(net184),
    .Y(_1820_));
 sg13g2_o21ai_1 _6159_ (.B1(_1820_),
    .Y(_1821_),
    .A1(net166),
    .A2(_1818_));
 sg13g2_a22oi_1 _6160_ (.Y(_1822_),
    .B1(net530),
    .B2(_1821_),
    .A2(net533),
    .A1(next_dm_addr_i_3_));
 sg13g2_o21ai_1 _6161_ (.B1(_1822_),
    .Y(_1823_),
    .A1(_0731_),
    .A2(_1817_));
 sg13g2_a221oi_1 _6162_ (.B2(net483),
    .C1(_1823_),
    .B1(_1815_),
    .A1(hartinfo_i_3_),
    .Y(_1824_),
    .A2(net527));
 sg13g2_a21oi_2 _6163_ (.B1(net405),
    .Y(_1825_),
    .A2(_1824_),
    .A1(_1814_));
 sg13g2_mux2_1 _6164_ (.A0(\i_dm_csrs.i_fifo.mem_q_39_ ),
    .A1(_1825_),
    .S(net478),
    .X(_0142_));
 sg13g2_mux2_1 _6165_ (.A0(\i_dm_csrs.i_fifo.mem_q_3_ ),
    .A1(_1795_),
    .S(net492),
    .X(_0143_));
 sg13g2_mux4_1 _6166_ (.S0(net149),
    .A0(\i_dm_csrs.progbuf_o_132_ ),
    .A1(\i_dm_csrs.progbuf_o_196_ ),
    .A2(\i_dm_csrs.progbuf_o_164_ ),
    .A3(\i_dm_csrs.progbuf_o_228_ ),
    .S1(net195),
    .X(_1826_));
 sg13g2_mux4_1 _6167_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_4_ ),
    .A1(\i_dm_csrs.progbuf_o_68_ ),
    .A2(\i_dm_csrs.progbuf_o_36_ ),
    .A3(\i_dm_csrs.progbuf_o_100_ ),
    .S1(net193),
    .X(_1827_));
 sg13g2_mux2_2 _6168_ (.A0(_1826_),
    .A1(_1827_),
    .S(net45),
    .X(_1828_));
 sg13g2_nand2_1 _6169_ (.Y(_1829_),
    .A(net582),
    .B(_1828_));
 sg13g2_mux2_1 _6170_ (.A0(\i_dm_csrs.sbdata_o_4_ ),
    .A1(\i_dm_csrs.sbdata_q_36_ ),
    .S(net172),
    .X(_1830_));
 sg13g2_and2_1 _6171_ (.A(data_csrs_mem_36_),
    .B(net163),
    .X(_1831_));
 sg13g2_a21oi_1 _6172_ (.A1(data_csrs_mem_4_),
    .A2(net591),
    .Y(_1832_),
    .B1(_1831_));
 sg13g2_nand2_1 _6173_ (.Y(_1833_),
    .A(net157),
    .B(\i_dm_csrs.sbaddr_q_36_ ));
 sg13g2_buf_2 fanout251 (.A(_3225_),
    .X(net251));
 sg13g2_nand3_1 _6175_ (.B(net601),
    .C(net48),
    .A(net182),
    .Y(_1835_));
 sg13g2_o21ai_1 _6176_ (.B1(_1835_),
    .Y(_1836_),
    .A1(net166),
    .A2(_1833_));
 sg13g2_a22oi_1 _6177_ (.Y(_1837_),
    .B1(net530),
    .B2(_1836_),
    .A2(net533),
    .A1(next_dm_addr_i_4_));
 sg13g2_o21ai_1 _6178_ (.B1(_1837_),
    .Y(_1838_),
    .A1(_0731_),
    .A2(_1832_));
 sg13g2_a221oi_1 _6179_ (.B2(net483),
    .C1(_1838_),
    .B1(_1830_),
    .A1(hartinfo_i_4_),
    .Y(_1839_),
    .A2(net527));
 sg13g2_a21oi_2 _6180_ (.B1(net405),
    .Y(_1840_),
    .A2(_1839_),
    .A1(_1829_));
 sg13g2_mux2_1 _6181_ (.A0(\i_dm_csrs.i_fifo.mem_q_40_ ),
    .A1(_1840_),
    .S(net479),
    .X(_0144_));
 sg13g2_mux4_1 _6182_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_133_ ),
    .A1(\i_dm_csrs.progbuf_o_197_ ),
    .A2(\i_dm_csrs.progbuf_o_165_ ),
    .A3(\i_dm_csrs.progbuf_o_229_ ),
    .S1(net195),
    .X(_1841_));
 sg13g2_mux4_1 _6183_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_5_ ),
    .A1(\i_dm_csrs.progbuf_o_69_ ),
    .A2(\i_dm_csrs.progbuf_o_37_ ),
    .A3(\i_dm_csrs.progbuf_o_101_ ),
    .S1(net193),
    .X(_1842_));
 sg13g2_mux2_1 _6184_ (.A0(_1841_),
    .A1(_1842_),
    .S(net45),
    .X(_1843_));
 sg13g2_nand2_1 _6185_ (.Y(_1844_),
    .A(net582),
    .B(_1843_));
 sg13g2_mux2_1 _6186_ (.A0(\i_dm_csrs.sbdata_o_5_ ),
    .A1(\i_dm_csrs.sbdata_q_37_ ),
    .S(net172),
    .X(_1845_));
 sg13g2_and2_1 _6187_ (.A(data_csrs_mem_37_),
    .B(net171),
    .X(_1846_));
 sg13g2_a21oi_1 _6188_ (.A1(data_csrs_mem_5_),
    .A2(net591),
    .Y(_1847_),
    .B1(_1846_));
 sg13g2_nand2_1 _6189_ (.Y(_1848_),
    .A(net156),
    .B(\i_dm_csrs.sbaddr_q_37_ ));
 sg13g2_buf_2 fanout250 (.A(_3225_),
    .X(net250));
 sg13g2_nand3_1 _6191_ (.B(net601),
    .C(master_add_o_5_),
    .A(net182),
    .Y(_1850_));
 sg13g2_o21ai_1 _6192_ (.B1(_1850_),
    .Y(_1851_),
    .A1(net166),
    .A2(_1848_));
 sg13g2_a22oi_1 _6193_ (.Y(_1852_),
    .B1(net530),
    .B2(_1851_),
    .A2(net533),
    .A1(next_dm_addr_i_5_));
 sg13g2_o21ai_1 _6194_ (.B1(_1852_),
    .Y(_1853_),
    .A1(_0731_),
    .A2(_1847_));
 sg13g2_a221oi_1 _6195_ (.B2(net483),
    .C1(_1853_),
    .B1(_1845_),
    .A1(hartinfo_i_5_),
    .Y(_1854_),
    .A2(net527));
 sg13g2_a21oi_2 _6196_ (.B1(net405),
    .Y(_1855_),
    .A2(_1854_),
    .A1(_1844_));
 sg13g2_mux2_1 _6197_ (.A0(\i_dm_csrs.i_fifo.mem_q_41_ ),
    .A1(_1855_),
    .S(net478),
    .X(_0145_));
 sg13g2_mux4_1 _6198_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_134_ ),
    .A1(\i_dm_csrs.progbuf_o_198_ ),
    .A2(\i_dm_csrs.progbuf_o_166_ ),
    .A3(\i_dm_csrs.progbuf_o_230_ ),
    .S1(net195),
    .X(_1856_));
 sg13g2_mux4_1 _6199_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_6_ ),
    .A1(\i_dm_csrs.progbuf_o_70_ ),
    .A2(\i_dm_csrs.progbuf_o_38_ ),
    .A3(\i_dm_csrs.progbuf_o_102_ ),
    .S1(net193),
    .X(_1857_));
 sg13g2_mux2_1 _6200_ (.A0(_1856_),
    .A1(_1857_),
    .S(net45),
    .X(_1858_));
 sg13g2_nand2_1 _6201_ (.Y(_1859_),
    .A(net582),
    .B(_1858_));
 sg13g2_mux2_1 _6202_ (.A0(\i_dm_csrs.sbdata_o_6_ ),
    .A1(\i_dm_csrs.sbdata_q_38_ ),
    .S(net172),
    .X(_1860_));
 sg13g2_and2_1 _6203_ (.A(data_csrs_mem_38_),
    .B(net171),
    .X(_1861_));
 sg13g2_a21oi_1 _6204_ (.A1(data_csrs_mem_6_),
    .A2(net591),
    .Y(_1862_),
    .B1(_1861_));
 sg13g2_nand2_1 _6205_ (.Y(_1863_),
    .A(net156),
    .B(\i_dm_csrs.sbaddr_q_38_ ));
 sg13g2_nand3_1 _6206_ (.B(net601),
    .C(master_add_o_6_),
    .A(net182),
    .Y(_1864_));
 sg13g2_o21ai_1 _6207_ (.B1(_1864_),
    .Y(_1865_),
    .A1(net166),
    .A2(_1863_));
 sg13g2_a22oi_1 _6208_ (.Y(_1866_),
    .B1(net530),
    .B2(_1865_),
    .A2(net533),
    .A1(next_dm_addr_i_6_));
 sg13g2_o21ai_1 _6209_ (.B1(_1866_),
    .Y(_1867_),
    .A1(_0731_),
    .A2(_1862_));
 sg13g2_a221oi_1 _6210_ (.B2(net483),
    .C1(_1867_),
    .B1(_1860_),
    .A1(hartinfo_i_6_),
    .Y(_1868_),
    .A2(net527));
 sg13g2_a21oi_2 _6211_ (.B1(net405),
    .Y(_1869_),
    .A2(_1868_),
    .A1(_1859_));
 sg13g2_mux2_1 _6212_ (.A0(\i_dm_csrs.i_fifo.mem_q_42_ ),
    .A1(_1869_),
    .S(net478),
    .X(_0146_));
 sg13g2_mux4_1 _6213_ (.S0(net150),
    .A0(\i_dm_csrs.progbuf_o_7_ ),
    .A1(\i_dm_csrs.progbuf_o_71_ ),
    .A2(\i_dm_csrs.progbuf_o_39_ ),
    .A3(\i_dm_csrs.progbuf_o_103_ ),
    .S1(net195),
    .X(_1870_));
 sg13g2_mux4_1 _6214_ (.S0(net148),
    .A0(\i_dm_csrs.progbuf_o_135_ ),
    .A1(\i_dm_csrs.progbuf_o_199_ ),
    .A2(\i_dm_csrs.progbuf_o_167_ ),
    .A3(\i_dm_csrs.progbuf_o_231_ ),
    .S1(net193),
    .X(_1871_));
 sg13g2_mux2_1 _6215_ (.A0(_1870_),
    .A1(_1871_),
    .S(net139),
    .X(_1872_));
 sg13g2_nand2_1 _6216_ (.Y(_1873_),
    .A(net582),
    .B(_1872_));
 sg13g2_mux2_1 _6217_ (.A0(\i_dm_csrs.sbdata_o_7_ ),
    .A1(\i_dm_csrs.sbdata_q_39_ ),
    .S(net172),
    .X(_1874_));
 sg13g2_a22oi_1 _6218_ (.Y(_1875_),
    .B1(net581),
    .B2(master_add_o_7_),
    .A2(net548),
    .A1(\i_dm_csrs.sbaddr_q_39_ ));
 sg13g2_mux2_1 _6219_ (.A0(data_csrs_mem_7_),
    .A1(data_csrs_mem_39_),
    .S(net171),
    .X(_1876_));
 sg13g2_nand3_1 _6220_ (.B(net133),
    .C(next_dm_addr_i_7_),
    .A(net142),
    .Y(_1877_));
 sg13g2_o21ai_1 _6221_ (.B1(_1877_),
    .Y(_1878_),
    .A1(net138),
    .A2(net132));
 sg13g2_nor2b_1 _6222_ (.A(_0595_),
    .B_N(net581),
    .Y(_1879_));
 sg13g2_a22oi_1 _6223_ (.Y(_1880_),
    .B1(_1878_),
    .B2(_1879_),
    .A2(_1876_),
    .A1(net539));
 sg13g2_o21ai_1 _6224_ (.B1(_1880_),
    .Y(_1881_),
    .A1(_1495_),
    .A2(_1875_));
 sg13g2_a221oi_1 _6225_ (.B2(net483),
    .C1(_1881_),
    .B1(_1874_),
    .A1(hartinfo_i_7_),
    .Y(_1882_),
    .A2(net527));
 sg13g2_a21oi_2 _6226_ (.B1(net405),
    .Y(_1883_),
    .A2(_1882_),
    .A1(_1873_));
 sg13g2_mux2_1 _6227_ (.A0(\i_dm_csrs.i_fifo.mem_q_43_ ),
    .A1(_1883_),
    .S(net481),
    .X(_0147_));
 sg13g2_buf_1 fanout249 (.A(net250),
    .X(net249));
 sg13g2_mux2_1 _6229_ (.A0(\i_dm_csrs.i_fifo.mem_q_44_ ),
    .A1(_1334_),
    .S(net479),
    .X(_0148_));
 sg13g2_mux2_1 _6230_ (.A0(\i_dm_csrs.i_fifo.mem_q_45_ ),
    .A1(_1351_),
    .S(net480),
    .X(_0149_));
 sg13g2_mux2_1 _6231_ (.A0(\i_dm_csrs.i_fifo.mem_q_46_ ),
    .A1(_1375_),
    .S(net481),
    .X(_0150_));
 sg13g2_mux2_1 _6232_ (.A0(\i_dm_csrs.i_fifo.mem_q_47_ ),
    .A1(_1396_),
    .S(net478),
    .X(_0151_));
 sg13g2_mux2_1 _6233_ (.A0(\i_dm_csrs.i_fifo.mem_q_48_ ),
    .A1(_1416_),
    .S(net482),
    .X(_0152_));
 sg13g2_mux2_1 _6234_ (.A0(\i_dm_csrs.i_fifo.mem_q_49_ ),
    .A1(_1431_),
    .S(net479),
    .X(_0153_));
 sg13g2_mux2_1 _6235_ (.A0(\i_dm_csrs.i_fifo.mem_q_4_ ),
    .A1(_1810_),
    .S(net491),
    .X(_0154_));
 sg13g2_mux2_1 _6236_ (.A0(\i_dm_csrs.i_fifo.mem_q_50_ ),
    .A1(_1452_),
    .S(net478),
    .X(_0155_));
 sg13g2_mux2_1 _6237_ (.A0(\i_dm_csrs.i_fifo.mem_q_51_ ),
    .A1(_1467_),
    .S(net482),
    .X(_0156_));
 sg13g2_mux2_1 _6238_ (.A0(\i_dm_csrs.i_fifo.mem_q_52_ ),
    .A1(_1489_),
    .S(net479),
    .X(_0157_));
 sg13g2_mux2_1 _6239_ (.A0(\i_dm_csrs.i_fifo.mem_q_53_ ),
    .A1(_1511_),
    .S(net481),
    .X(_0158_));
 sg13g2_buf_1 fanout248 (.A(net249),
    .X(net248));
 sg13g2_mux2_1 _6241_ (.A0(\i_dm_csrs.i_fifo.mem_q_54_ ),
    .A1(_1530_),
    .S(net479),
    .X(_0159_));
 sg13g2_mux2_1 _6242_ (.A0(\i_dm_csrs.i_fifo.mem_q_55_ ),
    .A1(_1549_),
    .S(net481),
    .X(_0160_));
 sg13g2_mux2_1 _6243_ (.A0(\i_dm_csrs.i_fifo.mem_q_56_ ),
    .A1(_1570_),
    .S(net482),
    .X(_0161_));
 sg13g2_mux2_1 _6244_ (.A0(\i_dm_csrs.i_fifo.mem_q_57_ ),
    .A1(_1589_),
    .S(net481),
    .X(_0162_));
 sg13g2_mux2_1 _6245_ (.A0(\i_dm_csrs.i_fifo.mem_q_58_ ),
    .A1(_1606_),
    .S(net478),
    .X(_0163_));
 sg13g2_mux2_1 _6246_ (.A0(\i_dm_csrs.i_fifo.mem_q_59_ ),
    .A1(_1624_),
    .S(net482),
    .X(_0164_));
 sg13g2_mux2_1 _6247_ (.A0(\i_dm_csrs.i_fifo.mem_q_5_ ),
    .A1(_1825_),
    .S(net488),
    .X(_0165_));
 sg13g2_mux2_1 _6248_ (.A0(\i_dm_csrs.i_fifo.mem_q_60_ ),
    .A1(_1640_),
    .S(net482),
    .X(_0166_));
 sg13g2_mux2_1 _6249_ (.A0(\i_dm_csrs.i_fifo.mem_q_61_ ),
    .A1(_1655_),
    .S(net481),
    .X(_0167_));
 sg13g2_mux2_1 _6250_ (.A0(\i_dm_csrs.i_fifo.mem_q_62_ ),
    .A1(_1671_),
    .S(net480),
    .X(_0168_));
 sg13g2_mux2_1 _6251_ (.A0(\i_dm_csrs.i_fifo.mem_q_63_ ),
    .A1(_1688_),
    .S(net480),
    .X(_0169_));
 sg13g2_mux2_1 _6252_ (.A0(\i_dm_csrs.i_fifo.mem_q_64_ ),
    .A1(_1726_),
    .S(net481),
    .X(_0170_));
 sg13g2_mux2_1 _6253_ (.A0(\i_dm_csrs.i_fifo.mem_q_65_ ),
    .A1(_1740_),
    .S(net478),
    .X(_0171_));
 sg13g2_mux2_1 _6254_ (.A0(\i_dm_csrs.i_fifo.mem_q_66_ ),
    .A1(_1757_),
    .S(net478),
    .X(_0172_));
 sg13g2_mux2_1 _6255_ (.A0(\i_dm_csrs.i_fifo.mem_q_67_ ),
    .A1(_1771_),
    .S(net479),
    .X(_0173_));
 sg13g2_mux2_1 _6256_ (.A0(\i_dm_csrs.i_fifo.mem_q_6_ ),
    .A1(_1840_),
    .S(net489),
    .X(_0174_));
 sg13g2_mux2_1 _6257_ (.A0(\i_dm_csrs.i_fifo.mem_q_7_ ),
    .A1(_1855_),
    .S(net488),
    .X(_0175_));
 sg13g2_mux2_1 _6258_ (.A0(\i_dm_csrs.i_fifo.mem_q_8_ ),
    .A1(_1869_),
    .S(net488),
    .X(_0176_));
 sg13g2_mux2_1 _6259_ (.A0(\i_dm_csrs.i_fifo.mem_q_9_ ),
    .A1(_1883_),
    .S(net491),
    .X(_0177_));
 sg13g2_nand2_2 _6260_ (.Y(_1886_),
    .A(dmi_resp_ready_i),
    .B(dmi_resp_valid_o));
 sg13g2_mux2_1 _6261_ (.A0(\i_dm_csrs.i_fifo.read_pointer_n ),
    .A1(net638),
    .S(_1886_),
    .X(_1887_));
 sg13g2_and2_1 _6262_ (.A(dmi_rst_ni),
    .B(_1887_),
    .X(_0178_));
 sg13g2_nand2b_1 _6263_ (.Y(_1888_),
    .B(dmi_resp_ready_i),
    .A_N(\i_dm_csrs.i_fifo.status_cnt_q_0_ ));
 sg13g2_a21oi_2 _6264_ (.B1(net44),
    .Y(_1889_),
    .A2(_1888_),
    .A1(\i_dm_csrs.i_fifo.status_cnt_q_1_ ));
 sg13g2_nor2b_1 _6265_ (.A(dmi_resp_ready_i),
    .B_N(\i_dm_csrs.i_fifo.status_cnt_q_0_ ),
    .Y(_1890_));
 sg13g2_and3_1 _6266_ (.X(_1891_),
    .A(\i_dm_csrs.i_fifo.status_cnt_q_1_ ),
    .B(net44),
    .C(_1890_));
 sg13g2_o21ai_1 _6267_ (.B1(dmi_rst_ni),
    .Y(_1892_),
    .A1(\i_dm_csrs.i_fifo.status_cnt_q_1_ ),
    .A2(_1890_));
 sg13g2_nor3_1 _6268_ (.A(_1889_),
    .B(_1891_),
    .C(_1892_),
    .Y(_0179_));
 sg13g2_a21o_1 _6269_ (.A2(_0612_),
    .A1(dmi_resp_ready_i),
    .B1(\i_dm_csrs.i_fifo.status_cnt_n_0_ ),
    .X(_1893_));
 sg13g2_and2_1 _6270_ (.A(\i_dm_csrs.i_fifo.status_cnt_q_1_ ),
    .B(dmi_resp_ready_i),
    .X(_1894_));
 sg13g2_a21oi_1 _6271_ (.A1(\i_dm_csrs.i_fifo.status_cnt_n_0_ ),
    .A2(_1894_),
    .Y(_1895_),
    .B1(_1890_));
 sg13g2_nand3b_1 _6272_ (.B(_0612_),
    .C(\i_dm_csrs.i_fifo.status_cnt_n_0_ ),
    .Y(_1896_),
    .A_N(_1894_));
 sg13g2_o21ai_1 _6273_ (.B1(_1896_),
    .Y(_1897_),
    .A1(net44),
    .A2(_1895_));
 sg13g2_a21oi_1 _6274_ (.A1(\i_dm_csrs.i_fifo.status_cnt_q_0_ ),
    .A2(_1893_),
    .Y(_1898_),
    .B1(_1897_));
 sg13g2_nor2b_1 _6275_ (.A(_1898_),
    .B_N(dmi_rst_ni),
    .Y(_0180_));
 sg13g2_a21oi_1 _6276_ (.A1(\i_dm_csrs.i_fifo.write_pointer_q ),
    .A2(_0598_),
    .Y(_1899_),
    .B1(net489));
 sg13g2_nor2b_1 _6277_ (.A(_1899_),
    .B_N(dmi_rst_ni),
    .Y(_0181_));
 sg13g2_inv_1 _6278_ (.Y(_1900_),
    .A(\i_dm_csrs.progbuf_o_0_ ));
 sg13g2_a21oi_2 _6279_ (.B1(net639),
    .Y(_1901_),
    .A2(net586),
    .A1(_0901_));
 sg13g2_nor2_1 _6280_ (.A(net640),
    .B(_1148_),
    .Y(_1902_));
 sg13g2_nor2_2 _6281_ (.A(_1901_),
    .B(_1902_),
    .Y(_1903_));
 sg13g2_buf_2 fanout247 (.A(net249),
    .X(net247));
 sg13g2_nand2_2 _6283_ (.Y(_1905_),
    .A(net83),
    .B(net589));
 sg13g2_nor3_2 _6284_ (.A(net147),
    .B(net140),
    .C(_1905_),
    .Y(_1906_));
 sg13g2_buf_2 fanout246 (.A(dmi_req_i_0_),
    .X(net246));
 sg13g2_buf_4 fanout245 (.X(net245),
    .A(dmi_req_i_0_));
 sg13g2_nand3_1 _6287_ (.B(net525),
    .C(net349),
    .A(net246),
    .Y(_1909_));
 sg13g2_o21ai_1 _6288_ (.B1(_1909_),
    .Y(_0182_),
    .A1(_1900_),
    .A2(net349));
 sg13g2_nand2_2 _6289_ (.Y(_1910_),
    .A(net83),
    .B(net166));
 sg13g2_nand2_1 _6290_ (.Y(_1911_),
    .A(net156),
    .B(net45));
 sg13g2_nor2_2 _6291_ (.A(_1910_),
    .B(_1911_),
    .Y(_1912_));
 sg13g2_nand2_1 _6292_ (.Y(_1913_),
    .A(net127),
    .B(net435));
 sg13g2_nor3_1 _6293_ (.A(net589),
    .B(net607),
    .C(net141),
    .Y(_1914_));
 sg13g2_inv_2 _6294_ (.Y(_1915_),
    .A(_1901_));
 sg13g2_o21ai_1 _6295_ (.B1(_1915_),
    .Y(_1916_),
    .A1(net640),
    .A2(_1914_));
 sg13g2_buf_2 fanout244 (.A(dmi_req_i_10_),
    .X(net244));
 sg13g2_buf_4 fanout243 (.X(net243),
    .A(dmi_req_i_10_));
 sg13g2_buf_1 fanout242 (.A(dmi_req_i_11_),
    .X(net242));
 sg13g2_nand2_2 _6299_ (.Y(_1920_),
    .A(\i_dm_csrs.progbuf_o_100_ ),
    .B(net263));
 sg13g2_o21ai_1 _6300_ (.B1(_1920_),
    .Y(_0183_),
    .A1(_1913_),
    .A2(net262));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(dmi_req_i_11_));
 sg13g2_nand2_1 _6302_ (.Y(_1922_),
    .A(net125),
    .B(net438));
 sg13g2_nand2_2 _6303_ (.Y(_1923_),
    .A(\i_dm_csrs.progbuf_o_101_ ),
    .B(net271));
 sg13g2_o21ai_1 _6304_ (.B1(_1923_),
    .Y(_0184_),
    .A1(net271),
    .A2(_1922_));
 sg13g2_nand2_1 _6305_ (.Y(_1924_),
    .A(net123),
    .B(net437));
 sg13g2_nand2_2 _6306_ (.Y(_1925_),
    .A(\i_dm_csrs.progbuf_o_102_ ),
    .B(net267));
 sg13g2_o21ai_1 _6307_ (.B1(_1925_),
    .Y(_0185_),
    .A1(net267),
    .A2(_1924_));
 sg13g2_nand2_1 _6308_ (.Y(_1926_),
    .A(net121),
    .B(net436));
 sg13g2_nand2_2 _6309_ (.Y(_1927_),
    .A(\i_dm_csrs.progbuf_o_103_ ),
    .B(net265));
 sg13g2_o21ai_1 _6310_ (.B1(_1927_),
    .Y(_0186_),
    .A1(net265),
    .A2(_1926_));
 sg13g2_buf_1 fanout240 (.A(dmi_req_i_12_),
    .X(net240));
 sg13g2_nand2_1 _6312_ (.Y(_1929_),
    .A(net119),
    .B(net436));
 sg13g2_nand2_2 _6313_ (.Y(_1930_),
    .A(\i_dm_csrs.progbuf_o_104_ ),
    .B(net266));
 sg13g2_o21ai_1 _6314_ (.B1(_1930_),
    .Y(_0187_),
    .A1(net266),
    .A2(_1929_));
 sg13g2_nand2_1 _6315_ (.Y(_1931_),
    .A(net117),
    .B(net439));
 sg13g2_nand2_2 _6316_ (.Y(_1932_),
    .A(\i_dm_csrs.progbuf_o_105_ ),
    .B(net272));
 sg13g2_o21ai_1 _6317_ (.B1(_1932_),
    .Y(_0188_),
    .A1(net272),
    .A2(_1931_));
 sg13g2_nand2_1 _6318_ (.Y(_1933_),
    .A(net244),
    .B(net438));
 sg13g2_nand2_2 _6319_ (.Y(_1934_),
    .A(\i_dm_csrs.progbuf_o_106_ ),
    .B(net270));
 sg13g2_o21ai_1 _6320_ (.B1(_1934_),
    .Y(_0189_),
    .A1(net270),
    .A2(_1933_));
 sg13g2_buf_8 fanout239 (.A(dmi_req_i_12_),
    .X(net239));
 sg13g2_nand2_1 _6322_ (.Y(_1936_),
    .A(net242),
    .B(net438));
 sg13g2_nand2_2 _6323_ (.Y(_1937_),
    .A(\i_dm_csrs.progbuf_o_107_ ),
    .B(net271));
 sg13g2_o21ai_1 _6324_ (.B1(_1937_),
    .Y(_0190_),
    .A1(net271),
    .A2(_1936_));
 sg13g2_buf_1 fanout238 (.A(dmi_req_i_14_),
    .X(net238));
 sg13g2_nand2_1 _6326_ (.Y(_1939_),
    .A(net240),
    .B(net435));
 sg13g2_buf_4 fanout237 (.X(net237),
    .A(dmi_req_i_14_));
 sg13g2_nand2_2 _6328_ (.Y(_1941_),
    .A(\i_dm_csrs.progbuf_o_108_ ),
    .B(net264));
 sg13g2_o21ai_1 _6329_ (.B1(_1941_),
    .Y(_0191_),
    .A1(net264),
    .A2(_1939_));
 sg13g2_buf_1 fanout236 (.A(dmi_req_i_15_),
    .X(net236));
 sg13g2_nand2_1 _6331_ (.Y(_1943_),
    .A(net800),
    .B(net435));
 sg13g2_nand2_2 _6332_ (.Y(_1944_),
    .A(\i_dm_csrs.progbuf_o_109_ ),
    .B(net263));
 sg13g2_o21ai_1 _6333_ (.B1(_1944_),
    .Y(_0192_),
    .A1(net262),
    .A2(_1943_));
 sg13g2_inv_1 _6334_ (.Y(_1945_),
    .A(\i_dm_csrs.progbuf_o_10_ ));
 sg13g2_nand3_1 _6335_ (.B(net524),
    .C(net347),
    .A(net244),
    .Y(_1946_));
 sg13g2_o21ai_1 _6336_ (.B1(_1946_),
    .Y(_0193_),
    .A1(_1945_),
    .A2(net347));
 sg13g2_buf_4 fanout235 (.X(net235),
    .A(dmi_req_i_15_));
 sg13g2_buf_1 fanout234 (.A(dmi_req_i_16_),
    .X(net234));
 sg13g2_nand2_1 _6339_ (.Y(_1949_),
    .A(net238),
    .B(net436));
 sg13g2_nand2_2 _6340_ (.Y(_1950_),
    .A(\i_dm_csrs.progbuf_o_110_ ),
    .B(net265));
 sg13g2_o21ai_1 _6341_ (.B1(_1950_),
    .Y(_0194_),
    .A1(net265),
    .A2(_1949_));
 sg13g2_buf_4 fanout233 (.X(net233),
    .A(dmi_req_i_16_));
 sg13g2_buf_2 fanout232 (.A(dmi_req_i_17_),
    .X(net232));
 sg13g2_nand2_1 _6344_ (.Y(_1953_),
    .A(net236),
    .B(net435));
 sg13g2_nand2_2 _6345_ (.Y(_1954_),
    .A(\i_dm_csrs.progbuf_o_111_ ),
    .B(net263));
 sg13g2_o21ai_1 _6346_ (.B1(_1954_),
    .Y(_0195_),
    .A1(net263),
    .A2(_1953_));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(dmi_req_i_17_));
 sg13g2_nand2_1 _6348_ (.Y(_1956_),
    .A(net234),
    .B(net439));
 sg13g2_nand2_2 _6349_ (.Y(_1957_),
    .A(\i_dm_csrs.progbuf_o_112_ ),
    .B(net270));
 sg13g2_o21ai_1 _6350_ (.B1(_1957_),
    .Y(_0196_),
    .A1(net270),
    .A2(_1956_));
 sg13g2_buf_1 fanout230 (.A(dmi_req_i_18_),
    .X(net230));
 sg13g2_nand2_1 _6352_ (.Y(_1959_),
    .A(net232),
    .B(net438));
 sg13g2_nand2_2 _6353_ (.Y(_1960_),
    .A(\i_dm_csrs.progbuf_o_113_ ),
    .B(net269));
 sg13g2_o21ai_1 _6354_ (.B1(_1960_),
    .Y(_0197_),
    .A1(net269),
    .A2(_1959_));
 sg13g2_buf_4 fanout229 (.X(net229),
    .A(dmi_req_i_18_));
 sg13g2_nand2_1 _6356_ (.Y(_1962_),
    .A(net230),
    .B(net438));
 sg13g2_nand2_2 _6357_ (.Y(_1963_),
    .A(\i_dm_csrs.progbuf_o_114_ ),
    .B(net269));
 sg13g2_o21ai_1 _6358_ (.B1(_1963_),
    .Y(_0198_),
    .A1(net269),
    .A2(_1962_));
 sg13g2_buf_2 fanout228 (.A(dmi_req_i_19_),
    .X(net228));
 sg13g2_nand2_1 _6360_ (.Y(_1965_),
    .A(net228),
    .B(net438));
 sg13g2_nand2_2 _6361_ (.Y(_1966_),
    .A(\i_dm_csrs.progbuf_o_115_ ),
    .B(net269));
 sg13g2_o21ai_1 _6362_ (.B1(_1966_),
    .Y(_0199_),
    .A1(net269),
    .A2(_1965_));
 sg13g2_buf_4 fanout227 (.X(net227),
    .A(dmi_req_i_19_));
 sg13g2_nand2_1 _6364_ (.Y(_1968_),
    .A(net224),
    .B(net435));
 sg13g2_nand2_2 _6365_ (.Y(_1969_),
    .A(\i_dm_csrs.progbuf_o_116_ ),
    .B(net262));
 sg13g2_o21ai_1 _6366_ (.B1(_1969_),
    .Y(_0200_),
    .A1(net262),
    .A2(_1968_));
 sg13g2_buf_1 fanout226 (.A(dmi_req_i_1_),
    .X(net226));
 sg13g2_nand2_1 _6368_ (.Y(_1971_),
    .A(net222),
    .B(net435));
 sg13g2_nand2_2 _6369_ (.Y(_1972_),
    .A(\i_dm_csrs.progbuf_o_117_ ),
    .B(net262));
 sg13g2_o21ai_1 _6370_ (.B1(_1972_),
    .Y(_0201_),
    .A1(net262),
    .A2(_1971_));
 sg13g2_buf_8 fanout225 (.A(dmi_req_i_1_),
    .X(net225));
 sg13g2_nand2_1 _6372_ (.Y(_1974_),
    .A(net220),
    .B(net437));
 sg13g2_buf_2 fanout224 (.A(dmi_req_i_20_),
    .X(net224));
 sg13g2_nand2_2 _6374_ (.Y(_1976_),
    .A(\i_dm_csrs.progbuf_o_118_ ),
    .B(net267));
 sg13g2_o21ai_1 _6375_ (.B1(_1976_),
    .Y(_0202_),
    .A1(net267),
    .A2(_1974_));
 sg13g2_buf_8 fanout223 (.A(dmi_req_i_20_),
    .X(net223));
 sg13g2_nand2_1 _6377_ (.Y(_1978_),
    .A(net799),
    .B(net436));
 sg13g2_nand2_2 _6378_ (.Y(_1979_),
    .A(\i_dm_csrs.progbuf_o_119_ ),
    .B(net266));
 sg13g2_o21ai_1 _6379_ (.B1(_1979_),
    .Y(_0203_),
    .A1(net266),
    .A2(_1978_));
 sg13g2_inv_1 _6380_ (.Y(_1980_),
    .A(\i_dm_csrs.progbuf_o_11_ ));
 sg13g2_nand3_1 _6381_ (.B(net524),
    .C(net348),
    .A(net242),
    .Y(_1981_));
 sg13g2_o21ai_1 _6382_ (.B1(_1981_),
    .Y(_0204_),
    .A1(_1980_),
    .A2(net348));
 sg13g2_buf_1 fanout222 (.A(dmi_req_i_21_),
    .X(net222));
 sg13g2_buf_4 fanout221 (.X(net221),
    .A(dmi_req_i_21_));
 sg13g2_nand2_1 _6385_ (.Y(_1984_),
    .A(net218),
    .B(net435));
 sg13g2_nand2_2 _6386_ (.Y(_1985_),
    .A(\i_dm_csrs.progbuf_o_120_ ),
    .B(net264));
 sg13g2_o21ai_1 _6387_ (.B1(_1985_),
    .Y(_0205_),
    .A1(net268),
    .A2(_1984_));
 sg13g2_buf_2 fanout220 (.A(dmi_req_i_22_),
    .X(net220));
 sg13g2_buf_4 fanout219 (.X(net219),
    .A(dmi_req_i_22_));
 sg13g2_nand2_1 _6390_ (.Y(_1988_),
    .A(net216),
    .B(net438));
 sg13g2_nand2_2 _6391_ (.Y(_1989_),
    .A(\i_dm_csrs.progbuf_o_121_ ),
    .B(net271));
 sg13g2_o21ai_1 _6392_ (.B1(_1989_),
    .Y(_0206_),
    .A1(net271),
    .A2(_1988_));
 sg13g2_buf_2 fanout218 (.A(dmi_req_i_24_),
    .X(net218));
 sg13g2_nand2_1 _6394_ (.Y(_1991_),
    .A(net214),
    .B(net435));
 sg13g2_nand2_2 _6395_ (.Y(_1992_),
    .A(\i_dm_csrs.progbuf_o_122_ ),
    .B(net262));
 sg13g2_o21ai_1 _6396_ (.B1(_1992_),
    .Y(_0207_),
    .A1(net262),
    .A2(_1991_));
 sg13g2_buf_4 fanout217 (.X(net217),
    .A(dmi_req_i_24_));
 sg13g2_nand2_1 _6398_ (.Y(_1994_),
    .A(net212),
    .B(net438));
 sg13g2_nand2_2 _6399_ (.Y(_1995_),
    .A(\i_dm_csrs.progbuf_o_123_ ),
    .B(net271));
 sg13g2_o21ai_1 _6400_ (.B1(_1995_),
    .Y(_0208_),
    .A1(net271),
    .A2(_1994_));
 sg13g2_nand2_1 _6401_ (.Y(_1996_),
    .A(net210),
    .B(net439));
 sg13g2_nand2_2 _6402_ (.Y(_1997_),
    .A(\i_dm_csrs.progbuf_o_124_ ),
    .B(net269));
 sg13g2_o21ai_1 _6403_ (.B1(_1997_),
    .Y(_0209_),
    .A1(net269),
    .A2(_1996_));
 sg13g2_buf_2 fanout216 (.A(dmi_req_i_25_),
    .X(net216));
 sg13g2_nand2_1 _6405_ (.Y(_1999_),
    .A(net208),
    .B(net437));
 sg13g2_nand2_2 _6406_ (.Y(_2000_),
    .A(\i_dm_csrs.progbuf_o_125_ ),
    .B(net264));
 sg13g2_o21ai_1 _6407_ (.B1(_2000_),
    .Y(_0210_),
    .A1(net268),
    .A2(_1999_));
 sg13g2_buf_4 fanout215 (.X(net215),
    .A(dmi_req_i_25_));
 sg13g2_nand2_1 _6409_ (.Y(_2002_),
    .A(net204),
    .B(net437));
 sg13g2_nand2_2 _6410_ (.Y(_2003_),
    .A(\i_dm_csrs.progbuf_o_126_ ),
    .B(net264));
 sg13g2_o21ai_1 _6411_ (.B1(_2003_),
    .Y(_0211_),
    .A1(net264),
    .A2(_2002_));
 sg13g2_buf_1 fanout214 (.A(dmi_req_i_26_),
    .X(net214));
 sg13g2_nand2_1 _6413_ (.Y(_2005_),
    .A(net202),
    .B(net436));
 sg13g2_nand2_2 _6414_ (.Y(_2006_),
    .A(\i_dm_csrs.progbuf_o_127_ ),
    .B(net266));
 sg13g2_o21ai_1 _6415_ (.B1(_2006_),
    .Y(_0212_),
    .A1(net266),
    .A2(_2005_));
 sg13g2_inv_1 _6416_ (.Y(_2007_),
    .A(\i_dm_csrs.progbuf_o_128_ ));
 sg13g2_and2_1 _6417_ (.A(net134),
    .B(_0602_),
    .X(_2008_));
 sg13g2_nor2_1 _6418_ (.A(net639),
    .B(_2008_),
    .Y(_2009_));
 sg13g2_nor2_2 _6419_ (.A(_1901_),
    .B(_2009_),
    .Y(_2010_));
 sg13g2_buf_4 fanout213 (.X(net213),
    .A(dmi_req_i_26_));
 sg13g2_nor2_2 _6421_ (.A(_0896_),
    .B(_1905_),
    .Y(_2012_));
 sg13g2_buf_2 fanout212 (.A(dmi_req_i_27_),
    .X(net212));
 sg13g2_buf_4 fanout211 (.X(net211),
    .A(dmi_req_i_27_));
 sg13g2_nand3_1 _6424_ (.B(net520),
    .C(net338),
    .A(net246),
    .Y(_2015_));
 sg13g2_o21ai_1 _6425_ (.B1(_2015_),
    .Y(_0213_),
    .A1(_2007_),
    .A2(net338));
 sg13g2_inv_1 _6426_ (.Y(_2016_),
    .A(\i_dm_csrs.progbuf_o_129_ ));
 sg13g2_nand3_1 _6427_ (.B(net517),
    .C(net331),
    .A(net226),
    .Y(_2017_));
 sg13g2_o21ai_1 _6428_ (.B1(_2017_),
    .Y(_0214_),
    .A1(_2016_),
    .A2(net331));
 sg13g2_inv_1 _6429_ (.Y(_2018_),
    .A(\i_dm_csrs.progbuf_o_12_ ));
 sg13g2_nand3_1 _6430_ (.B(net521),
    .C(net341),
    .A(net240),
    .Y(_2019_));
 sg13g2_o21ai_1 _6431_ (.B1(_2019_),
    .Y(_0215_),
    .A1(_2018_),
    .A2(net341));
 sg13g2_inv_1 _6432_ (.Y(_2020_),
    .A(\i_dm_csrs.progbuf_o_130_ ));
 sg13g2_nand3_1 _6433_ (.B(net517),
    .C(net333),
    .A(net206),
    .Y(_2021_));
 sg13g2_o21ai_1 _6434_ (.B1(_2021_),
    .Y(_0216_),
    .A1(_2020_),
    .A2(net333));
 sg13g2_inv_1 _6435_ (.Y(_2022_),
    .A(\i_dm_csrs.progbuf_o_131_ ));
 sg13g2_nand3_1 _6436_ (.B(net517),
    .C(net332),
    .A(net129),
    .Y(_2023_));
 sg13g2_o21ai_1 _6437_ (.B1(_2023_),
    .Y(_0217_),
    .A1(_2022_),
    .A2(net331));
 sg13g2_inv_1 _6438_ (.Y(_2024_),
    .A(\i_dm_csrs.progbuf_o_132_ ));
 sg13g2_nand3_1 _6439_ (.B(net516),
    .C(net329),
    .A(net127),
    .Y(_2025_));
 sg13g2_o21ai_1 _6440_ (.B1(_2025_),
    .Y(_0218_),
    .A1(_2024_),
    .A2(net328));
 sg13g2_inv_1 _6441_ (.Y(_2026_),
    .A(\i_dm_csrs.progbuf_o_133_ ));
 sg13g2_nand3_1 _6442_ (.B(net519),
    .C(net337),
    .A(net125),
    .Y(_2027_));
 sg13g2_o21ai_1 _6443_ (.B1(_2027_),
    .Y(_0219_),
    .A1(_2026_),
    .A2(net337));
 sg13g2_inv_1 _6444_ (.Y(_2028_),
    .A(\i_dm_csrs.progbuf_o_134_ ));
 sg13g2_nand3_1 _6445_ (.B(net517),
    .C(net333),
    .A(net123),
    .Y(_2029_));
 sg13g2_o21ai_1 _6446_ (.B1(_2029_),
    .Y(_0220_),
    .A1(_2028_),
    .A2(net334));
 sg13g2_inv_1 _6447_ (.Y(_2030_),
    .A(\i_dm_csrs.progbuf_o_135_ ));
 sg13g2_nand3_1 _6448_ (.B(net517),
    .C(net333),
    .A(net121),
    .Y(_2031_));
 sg13g2_o21ai_1 _6449_ (.B1(_2031_),
    .Y(_0221_),
    .A1(_2030_),
    .A2(net333));
 sg13g2_inv_1 _6450_ (.Y(_2032_),
    .A(\i_dm_csrs.progbuf_o_136_ ));
 sg13g2_buf_2 fanout210 (.A(dmi_req_i_28_),
    .X(net210));
 sg13g2_nand3_1 _6452_ (.B(net517),
    .C(net332),
    .A(net119),
    .Y(_2034_));
 sg13g2_o21ai_1 _6453_ (.B1(_2034_),
    .Y(_0222_),
    .A1(_2032_),
    .A2(net331));
 sg13g2_inv_1 _6454_ (.Y(_2035_),
    .A(\i_dm_csrs.progbuf_o_137_ ));
 sg13g2_nand3_1 _6455_ (.B(net520),
    .C(net338),
    .A(net117),
    .Y(_2036_));
 sg13g2_o21ai_1 _6456_ (.B1(_2036_),
    .Y(_0223_),
    .A1(_2035_),
    .A2(net338));
 sg13g2_inv_1 _6457_ (.Y(_2037_),
    .A(\i_dm_csrs.progbuf_o_138_ ));
 sg13g2_buf_4 fanout209 (.X(net209),
    .A(dmi_req_i_28_));
 sg13g2_buf_1 fanout208 (.A(dmi_req_i_29_),
    .X(net208));
 sg13g2_nand3_1 _6460_ (.B(net519),
    .C(net335),
    .A(net244),
    .Y(_2040_));
 sg13g2_o21ai_1 _6461_ (.B1(_2040_),
    .Y(_0224_),
    .A1(_2037_),
    .A2(net336));
 sg13g2_inv_1 _6462_ (.Y(_2041_),
    .A(\i_dm_csrs.progbuf_o_139_ ));
 sg13g2_nand3_1 _6463_ (.B(net519),
    .C(net337),
    .A(net242),
    .Y(_2042_));
 sg13g2_o21ai_1 _6464_ (.B1(_2042_),
    .Y(_0225_),
    .A1(_2041_),
    .A2(net337));
 sg13g2_inv_1 _6465_ (.Y(_2043_),
    .A(\i_dm_csrs.progbuf_o_13_ ));
 sg13g2_nand3_1 _6466_ (.B(net521),
    .C(net340),
    .A(net800),
    .Y(_2044_));
 sg13g2_o21ai_1 _6467_ (.B1(_2044_),
    .Y(_0226_),
    .A1(_2043_),
    .A2(net339));
 sg13g2_inv_1 _6468_ (.Y(_2045_),
    .A(\i_dm_csrs.progbuf_o_140_ ));
 sg13g2_nand3_1 _6469_ (.B(net516),
    .C(net330),
    .A(net240),
    .Y(_2046_));
 sg13g2_o21ai_1 _6470_ (.B1(_2046_),
    .Y(_0227_),
    .A1(_2045_),
    .A2(net330));
 sg13g2_inv_1 _6471_ (.Y(_2047_),
    .A(\i_dm_csrs.progbuf_o_141_ ));
 sg13g2_nand3_1 _6472_ (.B(net516),
    .C(net329),
    .A(net800),
    .Y(_2048_));
 sg13g2_o21ai_1 _6473_ (.B1(_2048_),
    .Y(_0228_),
    .A1(_2047_),
    .A2(net329));
 sg13g2_inv_1 _6474_ (.Y(_2049_),
    .A(\i_dm_csrs.progbuf_o_142_ ));
 sg13g2_nand3_1 _6475_ (.B(net517),
    .C(net331),
    .A(net238),
    .Y(_2050_));
 sg13g2_o21ai_1 _6476_ (.B1(_2050_),
    .Y(_0229_),
    .A1(_2049_),
    .A2(net331));
 sg13g2_inv_1 _6477_ (.Y(_2051_),
    .A(\i_dm_csrs.progbuf_o_143_ ));
 sg13g2_nand3_1 _6478_ (.B(net516),
    .C(net329),
    .A(net236),
    .Y(_2052_));
 sg13g2_o21ai_1 _6479_ (.B1(_2052_),
    .Y(_0230_),
    .A1(_2051_),
    .A2(net329));
 sg13g2_inv_1 _6480_ (.Y(_2053_),
    .A(\i_dm_csrs.progbuf_o_144_ ));
 sg13g2_nand3_1 _6481_ (.B(net519),
    .C(net335),
    .A(net234),
    .Y(_2054_));
 sg13g2_o21ai_1 _6482_ (.B1(_2054_),
    .Y(_0231_),
    .A1(_2053_),
    .A2(net336));
 sg13g2_inv_1 _6483_ (.Y(_2055_),
    .A(\i_dm_csrs.progbuf_o_145_ ));
 sg13g2_nand3_1 _6484_ (.B(net519),
    .C(net335),
    .A(net232),
    .Y(_2056_));
 sg13g2_o21ai_1 _6485_ (.B1(_2056_),
    .Y(_0232_),
    .A1(_2055_),
    .A2(net335));
 sg13g2_inv_1 _6486_ (.Y(_2057_),
    .A(\i_dm_csrs.progbuf_o_146_ ));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(dmi_req_i_29_));
 sg13g2_nand3_1 _6488_ (.B(net519),
    .C(net335),
    .A(net230),
    .Y(_2059_));
 sg13g2_o21ai_1 _6489_ (.B1(_2059_),
    .Y(_0233_),
    .A1(_2057_),
    .A2(net335));
 sg13g2_inv_1 _6490_ (.Y(_2060_),
    .A(\i_dm_csrs.progbuf_o_147_ ));
 sg13g2_nand3_1 _6491_ (.B(net519),
    .C(net336),
    .A(net228),
    .Y(_2061_));
 sg13g2_o21ai_1 _6492_ (.B1(_2061_),
    .Y(_0234_),
    .A1(_2060_),
    .A2(net336));
 sg13g2_inv_1 _6493_ (.Y(_2062_),
    .A(\i_dm_csrs.progbuf_o_148_ ));
 sg13g2_buf_1 fanout206 (.A(dmi_req_i_2_),
    .X(net206));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(dmi_req_i_2_));
 sg13g2_nand3_1 _6496_ (.B(net516),
    .C(net328),
    .A(net224),
    .Y(_2065_));
 sg13g2_o21ai_1 _6497_ (.B1(_2065_),
    .Y(_0235_),
    .A1(_2062_),
    .A2(net328));
 sg13g2_inv_1 _6498_ (.Y(_2066_),
    .A(\i_dm_csrs.progbuf_o_149_ ));
 sg13g2_nand3_1 _6499_ (.B(net516),
    .C(net328),
    .A(net222),
    .Y(_2067_));
 sg13g2_o21ai_1 _6500_ (.B1(_2067_),
    .Y(_0236_),
    .A1(_2066_),
    .A2(net328));
 sg13g2_inv_1 _6501_ (.Y(_2068_),
    .A(\i_dm_csrs.progbuf_o_14_ ));
 sg13g2_nand3_1 _6502_ (.B(net522),
    .C(net342),
    .A(net238),
    .Y(_2069_));
 sg13g2_o21ai_1 _6503_ (.B1(_2069_),
    .Y(_0237_),
    .A1(_2068_),
    .A2(net342));
 sg13g2_inv_1 _6504_ (.Y(_2070_),
    .A(\i_dm_csrs.progbuf_o_150_ ));
 sg13g2_nand3_1 _6505_ (.B(net518),
    .C(net334),
    .A(net220),
    .Y(_2071_));
 sg13g2_o21ai_1 _6506_ (.B1(_2071_),
    .Y(_0238_),
    .A1(_2070_),
    .A2(net334));
 sg13g2_inv_1 _6507_ (.Y(_2072_),
    .A(\i_dm_csrs.progbuf_o_151_ ));
 sg13g2_nand3_1 _6508_ (.B(net518),
    .C(net332),
    .A(net799),
    .Y(_2073_));
 sg13g2_o21ai_1 _6509_ (.B1(_2073_),
    .Y(_0239_),
    .A1(_2072_),
    .A2(net332));
 sg13g2_inv_1 _6510_ (.Y(_2074_),
    .A(\i_dm_csrs.progbuf_o_152_ ));
 sg13g2_nand3_1 _6511_ (.B(net518),
    .C(net330),
    .A(net218),
    .Y(_2075_));
 sg13g2_o21ai_1 _6512_ (.B1(_2075_),
    .Y(_0240_),
    .A1(_2074_),
    .A2(net330));
 sg13g2_inv_1 _6513_ (.Y(_2076_),
    .A(\i_dm_csrs.progbuf_o_153_ ));
 sg13g2_nand3_1 _6514_ (.B(net520),
    .C(net337),
    .A(net216),
    .Y(_2077_));
 sg13g2_o21ai_1 _6515_ (.B1(_2077_),
    .Y(_0241_),
    .A1(_2076_),
    .A2(net337));
 sg13g2_inv_1 _6516_ (.Y(_2078_),
    .A(\i_dm_csrs.progbuf_o_154_ ));
 sg13g2_nand3_1 _6517_ (.B(net516),
    .C(net328),
    .A(net214),
    .Y(_2079_));
 sg13g2_o21ai_1 _6518_ (.B1(_2079_),
    .Y(_0242_),
    .A1(_2078_),
    .A2(net328));
 sg13g2_inv_1 _6519_ (.Y(_2080_),
    .A(\i_dm_csrs.progbuf_o_155_ ));
 sg13g2_nand3_1 _6520_ (.B(net519),
    .C(net337),
    .A(net212),
    .Y(_2081_));
 sg13g2_o21ai_1 _6521_ (.B1(_2081_),
    .Y(_0243_),
    .A1(_2080_),
    .A2(net337));
 sg13g2_inv_1 _6522_ (.Y(_2082_),
    .A(\i_dm_csrs.progbuf_o_156_ ));
 sg13g2_nand3_1 _6523_ (.B(net520),
    .C(net335),
    .A(net210),
    .Y(_2083_));
 sg13g2_o21ai_1 _6524_ (.B1(_2083_),
    .Y(_0244_),
    .A1(_2082_),
    .A2(net335));
 sg13g2_inv_1 _6525_ (.Y(_2084_),
    .A(\i_dm_csrs.progbuf_o_157_ ));
 sg13g2_nand3_1 _6526_ (.B(net518),
    .C(net330),
    .A(net208),
    .Y(_2085_));
 sg13g2_o21ai_1 _6527_ (.B1(_2085_),
    .Y(_0245_),
    .A1(_2084_),
    .A2(net330));
 sg13g2_inv_1 _6528_ (.Y(_2086_),
    .A(\i_dm_csrs.progbuf_o_158_ ));
 sg13g2_nand3_1 _6529_ (.B(net516),
    .C(net328),
    .A(net204),
    .Y(_2087_));
 sg13g2_o21ai_1 _6530_ (.B1(_2087_),
    .Y(_0246_),
    .A1(_2086_),
    .A2(net329));
 sg13g2_inv_1 _6531_ (.Y(_2088_),
    .A(\i_dm_csrs.progbuf_o_159_ ));
 sg13g2_nand3_1 _6532_ (.B(net517),
    .C(net331),
    .A(net202),
    .Y(_2089_));
 sg13g2_o21ai_1 _6533_ (.B1(_2089_),
    .Y(_0247_),
    .A1(_2088_),
    .A2(net331));
 sg13g2_inv_1 _6534_ (.Y(_2090_),
    .A(\i_dm_csrs.progbuf_o_15_ ));
 sg13g2_nand3_1 _6535_ (.B(net521),
    .C(net340),
    .A(net236),
    .Y(_2091_));
 sg13g2_o21ai_1 _6536_ (.B1(_2091_),
    .Y(_0248_),
    .A1(_2090_),
    .A2(net339));
 sg13g2_nor2_2 _6537_ (.A(_0896_),
    .B(_1910_),
    .Y(_2092_));
 sg13g2_nand2_1 _6538_ (.Y(_2093_),
    .A(net246),
    .B(net477));
 sg13g2_o21ai_1 _6539_ (.B1(_1915_),
    .Y(_2094_),
    .A1(net639),
    .A2(_1326_));
 sg13g2_buf_2 fanout204 (.A(dmi_req_i_30_),
    .X(net204));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(dmi_req_i_30_));
 sg13g2_buf_1 fanout202 (.A(dmi_req_i_31_),
    .X(net202));
 sg13g2_nand2_2 _6543_ (.Y(_2098_),
    .A(\i_dm_csrs.progbuf_o_160_ ),
    .B(net261));
 sg13g2_o21ai_1 _6544_ (.B1(_2098_),
    .Y(_0249_),
    .A1(_2093_),
    .A2(net261));
 sg13g2_buf_8 fanout201 (.A(dmi_req_i_31_),
    .X(net201));
 sg13g2_nand2_1 _6546_ (.Y(_2100_),
    .A(net226),
    .B(net474));
 sg13g2_nand2_2 _6547_ (.Y(_2101_),
    .A(\i_dm_csrs.progbuf_o_161_ ),
    .B(net255));
 sg13g2_o21ai_1 _6548_ (.B1(_2101_),
    .Y(_0250_),
    .A1(net255),
    .A2(_2100_));
 sg13g2_nand2_1 _6549_ (.Y(_2102_),
    .A(net206),
    .B(net474));
 sg13g2_nand2_2 _6550_ (.Y(_2103_),
    .A(\i_dm_csrs.progbuf_o_162_ ),
    .B(net256));
 sg13g2_o21ai_1 _6551_ (.B1(_2103_),
    .Y(_0251_),
    .A1(net256),
    .A2(_2102_));
 sg13g2_nand2_1 _6552_ (.Y(_2104_),
    .A(net129),
    .B(net474));
 sg13g2_nand2_2 _6553_ (.Y(_2105_),
    .A(\i_dm_csrs.progbuf_o_163_ ),
    .B(net255));
 sg13g2_o21ai_1 _6554_ (.B1(_2105_),
    .Y(_0252_),
    .A1(net256),
    .A2(_2104_));
 sg13g2_nand2_1 _6555_ (.Y(_2106_),
    .A(net127),
    .B(net473));
 sg13g2_nand2_2 _6556_ (.Y(_2107_),
    .A(\i_dm_csrs.progbuf_o_164_ ),
    .B(net253));
 sg13g2_o21ai_1 _6557_ (.B1(_2107_),
    .Y(_0253_),
    .A1(net252),
    .A2(_2106_));
 sg13g2_nand2_1 _6558_ (.Y(_2108_),
    .A(net125),
    .B(net476));
 sg13g2_nand2_2 _6559_ (.Y(_2109_),
    .A(\i_dm_csrs.progbuf_o_165_ ),
    .B(net260));
 sg13g2_o21ai_1 _6560_ (.B1(_2109_),
    .Y(_0254_),
    .A1(net260),
    .A2(_2108_));
 sg13g2_nand2_1 _6561_ (.Y(_2110_),
    .A(net123),
    .B(net474));
 sg13g2_nand2_2 _6562_ (.Y(_2111_),
    .A(\i_dm_csrs.progbuf_o_166_ ),
    .B(net256));
 sg13g2_o21ai_1 _6563_ (.B1(_2111_),
    .Y(_0255_),
    .A1(net256),
    .A2(_2110_));
 sg13g2_nand2_1 _6564_ (.Y(_2112_),
    .A(net121),
    .B(net474));
 sg13g2_nand2_2 _6565_ (.Y(_2113_),
    .A(\i_dm_csrs.progbuf_o_167_ ),
    .B(net256));
 sg13g2_o21ai_1 _6566_ (.B1(_2113_),
    .Y(_0256_),
    .A1(net256),
    .A2(_2112_));
 sg13g2_nand2_1 _6567_ (.Y(_2114_),
    .A(net119),
    .B(net474));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(dmi_req_i_34_));
 sg13g2_nand2_1 _6569_ (.Y(_2116_),
    .A(\i_dm_csrs.progbuf_o_168_ ),
    .B(net257));
 sg13g2_o21ai_1 _6570_ (.B1(_2116_),
    .Y(_0257_),
    .A1(net255),
    .A2(_2114_));
 sg13g2_nand2_1 _6571_ (.Y(_2117_),
    .A(net117),
    .B(net477));
 sg13g2_nand2_2 _6572_ (.Y(_2118_),
    .A(\i_dm_csrs.progbuf_o_169_ ),
    .B(net261));
 sg13g2_o21ai_1 _6573_ (.B1(_2118_),
    .Y(_0258_),
    .A1(net261),
    .A2(_2117_));
 sg13g2_inv_1 _6574_ (.Y(_2119_),
    .A(\i_dm_csrs.progbuf_o_16_ ));
 sg13g2_nand3_1 _6575_ (.B(net524),
    .C(net347),
    .A(net234),
    .Y(_2120_));
 sg13g2_o21ai_1 _6576_ (.B1(_2120_),
    .Y(_0259_),
    .A1(_2119_),
    .A2(net347));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net200));
 sg13g2_nand2_1 _6578_ (.Y(_2122_),
    .A(net244),
    .B(net476));
 sg13g2_nand2_2 _6579_ (.Y(_2123_),
    .A(\i_dm_csrs.progbuf_o_170_ ),
    .B(net258));
 sg13g2_o21ai_1 _6580_ (.B1(_2123_),
    .Y(_0260_),
    .A1(net259),
    .A2(_2122_));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(net200));
 sg13g2_nand2_1 _6582_ (.Y(_2125_),
    .A(net242),
    .B(net476));
 sg13g2_nand2_2 _6583_ (.Y(_2126_),
    .A(\i_dm_csrs.progbuf_o_171_ ),
    .B(net260));
 sg13g2_o21ai_1 _6584_ (.B1(_2126_),
    .Y(_0261_),
    .A1(net260),
    .A2(_2125_));
 sg13g2_nand2_1 _6585_ (.Y(_2127_),
    .A(net240),
    .B(net473));
 sg13g2_nand2_2 _6586_ (.Y(_2128_),
    .A(\i_dm_csrs.progbuf_o_172_ ),
    .B(net254));
 sg13g2_o21ai_1 _6587_ (.B1(_2128_),
    .Y(_0262_),
    .A1(net254),
    .A2(_2127_));
 sg13g2_nand2_1 _6588_ (.Y(_2129_),
    .A(net800),
    .B(net473));
 sg13g2_nand2_2 _6589_ (.Y(_2130_),
    .A(\i_dm_csrs.progbuf_o_173_ ),
    .B(net253));
 sg13g2_o21ai_1 _6590_ (.B1(_2130_),
    .Y(_0263_),
    .A1(net253),
    .A2(_2129_));
 sg13g2_nand2_1 _6591_ (.Y(_2131_),
    .A(net238),
    .B(net474));
 sg13g2_nand2_2 _6592_ (.Y(_2132_),
    .A(\i_dm_csrs.progbuf_o_174_ ),
    .B(net255));
 sg13g2_o21ai_1 _6593_ (.B1(_2132_),
    .Y(_0264_),
    .A1(net255),
    .A2(_2131_));
 sg13g2_nand2_1 _6594_ (.Y(_2133_),
    .A(net236),
    .B(net473));
 sg13g2_nand2_2 _6595_ (.Y(_2134_),
    .A(\i_dm_csrs.progbuf_o_175_ ),
    .B(net253));
 sg13g2_o21ai_1 _6596_ (.B1(_2134_),
    .Y(_0265_),
    .A1(net253),
    .A2(_2133_));
 sg13g2_nand2_1 _6597_ (.Y(_2135_),
    .A(net234),
    .B(net477));
 sg13g2_nand2_2 _6598_ (.Y(_2136_),
    .A(\i_dm_csrs.progbuf_o_176_ ),
    .B(net258));
 sg13g2_o21ai_1 _6599_ (.B1(_2136_),
    .Y(_0266_),
    .A1(net259),
    .A2(_2135_));
 sg13g2_nand2_1 _6600_ (.Y(_2137_),
    .A(net232),
    .B(net476));
 sg13g2_nand2_2 _6601_ (.Y(_2138_),
    .A(\i_dm_csrs.progbuf_o_177_ ),
    .B(net258));
 sg13g2_o21ai_1 _6602_ (.B1(_2138_),
    .Y(_0267_),
    .A1(net258),
    .A2(_2137_));
 sg13g2_nand2_1 _6603_ (.Y(_2139_),
    .A(net230),
    .B(net476));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(net200));
 sg13g2_nand2_2 _6605_ (.Y(_2141_),
    .A(\i_dm_csrs.progbuf_o_178_ ),
    .B(net258));
 sg13g2_o21ai_1 _6606_ (.B1(_2141_),
    .Y(_0268_),
    .A1(net258),
    .A2(_2139_));
 sg13g2_nand2_1 _6607_ (.Y(_2142_),
    .A(net228),
    .B(net476));
 sg13g2_nand2_2 _6608_ (.Y(_2143_),
    .A(\i_dm_csrs.progbuf_o_179_ ),
    .B(net259));
 sg13g2_o21ai_1 _6609_ (.B1(_2143_),
    .Y(_0269_),
    .A1(net259),
    .A2(_2142_));
 sg13g2_inv_1 _6610_ (.Y(_2144_),
    .A(\i_dm_csrs.progbuf_o_17_ ));
 sg13g2_buf_8 fanout196 (.A(net200),
    .X(net196));
 sg13g2_nand3_1 _6612_ (.B(net524),
    .C(net346),
    .A(net232),
    .Y(_2146_));
 sg13g2_o21ai_1 _6613_ (.B1(_2146_),
    .Y(_0270_),
    .A1(_2144_),
    .A2(net346));
 sg13g2_buf_8 fanout195 (.A(net200),
    .X(net195));
 sg13g2_nand2_1 _6615_ (.Y(_2148_),
    .A(net224),
    .B(net473));
 sg13g2_nand2_2 _6616_ (.Y(_2149_),
    .A(\i_dm_csrs.progbuf_o_180_ ),
    .B(net252));
 sg13g2_o21ai_1 _6617_ (.B1(_2149_),
    .Y(_0271_),
    .A1(net252),
    .A2(_2148_));
 sg13g2_buf_8 fanout194 (.A(net200),
    .X(net194));
 sg13g2_nand2_1 _6619_ (.Y(_2151_),
    .A(net222),
    .B(net473));
 sg13g2_nand2_2 _6620_ (.Y(_2152_),
    .A(\i_dm_csrs.progbuf_o_181_ ),
    .B(net252));
 sg13g2_o21ai_1 _6621_ (.B1(_2152_),
    .Y(_0272_),
    .A1(net252),
    .A2(_2151_));
 sg13g2_nand2_1 _6622_ (.Y(_2153_),
    .A(net220),
    .B(net475));
 sg13g2_nand2_2 _6623_ (.Y(_2154_),
    .A(\i_dm_csrs.progbuf_o_182_ ),
    .B(net257));
 sg13g2_o21ai_1 _6624_ (.B1(_2154_),
    .Y(_0273_),
    .A1(net257),
    .A2(_2153_));
 sg13g2_nand2_1 _6625_ (.Y(_2155_),
    .A(net798),
    .B(net475));
 sg13g2_nand2_2 _6626_ (.Y(_2156_),
    .A(\i_dm_csrs.progbuf_o_183_ ),
    .B(net257));
 sg13g2_o21ai_1 _6627_ (.B1(_2156_),
    .Y(_0274_),
    .A1(net257),
    .A2(_2155_));
 sg13g2_nand2_1 _6628_ (.Y(_2157_),
    .A(net218),
    .B(net475));
 sg13g2_nand2_2 _6629_ (.Y(_2158_),
    .A(\i_dm_csrs.progbuf_o_184_ ),
    .B(net254));
 sg13g2_o21ai_1 _6630_ (.B1(_2158_),
    .Y(_0275_),
    .A1(net254),
    .A2(_2157_));
 sg13g2_nand2_1 _6631_ (.Y(_2159_),
    .A(net216),
    .B(net476));
 sg13g2_nand2_2 _6632_ (.Y(_2160_),
    .A(\i_dm_csrs.progbuf_o_185_ ),
    .B(net260));
 sg13g2_o21ai_1 _6633_ (.B1(_2160_),
    .Y(_0276_),
    .A1(net260),
    .A2(_2159_));
 sg13g2_nand2_1 _6634_ (.Y(_2161_),
    .A(net214),
    .B(net473));
 sg13g2_nand2_2 _6635_ (.Y(_2162_),
    .A(\i_dm_csrs.progbuf_o_186_ ),
    .B(net252));
 sg13g2_o21ai_1 _6636_ (.B1(_2162_),
    .Y(_0277_),
    .A1(net252),
    .A2(_2161_));
 sg13g2_nand2_1 _6637_ (.Y(_2163_),
    .A(net212),
    .B(net476));
 sg13g2_nand2_2 _6638_ (.Y(_2164_),
    .A(\i_dm_csrs.progbuf_o_187_ ),
    .B(net260));
 sg13g2_o21ai_1 _6639_ (.B1(_2164_),
    .Y(_0278_),
    .A1(net260),
    .A2(_2163_));
 sg13g2_nand2_1 _6640_ (.Y(_2165_),
    .A(net210),
    .B(net477));
 sg13g2_nand2_2 _6641_ (.Y(_2166_),
    .A(\i_dm_csrs.progbuf_o_188_ ),
    .B(net258));
 sg13g2_o21ai_1 _6642_ (.B1(_2166_),
    .Y(_0279_),
    .A1(net258),
    .A2(_2165_));
 sg13g2_nand2_1 _6643_ (.Y(_2167_),
    .A(net208),
    .B(net475));
 sg13g2_nand2_2 _6644_ (.Y(_2168_),
    .A(\i_dm_csrs.progbuf_o_189_ ),
    .B(net254));
 sg13g2_o21ai_1 _6645_ (.B1(_2168_),
    .Y(_0280_),
    .A1(net254),
    .A2(_2167_));
 sg13g2_inv_1 _6646_ (.Y(_2169_),
    .A(\i_dm_csrs.progbuf_o_18_ ));
 sg13g2_nand3_1 _6647_ (.B(net524),
    .C(net346),
    .A(net230),
    .Y(_2170_));
 sg13g2_o21ai_1 _6648_ (.B1(_2170_),
    .Y(_0281_),
    .A1(_2169_),
    .A2(net346));
 sg13g2_nand2_1 _6649_ (.Y(_2171_),
    .A(net204),
    .B(net473));
 sg13g2_nand2_2 _6650_ (.Y(_2172_),
    .A(\i_dm_csrs.progbuf_o_190_ ),
    .B(net252));
 sg13g2_o21ai_1 _6651_ (.B1(_2172_),
    .Y(_0282_),
    .A1(net253),
    .A2(_2171_));
 sg13g2_nand2_1 _6652_ (.Y(_2173_),
    .A(net202),
    .B(net474));
 sg13g2_nand2_2 _6653_ (.Y(_2174_),
    .A(\i_dm_csrs.progbuf_o_191_ ),
    .B(net255));
 sg13g2_o21ai_1 _6654_ (.B1(_2174_),
    .Y(_0283_),
    .A1(net255),
    .A2(_2173_));
 sg13g2_nand2_1 _6655_ (.Y(_2175_),
    .A(net156),
    .B(net137));
 sg13g2_nor2_2 _6656_ (.A(_2175_),
    .B(_1905_),
    .Y(_2176_));
 sg13g2_nand2_1 _6657_ (.Y(_2177_),
    .A(net246),
    .B(net472));
 sg13g2_a21oi_1 _6658_ (.A1(net141),
    .A2(net548),
    .Y(_2178_),
    .B1(net639));
 sg13g2_or2_2 _6659_ (.X(_2179_),
    .B(_2178_),
    .A(_1901_));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(net200));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(net200));
 sg13g2_buf_1 fanout191 (.A(dmi_req_i_34_),
    .X(net191));
 sg13g2_nand2_2 _6663_ (.Y(_2183_),
    .A(\i_dm_csrs.progbuf_o_192_ ),
    .B(net327));
 sg13g2_o21ai_1 _6664_ (.B1(_2183_),
    .Y(_0284_),
    .A1(_2177_),
    .A2(net323));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_nand2_1 _6666_ (.Y(_2185_),
    .A(net226),
    .B(net469));
 sg13g2_nand2_2 _6667_ (.Y(_2186_),
    .A(\i_dm_csrs.progbuf_o_193_ ),
    .B(net320));
 sg13g2_o21ai_1 _6668_ (.B1(_2186_),
    .Y(_0285_),
    .A1(net320),
    .A2(_2185_));
 sg13g2_nand2_1 _6669_ (.Y(_2187_),
    .A(net206),
    .B(net469));
 sg13g2_nand2_2 _6670_ (.Y(_2188_),
    .A(\i_dm_csrs.progbuf_o_194_ ),
    .B(net322));
 sg13g2_o21ai_1 _6671_ (.B1(_2188_),
    .Y(_0286_),
    .A1(net322),
    .A2(_2187_));
 sg13g2_nand2_1 _6672_ (.Y(_2189_),
    .A(net129),
    .B(net469));
 sg13g2_nand2_1 _6673_ (.Y(_2190_),
    .A(\i_dm_csrs.progbuf_o_195_ ),
    .B(net321));
 sg13g2_o21ai_1 _6674_ (.B1(_2190_),
    .Y(_0287_),
    .A1(net320),
    .A2(_2189_));
 sg13g2_nand2_1 _6675_ (.Y(_2191_),
    .A(net127),
    .B(net468));
 sg13g2_nand2_2 _6676_ (.Y(_2192_),
    .A(\i_dm_csrs.progbuf_o_196_ ),
    .B(net318));
 sg13g2_o21ai_1 _6677_ (.B1(_2192_),
    .Y(_0288_),
    .A1(net317),
    .A2(_2191_));
 sg13g2_nand2_1 _6678_ (.Y(_2193_),
    .A(net125),
    .B(net471));
 sg13g2_nand2_2 _6679_ (.Y(_2194_),
    .A(\i_dm_csrs.progbuf_o_197_ ),
    .B(net326));
 sg13g2_o21ai_1 _6680_ (.B1(_2194_),
    .Y(_0289_),
    .A1(net326),
    .A2(_2193_));
 sg13g2_nand2_1 _6681_ (.Y(_2195_),
    .A(net123),
    .B(net469));
 sg13g2_nand2_2 _6682_ (.Y(_2196_),
    .A(\i_dm_csrs.progbuf_o_198_ ),
    .B(net322));
 sg13g2_o21ai_1 _6683_ (.B1(_2196_),
    .Y(_0290_),
    .A1(net322),
    .A2(_2195_));
 sg13g2_nand2_1 _6684_ (.Y(_2197_),
    .A(net121),
    .B(net469));
 sg13g2_nand2_2 _6685_ (.Y(_2198_),
    .A(\i_dm_csrs.progbuf_o_199_ ),
    .B(net322));
 sg13g2_o21ai_1 _6686_ (.B1(_2198_),
    .Y(_0291_),
    .A1(net322),
    .A2(_2197_));
 sg13g2_inv_1 _6687_ (.Y(_2199_),
    .A(\i_dm_csrs.progbuf_o_19_ ));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(net191));
 sg13g2_buf_2 fanout188 (.A(net191),
    .X(net188));
 sg13g2_nand3_1 _6690_ (.B(net525),
    .C(net347),
    .A(net228),
    .Y(_2202_));
 sg13g2_o21ai_1 _6691_ (.B1(_2202_),
    .Y(_0292_),
    .A1(_2199_),
    .A2(net347));
 sg13g2_inv_1 _6692_ (.Y(_2203_),
    .A(\i_dm_csrs.progbuf_o_1_ ));
 sg13g2_nand3_1 _6693_ (.B(net522),
    .C(net342),
    .A(net226),
    .Y(_2204_));
 sg13g2_o21ai_1 _6694_ (.B1(_2204_),
    .Y(_0293_),
    .A1(_2203_),
    .A2(net342));
 sg13g2_nand2_1 _6695_ (.Y(_2205_),
    .A(net119),
    .B(net469));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(net191));
 sg13g2_nand2_1 _6697_ (.Y(_2207_),
    .A(\i_dm_csrs.progbuf_o_200_ ),
    .B(net321));
 sg13g2_o21ai_1 _6698_ (.B1(_2207_),
    .Y(_0294_),
    .A1(net320),
    .A2(_2205_));
 sg13g2_nand2_1 _6699_ (.Y(_2208_),
    .A(net117),
    .B(net472));
 sg13g2_nand2_2 _6700_ (.Y(_2209_),
    .A(\i_dm_csrs.progbuf_o_201_ ),
    .B(net327));
 sg13g2_o21ai_1 _6701_ (.B1(_2209_),
    .Y(_0295_),
    .A1(net327),
    .A2(_2208_));
 sg13g2_buf_1 fanout186 (.A(net189),
    .X(net186));
 sg13g2_nand2_1 _6703_ (.Y(_2211_),
    .A(net244),
    .B(net471));
 sg13g2_nand2_2 _6704_ (.Y(_2212_),
    .A(\i_dm_csrs.progbuf_o_202_ ),
    .B(net324));
 sg13g2_o21ai_1 _6705_ (.B1(_2212_),
    .Y(_0296_),
    .A1(net325),
    .A2(_2211_));
 sg13g2_buf_2 fanout185 (.A(net189),
    .X(net185));
 sg13g2_nand2_1 _6707_ (.Y(_2214_),
    .A(net242),
    .B(net471));
 sg13g2_nand2_2 _6708_ (.Y(_2215_),
    .A(\i_dm_csrs.progbuf_o_203_ ),
    .B(net326));
 sg13g2_o21ai_1 _6709_ (.B1(_2215_),
    .Y(_0297_),
    .A1(net326),
    .A2(_2214_));
 sg13g2_nand2_1 _6710_ (.Y(_2216_),
    .A(net240),
    .B(net468));
 sg13g2_nand2_2 _6711_ (.Y(_2217_),
    .A(\i_dm_csrs.progbuf_o_204_ ),
    .B(net319));
 sg13g2_o21ai_1 _6712_ (.B1(_2217_),
    .Y(_0298_),
    .A1(net319),
    .A2(_2216_));
 sg13g2_nand2_1 _6713_ (.Y(_2218_),
    .A(net800),
    .B(net468));
 sg13g2_nand2_2 _6714_ (.Y(_2219_),
    .A(\i_dm_csrs.progbuf_o_205_ ),
    .B(net318));
 sg13g2_o21ai_1 _6715_ (.B1(_2219_),
    .Y(_0299_),
    .A1(net318),
    .A2(_2218_));
 sg13g2_nand2_1 _6716_ (.Y(_2220_),
    .A(net238),
    .B(net469));
 sg13g2_nand2_2 _6717_ (.Y(_2221_),
    .A(\i_dm_csrs.progbuf_o_206_ ),
    .B(net320));
 sg13g2_o21ai_1 _6718_ (.B1(_2221_),
    .Y(_0300_),
    .A1(net320),
    .A2(_2220_));
 sg13g2_nand2_1 _6719_ (.Y(_2222_),
    .A(net236),
    .B(net468));
 sg13g2_nand2_2 _6720_ (.Y(_2223_),
    .A(\i_dm_csrs.progbuf_o_207_ ),
    .B(net318));
 sg13g2_o21ai_1 _6721_ (.B1(_2223_),
    .Y(_0301_),
    .A1(net318),
    .A2(_2222_));
 sg13g2_nand2_1 _6722_ (.Y(_2224_),
    .A(net234),
    .B(net472));
 sg13g2_nand2_2 _6723_ (.Y(_2225_),
    .A(\i_dm_csrs.progbuf_o_208_ ),
    .B(net324));
 sg13g2_o21ai_1 _6724_ (.B1(_2225_),
    .Y(_0302_),
    .A1(net325),
    .A2(_2224_));
 sg13g2_nand2_1 _6725_ (.Y(_2226_),
    .A(net232),
    .B(net471));
 sg13g2_nand2_2 _6726_ (.Y(_2227_),
    .A(\i_dm_csrs.progbuf_o_209_ ),
    .B(net324));
 sg13g2_o21ai_1 _6727_ (.B1(_2227_),
    .Y(_0303_),
    .A1(net324),
    .A2(_2226_));
 sg13g2_inv_1 _6728_ (.Y(_2228_),
    .A(\i_dm_csrs.progbuf_o_20_ ));
 sg13g2_nand3_1 _6729_ (.B(net521),
    .C(net339),
    .A(net224),
    .Y(_2229_));
 sg13g2_o21ai_1 _6730_ (.B1(_2229_),
    .Y(_0304_),
    .A1(_2228_),
    .A2(net339));
 sg13g2_nand2_1 _6731_ (.Y(_2230_),
    .A(net230),
    .B(net471));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net189));
 sg13g2_nand2_2 _6733_ (.Y(_2232_),
    .A(\i_dm_csrs.progbuf_o_210_ ),
    .B(net324));
 sg13g2_o21ai_1 _6734_ (.B1(_2232_),
    .Y(_0305_),
    .A1(net324),
    .A2(_2230_));
 sg13g2_nand2_1 _6735_ (.Y(_2233_),
    .A(net228),
    .B(net471));
 sg13g2_nand2_2 _6736_ (.Y(_2234_),
    .A(\i_dm_csrs.progbuf_o_211_ ),
    .B(net325));
 sg13g2_o21ai_1 _6737_ (.B1(_2234_),
    .Y(_0306_),
    .A1(net325),
    .A2(_2233_));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(net189));
 sg13g2_nand2_1 _6739_ (.Y(_2236_),
    .A(net224),
    .B(net468));
 sg13g2_nand2_2 _6740_ (.Y(_2237_),
    .A(\i_dm_csrs.progbuf_o_212_ ),
    .B(net317));
 sg13g2_o21ai_1 _6741_ (.B1(_2237_),
    .Y(_0307_),
    .A1(net317),
    .A2(_2236_));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net189));
 sg13g2_nand2_1 _6743_ (.Y(_2239_),
    .A(net222),
    .B(net468));
 sg13g2_nand2_2 _6744_ (.Y(_2240_),
    .A(\i_dm_csrs.progbuf_o_213_ ),
    .B(net317));
 sg13g2_o21ai_1 _6745_ (.B1(_2240_),
    .Y(_0308_),
    .A1(net317),
    .A2(_2239_));
 sg13g2_nand2_1 _6746_ (.Y(_2241_),
    .A(net220),
    .B(net470));
 sg13g2_nand2_2 _6747_ (.Y(_2242_),
    .A(\i_dm_csrs.progbuf_o_214_ ),
    .B(net323));
 sg13g2_o21ai_1 _6748_ (.B1(_2242_),
    .Y(_0309_),
    .A1(net323),
    .A2(_2241_));
 sg13g2_nand2_1 _6749_ (.Y(_2243_),
    .A(net798),
    .B(net470));
 sg13g2_nand2_2 _6750_ (.Y(_2244_),
    .A(\i_dm_csrs.progbuf_o_215_ ),
    .B(net321));
 sg13g2_o21ai_1 _6751_ (.B1(_2244_),
    .Y(_0310_),
    .A1(net321),
    .A2(_2243_));
 sg13g2_nand2_1 _6752_ (.Y(_2245_),
    .A(net218),
    .B(net470));
 sg13g2_nand2_2 _6753_ (.Y(_2246_),
    .A(\i_dm_csrs.progbuf_o_216_ ),
    .B(net319));
 sg13g2_o21ai_1 _6754_ (.B1(_2246_),
    .Y(_0311_),
    .A1(net319),
    .A2(_2245_));
 sg13g2_nand2_1 _6755_ (.Y(_2247_),
    .A(net216),
    .B(net471));
 sg13g2_nand2_2 _6756_ (.Y(_2248_),
    .A(\i_dm_csrs.progbuf_o_217_ ),
    .B(net326));
 sg13g2_o21ai_1 _6757_ (.B1(_2248_),
    .Y(_0312_),
    .A1(net326),
    .A2(_2247_));
 sg13g2_nand2_1 _6758_ (.Y(_2249_),
    .A(net214),
    .B(net468));
 sg13g2_nand2_2 _6759_ (.Y(_2250_),
    .A(\i_dm_csrs.progbuf_o_218_ ),
    .B(net317));
 sg13g2_o21ai_1 _6760_ (.B1(_2250_),
    .Y(_0313_),
    .A1(net317),
    .A2(_2249_));
 sg13g2_nand2_1 _6761_ (.Y(_2251_),
    .A(net212),
    .B(net471));
 sg13g2_nand2_2 _6762_ (.Y(_2252_),
    .A(\i_dm_csrs.progbuf_o_219_ ),
    .B(net326));
 sg13g2_o21ai_1 _6763_ (.B1(_2252_),
    .Y(_0314_),
    .A1(net326),
    .A2(_2251_));
 sg13g2_inv_1 _6764_ (.Y(_2253_),
    .A(\i_dm_csrs.progbuf_o_21_ ));
 sg13g2_nand3_1 _6765_ (.B(net521),
    .C(net339),
    .A(net222),
    .Y(_2254_));
 sg13g2_o21ai_1 _6766_ (.B1(_2254_),
    .Y(_0315_),
    .A1(_2253_),
    .A2(net339));
 sg13g2_nand2_1 _6767_ (.Y(_2255_),
    .A(net210),
    .B(net472));
 sg13g2_nand2_2 _6768_ (.Y(_2256_),
    .A(\i_dm_csrs.progbuf_o_220_ ),
    .B(net324));
 sg13g2_o21ai_1 _6769_ (.B1(_2256_),
    .Y(_0316_),
    .A1(net324),
    .A2(_2255_));
 sg13g2_nand2_1 _6770_ (.Y(_2257_),
    .A(net208),
    .B(net470));
 sg13g2_nand2_2 _6771_ (.Y(_2258_),
    .A(\i_dm_csrs.progbuf_o_221_ ),
    .B(net319));
 sg13g2_o21ai_1 _6772_ (.B1(_2258_),
    .Y(_0317_),
    .A1(net319),
    .A2(_2257_));
 sg13g2_nand2_1 _6773_ (.Y(_2259_),
    .A(net204),
    .B(net468));
 sg13g2_nand2_2 _6774_ (.Y(_2260_),
    .A(\i_dm_csrs.progbuf_o_222_ ),
    .B(net317));
 sg13g2_o21ai_1 _6775_ (.B1(_2260_),
    .Y(_0318_),
    .A1(net318),
    .A2(_2259_));
 sg13g2_nand2_1 _6776_ (.Y(_2261_),
    .A(net202),
    .B(net469));
 sg13g2_nand2_2 _6777_ (.Y(_2262_),
    .A(\i_dm_csrs.progbuf_o_223_ ),
    .B(net320));
 sg13g2_o21ai_1 _6778_ (.B1(_2262_),
    .Y(_0319_),
    .A1(net320),
    .A2(_2261_));
 sg13g2_inv_1 _6779_ (.Y(_2263_),
    .A(\i_dm_csrs.progbuf_o_224_ ));
 sg13g2_a21oi_2 _6780_ (.B1(_1901_),
    .Y(_2264_),
    .A2(_0621_),
    .A1(_0893_));
 sg13g2_buf_2 fanout181 (.A(net190),
    .X(net181));
 sg13g2_nor2_2 _6782_ (.A(_2175_),
    .B(_1910_),
    .Y(_2266_));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net190));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(net190));
 sg13g2_nand3_1 _6785_ (.B(net467),
    .C(net311),
    .A(net246),
    .Y(_2269_));
 sg13g2_o21ai_1 _6786_ (.B1(_2269_),
    .Y(_0320_),
    .A1(_2263_),
    .A2(net316));
 sg13g2_inv_1 _6787_ (.Y(_2270_),
    .A(\i_dm_csrs.progbuf_o_225_ ));
 sg13g2_nand3_1 _6788_ (.B(net464),
    .C(net309),
    .A(net226),
    .Y(_2271_));
 sg13g2_o21ai_1 _6789_ (.B1(_2271_),
    .Y(_0321_),
    .A1(_2270_),
    .A2(net309));
 sg13g2_inv_1 _6790_ (.Y(_2272_),
    .A(\i_dm_csrs.progbuf_o_226_ ));
 sg13g2_nand3_1 _6791_ (.B(net464),
    .C(net308),
    .A(net206),
    .Y(_2273_));
 sg13g2_o21ai_1 _6792_ (.B1(_2273_),
    .Y(_0322_),
    .A1(_2272_),
    .A2(net308));
 sg13g2_inv_1 _6793_ (.Y(_2274_),
    .A(\i_dm_csrs.progbuf_o_227_ ));
 sg13g2_nand3_1 _6794_ (.B(net464),
    .C(net310),
    .A(net129),
    .Y(_2275_));
 sg13g2_o21ai_1 _6795_ (.B1(_2275_),
    .Y(_0323_),
    .A1(_2274_),
    .A2(net308));
 sg13g2_inv_1 _6796_ (.Y(_2276_),
    .A(\i_dm_csrs.progbuf_o_228_ ));
 sg13g2_nand3_1 _6797_ (.B(net463),
    .C(net306),
    .A(net127),
    .Y(_2277_));
 sg13g2_o21ai_1 _6798_ (.B1(_2277_),
    .Y(_0324_),
    .A1(_2276_),
    .A2(net305));
 sg13g2_inv_1 _6799_ (.Y(_2278_),
    .A(\i_dm_csrs.progbuf_o_229_ ));
 sg13g2_nand3_1 _6800_ (.B(net466),
    .C(net315),
    .A(net125),
    .Y(_2279_));
 sg13g2_o21ai_1 _6801_ (.B1(_2279_),
    .Y(_0325_),
    .A1(_2278_),
    .A2(net315));
 sg13g2_inv_1 _6802_ (.Y(_2280_),
    .A(\i_dm_csrs.progbuf_o_22_ ));
 sg13g2_nand3_1 _6803_ (.B(net522),
    .C(net344),
    .A(net220),
    .Y(_2281_));
 sg13g2_o21ai_1 _6804_ (.B1(_2281_),
    .Y(_0326_),
    .A1(_2280_),
    .A2(net344));
 sg13g2_inv_1 _6805_ (.Y(_2282_),
    .A(\i_dm_csrs.progbuf_o_230_ ));
 sg13g2_nand3_1 _6806_ (.B(net464),
    .C(net308),
    .A(net123),
    .Y(_2283_));
 sg13g2_o21ai_1 _6807_ (.B1(_2283_),
    .Y(_0327_),
    .A1(_2282_),
    .A2(net308));
 sg13g2_inv_1 _6808_ (.Y(_2284_),
    .A(\i_dm_csrs.progbuf_o_231_ ));
 sg13g2_nand3_1 _6809_ (.B(net464),
    .C(net308),
    .A(net121),
    .Y(_2285_));
 sg13g2_o21ai_1 _6810_ (.B1(_2285_),
    .Y(_0328_),
    .A1(_2284_),
    .A2(net308));
 sg13g2_inv_1 _6811_ (.Y(_2286_),
    .A(\i_dm_csrs.progbuf_o_232_ ));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(net190));
 sg13g2_nand3_1 _6813_ (.B(net464),
    .C(net309),
    .A(net119),
    .Y(_2288_));
 sg13g2_o21ai_1 _6814_ (.B1(_2288_),
    .Y(_0329_),
    .A1(_2286_),
    .A2(net309));
 sg13g2_inv_1 _6815_ (.Y(_2289_),
    .A(\i_dm_csrs.progbuf_o_233_ ));
 sg13g2_nand3_1 _6816_ (.B(net467),
    .C(net316),
    .A(net117),
    .Y(_2290_));
 sg13g2_o21ai_1 _6817_ (.B1(_2290_),
    .Y(_0330_),
    .A1(_2289_),
    .A2(net316));
 sg13g2_inv_1 _6818_ (.Y(_2291_),
    .A(\i_dm_csrs.progbuf_o_234_ ));
 sg13g2_buf_2 fanout177 (.A(net190),
    .X(net177));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(net187));
 sg13g2_nand3_1 _6821_ (.B(net466),
    .C(net314),
    .A(net243),
    .Y(_2294_));
 sg13g2_o21ai_1 _6822_ (.B1(_2294_),
    .Y(_0331_),
    .A1(_2291_),
    .A2(net314));
 sg13g2_inv_1 _6823_ (.Y(_2295_),
    .A(\i_dm_csrs.progbuf_o_235_ ));
 sg13g2_nand3_1 _6824_ (.B(net465),
    .C(net307),
    .A(net241),
    .Y(_2296_));
 sg13g2_o21ai_1 _6825_ (.B1(_2296_),
    .Y(_0332_),
    .A1(_2295_),
    .A2(net307));
 sg13g2_inv_1 _6826_ (.Y(_2297_),
    .A(\i_dm_csrs.progbuf_o_236_ ));
 sg13g2_nand3_1 _6827_ (.B(net463),
    .C(net307),
    .A(net240),
    .Y(_2298_));
 sg13g2_o21ai_1 _6828_ (.B1(_2298_),
    .Y(_0333_),
    .A1(_2297_),
    .A2(net307));
 sg13g2_inv_1 _6829_ (.Y(_2299_),
    .A(\i_dm_csrs.progbuf_o_237_ ));
 sg13g2_nand3_1 _6830_ (.B(net463),
    .C(net306),
    .A(net800),
    .Y(_2300_));
 sg13g2_o21ai_1 _6831_ (.B1(_2300_),
    .Y(_0334_),
    .A1(_2299_),
    .A2(net306));
 sg13g2_inv_1 _6832_ (.Y(_2301_),
    .A(\i_dm_csrs.progbuf_o_238_ ));
 sg13g2_nand3_1 _6833_ (.B(net464),
    .C(net308),
    .A(net238),
    .Y(_2302_));
 sg13g2_o21ai_1 _6834_ (.B1(_2302_),
    .Y(_0335_),
    .A1(_2301_),
    .A2(net309));
 sg13g2_inv_1 _6835_ (.Y(_2303_),
    .A(\i_dm_csrs.progbuf_o_239_ ));
 sg13g2_nand3_1 _6836_ (.B(net463),
    .C(net306),
    .A(net236),
    .Y(_2304_));
 sg13g2_o21ai_1 _6837_ (.B1(_2304_),
    .Y(_0336_),
    .A1(_2303_),
    .A2(net306));
 sg13g2_inv_1 _6838_ (.Y(_2305_),
    .A(\i_dm_csrs.progbuf_o_23_ ));
 sg13g2_nand3_1 _6839_ (.B(net522),
    .C(net343),
    .A(net798),
    .Y(_2306_));
 sg13g2_o21ai_1 _6840_ (.B1(_2306_),
    .Y(_0337_),
    .A1(_2305_),
    .A2(net343));
 sg13g2_inv_1 _6841_ (.Y(_2307_),
    .A(\i_dm_csrs.progbuf_o_240_ ));
 sg13g2_nand3_1 _6842_ (.B(net466),
    .C(net314),
    .A(net234),
    .Y(_2308_));
 sg13g2_o21ai_1 _6843_ (.B1(_2308_),
    .Y(_0338_),
    .A1(_2307_),
    .A2(net314));
 sg13g2_inv_1 _6844_ (.Y(_2309_),
    .A(\i_dm_csrs.progbuf_o_241_ ));
 sg13g2_nand3_1 _6845_ (.B(net466),
    .C(net313),
    .A(net232),
    .Y(_2310_));
 sg13g2_o21ai_1 _6846_ (.B1(_2310_),
    .Y(_0339_),
    .A1(_2309_),
    .A2(net313));
 sg13g2_inv_1 _6847_ (.Y(_2311_),
    .A(\i_dm_csrs.progbuf_o_242_ ));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net187));
 sg13g2_nand3_1 _6849_ (.B(net466),
    .C(net313),
    .A(net230),
    .Y(_2313_));
 sg13g2_o21ai_1 _6850_ (.B1(_2313_),
    .Y(_0340_),
    .A1(_2311_),
    .A2(net313));
 sg13g2_inv_1 _6851_ (.Y(_2314_),
    .A(\i_dm_csrs.progbuf_o_243_ ));
 sg13g2_nand3_1 _6852_ (.B(net466),
    .C(net313),
    .A(net228),
    .Y(_2315_));
 sg13g2_o21ai_1 _6853_ (.B1(_2315_),
    .Y(_0341_),
    .A1(_2314_),
    .A2(net313));
 sg13g2_inv_1 _6854_ (.Y(_2316_),
    .A(\i_dm_csrs.progbuf_o_244_ ));
 sg13g2_buf_4 fanout174 (.X(net174),
    .A(net187));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(net187));
 sg13g2_nand3_1 _6857_ (.B(net463),
    .C(net305),
    .A(net224),
    .Y(_2319_));
 sg13g2_o21ai_1 _6858_ (.B1(_2319_),
    .Y(_0342_),
    .A1(_2316_),
    .A2(net305));
 sg13g2_inv_1 _6859_ (.Y(_2320_),
    .A(\i_dm_csrs.progbuf_o_245_ ));
 sg13g2_nand3_1 _6860_ (.B(net463),
    .C(net305),
    .A(net221),
    .Y(_2321_));
 sg13g2_o21ai_1 _6861_ (.B1(_2321_),
    .Y(_0343_),
    .A1(_2320_),
    .A2(net305));
 sg13g2_inv_1 _6862_ (.Y(_2322_),
    .A(\i_dm_csrs.progbuf_o_246_ ));
 sg13g2_nand3_1 _6863_ (.B(net465),
    .C(net311),
    .A(net220),
    .Y(_2323_));
 sg13g2_o21ai_1 _6864_ (.B1(_2323_),
    .Y(_0344_),
    .A1(_2322_),
    .A2(net311));
 sg13g2_inv_1 _6865_ (.Y(_2324_),
    .A(\i_dm_csrs.progbuf_o_247_ ));
 sg13g2_nand3_1 _6866_ (.B(net465),
    .C(net309),
    .A(net798),
    .Y(_2325_));
 sg13g2_o21ai_1 _6867_ (.B1(_2325_),
    .Y(_0345_),
    .A1(_2324_),
    .A2(net310));
 sg13g2_inv_1 _6868_ (.Y(_2326_),
    .A(\i_dm_csrs.progbuf_o_248_ ));
 sg13g2_nand3_1 _6869_ (.B(net465),
    .C(net307),
    .A(net218),
    .Y(_2327_));
 sg13g2_o21ai_1 _6870_ (.B1(_2327_),
    .Y(_0346_),
    .A1(_2326_),
    .A2(net312));
 sg13g2_inv_1 _6871_ (.Y(_2328_),
    .A(\i_dm_csrs.progbuf_o_249_ ));
 sg13g2_nand3_1 _6872_ (.B(net466),
    .C(net315),
    .A(net216),
    .Y(_2329_));
 sg13g2_o21ai_1 _6873_ (.B1(_2329_),
    .Y(_0347_),
    .A1(_2328_),
    .A2(net315));
 sg13g2_inv_1 _6874_ (.Y(_2330_),
    .A(\i_dm_csrs.progbuf_o_24_ ));
 sg13g2_nand3_1 _6875_ (.B(net521),
    .C(net341),
    .A(net218),
    .Y(_2331_));
 sg13g2_o21ai_1 _6876_ (.B1(_2331_),
    .Y(_0348_),
    .A1(_2330_),
    .A2(net341));
 sg13g2_inv_1 _6877_ (.Y(_2332_),
    .A(\i_dm_csrs.progbuf_o_250_ ));
 sg13g2_nand3_1 _6878_ (.B(net463),
    .C(net305),
    .A(net214),
    .Y(_2333_));
 sg13g2_o21ai_1 _6879_ (.B1(_2333_),
    .Y(_0349_),
    .A1(_2332_),
    .A2(net305));
 sg13g2_inv_1 _6880_ (.Y(_2334_),
    .A(\i_dm_csrs.progbuf_o_251_ ));
 sg13g2_nand3_1 _6881_ (.B(net466),
    .C(net315),
    .A(net212),
    .Y(_2335_));
 sg13g2_o21ai_1 _6882_ (.B1(_2335_),
    .Y(_0350_),
    .A1(_2334_),
    .A2(net315));
 sg13g2_inv_1 _6883_ (.Y(_2336_),
    .A(\i_dm_csrs.progbuf_o_252_ ));
 sg13g2_nand3_1 _6884_ (.B(net467),
    .C(net313),
    .A(net210),
    .Y(_2337_));
 sg13g2_o21ai_1 _6885_ (.B1(_2337_),
    .Y(_0351_),
    .A1(_2336_),
    .A2(net313));
 sg13g2_inv_1 _6886_ (.Y(_2338_),
    .A(\i_dm_csrs.progbuf_o_253_ ));
 sg13g2_nand3_1 _6887_ (.B(net465),
    .C(net307),
    .A(net208),
    .Y(_2339_));
 sg13g2_o21ai_1 _6888_ (.B1(_2339_),
    .Y(_0352_),
    .A1(_2338_),
    .A2(net312));
 sg13g2_inv_1 _6889_ (.Y(_2340_),
    .A(\i_dm_csrs.progbuf_o_254_ ));
 sg13g2_nand3_1 _6890_ (.B(net463),
    .C(net305),
    .A(net204),
    .Y(_2341_));
 sg13g2_o21ai_1 _6891_ (.B1(_2341_),
    .Y(_0353_),
    .A1(_2340_),
    .A2(net306));
 sg13g2_inv_1 _6892_ (.Y(_2342_),
    .A(\i_dm_csrs.progbuf_o_255_ ));
 sg13g2_nand3_1 _6893_ (.B(net464),
    .C(net309),
    .A(net202),
    .Y(_2343_));
 sg13g2_o21ai_1 _6894_ (.B1(_2343_),
    .Y(_0354_),
    .A1(_2342_),
    .A2(net309));
 sg13g2_inv_1 _6895_ (.Y(_2344_),
    .A(\i_dm_csrs.progbuf_o_25_ ));
 sg13g2_nand3_1 _6896_ (.B(net524),
    .C(net348),
    .A(net216),
    .Y(_2345_));
 sg13g2_o21ai_1 _6897_ (.B1(_2345_),
    .Y(_0355_),
    .A1(_2344_),
    .A2(net348));
 sg13g2_inv_1 _6898_ (.Y(_2346_),
    .A(\i_dm_csrs.progbuf_o_26_ ));
 sg13g2_buf_4 fanout172 (.X(net172),
    .A(net187));
 sg13g2_nand3_1 _6900_ (.B(net521),
    .C(net339),
    .A(net214),
    .Y(_2348_));
 sg13g2_o21ai_1 _6901_ (.B1(_2348_),
    .Y(_0356_),
    .A1(_2346_),
    .A2(net339));
 sg13g2_inv_1 _6902_ (.Y(_2349_),
    .A(\i_dm_csrs.progbuf_o_27_ ));
 sg13g2_nand3_1 _6903_ (.B(net524),
    .C(net346),
    .A(net212),
    .Y(_2350_));
 sg13g2_o21ai_1 _6904_ (.B1(_2350_),
    .Y(_0357_),
    .A1(_2349_),
    .A2(net346));
 sg13g2_inv_1 _6905_ (.Y(_2351_),
    .A(\i_dm_csrs.progbuf_o_28_ ));
 sg13g2_buf_4 fanout171 (.X(net171),
    .A(net187));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(net187));
 sg13g2_nand3_1 _6908_ (.B(net525),
    .C(net346),
    .A(net210),
    .Y(_2354_));
 sg13g2_o21ai_1 _6909_ (.B1(_2354_),
    .Y(_0358_),
    .A1(_2351_),
    .A2(net346));
 sg13g2_inv_1 _6910_ (.Y(_2355_),
    .A(\i_dm_csrs.progbuf_o_29_ ));
 sg13g2_nand3_1 _6911_ (.B(net523),
    .C(net341),
    .A(net207),
    .Y(_2356_));
 sg13g2_o21ai_1 _6912_ (.B1(_2356_),
    .Y(_0359_),
    .A1(_2355_),
    .A2(net345));
 sg13g2_inv_1 _6913_ (.Y(_2357_),
    .A(\i_dm_csrs.progbuf_o_2_ ));
 sg13g2_nand3_1 _6914_ (.B(net522),
    .C(net343),
    .A(net206),
    .Y(_2358_));
 sg13g2_o21ai_1 _6915_ (.B1(_2358_),
    .Y(_0360_),
    .A1(_2357_),
    .A2(net343));
 sg13g2_inv_1 _6916_ (.Y(_2359_),
    .A(\i_dm_csrs.progbuf_o_30_ ));
 sg13g2_nand3_1 _6917_ (.B(net523),
    .C(net341),
    .A(net204),
    .Y(_2360_));
 sg13g2_o21ai_1 _6918_ (.B1(_2360_),
    .Y(_0361_),
    .A1(_2359_),
    .A2(net345));
 sg13g2_inv_1 _6919_ (.Y(_2361_),
    .A(\i_dm_csrs.progbuf_o_31_ ));
 sg13g2_nand3_1 _6920_ (.B(net522),
    .C(net342),
    .A(net201),
    .Y(_2362_));
 sg13g2_o21ai_1 _6921_ (.B1(_2362_),
    .Y(_0362_),
    .A1(_2361_),
    .A2(net342));
 sg13g2_inv_1 _6922_ (.Y(_2363_),
    .A(\i_dm_csrs.progbuf_o_32_ ));
 sg13g2_and2_2 _6923_ (.A(net45),
    .B(net581),
    .X(_2364_));
 sg13g2_nor2_1 _6924_ (.A(net639),
    .B(_2364_),
    .Y(_2365_));
 sg13g2_nor2_2 _6925_ (.A(_1901_),
    .B(_2365_),
    .Y(_2366_));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(net187));
 sg13g2_nor3_2 _6927_ (.A(net147),
    .B(net141),
    .C(_1910_),
    .Y(_2368_));
 sg13g2_buf_2 fanout168 (.A(net188),
    .X(net168));
 sg13g2_buf_2 fanout167 (.A(net188),
    .X(net167));
 sg13g2_nand3_1 _6930_ (.B(net462),
    .C(net304),
    .A(net245),
    .Y(_2371_));
 sg13g2_o21ai_1 _6931_ (.B1(_2371_),
    .Y(_0363_),
    .A1(_2363_),
    .A2(net304));
 sg13g2_inv_1 _6932_ (.Y(_2372_),
    .A(\i_dm_csrs.progbuf_o_33_ ));
 sg13g2_nand3_1 _6933_ (.B(net459),
    .C(net298),
    .A(net225),
    .Y(_2373_));
 sg13g2_o21ai_1 _6934_ (.B1(_2373_),
    .Y(_0364_),
    .A1(_2372_),
    .A2(net298));
 sg13g2_inv_1 _6935_ (.Y(_2374_),
    .A(\i_dm_csrs.progbuf_o_34_ ));
 sg13g2_nand3_1 _6936_ (.B(net459),
    .C(net297),
    .A(net205),
    .Y(_2375_));
 sg13g2_o21ai_1 _6937_ (.B1(_2375_),
    .Y(_0365_),
    .A1(_2374_),
    .A2(net297));
 sg13g2_inv_1 _6938_ (.Y(_2376_),
    .A(\i_dm_csrs.progbuf_o_35_ ));
 sg13g2_nand3_1 _6939_ (.B(net459),
    .C(net297),
    .A(net129),
    .Y(_2377_));
 sg13g2_o21ai_1 _6940_ (.B1(_2377_),
    .Y(_0366_),
    .A1(_2376_),
    .A2(net297));
 sg13g2_inv_1 _6941_ (.Y(_2378_),
    .A(\i_dm_csrs.progbuf_o_36_ ));
 sg13g2_nand3_1 _6942_ (.B(net457),
    .C(net294),
    .A(net126),
    .Y(_2379_));
 sg13g2_o21ai_1 _6943_ (.B1(_2379_),
    .Y(_0367_),
    .A1(_2378_),
    .A2(net294));
 sg13g2_inv_1 _6944_ (.Y(_2380_),
    .A(\i_dm_csrs.progbuf_o_37_ ));
 sg13g2_nand3_1 _6945_ (.B(net461),
    .C(net303),
    .A(net124),
    .Y(_2381_));
 sg13g2_o21ai_1 _6946_ (.B1(_2381_),
    .Y(_0368_),
    .A1(_2380_),
    .A2(net303));
 sg13g2_inv_1 _6947_ (.Y(_2382_),
    .A(\i_dm_csrs.progbuf_o_38_ ));
 sg13g2_nand3_1 _6948_ (.B(net457),
    .C(net296),
    .A(net122),
    .Y(_2383_));
 sg13g2_o21ai_1 _6949_ (.B1(_2383_),
    .Y(_0369_),
    .A1(_2382_),
    .A2(net296));
 sg13g2_inv_1 _6950_ (.Y(_2384_),
    .A(\i_dm_csrs.progbuf_o_39_ ));
 sg13g2_nand3_1 _6951_ (.B(net459),
    .C(net297),
    .A(net120),
    .Y(_2385_));
 sg13g2_o21ai_1 _6952_ (.B1(_2385_),
    .Y(_0370_),
    .A1(_2384_),
    .A2(net297));
 sg13g2_inv_1 _6953_ (.Y(_2386_),
    .A(\i_dm_csrs.progbuf_o_3_ ));
 sg13g2_nand3_1 _6954_ (.B(net523),
    .C(net344),
    .A(net128),
    .Y(_2387_));
 sg13g2_o21ai_1 _6955_ (.B1(_2387_),
    .Y(_0371_),
    .A1(_2386_),
    .A2(net344));
 sg13g2_inv_1 _6956_ (.Y(_2388_),
    .A(\i_dm_csrs.progbuf_o_40_ ));
 sg13g2_buf_4 fanout166 (.X(net166),
    .A(net188));
 sg13g2_nand3_1 _6958_ (.B(net459),
    .C(net298),
    .A(net119),
    .Y(_2390_));
 sg13g2_o21ai_1 _6959_ (.B1(_2390_),
    .Y(_0372_),
    .A1(_2388_),
    .A2(net298));
 sg13g2_inv_1 _6960_ (.Y(_2391_),
    .A(\i_dm_csrs.progbuf_o_41_ ));
 sg13g2_nand3_1 _6961_ (.B(net462),
    .C(net304),
    .A(net116),
    .Y(_2392_));
 sg13g2_o21ai_1 _6962_ (.B1(_2392_),
    .Y(_0373_),
    .A1(_2391_),
    .A2(net304));
 sg13g2_inv_1 _6963_ (.Y(_2393_),
    .A(\i_dm_csrs.progbuf_o_42_ ));
 sg13g2_buf_2 fanout165 (.A(net188),
    .X(net165));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(net188));
 sg13g2_nand3_1 _6966_ (.B(net461),
    .C(net302),
    .A(net243),
    .Y(_2396_));
 sg13g2_o21ai_1 _6967_ (.B1(_2396_),
    .Y(_0374_),
    .A1(_2393_),
    .A2(net302));
 sg13g2_inv_1 _6968_ (.Y(_2397_),
    .A(\i_dm_csrs.progbuf_o_43_ ));
 sg13g2_nand3_1 _6969_ (.B(net458),
    .C(net303),
    .A(net241),
    .Y(_2398_));
 sg13g2_o21ai_1 _6970_ (.B1(_2398_),
    .Y(_0375_),
    .A1(_2397_),
    .A2(net295));
 sg13g2_inv_1 _6971_ (.Y(_2399_),
    .A(\i_dm_csrs.progbuf_o_44_ ));
 sg13g2_nand3_1 _6972_ (.B(net458),
    .C(net295),
    .A(net239),
    .Y(_2400_));
 sg13g2_o21ai_1 _6973_ (.B1(_2400_),
    .Y(_0376_),
    .A1(_2399_),
    .A2(net295));
 sg13g2_inv_1 _6974_ (.Y(_2401_),
    .A(\i_dm_csrs.progbuf_o_45_ ));
 sg13g2_nand3_1 _6975_ (.B(net457),
    .C(net293),
    .A(net800),
    .Y(_2402_));
 sg13g2_o21ai_1 _6976_ (.B1(_2402_),
    .Y(_0377_),
    .A1(_2401_),
    .A2(net293));
 sg13g2_inv_1 _6977_ (.Y(_2403_),
    .A(\i_dm_csrs.progbuf_o_46_ ));
 sg13g2_nand3_1 _6978_ (.B(net459),
    .C(net297),
    .A(net237),
    .Y(_2404_));
 sg13g2_o21ai_1 _6979_ (.B1(_2404_),
    .Y(_0378_),
    .A1(_2403_),
    .A2(net297));
 sg13g2_inv_1 _6980_ (.Y(_2405_),
    .A(\i_dm_csrs.progbuf_o_47_ ));
 sg13g2_nand3_1 _6981_ (.B(net457),
    .C(net294),
    .A(net235),
    .Y(_2406_));
 sg13g2_o21ai_1 _6982_ (.B1(_2406_),
    .Y(_0379_),
    .A1(_2405_),
    .A2(net294));
 sg13g2_inv_1 _6983_ (.Y(_2407_),
    .A(\i_dm_csrs.progbuf_o_48_ ));
 sg13g2_nand3_1 _6984_ (.B(net461),
    .C(net302),
    .A(net233),
    .Y(_2408_));
 sg13g2_o21ai_1 _6985_ (.B1(_2408_),
    .Y(_0380_),
    .A1(_2407_),
    .A2(net302));
 sg13g2_inv_1 _6986_ (.Y(_2409_),
    .A(\i_dm_csrs.progbuf_o_49_ ));
 sg13g2_nand3_1 _6987_ (.B(net461),
    .C(net301),
    .A(net231),
    .Y(_2410_));
 sg13g2_o21ai_1 _6988_ (.B1(_2410_),
    .Y(_0381_),
    .A1(_2409_),
    .A2(net301));
 sg13g2_inv_1 _6989_ (.Y(_2411_),
    .A(\i_dm_csrs.progbuf_o_4_ ));
 sg13g2_nand3_1 _6990_ (.B(net521),
    .C(net340),
    .A(net126),
    .Y(_2412_));
 sg13g2_o21ai_1 _6991_ (.B1(_2412_),
    .Y(_0382_),
    .A1(_2411_),
    .A2(net340));
 sg13g2_inv_1 _6992_ (.Y(_2413_),
    .A(\i_dm_csrs.progbuf_o_50_ ));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(net188));
 sg13g2_nand3_1 _6994_ (.B(net461),
    .C(net301),
    .A(net229),
    .Y(_2415_));
 sg13g2_o21ai_1 _6995_ (.B1(_2415_),
    .Y(_0383_),
    .A1(_2413_),
    .A2(net301));
 sg13g2_inv_1 _6996_ (.Y(_2416_),
    .A(\i_dm_csrs.progbuf_o_51_ ));
 sg13g2_nand3_1 _6997_ (.B(net461),
    .C(net302),
    .A(net227),
    .Y(_2417_));
 sg13g2_o21ai_1 _6998_ (.B1(_2417_),
    .Y(_0384_),
    .A1(_2416_),
    .A2(net301));
 sg13g2_inv_1 _6999_ (.Y(_2418_),
    .A(\i_dm_csrs.progbuf_o_52_ ));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(net188));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(net188));
 sg13g2_nand3_1 _7002_ (.B(net457),
    .C(net293),
    .A(net223),
    .Y(_2421_));
 sg13g2_o21ai_1 _7003_ (.B1(_2421_),
    .Y(_0385_),
    .A1(_2418_),
    .A2(net293));
 sg13g2_inv_1 _7004_ (.Y(_2422_),
    .A(\i_dm_csrs.progbuf_o_53_ ));
 sg13g2_nand3_1 _7005_ (.B(net457),
    .C(net293),
    .A(net221),
    .Y(_2423_));
 sg13g2_o21ai_1 _7006_ (.B1(_2423_),
    .Y(_0386_),
    .A1(_2422_),
    .A2(net293));
 sg13g2_inv_1 _7007_ (.Y(_2424_),
    .A(\i_dm_csrs.progbuf_o_54_ ));
 sg13g2_nand3_1 _7008_ (.B(net460),
    .C(net299),
    .A(net219),
    .Y(_2425_));
 sg13g2_o21ai_1 _7009_ (.B1(_2425_),
    .Y(_0387_),
    .A1(_2424_),
    .A2(net299));
 sg13g2_inv_1 _7010_ (.Y(_2426_),
    .A(\i_dm_csrs.progbuf_o_55_ ));
 sg13g2_nand3_1 _7011_ (.B(net459),
    .C(net298),
    .A(net798),
    .Y(_2427_));
 sg13g2_o21ai_1 _7012_ (.B1(_2427_),
    .Y(_0388_),
    .A1(_2426_),
    .A2(net298));
 sg13g2_inv_1 _7013_ (.Y(_2428_),
    .A(\i_dm_csrs.progbuf_o_56_ ));
 sg13g2_nand3_1 _7014_ (.B(net458),
    .C(net295),
    .A(net217),
    .Y(_2429_));
 sg13g2_o21ai_1 _7015_ (.B1(_2429_),
    .Y(_0389_),
    .A1(_2428_),
    .A2(net296));
 sg13g2_inv_1 _7016_ (.Y(_2430_),
    .A(\i_dm_csrs.progbuf_o_57_ ));
 sg13g2_nand3_1 _7017_ (.B(net461),
    .C(net303),
    .A(net215),
    .Y(_2431_));
 sg13g2_o21ai_1 _7018_ (.B1(_2431_),
    .Y(_0390_),
    .A1(_2430_),
    .A2(net303));
 sg13g2_inv_1 _7019_ (.Y(_2432_),
    .A(\i_dm_csrs.progbuf_o_58_ ));
 sg13g2_nand3_1 _7020_ (.B(net457),
    .C(net293),
    .A(net213),
    .Y(_2433_));
 sg13g2_o21ai_1 _7021_ (.B1(_2433_),
    .Y(_0391_),
    .A1(_2432_),
    .A2(net293));
 sg13g2_inv_1 _7022_ (.Y(_2434_),
    .A(\i_dm_csrs.progbuf_o_59_ ));
 sg13g2_nand3_1 _7023_ (.B(net461),
    .C(net303),
    .A(net211),
    .Y(_2435_));
 sg13g2_o21ai_1 _7024_ (.B1(_2435_),
    .Y(_0392_),
    .A1(_2434_),
    .A2(net301));
 sg13g2_inv_1 _7025_ (.Y(_2436_),
    .A(\i_dm_csrs.progbuf_o_5_ ));
 sg13g2_nand3_1 _7026_ (.B(net524),
    .C(net348),
    .A(net124),
    .Y(_2437_));
 sg13g2_o21ai_1 _7027_ (.B1(_2437_),
    .Y(_0393_),
    .A1(_2436_),
    .A2(net348));
 sg13g2_inv_1 _7028_ (.Y(_2438_),
    .A(\i_dm_csrs.progbuf_o_60_ ));
 sg13g2_nand3_1 _7029_ (.B(net462),
    .C(net301),
    .A(net209),
    .Y(_2439_));
 sg13g2_o21ai_1 _7030_ (.B1(_2439_),
    .Y(_0394_),
    .A1(_2438_),
    .A2(net301));
 sg13g2_inv_1 _7031_ (.Y(_2440_),
    .A(\i_dm_csrs.progbuf_o_61_ ));
 sg13g2_nand3_1 _7032_ (.B(net458),
    .C(net295),
    .A(net207),
    .Y(_2441_));
 sg13g2_o21ai_1 _7033_ (.B1(_2441_),
    .Y(_0395_),
    .A1(_2440_),
    .A2(net295));
 sg13g2_inv_1 _7034_ (.Y(_2442_),
    .A(\i_dm_csrs.progbuf_o_62_ ));
 sg13g2_nand3_1 _7035_ (.B(net457),
    .C(net295),
    .A(net203),
    .Y(_2443_));
 sg13g2_o21ai_1 _7036_ (.B1(_2443_),
    .Y(_0396_),
    .A1(_2442_),
    .A2(net295));
 sg13g2_inv_1 _7037_ (.Y(_2444_),
    .A(\i_dm_csrs.progbuf_o_63_ ));
 sg13g2_nand3_1 _7038_ (.B(net459),
    .C(net298),
    .A(net201),
    .Y(_2445_));
 sg13g2_o21ai_1 _7039_ (.B1(_2445_),
    .Y(_0397_),
    .A1(_2444_),
    .A2(net298));
 sg13g2_inv_1 _7040_ (.Y(_2446_),
    .A(\i_dm_csrs.progbuf_o_64_ ));
 sg13g2_nor3_1 _7041_ (.A(net176),
    .B(net607),
    .C(net141),
    .Y(_2447_));
 sg13g2_nor2_1 _7042_ (.A(net639),
    .B(_2447_),
    .Y(_2448_));
 sg13g2_nor2_2 _7043_ (.A(_1901_),
    .B(_2448_),
    .Y(_2449_));
 sg13g2_buf_2 fanout160 (.A(dmi_req_i_35_),
    .X(net160));
 sg13g2_nor2_2 _7045_ (.A(_1905_),
    .B(_1911_),
    .Y(_2451_));
 sg13g2_buf_4 fanout159 (.X(net159),
    .A(net160));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(net160));
 sg13g2_nand3_1 _7048_ (.B(net434),
    .C(net292),
    .A(net245),
    .Y(_2454_));
 sg13g2_o21ai_1 _7049_ (.B1(_2454_),
    .Y(_0398_),
    .A1(_2446_),
    .A2(net292));
 sg13g2_inv_1 _7050_ (.Y(_2455_),
    .A(\i_dm_csrs.progbuf_o_65_ ));
 sg13g2_nand3_1 _7051_ (.B(net431),
    .C(net286),
    .A(net225),
    .Y(_2456_));
 sg13g2_o21ai_1 _7052_ (.B1(_2456_),
    .Y(_0399_),
    .A1(_2455_),
    .A2(net286));
 sg13g2_inv_1 _7053_ (.Y(_2457_),
    .A(\i_dm_csrs.progbuf_o_66_ ));
 sg13g2_nand3_1 _7054_ (.B(net431),
    .C(net287),
    .A(net205),
    .Y(_2458_));
 sg13g2_o21ai_1 _7055_ (.B1(_2458_),
    .Y(_0400_),
    .A1(_2457_),
    .A2(net287));
 sg13g2_inv_1 _7056_ (.Y(_2459_),
    .A(\i_dm_csrs.progbuf_o_67_ ));
 sg13g2_nand3_1 _7057_ (.B(net432),
    .C(net288),
    .A(net128),
    .Y(_2460_));
 sg13g2_o21ai_1 _7058_ (.B1(_2460_),
    .Y(_0401_),
    .A1(_2459_),
    .A2(net288));
 sg13g2_inv_1 _7059_ (.Y(_2461_),
    .A(\i_dm_csrs.progbuf_o_68_ ));
 sg13g2_nand3_1 _7060_ (.B(net430),
    .C(net283),
    .A(net126),
    .Y(_2462_));
 sg13g2_o21ai_1 _7061_ (.B1(_2462_),
    .Y(_0402_),
    .A1(_2461_),
    .A2(net283));
 sg13g2_inv_1 _7062_ (.Y(_2463_),
    .A(\i_dm_csrs.progbuf_o_69_ ));
 sg13g2_nand3_1 _7063_ (.B(net433),
    .C(net291),
    .A(net124),
    .Y(_2464_));
 sg13g2_o21ai_1 _7064_ (.B1(_2464_),
    .Y(_0403_),
    .A1(_2463_),
    .A2(net291));
 sg13g2_inv_1 _7065_ (.Y(_2465_),
    .A(\i_dm_csrs.progbuf_o_6_ ));
 sg13g2_nand3_1 _7066_ (.B(net523),
    .C(net344),
    .A(net122),
    .Y(_2466_));
 sg13g2_o21ai_1 _7067_ (.B1(_2466_),
    .Y(_0404_),
    .A1(_2465_),
    .A2(net344));
 sg13g2_inv_1 _7068_ (.Y(_2467_),
    .A(\i_dm_csrs.progbuf_o_70_ ));
 sg13g2_nand3_1 _7069_ (.B(net431),
    .C(net288),
    .A(net122),
    .Y(_2468_));
 sg13g2_o21ai_1 _7070_ (.B1(_2468_),
    .Y(_0405_),
    .A1(_2467_),
    .A2(net288));
 sg13g2_inv_1 _7071_ (.Y(_2469_),
    .A(\i_dm_csrs.progbuf_o_71_ ));
 sg13g2_nand3_1 _7072_ (.B(net431),
    .C(net287),
    .A(net120),
    .Y(_2470_));
 sg13g2_o21ai_1 _7073_ (.B1(_2470_),
    .Y(_0406_),
    .A1(_2469_),
    .A2(net287));
 sg13g2_inv_1 _7074_ (.Y(_2471_),
    .A(\i_dm_csrs.progbuf_o_72_ ));
 sg13g2_buf_2 fanout157 (.A(net159),
    .X(net157));
 sg13g2_nand3_1 _7076_ (.B(net431),
    .C(net287),
    .A(net118),
    .Y(_2473_));
 sg13g2_o21ai_1 _7077_ (.B1(_2473_),
    .Y(_0407_),
    .A1(_2471_),
    .A2(net287));
 sg13g2_inv_1 _7078_ (.Y(_2474_),
    .A(\i_dm_csrs.progbuf_o_73_ ));
 sg13g2_nand3_1 _7079_ (.B(net434),
    .C(net292),
    .A(net116),
    .Y(_2475_));
 sg13g2_o21ai_1 _7080_ (.B1(_2475_),
    .Y(_0408_),
    .A1(_2474_),
    .A2(net292));
 sg13g2_inv_1 _7081_ (.Y(_2476_),
    .A(\i_dm_csrs.progbuf_o_74_ ));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net159));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(net159));
 sg13g2_nand3_1 _7084_ (.B(net433),
    .C(net290),
    .A(net243),
    .Y(_2479_));
 sg13g2_o21ai_1 _7085_ (.B1(_2479_),
    .Y(_0409_),
    .A1(_2476_),
    .A2(net290));
 sg13g2_inv_1 _7086_ (.Y(_2480_),
    .A(\i_dm_csrs.progbuf_o_75_ ));
 sg13g2_nand3_1 _7087_ (.B(net433),
    .C(net291),
    .A(net241),
    .Y(_2481_));
 sg13g2_o21ai_1 _7088_ (.B1(_2481_),
    .Y(_0410_),
    .A1(_2480_),
    .A2(net291));
 sg13g2_inv_1 _7089_ (.Y(_2482_),
    .A(\i_dm_csrs.progbuf_o_76_ ));
 sg13g2_nand3_1 _7090_ (.B(net430),
    .C(net284),
    .A(net239),
    .Y(_2483_));
 sg13g2_o21ai_1 _7091_ (.B1(_2483_),
    .Y(_0411_),
    .A1(_2482_),
    .A2(net284));
 sg13g2_inv_1 _7092_ (.Y(_2484_),
    .A(\i_dm_csrs.progbuf_o_77_ ));
 sg13g2_nand3_1 _7093_ (.B(net430),
    .C(net285),
    .A(net800),
    .Y(_2485_));
 sg13g2_o21ai_1 _7094_ (.B1(_2485_),
    .Y(_0412_),
    .A1(_2484_),
    .A2(net285));
 sg13g2_inv_1 _7095_ (.Y(_2486_),
    .A(\i_dm_csrs.progbuf_o_78_ ));
 sg13g2_nand3_1 _7096_ (.B(net431),
    .C(net286),
    .A(net237),
    .Y(_2487_));
 sg13g2_o21ai_1 _7097_ (.B1(_2487_),
    .Y(_0413_),
    .A1(_2486_),
    .A2(net286));
 sg13g2_inv_1 _7098_ (.Y(_2488_),
    .A(\i_dm_csrs.progbuf_o_79_ ));
 sg13g2_nand3_1 _7099_ (.B(net430),
    .C(net283),
    .A(net235),
    .Y(_2489_));
 sg13g2_o21ai_1 _7100_ (.B1(_2489_),
    .Y(_0414_),
    .A1(_2488_),
    .A2(net285));
 sg13g2_inv_1 _7101_ (.Y(_2490_),
    .A(\i_dm_csrs.progbuf_o_7_ ));
 sg13g2_nand3_1 _7102_ (.B(net522),
    .C(net343),
    .A(net120),
    .Y(_2491_));
 sg13g2_o21ai_1 _7103_ (.B1(_2491_),
    .Y(_0415_),
    .A1(_2490_),
    .A2(net343));
 sg13g2_inv_1 _7104_ (.Y(_2492_),
    .A(\i_dm_csrs.progbuf_o_80_ ));
 sg13g2_nand3_1 _7105_ (.B(net433),
    .C(net290),
    .A(net233),
    .Y(_2493_));
 sg13g2_o21ai_1 _7106_ (.B1(_2493_),
    .Y(_0416_),
    .A1(_2492_),
    .A2(net290));
 sg13g2_inv_1 _7107_ (.Y(_2494_),
    .A(\i_dm_csrs.progbuf_o_81_ ));
 sg13g2_nand3_1 _7108_ (.B(net433),
    .C(net289),
    .A(net231),
    .Y(_2495_));
 sg13g2_o21ai_1 _7109_ (.B1(_2495_),
    .Y(_0417_),
    .A1(_2494_),
    .A2(net289));
 sg13g2_inv_1 _7110_ (.Y(_2496_),
    .A(\i_dm_csrs.progbuf_o_82_ ));
 sg13g2_buf_8 fanout154 (.A(net158),
    .X(net154));
 sg13g2_nand3_1 _7112_ (.B(net433),
    .C(net289),
    .A(net229),
    .Y(_2498_));
 sg13g2_o21ai_1 _7113_ (.B1(_2498_),
    .Y(_0418_),
    .A1(_2496_),
    .A2(net289));
 sg13g2_inv_1 _7114_ (.Y(_2499_),
    .A(\i_dm_csrs.progbuf_o_83_ ));
 sg13g2_nand3_1 _7115_ (.B(net433),
    .C(net290),
    .A(net227),
    .Y(_2500_));
 sg13g2_o21ai_1 _7116_ (.B1(_2500_),
    .Y(_0419_),
    .A1(_2499_),
    .A2(net290));
 sg13g2_inv_1 _7117_ (.Y(_2501_),
    .A(\i_dm_csrs.progbuf_o_84_ ));
 sg13g2_buf_8 fanout153 (.A(net158),
    .X(net153));
 sg13g2_buf_8 fanout152 (.A(net158),
    .X(net152));
 sg13g2_nand3_1 _7120_ (.B(net430),
    .C(net283),
    .A(net223),
    .Y(_2504_));
 sg13g2_o21ai_1 _7121_ (.B1(_2504_),
    .Y(_0420_),
    .A1(_2501_),
    .A2(net283));
 sg13g2_inv_1 _7122_ (.Y(_2505_),
    .A(\i_dm_csrs.progbuf_o_85_ ));
 sg13g2_nand3_1 _7123_ (.B(net430),
    .C(net283),
    .A(net221),
    .Y(_2506_));
 sg13g2_o21ai_1 _7124_ (.B1(_2506_),
    .Y(_0421_),
    .A1(_2505_),
    .A2(net284));
 sg13g2_inv_1 _7125_ (.Y(_2507_),
    .A(\i_dm_csrs.progbuf_o_86_ ));
 sg13g2_nand3_1 _7126_ (.B(net432),
    .C(net288),
    .A(net219),
    .Y(_2508_));
 sg13g2_o21ai_1 _7127_ (.B1(_2508_),
    .Y(_0422_),
    .A1(_2507_),
    .A2(net288));
 sg13g2_inv_1 _7128_ (.Y(_2509_),
    .A(\i_dm_csrs.progbuf_o_87_ ));
 sg13g2_nand3_1 _7129_ (.B(net431),
    .C(net286),
    .A(net798),
    .Y(_2510_));
 sg13g2_o21ai_1 _7130_ (.B1(_2510_),
    .Y(_0423_),
    .A1(_2509_),
    .A2(net286));
 sg13g2_inv_1 _7131_ (.Y(_2511_),
    .A(\i_dm_csrs.progbuf_o_88_ ));
 sg13g2_nand3_1 _7132_ (.B(net432),
    .C(net284),
    .A(net217),
    .Y(_2512_));
 sg13g2_o21ai_1 _7133_ (.B1(_2512_),
    .Y(_0424_),
    .A1(_2511_),
    .A2(net284));
 sg13g2_inv_1 _7134_ (.Y(_2513_),
    .A(\i_dm_csrs.progbuf_o_89_ ));
 sg13g2_nand3_1 _7135_ (.B(net433),
    .C(net291),
    .A(net215),
    .Y(_2514_));
 sg13g2_o21ai_1 _7136_ (.B1(_2514_),
    .Y(_0425_),
    .A1(_2513_),
    .A2(net291));
 sg13g2_inv_1 _7137_ (.Y(_2515_),
    .A(\i_dm_csrs.progbuf_o_8_ ));
 sg13g2_nand3_1 _7138_ (.B(net522),
    .C(net342),
    .A(net118),
    .Y(_2516_));
 sg13g2_o21ai_1 _7139_ (.B1(_2516_),
    .Y(_0426_),
    .A1(_2515_),
    .A2(net342));
 sg13g2_inv_1 _7140_ (.Y(_2517_),
    .A(\i_dm_csrs.progbuf_o_90_ ));
 sg13g2_nand3_1 _7141_ (.B(net430),
    .C(net283),
    .A(net213),
    .Y(_2518_));
 sg13g2_o21ai_1 _7142_ (.B1(_2518_),
    .Y(_0427_),
    .A1(_2517_),
    .A2(net283));
 sg13g2_inv_1 _7143_ (.Y(_2519_),
    .A(\i_dm_csrs.progbuf_o_91_ ));
 sg13g2_nand3_1 _7144_ (.B(net434),
    .C(net289),
    .A(net211),
    .Y(_2520_));
 sg13g2_o21ai_1 _7145_ (.B1(_2520_),
    .Y(_0428_),
    .A1(_2519_),
    .A2(net289));
 sg13g2_inv_1 _7146_ (.Y(_2521_),
    .A(\i_dm_csrs.progbuf_o_92_ ));
 sg13g2_nand3_1 _7147_ (.B(net434),
    .C(net289),
    .A(net209),
    .Y(_2522_));
 sg13g2_o21ai_1 _7148_ (.B1(_2522_),
    .Y(_0429_),
    .A1(_2521_),
    .A2(net289));
 sg13g2_inv_1 _7149_ (.Y(_2523_),
    .A(\i_dm_csrs.progbuf_o_93_ ));
 sg13g2_nand3_1 _7150_ (.B(net432),
    .C(net284),
    .A(net207),
    .Y(_2524_));
 sg13g2_o21ai_1 _7151_ (.B1(_2524_),
    .Y(_0430_),
    .A1(_2523_),
    .A2(net284));
 sg13g2_inv_1 _7152_ (.Y(_2525_),
    .A(\i_dm_csrs.progbuf_o_94_ ));
 sg13g2_nand3_1 _7153_ (.B(net430),
    .C(net284),
    .A(net203),
    .Y(_2526_));
 sg13g2_o21ai_1 _7154_ (.B1(_2526_),
    .Y(_0431_),
    .A1(_2525_),
    .A2(net285));
 sg13g2_inv_1 _7155_ (.Y(_2527_),
    .A(\i_dm_csrs.progbuf_o_95_ ));
 sg13g2_nand3_1 _7156_ (.B(net431),
    .C(net286),
    .A(net201),
    .Y(_2528_));
 sg13g2_o21ai_1 _7157_ (.B1(_2528_),
    .Y(_0432_),
    .A1(_2527_),
    .A2(net286));
 sg13g2_nand2_1 _7158_ (.Y(_2529_),
    .A(net245),
    .B(net439));
 sg13g2_nand2_2 _7159_ (.Y(_2530_),
    .A(\i_dm_csrs.progbuf_o_96_ ),
    .B(net272));
 sg13g2_o21ai_1 _7160_ (.B1(_2530_),
    .Y(_0433_),
    .A1(net272),
    .A2(_2529_));
 sg13g2_nand2_1 _7161_ (.Y(_2531_),
    .A(net225),
    .B(net436));
 sg13g2_nand2_2 _7162_ (.Y(_2532_),
    .A(\i_dm_csrs.progbuf_o_97_ ),
    .B(net266));
 sg13g2_o21ai_1 _7163_ (.B1(_2532_),
    .Y(_0434_),
    .A1(net266),
    .A2(_2531_));
 sg13g2_nand2_1 _7164_ (.Y(_2533_),
    .A(net205),
    .B(net436));
 sg13g2_nand2_2 _7165_ (.Y(_2534_),
    .A(\i_dm_csrs.progbuf_o_98_ ),
    .B(net265));
 sg13g2_o21ai_1 _7166_ (.B1(_2534_),
    .Y(_0435_),
    .A1(net265),
    .A2(_2533_));
 sg13g2_nand2_1 _7167_ (.Y(_2535_),
    .A(net128),
    .B(net436));
 sg13g2_nand2_2 _7168_ (.Y(_2536_),
    .A(\i_dm_csrs.progbuf_o_99_ ),
    .B(net265));
 sg13g2_o21ai_1 _7169_ (.B1(_2536_),
    .Y(_0436_),
    .A1(net265),
    .A2(_2535_));
 sg13g2_inv_1 _7170_ (.Y(_2537_),
    .A(\i_dm_csrs.progbuf_o_9_ ));
 sg13g2_nand3_1 _7171_ (.B(net525),
    .C(net349),
    .A(net116),
    .Y(_2538_));
 sg13g2_o21ai_1 _7172_ (.B1(_2538_),
    .Y(_0437_),
    .A1(_2537_),
    .A2(net349));
 sg13g2_buf_8 fanout151 (.A(net158),
    .X(net151));
 sg13g2_nand4_1 _7174_ (.B(_1148_),
    .C(net42),
    .A(_0599_),
    .Y(_2540_),
    .D(net41));
 sg13g2_and2_2 _7175_ (.A(_0893_),
    .B(_2540_),
    .X(_2541_));
 sg13g2_buf_8 fanout150 (.A(net158),
    .X(net150));
 sg13g2_a21oi_1 _7177_ (.A1(_1148_),
    .A2(net41),
    .Y(_2543_),
    .B1(net640));
 sg13g2_nand3_1 _7178_ (.B(net42),
    .C(net525),
    .A(_0599_),
    .Y(_2544_));
 sg13g2_nor2_2 _7179_ (.A(_2543_),
    .B(_2544_),
    .Y(_2545_));
 sg13g2_and2_2 _7180_ (.A(net41),
    .B(_2545_),
    .X(_2546_));
 sg13g2_a22oi_1 _7181_ (.Y(_2547_),
    .B1(_2546_),
    .B2(net231),
    .A2(net428),
    .A1(net633));
 sg13g2_inv_1 _7182_ (.Y(_0438_),
    .A(_2547_));
 sg13g2_nand3_1 _7183_ (.B(_0602_),
    .C(net530),
    .A(_0599_),
    .Y(_2548_));
 sg13g2_nand2_1 _7184_ (.Y(_2549_),
    .A(net229),
    .B(net41));
 sg13g2_o21ai_1 _7185_ (.B1(net95),
    .Y(_2550_),
    .A1(_2548_),
    .A2(_2549_));
 sg13g2_nand2_2 _7186_ (.Y(_2551_),
    .A(_0001_),
    .B(net428));
 sg13g2_o21ai_1 _7187_ (.B1(_2551_),
    .Y(_0439_),
    .A1(net428),
    .A2(_2550_));
 sg13g2_a22oi_1 _7188_ (.Y(_2552_),
    .B1(_2546_),
    .B2(net227),
    .A2(net428),
    .A1(net628));
 sg13g2_inv_1 _7189_ (.Y(_0440_),
    .A(_2552_));
 sg13g2_nor4_2 _7190_ (.A(\i_dm_csrs.sbcs_q_22_ ),
    .B(_0614_),
    .C(_1279_),
    .Y(_2553_),
    .D(_1315_));
 sg13g2_nand2_2 _7191_ (.Y(_2554_),
    .A(_2364_),
    .B(_2553_));
 sg13g2_buf_8 fanout149 (.A(net158),
    .X(net149));
 sg13g2_buf_8 fanout148 (.A(net158),
    .X(net148));
 sg13g2_inv_1 _7194_ (.Y(_2557_),
    .A(net77));
 sg13g2_nand2_2 _7195_ (.Y(_2558_),
    .A(_1517_),
    .B(_1536_));
 sg13g2_nor3_1 _7196_ (.A(\i_dm_sba.state_q_2_ ),
    .B(\i_dm_sba.state_q_0__$_NOT__A_Y ),
    .C(\i_dm_sba.state_q_1__$_NOT__A_Y ),
    .Y(_2559_));
 sg13g2_nor3_1 _7197_ (.A(\i_dm_csrs.sbbusy_i_$_OR__Y_A_$_OR__A_B ),
    .B(\i_dm_sba.state_q_0_ ),
    .C(\i_dm_sba.state_q_1_ ),
    .Y(_2560_));
 sg13g2_nor2_1 _7198_ (.A(_2559_),
    .B(_2560_),
    .Y(_2561_));
 sg13g2_buf_4 fanout147 (.X(net147),
    .A(net158));
 sg13g2_nor2b_2 _7200_ (.A(_2561_),
    .B_N(net795),
    .Y(_2563_));
 sg13g2_nand2_1 _7201_ (.Y(_2564_),
    .A(\i_dm_csrs.sbautoincrement_o ),
    .B(_2563_));
 sg13g2_nor3_1 _7202_ (.A(net546),
    .B(_2558_),
    .C(net427),
    .Y(_2565_));
 sg13g2_xnor2_1 _7203_ (.Y(_2566_),
    .A(master_add_o_0_),
    .B(_2565_));
 sg13g2_buf_8 fanout146 (.A(net159),
    .X(net146));
 sg13g2_nand2_2 _7205_ (.Y(_2568_),
    .A(_2566_),
    .B(net404));
 sg13g2_o21ai_1 _7206_ (.B1(_2568_),
    .Y(_2569_),
    .A1(net245),
    .A2(net404));
 sg13g2_nor2_1 _7207_ (.A(net598),
    .B(_2569_),
    .Y(\master_add_o[0]_reg_D ));
 sg13g2_inv_1 _7208_ (.Y(_2570_),
    .A(master_add_o_6_));
 sg13g2_a21oi_1 _7209_ (.A1(net48),
    .A2(net79),
    .Y(_2571_),
    .B1(master_add_o_5_));
 sg13g2_nand2b_1 _7210_ (.Y(_2572_),
    .B(net631),
    .A_N(_2571_));
 sg13g2_and2_1 _7211_ (.A(net48),
    .B(master_add_o_5_),
    .X(_2573_));
 sg13g2_nand2_1 _7212_ (.Y(_2574_),
    .A(net78),
    .B(_2573_));
 sg13g2_nand2b_2 _7213_ (.Y(_2575_),
    .B(\i_dm_csrs.sbaccess_o_2_ ),
    .A_N(net629));
 sg13g2_a221oi_1 _7214_ (.B2(_2574_),
    .C1(_2575_),
    .B1(_2572_),
    .A1(_2570_),
    .Y(_2576_),
    .A2(net546));
 sg13g2_buf_8 fanout145 (.A(net159),
    .X(net145));
 sg13g2_a21o_1 _7216_ (.A2(\i_dm_sba.sbaccess_mask_3__$_AND__B_A_$_AND__Y_A ),
    .A1(master_add_o_6_),
    .B1(master_add_o_7_),
    .X(_2578_));
 sg13g2_o21ai_1 _7217_ (.B1(net631),
    .Y(_2579_),
    .A1(_2576_),
    .A2(_2578_));
 sg13g2_and2_1 _7218_ (.A(master_add_o_6_),
    .B(master_add_o_7_),
    .X(_2580_));
 sg13g2_nand2_1 _7219_ (.Y(_2581_),
    .A(net78),
    .B(_2580_));
 sg13g2_nand2_1 _7220_ (.Y(_2582_),
    .A(net629),
    .B(\i_dm_csrs.sbaccess_o_2_ ));
 sg13g2_a21o_1 _7221_ (.A2(_2581_),
    .A1(_2579_),
    .B1(_2582_),
    .X(_2583_));
 sg13g2_o21ai_1 _7222_ (.B1(master_add_o_3_),
    .Y(_2584_),
    .A1(net50),
    .A2(net77));
 sg13g2_nand2b_1 _7223_ (.Y(_2585_),
    .B(net630),
    .A_N(net628));
 sg13g2_nand2_2 _7224_ (.Y(_2586_),
    .A(net50),
    .B(master_add_o_3_));
 sg13g2_nor3_2 _7225_ (.A(net50),
    .B(master_add_o_3_),
    .C(net79),
    .Y(_2587_));
 sg13g2_a221oi_1 _7226_ (.B2(_2586_),
    .C1(_2587_),
    .B1(_2585_),
    .A1(_1496_),
    .Y(_2588_),
    .A2(_2584_));
 sg13g2_nor2_2 _7227_ (.A(net629),
    .B(\i_dm_csrs.sbaccess_o_2_ ),
    .Y(_2589_));
 sg13g2_a21oi_1 _7228_ (.A1(net51),
    .A2(net79),
    .Y(_2590_),
    .B1(master_add_o_1_));
 sg13g2_nand3_1 _7229_ (.B(master_add_o_1_),
    .C(net77),
    .A(net51),
    .Y(_2591_));
 sg13g2_o21ai_1 _7230_ (.B1(_2591_),
    .Y(_2592_),
    .A1(_1496_),
    .A2(_2590_));
 sg13g2_a22oi_1 _7231_ (.Y(_2593_),
    .B1(net77),
    .B2(net50),
    .A2(master_add_o_3_),
    .A1(net631));
 sg13g2_nor2_1 _7232_ (.A(_2585_),
    .B(_2593_),
    .Y(_2594_));
 sg13g2_a21o_1 _7233_ (.A2(_2592_),
    .A1(_2589_),
    .B1(_2594_),
    .X(_2595_));
 sg13g2_and2_1 _7234_ (.A(_2588_),
    .B(_2595_),
    .X(_2596_));
 sg13g2_xor2_1 _7235_ (.B(net79),
    .A(net48),
    .X(_2597_));
 sg13g2_nor2b_1 _7236_ (.A(master_add_o_5_),
    .B_N(net631),
    .Y(_2598_));
 sg13g2_nor2b_1 _7237_ (.A(net631),
    .B_N(net77),
    .Y(_2599_));
 sg13g2_nor2b_1 _7238_ (.A(master_add_o_4_),
    .B_N(master_add_o_5_),
    .Y(_2600_));
 sg13g2_a22oi_1 _7239_ (.Y(_2601_),
    .B1(_2599_),
    .B2(_2600_),
    .A2(_2598_),
    .A1(_2597_));
 sg13g2_nor2_1 _7240_ (.A(net631),
    .B(net77),
    .Y(_2602_));
 sg13g2_o21ai_1 _7241_ (.B1(_2573_),
    .Y(_2603_),
    .A1(_2575_),
    .A2(_2602_));
 sg13g2_o21ai_1 _7242_ (.B1(_2603_),
    .Y(_2604_),
    .A1(_2575_),
    .A2(_2601_));
 sg13g2_nand2_1 _7243_ (.Y(_2605_),
    .A(master_add_o_6_),
    .B(master_add_o_7_));
 sg13g2_nor2_1 _7244_ (.A(net631),
    .B(master_add_o_7_),
    .Y(_2606_));
 sg13g2_a221oi_1 _7245_ (.B2(_2605_),
    .C1(_2606_),
    .B1(_2582_),
    .A1(_2570_),
    .Y(_2607_),
    .A2(net546));
 sg13g2_and2_1 _7246_ (.A(_2604_),
    .B(_2607_),
    .X(_2608_));
 sg13g2_a21oi_1 _7247_ (.A1(_2572_),
    .A2(_2574_),
    .Y(_2609_),
    .B1(_2575_));
 sg13g2_a22oi_1 _7248_ (.Y(_2610_),
    .B1(_2609_),
    .B2(_2580_),
    .A2(_2608_),
    .A1(_2596_));
 sg13g2_a21oi_1 _7249_ (.A1(_2583_),
    .A2(_2610_),
    .Y(_2611_),
    .B1(net427));
 sg13g2_buf_4 fanout144 (.X(net144),
    .A(net159));
 sg13g2_nand3_1 _7251_ (.B(master_add_o_9_),
    .C(net279),
    .A(master_add_o_8_),
    .Y(_2613_));
 sg13g2_xor2_1 _7252_ (.B(_2613_),
    .A(master_add_o_10_),
    .X(_2614_));
 sg13g2_buf_2 fanout143 (.A(net159),
    .X(net143));
 sg13g2_nor2_1 _7254_ (.A(net243),
    .B(net394),
    .Y(_2616_));
 sg13g2_a21oi_1 _7255_ (.A1(net396),
    .A2(_2614_),
    .Y(_2617_),
    .B1(_2616_));
 sg13g2_and2_1 _7256_ (.A(net81),
    .B(_2617_),
    .X(\master_add_o[10]_reg_D ));
 sg13g2_buf_2 fanout142 (.A(dmi_req_i_36_),
    .X(net142));
 sg13g2_and3_1 _7258_ (.X(_2619_),
    .A(master_add_o_8_),
    .B(master_add_o_9_),
    .C(master_add_o_10_));
 sg13g2_nand2_2 _7259_ (.Y(_2620_),
    .A(net279),
    .B(_2619_));
 sg13g2_xor2_1 _7260_ (.B(_2620_),
    .A(master_add_o_11_),
    .X(_2621_));
 sg13g2_nor2_1 _7261_ (.A(net241),
    .B(net394),
    .Y(_2622_));
 sg13g2_a21oi_1 _7262_ (.A1(net394),
    .A2(_2621_),
    .Y(_2623_),
    .B1(_2622_));
 sg13g2_and2_1 _7263_ (.A(net81),
    .B(_2623_),
    .X(\master_add_o[11]_reg_D ));
 sg13g2_nand3_1 _7264_ (.B(net279),
    .C(_2619_),
    .A(master_add_o_11_),
    .Y(_2624_));
 sg13g2_xor2_1 _7265_ (.B(_2624_),
    .A(master_add_o_12_),
    .X(_2625_));
 sg13g2_nor2_1 _7266_ (.A(net239),
    .B(net394),
    .Y(_2626_));
 sg13g2_a21oi_1 _7267_ (.A1(net396),
    .A2(_2625_),
    .Y(_2627_),
    .B1(_2626_));
 sg13g2_and2_1 _7268_ (.A(net81),
    .B(_2627_),
    .X(\master_add_o[12]_reg_D ));
 sg13g2_and3_1 _7269_ (.X(_2628_),
    .A(master_add_o_11_),
    .B(master_add_o_12_),
    .C(_2619_));
 sg13g2_nand2_2 _7270_ (.Y(_2629_),
    .A(net279),
    .B(_2628_));
 sg13g2_xor2_1 _7271_ (.B(_2629_),
    .A(master_add_o_13_),
    .X(_2630_));
 sg13g2_nor2_1 _7272_ (.A(net802),
    .B(net396),
    .Y(_2631_));
 sg13g2_a21oi_1 _7273_ (.A1(net396),
    .A2(_2630_),
    .Y(_2632_),
    .B1(_2631_));
 sg13g2_and2_1 _7274_ (.A(net81),
    .B(_2632_),
    .X(\master_add_o[13]_reg_D ));
 sg13g2_nand3_1 _7275_ (.B(net279),
    .C(_2628_),
    .A(master_add_o_13_),
    .Y(_2633_));
 sg13g2_xor2_1 _7276_ (.B(_2633_),
    .A(master_add_o_14_),
    .X(_2634_));
 sg13g2_nor2_1 _7277_ (.A(net237),
    .B(net396),
    .Y(_2635_));
 sg13g2_a21oi_1 _7278_ (.A1(net396),
    .A2(_2634_),
    .Y(_2636_),
    .B1(_2635_));
 sg13g2_and2_1 _7279_ (.A(net81),
    .B(_2636_),
    .X(\master_add_o[14]_reg_D ));
 sg13g2_and3_2 _7280_ (.X(_2637_),
    .A(master_add_o_13_),
    .B(master_add_o_14_),
    .C(_2628_));
 sg13g2_nand2_2 _7281_ (.Y(_2638_),
    .A(net279),
    .B(_2637_));
 sg13g2_xor2_1 _7282_ (.B(_2638_),
    .A(master_add_o_15_),
    .X(_2639_));
 sg13g2_nor2_1 _7283_ (.A(net235),
    .B(net394),
    .Y(_2640_));
 sg13g2_a21oi_1 _7284_ (.A1(net394),
    .A2(_2639_),
    .Y(_2641_),
    .B1(_2640_));
 sg13g2_and2_1 _7285_ (.A(net81),
    .B(_2641_),
    .X(\master_add_o[15]_reg_D ));
 sg13g2_buf_2 fanout141 (.A(net797),
    .X(net141));
 sg13g2_buf_4 fanout140 (.X(net140),
    .A(net797));
 sg13g2_nand3_1 _7288_ (.B(net279),
    .C(_2637_),
    .A(master_add_o_15_),
    .Y(_2644_));
 sg13g2_xor2_1 _7289_ (.B(_2644_),
    .A(master_add_o_16_),
    .X(_2645_));
 sg13g2_nor2_1 _7290_ (.A(net233),
    .B(net394),
    .Y(_2646_));
 sg13g2_a21oi_1 _7291_ (.A1(net395),
    .A2(_2645_),
    .Y(_2647_),
    .B1(_2646_));
 sg13g2_and2_1 _7292_ (.A(net83),
    .B(_2647_),
    .X(\master_add_o[16]_reg_D ));
 sg13g2_and2_1 _7293_ (.A(master_add_o_15_),
    .B(master_add_o_16_),
    .X(_2648_));
 sg13g2_nand3_1 _7294_ (.B(_2637_),
    .C(_2648_),
    .A(net279),
    .Y(_2649_));
 sg13g2_xor2_1 _7295_ (.B(_2649_),
    .A(master_add_o_17_),
    .X(_2650_));
 sg13g2_nor2_1 _7296_ (.A(net231),
    .B(net394),
    .Y(_2651_));
 sg13g2_a21oi_1 _7297_ (.A1(net395),
    .A2(_2650_),
    .Y(_2652_),
    .B1(_2651_));
 sg13g2_and2_1 _7298_ (.A(net83),
    .B(_2652_),
    .X(\master_add_o[17]_reg_D ));
 sg13g2_nand4_1 _7299_ (.B(net282),
    .C(_2637_),
    .A(master_add_o_17_),
    .Y(_2653_),
    .D(_2648_));
 sg13g2_xor2_1 _7300_ (.B(_2653_),
    .A(master_add_o_18_),
    .X(_2654_));
 sg13g2_nor2_1 _7301_ (.A(net229),
    .B(net395),
    .Y(_2655_));
 sg13g2_a21oi_1 _7302_ (.A1(net395),
    .A2(_2654_),
    .Y(_2656_),
    .B1(_2655_));
 sg13g2_and2_1 _7303_ (.A(net82),
    .B(_2656_),
    .X(\master_add_o[18]_reg_D ));
 sg13g2_and4_1 _7304_ (.A(master_add_o_17_),
    .B(master_add_o_18_),
    .C(_2637_),
    .D(_2648_),
    .X(_2657_));
 sg13g2_buf_8 fanout139 (.A(net797),
    .X(net139));
 sg13g2_nand2_2 _7306_ (.Y(_2659_),
    .A(net281),
    .B(net456));
 sg13g2_xor2_1 _7307_ (.B(_2659_),
    .A(master_add_o_19_),
    .X(_2660_));
 sg13g2_nor2_1 _7308_ (.A(net227),
    .B(net401),
    .Y(_2661_));
 sg13g2_a21oi_1 _7309_ (.A1(net401),
    .A2(_2660_),
    .Y(_2662_),
    .B1(_2661_));
 sg13g2_and2_1 _7310_ (.A(net82),
    .B(_2662_),
    .X(\master_add_o[19]_reg_D ));
 sg13g2_nand2_2 _7311_ (.Y(_2663_),
    .A(net51),
    .B(net77));
 sg13g2_xnor2_1 _7312_ (.Y(_2664_),
    .A(_1496_),
    .B(_2663_));
 sg13g2_nor3_2 _7313_ (.A(_2558_),
    .B(net427),
    .C(_2664_),
    .Y(_2665_));
 sg13g2_xnor2_1 _7314_ (.Y(_2666_),
    .A(master_add_o_1_),
    .B(_2665_));
 sg13g2_nand2_2 _7315_ (.Y(_2667_),
    .A(net404),
    .B(_2666_));
 sg13g2_o21ai_1 _7316_ (.B1(_2667_),
    .Y(_2668_),
    .A1(net225),
    .A2(net404));
 sg13g2_nor2_1 _7317_ (.A(net598),
    .B(_2668_),
    .Y(\master_add_o[1]_reg_D ));
 sg13g2_nand3_1 _7318_ (.B(net280),
    .C(net456),
    .A(master_add_o_19_),
    .Y(_2669_));
 sg13g2_xor2_1 _7319_ (.B(_2669_),
    .A(master_add_o_20_),
    .X(_2670_));
 sg13g2_buf_8 fanout138 (.A(net797),
    .X(net138));
 sg13g2_nor2_1 _7321_ (.A(net223),
    .B(net399),
    .Y(_2672_));
 sg13g2_a21oi_1 _7322_ (.A1(net400),
    .A2(_2670_),
    .Y(_2673_),
    .B1(_2672_));
 sg13g2_and2_1 _7323_ (.A(net82),
    .B(_2673_),
    .X(\master_add_o[20]_reg_D ));
 sg13g2_nand4_1 _7324_ (.B(master_add_o_20_),
    .C(net280),
    .A(master_add_o_19_),
    .Y(_2674_),
    .D(net455));
 sg13g2_xor2_1 _7325_ (.B(_2674_),
    .A(master_add_o_21_),
    .X(_2675_));
 sg13g2_nor2_1 _7326_ (.A(net221),
    .B(net399),
    .Y(_2676_));
 sg13g2_a21oi_1 _7327_ (.A1(net399),
    .A2(_2675_),
    .Y(_2677_),
    .B1(_2676_));
 sg13g2_and2_1 _7328_ (.A(net82),
    .B(_2677_),
    .X(\master_add_o[21]_reg_D ));
 sg13g2_and3_1 _7329_ (.X(_2678_),
    .A(master_add_o_19_),
    .B(master_add_o_20_),
    .C(master_add_o_21_));
 sg13g2_nand3_1 _7330_ (.B(net456),
    .C(_2678_),
    .A(net281),
    .Y(_2679_));
 sg13g2_xor2_1 _7331_ (.B(_2679_),
    .A(master_add_o_22_),
    .X(_2680_));
 sg13g2_nor2_1 _7332_ (.A(net219),
    .B(net400),
    .Y(_2681_));
 sg13g2_a21oi_1 _7333_ (.A1(net400),
    .A2(_2680_),
    .Y(_2682_),
    .B1(_2681_));
 sg13g2_and2_1 _7334_ (.A(net82),
    .B(_2682_),
    .X(\master_add_o[22]_reg_D ));
 sg13g2_nand4_1 _7335_ (.B(net280),
    .C(net456),
    .A(master_add_o_22_),
    .Y(_2683_),
    .D(_2678_));
 sg13g2_xor2_1 _7336_ (.B(_2683_),
    .A(master_add_o_23_),
    .X(_2684_));
 sg13g2_nor2_1 _7337_ (.A(net799),
    .B(net399),
    .Y(_2685_));
 sg13g2_a21oi_1 _7338_ (.A1(net400),
    .A2(_2684_),
    .Y(_2686_),
    .B1(_2685_));
 sg13g2_and2_1 _7339_ (.A(net82),
    .B(_2686_),
    .X(\master_add_o[23]_reg_D ));
 sg13g2_and2_1 _7340_ (.A(master_add_o_22_),
    .B(master_add_o_23_),
    .X(_2687_));
 sg13g2_nand4_1 _7341_ (.B(net456),
    .C(_2678_),
    .A(net280),
    .Y(_2688_),
    .D(_2687_));
 sg13g2_xor2_1 _7342_ (.B(_2688_),
    .A(master_add_o_24_),
    .X(_2689_));
 sg13g2_nor2_1 _7343_ (.A(net217),
    .B(net399),
    .Y(_2690_));
 sg13g2_a21oi_1 _7344_ (.A1(net399),
    .A2(_2689_),
    .Y(_2691_),
    .B1(_2690_));
 sg13g2_and2_1 _7345_ (.A(net82),
    .B(_2691_),
    .X(\master_add_o[24]_reg_D ));
 sg13g2_and3_2 _7346_ (.X(_2692_),
    .A(master_add_o_24_),
    .B(_2678_),
    .C(_2687_));
 sg13g2_nand3_1 _7347_ (.B(net455),
    .C(_2692_),
    .A(net281),
    .Y(_2693_));
 sg13g2_xor2_1 _7348_ (.B(_2693_),
    .A(master_add_o_25_),
    .X(_2694_));
 sg13g2_nor2_1 _7349_ (.A(net215),
    .B(net402),
    .Y(_2695_));
 sg13g2_a21oi_1 _7350_ (.A1(net401),
    .A2(_2694_),
    .Y(_2696_),
    .B1(_2695_));
 sg13g2_and2_1 _7351_ (.A(net82),
    .B(_2696_),
    .X(\master_add_o[25]_reg_D ));
 sg13g2_buf_8 fanout137 (.A(net797),
    .X(net137));
 sg13g2_nand4_1 _7353_ (.B(net281),
    .C(net455),
    .A(master_add_o_25_),
    .Y(_2698_),
    .D(_2692_));
 sg13g2_xor2_1 _7354_ (.B(_2698_),
    .A(master_add_o_26_),
    .X(_2699_));
 sg13g2_nor2_1 _7355_ (.A(net213),
    .B(net402),
    .Y(_2700_));
 sg13g2_a21oi_1 _7356_ (.A1(net402),
    .A2(_2699_),
    .Y(_2701_),
    .B1(_2700_));
 sg13g2_and2_1 _7357_ (.A(net80),
    .B(_2701_),
    .X(\master_add_o[26]_reg_D ));
 sg13g2_and2_1 _7358_ (.A(master_add_o_25_),
    .B(master_add_o_26_),
    .X(_2702_));
 sg13g2_nand4_1 _7359_ (.B(net455),
    .C(_2692_),
    .A(net280),
    .Y(_2703_),
    .D(_2702_));
 sg13g2_xor2_1 _7360_ (.B(_2703_),
    .A(master_add_o_27_),
    .X(_2704_));
 sg13g2_nor2_1 _7361_ (.A(net211),
    .B(net401),
    .Y(_2705_));
 sg13g2_a21oi_1 _7362_ (.A1(net401),
    .A2(_2704_),
    .Y(_2706_),
    .B1(_2705_));
 sg13g2_and2_1 _7363_ (.A(net80),
    .B(_2706_),
    .X(\master_add_o[27]_reg_D ));
 sg13g2_and2_1 _7364_ (.A(master_add_o_27_),
    .B(_2702_),
    .X(_2707_));
 sg13g2_nand4_1 _7365_ (.B(net455),
    .C(_2692_),
    .A(net280),
    .Y(_2708_),
    .D(_2707_));
 sg13g2_xor2_1 _7366_ (.B(_2708_),
    .A(master_add_o_28_),
    .X(_2709_));
 sg13g2_nor2_1 _7367_ (.A(net209),
    .B(net401),
    .Y(_2710_));
 sg13g2_a21oi_1 _7368_ (.A1(net401),
    .A2(_2709_),
    .Y(_2711_),
    .B1(_2710_));
 sg13g2_and2_1 _7369_ (.A(net80),
    .B(_2711_),
    .X(\master_add_o[28]_reg_D ));
 sg13g2_and2_1 _7370_ (.A(master_add_o_28_),
    .B(_2707_),
    .X(_2712_));
 sg13g2_nand4_1 _7371_ (.B(net455),
    .C(_2692_),
    .A(net280),
    .Y(_2713_),
    .D(_2712_));
 sg13g2_xor2_1 _7372_ (.B(_2713_),
    .A(master_add_o_29_),
    .X(_2714_));
 sg13g2_nor2_1 _7373_ (.A(net207),
    .B(net403),
    .Y(_2715_));
 sg13g2_a21oi_1 _7374_ (.A1(net403),
    .A2(_2714_),
    .Y(_2716_),
    .B1(_2715_));
 sg13g2_and2_1 _7375_ (.A(net80),
    .B(_2716_),
    .X(\master_add_o[29]_reg_D ));
 sg13g2_nor2_1 _7376_ (.A(_1517_),
    .B(net628),
    .Y(_2717_));
 sg13g2_a22oi_1 _7377_ (.Y(_2718_),
    .B1(_2592_),
    .B2(_2589_),
    .A2(_2717_),
    .A1(net78));
 sg13g2_nor2_1 _7378_ (.A(_2564_),
    .B(_2718_),
    .Y(_2719_));
 sg13g2_xnor2_1 _7379_ (.Y(_2720_),
    .A(net50),
    .B(_2719_));
 sg13g2_nand2_2 _7380_ (.Y(_2721_),
    .A(net398),
    .B(_2720_));
 sg13g2_o21ai_1 _7381_ (.B1(_2721_),
    .Y(_2722_),
    .A1(net205),
    .A2(net398));
 sg13g2_nor2_1 _7382_ (.A(net598),
    .B(_2722_),
    .Y(\master_add_o[2]_reg_D ));
 sg13g2_and3_1 _7383_ (.X(_2723_),
    .A(master_add_o_29_),
    .B(_2692_),
    .C(_2712_));
 sg13g2_nand3_1 _7384_ (.B(net455),
    .C(_2723_),
    .A(net282),
    .Y(_2724_));
 sg13g2_xor2_1 _7385_ (.B(_2724_),
    .A(master_add_o_30_),
    .X(_2725_));
 sg13g2_nor2_1 _7386_ (.A(net203),
    .B(net403),
    .Y(_2726_));
 sg13g2_a21oi_1 _7387_ (.A1(net403),
    .A2(_2725_),
    .Y(_2727_),
    .B1(_2726_));
 sg13g2_and2_1 _7388_ (.A(net80),
    .B(_2727_),
    .X(\master_add_o[30]_reg_D ));
 sg13g2_nand4_1 _7389_ (.B(net282),
    .C(net455),
    .A(master_add_o_30_),
    .Y(_2728_),
    .D(_2723_));
 sg13g2_xor2_1 _7390_ (.B(_2728_),
    .A(master_add_o_31_),
    .X(_2729_));
 sg13g2_nor2_1 _7391_ (.A(net201),
    .B(net403),
    .Y(_2730_));
 sg13g2_a21oi_1 _7392_ (.A1(net403),
    .A2(_2729_),
    .Y(_2731_),
    .B1(_2730_));
 sg13g2_and2_1 _7393_ (.A(net80),
    .B(_2731_),
    .X(\master_add_o[31]_reg_D ));
 sg13g2_nand2_2 _7394_ (.Y(_2732_),
    .A(_2447_),
    .B(net803));
 sg13g2_buf_8 fanout136 (.A(net797),
    .X(net136));
 sg13g2_nor2_2 _7396_ (.A(_0606_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_32__reg_D ));
 sg13g2_nor2_2 _7397_ (.A(_0655_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_33__reg_D ));
 sg13g2_nor2_2 _7398_ (.A(_0679_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_34__reg_D ));
 sg13g2_nor2_2 _7399_ (.A(_0687_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_35__reg_D ));
 sg13g2_nor2_2 _7400_ (.A(_0690_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_36__reg_D ));
 sg13g2_nor2_2 _7401_ (.A(_0693_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_37__reg_D ));
 sg13g2_nor2_2 _7402_ (.A(_0696_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_38__reg_D ));
 sg13g2_nor2_2 _7403_ (.A(_0699_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_39__reg_D ));
 sg13g2_nand2b_1 _7404_ (.Y(_2734_),
    .B(net50),
    .A_N(_2718_));
 sg13g2_nand2_1 _7405_ (.Y(_2735_),
    .A(net632),
    .B(_2717_));
 sg13g2_xnor2_1 _7406_ (.Y(_2736_),
    .A(_2734_),
    .B(_2735_));
 sg13g2_nor2_1 _7407_ (.A(_2564_),
    .B(_2736_),
    .Y(_2737_));
 sg13g2_xnor2_1 _7408_ (.Y(_2738_),
    .A(master_add_o_3_),
    .B(_2737_));
 sg13g2_nand2_2 _7409_ (.Y(_2739_),
    .A(net404),
    .B(_2738_));
 sg13g2_o21ai_1 _7410_ (.B1(_2739_),
    .Y(_2740_),
    .A1(net128),
    .A2(net404));
 sg13g2_nor2_1 _7411_ (.A(net598),
    .B(_2740_),
    .Y(\master_add_o[3]_reg_D ));
 sg13g2_nor2_2 _7412_ (.A(_0701_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_40__reg_D ));
 sg13g2_nor2_2 _7413_ (.A(_0703_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_41__reg_D ));
 sg13g2_buf_4 fanout135 (.X(net135),
    .A(net797));
 sg13g2_nor2_2 _7415_ (.A(_0631_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_42__reg_D ));
 sg13g2_nor2_2 _7416_ (.A(_0633_),
    .B(net389),
    .Y(\i_dm_csrs.sbaddr_q_43__reg_D ));
 sg13g2_nor2_2 _7417_ (.A(_0635_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_44__reg_D ));
 sg13g2_nand2_1 _7418_ (.Y(_2742_),
    .A(net85),
    .B(net802));
 sg13g2_nor2_2 _7419_ (.A(net392),
    .B(_2742_),
    .Y(\i_dm_csrs.sbaddr_q_45__reg_D ));
 sg13g2_nor2_2 _7420_ (.A(_0638_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_46__reg_D ));
 sg13g2_nor2_2 _7421_ (.A(_0640_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_47__reg_D ));
 sg13g2_nor2_2 _7422_ (.A(_0643_),
    .B(net390),
    .Y(\i_dm_csrs.sbaddr_q_48__reg_D ));
 sg13g2_nor2_2 _7423_ (.A(_0646_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_49__reg_D ));
 sg13g2_nor2_1 _7424_ (.A(net546),
    .B(_2575_),
    .Y(_2743_));
 sg13g2_xnor2_1 _7425_ (.Y(_2744_),
    .A(_2596_),
    .B(_2743_));
 sg13g2_nor2_1 _7426_ (.A(net427),
    .B(_2744_),
    .Y(_2745_));
 sg13g2_xnor2_1 _7427_ (.Y(_2746_),
    .A(master_add_o_4_),
    .B(_2745_));
 sg13g2_nand2_1 _7428_ (.Y(_2747_),
    .A(net397),
    .B(_2746_));
 sg13g2_o21ai_1 _7429_ (.B1(_2747_),
    .Y(_2748_),
    .A1(net126),
    .A2(net397));
 sg13g2_nor2_1 _7430_ (.A(net598),
    .B(_2748_),
    .Y(\master_add_o[4]_reg_D ));
 sg13g2_nor2_2 _7431_ (.A(_0648_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_50__reg_D ));
 sg13g2_nor2_2 _7432_ (.A(_0650_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_51__reg_D ));
 sg13g2_nor2_2 _7433_ (.A(_0658_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_52__reg_D ));
 sg13g2_buf_2 fanout134 (.A(net797),
    .X(net134));
 sg13g2_nor2_2 _7435_ (.A(_0660_),
    .B(net393),
    .Y(\i_dm_csrs.sbaddr_q_53__reg_D ));
 sg13g2_nor2_2 _7436_ (.A(_0662_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_54__reg_D ));
 sg13g2_nor2_2 _7437_ (.A(_1163_),
    .B(net393),
    .Y(\i_dm_csrs.sbaddr_q_55__reg_D ));
 sg13g2_nor2_2 _7438_ (.A(_0665_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_56__reg_D ));
 sg13g2_nor2_2 _7439_ (.A(_0667_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_57__reg_D ));
 sg13g2_nor2_2 _7440_ (.A(_0669_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_58__reg_D ));
 sg13g2_nor2_2 _7441_ (.A(_0671_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_59__reg_D ));
 sg13g2_or2_1 _7442_ (.X(_2750_),
    .B(net396),
    .A(net124));
 sg13g2_nor2_1 _7443_ (.A(net629),
    .B(_1536_),
    .Y(_2751_));
 sg13g2_nand3_1 _7444_ (.B(_2588_),
    .C(_2595_),
    .A(net48),
    .Y(_2752_));
 sg13g2_a21oi_1 _7445_ (.A1(_2588_),
    .A2(_2595_),
    .Y(_2753_),
    .B1(net48));
 sg13g2_a21oi_1 _7446_ (.A1(net546),
    .A2(_2752_),
    .Y(_2754_),
    .B1(_2753_));
 sg13g2_nand2b_1 _7447_ (.Y(_2755_),
    .B(_2599_),
    .A_N(_2753_));
 sg13g2_o21ai_1 _7448_ (.B1(_2755_),
    .Y(_2756_),
    .A1(_1496_),
    .A2(_2754_));
 sg13g2_a21oi_1 _7449_ (.A1(net631),
    .A2(_2751_),
    .Y(_2757_),
    .B1(_2752_));
 sg13g2_a21oi_2 _7450_ (.B1(_2757_),
    .Y(_2758_),
    .A2(_2756_),
    .A1(_2751_));
 sg13g2_or3_1 _7451_ (.A(master_add_o_5_),
    .B(net427),
    .C(_2758_),
    .X(_2759_));
 sg13g2_o21ai_1 _7452_ (.B1(master_add_o_5_),
    .Y(_2760_),
    .A1(net427),
    .A2(_2758_));
 sg13g2_nand3_1 _7453_ (.B(_2759_),
    .C(_2760_),
    .A(net397),
    .Y(_2761_));
 sg13g2_and3_1 _7454_ (.X(\master_add_o[5]_reg_D ),
    .A(net81),
    .B(_2750_),
    .C(_2761_));
 sg13g2_nor2_2 _7455_ (.A(_0673_),
    .B(net393),
    .Y(\i_dm_csrs.sbaddr_q_60__reg_D ));
 sg13g2_nor2_2 _7456_ (.A(_0675_),
    .B(net392),
    .Y(\i_dm_csrs.sbaddr_q_61__reg_D ));
 sg13g2_nor2_2 _7457_ (.A(_0682_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_62__reg_D ));
 sg13g2_nor2_2 _7458_ (.A(_0684_),
    .B(net391),
    .Y(\i_dm_csrs.sbaddr_q_63__reg_D ));
 sg13g2_nand3_1 _7459_ (.B(_2588_),
    .C(_2595_),
    .A(_2604_),
    .Y(_2762_));
 sg13g2_nor4_2 _7460_ (.A(_1517_),
    .B(_1536_),
    .C(net546),
    .Y(_2763_),
    .D(_2762_));
 sg13g2_and2_1 _7461_ (.A(\i_dm_csrs.sbautoincrement_o ),
    .B(_2563_),
    .X(_2764_));
 sg13g2_nand3_1 _7462_ (.B(net628),
    .C(net77),
    .A(net629),
    .Y(_2765_));
 sg13g2_nand3b_1 _7463_ (.B(_2765_),
    .C(_2762_),
    .Y(_2766_),
    .A_N(_2609_));
 sg13g2_nand3b_1 _7464_ (.B(_2764_),
    .C(_2766_),
    .Y(_2767_),
    .A_N(_2763_));
 sg13g2_xnor2_1 _7465_ (.Y(_2768_),
    .A(_2570_),
    .B(_2767_));
 sg13g2_nor2_1 _7466_ (.A(net122),
    .B(net395),
    .Y(_2769_));
 sg13g2_a21oi_1 _7467_ (.A1(net398),
    .A2(_2768_),
    .Y(_2770_),
    .B1(_2769_));
 sg13g2_and2_1 _7468_ (.A(net80),
    .B(_2770_),
    .X(\master_add_o[6]_reg_D ));
 sg13g2_or2_1 _7469_ (.X(_2771_),
    .B(net396),
    .A(net120));
 sg13g2_nand3_1 _7470_ (.B(net630),
    .C(net628),
    .A(net633),
    .Y(_2772_));
 sg13g2_a21oi_1 _7471_ (.A1(master_add_o_6_),
    .A2(_2766_),
    .Y(_2773_),
    .B1(_2763_));
 sg13g2_xnor2_1 _7472_ (.Y(_2774_),
    .A(_2772_),
    .B(_2773_));
 sg13g2_or3_1 _7473_ (.A(master_add_o_7_),
    .B(net427),
    .C(_2774_),
    .X(_2775_));
 sg13g2_o21ai_1 _7474_ (.B1(master_add_o_7_),
    .Y(_2776_),
    .A1(net427),
    .A2(_2774_));
 sg13g2_nand3_1 _7475_ (.B(_2775_),
    .C(_2776_),
    .A(net397),
    .Y(_2777_));
 sg13g2_and3_1 _7476_ (.X(\master_add_o[7]_reg_D ),
    .A(net81),
    .B(_2771_),
    .C(_2777_));
 sg13g2_xnor2_1 _7477_ (.Y(_2778_),
    .A(master_add_o_8_),
    .B(net280));
 sg13g2_nand2_1 _7478_ (.Y(_2779_),
    .A(net399),
    .B(_2778_));
 sg13g2_o21ai_1 _7479_ (.B1(_2779_),
    .Y(_2780_),
    .A1(net118),
    .A2(net399));
 sg13g2_nor2_1 _7480_ (.A(net598),
    .B(_2780_),
    .Y(\master_add_o[8]_reg_D ));
 sg13g2_nand2_2 _7481_ (.Y(_2781_),
    .A(master_add_o_8_),
    .B(net281));
 sg13g2_xor2_1 _7482_ (.B(_2781_),
    .A(master_add_o_9_),
    .X(_2782_));
 sg13g2_nor2_1 _7483_ (.A(net116),
    .B(net401),
    .Y(_2783_));
 sg13g2_a21oi_1 _7484_ (.A1(net404),
    .A2(_2782_),
    .Y(_2784_),
    .B1(_2783_));
 sg13g2_and2_1 _7485_ (.A(net80),
    .B(_2784_),
    .X(\master_add_o[9]_reg_D ));
 sg13g2_a22oi_1 _7486_ (.Y(_2785_),
    .B1(_2546_),
    .B2(net233),
    .A2(net428),
    .A1(\i_dm_csrs.sbautoincrement_o ));
 sg13g2_inv_1 _7487_ (.Y(_0441_),
    .A(_2785_));
 sg13g2_a21oi_1 _7488_ (.A1(net141),
    .A2(_1169_),
    .Y(_2786_),
    .B1(_0611_));
 sg13g2_nand2_1 _7489_ (.Y(_2787_),
    .A(_0611_),
    .B(_1271_));
 sg13g2_o21ai_1 _7490_ (.B1(_2787_),
    .Y(_2788_),
    .A1(net147),
    .A2(_2786_));
 sg13g2_a21oi_1 _7491_ (.A1(\i_dm_csrs.sbcs_q_22_ ),
    .A2(_0614_),
    .Y(_2789_),
    .B1(_1315_));
 sg13g2_nor3_1 _7492_ (.A(_0598_),
    .B(_1279_),
    .C(_2789_),
    .Y(_2790_));
 sg13g2_nand4_1 _7493_ (.B(_0599_),
    .C(_0602_),
    .A(net219),
    .Y(_2791_),
    .D(net532));
 sg13g2_a22oi_1 _7494_ (.Y(_2792_),
    .B1(_2791_),
    .B2(\i_dm_csrs.sbcs_q_22_ ),
    .A2(_2790_),
    .A1(_2788_));
 sg13g2_nor2_1 _7495_ (.A(net597),
    .B(_2792_),
    .Y(\i_dm_csrs.sbcs_q_22__reg_D ));
 sg13g2_nor2_1 _7496_ (.A(_2570_),
    .B(net78),
    .Y(_2793_));
 sg13g2_or2_1 _7497_ (.X(_2794_),
    .B(master_add_o_5_),
    .A(net48));
 sg13g2_o21ai_1 _7498_ (.B1(net629),
    .Y(_2795_),
    .A1(_2793_),
    .A2(_2794_));
 sg13g2_nor2b_1 _7499_ (.A(\i_dm_sba.sbaccess_mask_3__$_AND__B_A_$_AND__Y_A ),
    .B_N(net48),
    .Y(_2796_));
 sg13g2_or2_1 _7500_ (.X(_2797_),
    .B(master_add_o_1_),
    .A(net51));
 sg13g2_nor4_1 _7501_ (.A(net50),
    .B(master_add_o_3_),
    .C(_2796_),
    .D(_2797_),
    .Y(_2798_));
 sg13g2_a21o_1 _7502_ (.A2(master_add_o_2_),
    .A1(net629),
    .B1(net51),
    .X(_2799_));
 sg13g2_a221oi_1 _7503_ (.B2(net629),
    .C1(net628),
    .B1(_2797_),
    .A1(net546),
    .Y(_2800_),
    .A2(_2799_));
 sg13g2_a21oi_2 _7504_ (.B1(_2800_),
    .Y(_2801_),
    .A2(_2798_),
    .A1(_2795_));
 sg13g2_nand2_1 _7505_ (.Y(_2802_),
    .A(_1315_),
    .B(_2801_));
 sg13g2_nand2_1 _7506_ (.Y(_2803_),
    .A(net630),
    .B(\i_dm_sba.sbaccess_mask_3_ ));
 sg13g2_mux2_1 _7507_ (.A0(net79),
    .A1(_1536_),
    .S(_2803_),
    .X(_2804_));
 sg13g2_nor2_1 _7508_ (.A(net41),
    .B(_2804_),
    .Y(_2805_));
 sg13g2_nor2b_1 _7509_ (.A(_2805_),
    .B_N(_2563_),
    .Y(_2806_));
 sg13g2_nand2_1 _7510_ (.Y(_2807_),
    .A(master_r_other_err_i),
    .B(_2806_));
 sg13g2_buf_2 fanout133 (.A(dmi_req_i_37_),
    .X(net133));
 sg13g2_a21oi_1 _7512_ (.A1(_2802_),
    .A2(_2807_),
    .Y(_2809_),
    .B1(net599));
 sg13g2_inv_2 _7513_ (.Y(_2810_),
    .A(_2801_));
 sg13g2_a21oi_2 _7514_ (.B1(net41),
    .Y(_2811_),
    .A2(_2804_),
    .A1(_2810_));
 sg13g2_o21ai_1 _7515_ (.B1(_2563_),
    .Y(_2812_),
    .A1(master_r_err_i),
    .A2(master_r_other_err_i));
 sg13g2_inv_1 _7516_ (.Y(_2813_),
    .A(_2812_));
 sg13g2_nor3_1 _7517_ (.A(net239),
    .B(net237),
    .C(net802),
    .Y(_2814_));
 sg13g2_nor2_1 _7518_ (.A(_2540_),
    .B(_2814_),
    .Y(_2815_));
 sg13g2_nor4_2 _7519_ (.A(\ndmreset_o_reg_E_$_AND__Y_B_$_OR__Y_A ),
    .B(_2811_),
    .C(_2813_),
    .Y(_2816_),
    .D(_2815_));
 sg13g2_mux2_1 _7520_ (.A0(_2809_),
    .A1(\i_dm_csrs.sbcs_q_12_ ),
    .S(_2816_),
    .X(_0442_));
 sg13g2_o21ai_1 _7521_ (.B1(_2806_),
    .Y(_2817_),
    .A1(master_r_err_i),
    .A2(master_r_other_err_i));
 sg13g2_a21oi_1 _7522_ (.A1(_2802_),
    .A2(_2817_),
    .Y(_2818_),
    .B1(net599));
 sg13g2_mux2_1 _7523_ (.A0(_2818_),
    .A1(\i_dm_csrs.sbcs_q_13_ ),
    .S(_2816_),
    .X(_0443_));
 sg13g2_a21o_1 _7524_ (.A2(_2563_),
    .A1(master_r_other_err_i),
    .B1(_2805_),
    .X(_2819_));
 sg13g2_nand3_1 _7525_ (.B(_2802_),
    .C(_2819_),
    .A(net98),
    .Y(_2820_));
 sg13g2_nand2_1 _7526_ (.Y(_2821_),
    .A(\i_dm_csrs.sbcs_q_14_ ),
    .B(_2816_));
 sg13g2_o21ai_1 _7527_ (.B1(_2821_),
    .Y(_0444_),
    .A1(_2816_),
    .A2(_2820_));
 sg13g2_nor2_2 _7528_ (.A(net598),
    .B(_1255_),
    .Y(\i_dm_csrs.sbcs_q_21__reg_D ));
 sg13g2_a22oi_1 _7529_ (.Y(_2822_),
    .B1(_2545_),
    .B2(net799),
    .A2(net429),
    .A1(\i_dm_csrs.sbcs_q_23_ ));
 sg13g2_inv_1 _7530_ (.Y(_0445_),
    .A(_2822_));
 sg13g2_a22oi_1 _7531_ (.Y(_2823_),
    .B1(_2545_),
    .B2(net217),
    .A2(net429),
    .A1(\i_dm_csrs.sbcs_q_24_ ));
 sg13g2_inv_1 _7532_ (.Y(_0446_),
    .A(_2823_));
 sg13g2_a22oi_1 _7533_ (.Y(_2824_),
    .B1(_2545_),
    .B2(net215),
    .A2(net429),
    .A1(\i_dm_csrs.sbcs_q_25_ ));
 sg13g2_inv_1 _7534_ (.Y(_0447_),
    .A(_2824_));
 sg13g2_a22oi_1 _7535_ (.Y(_2825_),
    .B1(_2545_),
    .B2(net213),
    .A2(net429),
    .A1(\i_dm_csrs.sbcs_q_26_ ));
 sg13g2_inv_1 _7536_ (.Y(_0448_),
    .A(_2825_));
 sg13g2_a22oi_1 _7537_ (.Y(_2826_),
    .B1(_2545_),
    .B2(net211),
    .A2(net429),
    .A1(\i_dm_csrs.sbcs_q_27_ ));
 sg13g2_inv_1 _7538_ (.Y(_0449_),
    .A(_2826_));
 sg13g2_a22oi_1 _7539_ (.Y(_2827_),
    .B1(_2545_),
    .B2(net209),
    .A2(net428),
    .A1(\i_dm_csrs.sbcs_q_28_ ));
 sg13g2_inv_1 _7540_ (.Y(_0450_),
    .A(_2827_));
 sg13g2_or2_1 _7541_ (.X(_2828_),
    .B(net639),
    .A(net791));
 sg13g2_a21oi_2 _7542_ (.B1(_2828_),
    .Y(_2829_),
    .A2(net803),
    .A1(_2008_));
 sg13g2_buf_2 fanout132 (.A(dmi_req_i_37_),
    .X(net132));
 sg13g2_buf_1 fanout131 (.A(dmi_req_i_39_),
    .X(net131));
 sg13g2_buf_2 fanout130 (.A(dmi_req_i_39_),
    .X(net130));
 sg13g2_inv_1 _7546_ (.Y(_2833_),
    .A(master_add_o_1_));
 sg13g2_nor2_1 _7547_ (.A(_2833_),
    .B(_2558_),
    .Y(_2834_));
 sg13g2_nand2_1 _7548_ (.Y(_2835_),
    .A(master_add_o_1_),
    .B(_2589_));
 sg13g2_buf_1 fanout129 (.A(dmi_req_i_3_),
    .X(net129));
 sg13g2_and2_1 _7550_ (.A(master_r_rdata_i_0_),
    .B(net506),
    .X(_2837_));
 sg13g2_a21oi_1 _7551_ (.A1(master_r_rdata_i_16_),
    .A2(net451),
    .Y(_2838_),
    .B1(_2837_));
 sg13g2_nand3_1 _7552_ (.B(net78),
    .C(_2589_),
    .A(net51),
    .Y(_2839_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(dmi_req_i_3_));
 sg13g2_mux2_1 _7554_ (.A0(master_r_rdata_i_24_),
    .A1(master_r_rdata_i_8_),
    .S(net506),
    .X(_2841_));
 sg13g2_nor2_1 _7555_ (.A(_2841_),
    .B(net502),
    .Y(_2842_));
 sg13g2_a21oi_2 _7556_ (.B1(_2842_),
    .Y(_2843_),
    .A2(net502),
    .A1(_2838_));
 sg13g2_buf_1 fanout127 (.A(dmi_req_i_4_),
    .X(net127));
 sg13g2_nor2b_1 _7558_ (.A(net791),
    .B_N(net245),
    .Y(_2845_));
 sg13g2_a21oi_2 _7559_ (.B1(_2845_),
    .Y(_2846_),
    .A2(_2843_),
    .A1(net791));
 sg13g2_buf_8 fanout126 (.A(dmi_req_i_4_),
    .X(net126));
 sg13g2_nor3_2 _7561_ (.A(net596),
    .B(_2846_),
    .C(net22),
    .Y(_2848_));
 sg13g2_a21o_1 _7562_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_0_ ),
    .B1(_2848_),
    .X(_0451_));
 sg13g2_buf_1 fanout125 (.A(dmi_req_i_5_),
    .X(net125));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(dmi_req_i_5_));
 sg13g2_buf_1 fanout123 (.A(dmi_req_i_6_),
    .X(net123));
 sg13g2_mux2_1 _7566_ (.A0(master_r_rdata_i_26_),
    .A1(master_r_rdata_i_10_),
    .S(net508),
    .X(_2852_));
 sg13g2_nand2_2 _7567_ (.Y(_2853_),
    .A(net502),
    .B(_2852_));
 sg13g2_buf_4 fanout122 (.X(net122),
    .A(dmi_req_i_6_));
 sg13g2_buf_1 fanout121 (.A(dmi_req_i_7_),
    .X(net121));
 sg13g2_nor2_2 _7570_ (.A(_2558_),
    .B(_2663_),
    .Y(_2856_));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(dmi_req_i_7_));
 sg13g2_nand3_1 _7572_ (.B(net506),
    .C(net443),
    .A(master_r_rdata_i_18_),
    .Y(_2858_));
 sg13g2_nand3_1 _7573_ (.B(_2853_),
    .C(_2858_),
    .A(net780),
    .Y(_2859_));
 sg13g2_o21ai_1 _7574_ (.B1(_2859_),
    .Y(_2860_),
    .A1(net243),
    .A2(net785));
 sg13g2_nor3_2 _7575_ (.A(net594),
    .B(net20),
    .C(_2860_),
    .Y(_2861_));
 sg13g2_a21o_1 _7576_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_10_ ),
    .B1(_2861_),
    .X(_0452_));
 sg13g2_buf_2 fanout119 (.A(dmi_req_i_8_),
    .X(net119));
 sg13g2_mux2_1 _7578_ (.A0(master_r_rdata_i_27_),
    .A1(master_r_rdata_i_11_),
    .S(net507),
    .X(_2863_));
 sg13g2_nand2_1 _7579_ (.Y(_2864_),
    .A(net504),
    .B(_2863_));
 sg13g2_nand3_1 _7580_ (.B(net507),
    .C(net442),
    .A(master_r_rdata_i_19_),
    .Y(_2865_));
 sg13g2_nand3_1 _7581_ (.B(_2864_),
    .C(_2865_),
    .A(net781),
    .Y(_2866_));
 sg13g2_o21ai_1 _7582_ (.B1(_2866_),
    .Y(_2867_),
    .A1(net241),
    .A2(net781));
 sg13g2_nor3_2 _7583_ (.A(net595),
    .B(net19),
    .C(_2867_),
    .Y(_2868_));
 sg13g2_a21o_1 _7584_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_11_ ),
    .B1(_2868_),
    .X(_0453_));
 sg13g2_mux2_1 _7585_ (.A0(master_r_rdata_i_28_),
    .A1(master_r_rdata_i_12_),
    .S(net508),
    .X(_2869_));
 sg13g2_nand2_2 _7586_ (.Y(_2870_),
    .A(net504),
    .B(_2869_));
 sg13g2_nand3_1 _7587_ (.B(net508),
    .C(net442),
    .A(master_r_rdata_i_20_),
    .Y(_2871_));
 sg13g2_nand3_1 _7588_ (.B(_2870_),
    .C(_2871_),
    .A(net781),
    .Y(_2872_));
 sg13g2_o21ai_1 _7589_ (.B1(_2872_),
    .Y(_2873_),
    .A1(net239),
    .A2(net781));
 sg13g2_nor3_2 _7590_ (.A(net595),
    .B(net19),
    .C(_2873_),
    .Y(_2874_));
 sg13g2_a21o_1 _7591_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_12_ ),
    .B1(_2874_),
    .X(_0454_));
 sg13g2_mux2_1 _7592_ (.A0(master_r_rdata_i_29_),
    .A1(master_r_rdata_i_13_),
    .S(net506),
    .X(_2875_));
 sg13g2_nand2_2 _7593_ (.Y(_2876_),
    .A(net502),
    .B(_2875_));
 sg13g2_nand3_1 _7594_ (.B(net509),
    .C(net443),
    .A(master_r_rdata_i_21_),
    .Y(_2877_));
 sg13g2_nand3_1 _7595_ (.B(_2876_),
    .C(_2877_),
    .A(net780),
    .Y(_2878_));
 sg13g2_o21ai_1 _7596_ (.B1(_2878_),
    .Y(_2879_),
    .A1(net801),
    .A2(net780));
 sg13g2_nor3_2 _7597_ (.A(net594),
    .B(net19),
    .C(_2879_),
    .Y(_2880_));
 sg13g2_a21o_1 _7598_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_13_ ),
    .B1(_2880_),
    .X(_0455_));
 sg13g2_buf_4 fanout118 (.X(net118),
    .A(dmi_req_i_8_));
 sg13g2_mux2_1 _7600_ (.A0(master_r_rdata_i_30_),
    .A1(master_r_rdata_i_14_),
    .S(net507),
    .X(_2882_));
 sg13g2_nand2_2 _7601_ (.Y(_2883_),
    .A(net504),
    .B(_2882_));
 sg13g2_nand3_1 _7602_ (.B(net509),
    .C(net443),
    .A(master_r_rdata_i_22_),
    .Y(_2884_));
 sg13g2_nand3_1 _7603_ (.B(_2883_),
    .C(_2884_),
    .A(net780),
    .Y(_2885_));
 sg13g2_o21ai_1 _7604_ (.B1(_2885_),
    .Y(_2886_),
    .A1(net237),
    .A2(net787));
 sg13g2_nor3_2 _7605_ (.A(net594),
    .B(net19),
    .C(_2886_),
    .Y(_2887_));
 sg13g2_a21o_1 _7606_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_14_ ),
    .B1(_2887_),
    .X(_0456_));
 sg13g2_mux2_1 _7607_ (.A0(master_r_rdata_i_31_),
    .A1(master_r_rdata_i_15_),
    .S(net507),
    .X(_2888_));
 sg13g2_nand2_2 _7608_ (.Y(_2889_),
    .A(net503),
    .B(_2888_));
 sg13g2_nand3_1 _7609_ (.B(net507),
    .C(net442),
    .A(master_r_rdata_i_23_),
    .Y(_2890_));
 sg13g2_nand3_1 _7610_ (.B(_2889_),
    .C(_2890_),
    .A(net781),
    .Y(_2891_));
 sg13g2_o21ai_1 _7611_ (.B1(_2891_),
    .Y(_2892_),
    .A1(net235),
    .A2(net786));
 sg13g2_nor3_2 _7612_ (.A(net594),
    .B(net19),
    .C(_2892_),
    .Y(_2893_));
 sg13g2_a21o_1 _7613_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_15_ ),
    .B1(_2893_),
    .X(_0457_));
 sg13g2_nand2b_1 _7614_ (.Y(_2894_),
    .B(net233),
    .A_N(net784));
 sg13g2_buf_2 fanout117 (.A(dmi_req_i_9_),
    .X(net117));
 sg13g2_buf_4 fanout116 (.X(net116),
    .A(dmi_req_i_9_));
 sg13g2_mux2_1 _7617_ (.A0(master_r_rdata_i_16_),
    .A1(master_r_rdata_i_24_),
    .S(net443),
    .X(_2897_));
 sg13g2_nand3_1 _7618_ (.B(net510),
    .C(_2897_),
    .A(net784),
    .Y(_2898_));
 sg13g2_a21oi_1 _7619_ (.A1(_2894_),
    .A2(_2898_),
    .Y(_2899_),
    .B1(net593));
 sg13g2_buf_2 fanout115 (.A(slave_addr_i_3_),
    .X(net115));
 sg13g2_mux2_1 _7621_ (.A0(_2899_),
    .A1(\i_dm_csrs.sbdata_o_16_ ),
    .S(net20),
    .X(_0458_));
 sg13g2_nand2b_1 _7622_ (.Y(_2901_),
    .B(net231),
    .A_N(net782));
 sg13g2_mux2_1 _7623_ (.A0(master_r_rdata_i_17_),
    .A1(master_r_rdata_i_25_),
    .S(net442),
    .X(_2902_));
 sg13g2_nand3_1 _7624_ (.B(net510),
    .C(_2902_),
    .A(net782),
    .Y(_2903_));
 sg13g2_a21oi_1 _7625_ (.A1(_2901_),
    .A2(_2903_),
    .Y(_2904_),
    .B1(net592));
 sg13g2_mux2_1 _7626_ (.A0(_2904_),
    .A1(\i_dm_csrs.sbdata_o_17_ ),
    .S(net20),
    .X(_0459_));
 sg13g2_nand2b_1 _7627_ (.Y(_2905_),
    .B(net229),
    .A_N(net784));
 sg13g2_mux2_1 _7628_ (.A0(master_r_rdata_i_18_),
    .A1(master_r_rdata_i_26_),
    .S(net443),
    .X(_2906_));
 sg13g2_nand3_1 _7629_ (.B(net506),
    .C(_2906_),
    .A(net780),
    .Y(_2907_));
 sg13g2_a21oi_1 _7630_ (.A1(_2905_),
    .A2(_2907_),
    .Y(_2908_),
    .B1(net593));
 sg13g2_mux2_1 _7631_ (.A0(_2908_),
    .A1(\i_dm_csrs.sbdata_o_18_ ),
    .S(net20),
    .X(_0460_));
 sg13g2_nand2b_1 _7632_ (.Y(_2909_),
    .B(net227),
    .A_N(net782));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(net115));
 sg13g2_mux2_1 _7634_ (.A0(master_r_rdata_i_19_),
    .A1(master_r_rdata_i_27_),
    .S(net443),
    .X(_2911_));
 sg13g2_nand3_1 _7635_ (.B(net510),
    .C(_2911_),
    .A(net782),
    .Y(_2912_));
 sg13g2_a21oi_1 _7636_ (.A1(_2909_),
    .A2(_2912_),
    .Y(_2913_),
    .B1(net592));
 sg13g2_mux2_1 _7637_ (.A0(_2913_),
    .A1(\i_dm_csrs.sbdata_o_19_ ),
    .S(net20),
    .X(_0461_));
 sg13g2_buf_8 fanout113 (.A(net115),
    .X(net113));
 sg13g2_buf_8 fanout112 (.A(net115),
    .X(net112));
 sg13g2_and2_1 _7640_ (.A(master_r_rdata_i_1_),
    .B(net507),
    .X(_2916_));
 sg13g2_a21oi_1 _7641_ (.A1(master_r_rdata_i_17_),
    .A2(net451),
    .Y(_2917_),
    .B1(_2916_));
 sg13g2_mux2_1 _7642_ (.A0(master_r_rdata_i_25_),
    .A1(master_r_rdata_i_9_),
    .S(net508),
    .X(_2918_));
 sg13g2_nor2_2 _7643_ (.A(net503),
    .B(_2918_),
    .Y(_2919_));
 sg13g2_a21oi_2 _7644_ (.B1(_2919_),
    .Y(_2920_),
    .A2(_2917_),
    .A1(net503));
 sg13g2_nor2b_1 _7645_ (.A(net786),
    .B_N(net225),
    .Y(_2921_));
 sg13g2_a21oi_1 _7646_ (.A1(net787),
    .A2(_2920_),
    .Y(_2922_),
    .B1(_2921_));
 sg13g2_nor3_2 _7647_ (.A(net594),
    .B(net19),
    .C(_2922_),
    .Y(_2923_));
 sg13g2_a21o_1 _7648_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_1_ ),
    .B1(_2923_),
    .X(_0462_));
 sg13g2_nand2b_1 _7649_ (.Y(_2924_),
    .B(net223),
    .A_N(net782));
 sg13g2_buf_4 fanout111 (.X(net111),
    .A(slave_addr_i_3_));
 sg13g2_mux2_1 _7651_ (.A0(master_r_rdata_i_20_),
    .A1(master_r_rdata_i_28_),
    .S(net442),
    .X(_2926_));
 sg13g2_nand3_1 _7652_ (.B(net510),
    .C(_2926_),
    .A(net782),
    .Y(_2927_));
 sg13g2_a21oi_2 _7653_ (.B1(net592),
    .Y(_2928_),
    .A2(_2927_),
    .A1(_2924_));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110));
 sg13g2_mux2_1 _7655_ (.A0(_2928_),
    .A1(\i_dm_csrs.sbdata_o_20_ ),
    .S(net21),
    .X(_0463_));
 sg13g2_nand2b_1 _7656_ (.Y(_2930_),
    .B(net221),
    .A_N(net782));
 sg13g2_mux2_1 _7657_ (.A0(master_r_rdata_i_21_),
    .A1(master_r_rdata_i_29_),
    .S(net442),
    .X(_2931_));
 sg13g2_nand3_1 _7658_ (.B(net509),
    .C(_2931_),
    .A(net781),
    .Y(_2932_));
 sg13g2_a21oi_2 _7659_ (.B1(net592),
    .Y(_2933_),
    .A2(_2932_),
    .A1(_2930_));
 sg13g2_mux2_1 _7660_ (.A0(_2933_),
    .A1(\i_dm_csrs.sbdata_o_21_ ),
    .S(net21),
    .X(_0464_));
 sg13g2_buf_2 fanout109 (.A(slave_addr_i_3_),
    .X(net109));
 sg13g2_nand2b_1 _7662_ (.Y(_2935_),
    .B(net219),
    .A_N(net786));
 sg13g2_mux2_1 _7663_ (.A0(master_r_rdata_i_22_),
    .A1(master_r_rdata_i_30_),
    .S(net442),
    .X(_2936_));
 sg13g2_nand3_1 _7664_ (.B(net515),
    .C(_2936_),
    .A(net786),
    .Y(_2937_));
 sg13g2_a21oi_1 _7665_ (.A1(_2935_),
    .A2(_2937_),
    .Y(_2938_),
    .B1(net594));
 sg13g2_mux2_1 _7666_ (.A0(_2938_),
    .A1(\i_dm_csrs.sbdata_o_22_ ),
    .S(net21),
    .X(_0465_));
 sg13g2_nand2b_1 _7667_ (.Y(_2939_),
    .B(net799),
    .A_N(net787));
 sg13g2_mux2_1 _7668_ (.A0(master_r_rdata_i_23_),
    .A1(master_r_rdata_i_31_),
    .S(net450),
    .X(_2940_));
 sg13g2_nand3_1 _7669_ (.B(net515),
    .C(_2940_),
    .A(net787),
    .Y(_2941_));
 sg13g2_a21oi_1 _7670_ (.A1(_2939_),
    .A2(_2941_),
    .Y(_2942_),
    .B1(net594));
 sg13g2_mux2_1 _7671_ (.A0(_2942_),
    .A1(\i_dm_csrs.sbdata_o_23_ ),
    .S(net21),
    .X(_0466_));
 sg13g2_nand2b_1 _7672_ (.Y(_2943_),
    .B(net217),
    .A_N(net783));
 sg13g2_nor2_2 _7673_ (.A(net454),
    .B(net450),
    .Y(_2944_));
 sg13g2_buf_8 fanout108 (.A(net111),
    .X(net108));
 sg13g2_nand3_1 _7675_ (.B(master_r_rdata_i_24_),
    .C(net425),
    .A(net783),
    .Y(_2946_));
 sg13g2_a21oi_1 _7676_ (.A1(_2943_),
    .A2(_2946_),
    .Y(_2947_),
    .B1(net593));
 sg13g2_mux2_1 _7677_ (.A0(_2947_),
    .A1(\i_dm_csrs.sbdata_o_24_ ),
    .S(net21),
    .X(_0467_));
 sg13g2_nand2b_1 _7678_ (.Y(_2948_),
    .B(net215),
    .A_N(net783));
 sg13g2_nand3_1 _7679_ (.B(master_r_rdata_i_25_),
    .C(net425),
    .A(net783),
    .Y(_2949_));
 sg13g2_a21oi_1 _7680_ (.A1(_2948_),
    .A2(_2949_),
    .Y(_2950_),
    .B1(net592));
 sg13g2_mux2_1 _7681_ (.A0(_2950_),
    .A1(\i_dm_csrs.sbdata_o_25_ ),
    .S(net21),
    .X(_0468_));
 sg13g2_nand2b_1 _7682_ (.Y(_2951_),
    .B(net213),
    .A_N(net786));
 sg13g2_nand3_1 _7683_ (.B(master_r_rdata_i_26_),
    .C(net425),
    .A(net783),
    .Y(_2952_));
 sg13g2_a21oi_1 _7684_ (.A1(_2951_),
    .A2(_2952_),
    .Y(_2953_),
    .B1(net592));
 sg13g2_mux2_1 _7685_ (.A0(_2953_),
    .A1(\i_dm_csrs.sbdata_o_26_ ),
    .S(net21),
    .X(_0469_));
 sg13g2_nand2b_1 _7686_ (.Y(_2954_),
    .B(net211),
    .A_N(net785));
 sg13g2_nand3_1 _7687_ (.B(master_r_rdata_i_27_),
    .C(net425),
    .A(net785),
    .Y(_2955_));
 sg13g2_a21oi_1 _7688_ (.A1(_2954_),
    .A2(_2955_),
    .Y(_2956_),
    .B1(net593));
 sg13g2_mux2_1 _7689_ (.A0(_2956_),
    .A1(\i_dm_csrs.sbdata_o_27_ ),
    .S(net20),
    .X(_0470_));
 sg13g2_nand2b_1 _7690_ (.Y(_2957_),
    .B(net209),
    .A_N(net783));
 sg13g2_nand3_1 _7691_ (.B(master_r_rdata_i_28_),
    .C(net425),
    .A(net782),
    .Y(_2958_));
 sg13g2_a21oi_1 _7692_ (.A1(_2957_),
    .A2(_2958_),
    .Y(_2959_),
    .B1(net592));
 sg13g2_mux2_1 _7693_ (.A0(_2959_),
    .A1(\i_dm_csrs.sbdata_o_28_ ),
    .S(net20),
    .X(_0471_));
 sg13g2_nand2b_1 _7694_ (.Y(_2960_),
    .B(net207),
    .A_N(net785));
 sg13g2_nand3_1 _7695_ (.B(master_r_rdata_i_29_),
    .C(net425),
    .A(net785),
    .Y(_2961_));
 sg13g2_a21oi_1 _7696_ (.A1(_2960_),
    .A2(_2961_),
    .Y(_2962_),
    .B1(net592));
 sg13g2_mux2_1 _7697_ (.A0(_2962_),
    .A1(\i_dm_csrs.sbdata_o_29_ ),
    .S(net20),
    .X(_0472_));
 sg13g2_and2_1 _7698_ (.A(master_r_rdata_i_2_),
    .B(net506),
    .X(_2963_));
 sg13g2_a21oi_1 _7699_ (.A1(master_r_rdata_i_18_),
    .A2(net451),
    .Y(_2964_),
    .B1(_2963_));
 sg13g2_nor2_2 _7700_ (.A(net502),
    .B(_2852_),
    .Y(_2965_));
 sg13g2_a21oi_2 _7701_ (.B1(_2965_),
    .Y(_2966_),
    .A2(_2964_),
    .A1(net502));
 sg13g2_nor2b_1 _7702_ (.A(net788),
    .B_N(net205),
    .Y(_2967_));
 sg13g2_a21oi_2 _7703_ (.B1(_2967_),
    .Y(_2968_),
    .A2(_2966_),
    .A1(net788));
 sg13g2_nor3_2 _7704_ (.A(net596),
    .B(net18),
    .C(_2968_),
    .Y(_2969_));
 sg13g2_a21o_1 _7705_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_2_ ),
    .B1(_2969_),
    .X(_0473_));
 sg13g2_nand2b_1 _7706_ (.Y(_2970_),
    .B(net203),
    .A_N(net785));
 sg13g2_nand3_1 _7707_ (.B(master_r_rdata_i_30_),
    .C(net425),
    .A(net785),
    .Y(_2971_));
 sg13g2_a21oi_1 _7708_ (.A1(_2970_),
    .A2(_2971_),
    .Y(_2972_),
    .B1(net593));
 sg13g2_mux2_1 _7709_ (.A0(_2972_),
    .A1(\i_dm_csrs.sbdata_o_30_ ),
    .S(net19),
    .X(_0474_));
 sg13g2_nand2b_1 _7710_ (.Y(_2973_),
    .B(net201),
    .A_N(net787));
 sg13g2_nand3_1 _7711_ (.B(master_r_rdata_i_31_),
    .C(net425),
    .A(net786),
    .Y(_2974_));
 sg13g2_a21oi_1 _7712_ (.A1(_2973_),
    .A2(_2974_),
    .Y(_2975_),
    .B1(net594));
 sg13g2_mux2_1 _7713_ (.A0(_2975_),
    .A1(\i_dm_csrs.sbdata_o_31_ ),
    .S(net19),
    .X(_0475_));
 sg13g2_and2_1 _7714_ (.A(master_r_rdata_i_3_),
    .B(net507),
    .X(_2976_));
 sg13g2_a21oi_1 _7715_ (.A1(master_r_rdata_i_19_),
    .A2(net451),
    .Y(_2977_),
    .B1(_2976_));
 sg13g2_nor2_1 _7716_ (.A(net504),
    .B(_2863_),
    .Y(_2978_));
 sg13g2_a21oi_2 _7717_ (.B1(_2978_),
    .Y(_2979_),
    .A2(_2977_),
    .A1(net503));
 sg13g2_nor2b_1 _7718_ (.A(net788),
    .B_N(net128),
    .Y(_2980_));
 sg13g2_a21oi_1 _7719_ (.A1(net788),
    .A2(_2979_),
    .Y(_2981_),
    .B1(_2980_));
 sg13g2_nor3_2 _7720_ (.A(net597),
    .B(net18),
    .C(_2981_),
    .Y(_2982_));
 sg13g2_a21o_1 _7721_ (.A2(net22),
    .A1(\i_dm_csrs.sbdata_o_3_ ),
    .B1(_2982_),
    .X(_0476_));
 sg13g2_and2_1 _7722_ (.A(master_r_rdata_i_4_),
    .B(net508),
    .X(_2983_));
 sg13g2_a21oi_1 _7723_ (.A1(master_r_rdata_i_20_),
    .A2(net451),
    .Y(_2984_),
    .B1(_2983_));
 sg13g2_nor2_2 _7724_ (.A(net503),
    .B(_2869_),
    .Y(_2985_));
 sg13g2_a21oi_2 _7725_ (.B1(_2985_),
    .Y(_2986_),
    .A2(_2984_),
    .A1(net503));
 sg13g2_nor2b_1 _7726_ (.A(net786),
    .B_N(net126),
    .Y(_2987_));
 sg13g2_a21oi_2 _7727_ (.B1(_2987_),
    .Y(_2988_),
    .A2(_2986_),
    .A1(net786));
 sg13g2_nor3_2 _7728_ (.A(net596),
    .B(net18),
    .C(_2988_),
    .Y(_2989_));
 sg13g2_a21o_1 _7729_ (.A2(net24),
    .A1(\i_dm_csrs.sbdata_o_4_ ),
    .B1(_2989_),
    .X(_0477_));
 sg13g2_and2_1 _7730_ (.A(master_r_rdata_i_5_),
    .B(net506),
    .X(_2990_));
 sg13g2_a21oi_1 _7731_ (.A1(master_r_rdata_i_21_),
    .A2(net451),
    .Y(_2991_),
    .B1(_2990_));
 sg13g2_nor2_1 _7732_ (.A(net505),
    .B(_2875_),
    .Y(_2992_));
 sg13g2_a21oi_2 _7733_ (.B1(_2992_),
    .Y(_2993_),
    .A2(_2991_),
    .A1(net502));
 sg13g2_nor2b_1 _7734_ (.A(net780),
    .B_N(net124),
    .Y(_2994_));
 sg13g2_a21oi_2 _7735_ (.B1(_2994_),
    .Y(_2995_),
    .A2(_2993_),
    .A1(net780));
 sg13g2_nor3_2 _7736_ (.A(net596),
    .B(net18),
    .C(_2995_),
    .Y(_2996_));
 sg13g2_a21o_1 _7737_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_5_ ),
    .B1(_2996_),
    .X(_0478_));
 sg13g2_and2_1 _7738_ (.A(master_r_rdata_i_6_),
    .B(net507),
    .X(_2997_));
 sg13g2_a21oi_1 _7739_ (.A1(master_r_rdata_i_22_),
    .A2(net451),
    .Y(_2998_),
    .B1(_2997_));
 sg13g2_nor2_2 _7740_ (.A(net504),
    .B(_2882_),
    .Y(_2999_));
 sg13g2_a21oi_2 _7741_ (.B1(_2999_),
    .Y(_3000_),
    .A2(_2998_),
    .A1(net504));
 sg13g2_nor2b_1 _7742_ (.A(net785),
    .B_N(net122),
    .Y(_3001_));
 sg13g2_a21oi_2 _7743_ (.B1(_3001_),
    .Y(_3002_),
    .A2(_3000_),
    .A1(net787));
 sg13g2_nor3_2 _7744_ (.A(net596),
    .B(net18),
    .C(_3002_),
    .Y(_3003_));
 sg13g2_a21o_1 _7745_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_6_ ),
    .B1(_3003_),
    .X(_0479_));
 sg13g2_and2_1 _7746_ (.A(master_r_rdata_i_7_),
    .B(net508),
    .X(_3004_));
 sg13g2_a21oi_1 _7747_ (.A1(master_r_rdata_i_23_),
    .A2(net451),
    .Y(_3005_),
    .B1(_3004_));
 sg13g2_nor2_2 _7748_ (.A(net503),
    .B(_2888_),
    .Y(_3006_));
 sg13g2_a21oi_2 _7749_ (.B1(_3006_),
    .Y(_3007_),
    .A2(_3005_),
    .A1(net503));
 sg13g2_nor2b_1 _7750_ (.A(net788),
    .B_N(net120),
    .Y(_3008_));
 sg13g2_a21oi_2 _7751_ (.B1(_3008_),
    .Y(_3009_),
    .A2(_3007_),
    .A1(net788));
 sg13g2_nor3_2 _7752_ (.A(net596),
    .B(net18),
    .C(_3009_),
    .Y(_3010_));
 sg13g2_a21o_1 _7753_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_7_ ),
    .B1(_3010_),
    .X(_0480_));
 sg13g2_nand2_2 _7754_ (.Y(_3011_),
    .A(_2841_),
    .B(net502));
 sg13g2_nand3_1 _7755_ (.B(net506),
    .C(net443),
    .A(master_r_rdata_i_16_),
    .Y(_3012_));
 sg13g2_nand3_1 _7756_ (.B(_3011_),
    .C(_3012_),
    .A(net780),
    .Y(_3013_));
 sg13g2_o21ai_1 _7757_ (.B1(_3013_),
    .Y(_3014_),
    .A1(net118),
    .A2(net789));
 sg13g2_nor3_2 _7758_ (.A(net596),
    .B(net18),
    .C(_3014_),
    .Y(_3015_));
 sg13g2_a21o_1 _7759_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_8_ ),
    .B1(_3015_),
    .X(_0481_));
 sg13g2_nand2_2 _7760_ (.Y(_3016_),
    .A(net504),
    .B(_2918_));
 sg13g2_nand3_1 _7761_ (.B(net508),
    .C(net442),
    .A(master_r_rdata_i_17_),
    .Y(_3017_));
 sg13g2_nand3_1 _7762_ (.B(_3016_),
    .C(_3017_),
    .A(net781),
    .Y(_3018_));
 sg13g2_o21ai_1 _7763_ (.B1(_3018_),
    .Y(_3019_),
    .A1(net116),
    .A2(net788));
 sg13g2_nor3_2 _7764_ (.A(net596),
    .B(net18),
    .C(_3019_),
    .Y(_3020_));
 sg13g2_a21o_1 _7765_ (.A2(net23),
    .A1(\i_dm_csrs.sbdata_o_9_ ),
    .B1(_3020_),
    .X(_0482_));
 sg13g2_a21oi_2 _7766_ (.B1(_2828_),
    .Y(_3021_),
    .A2(net803),
    .A1(_1326_));
 sg13g2_buf_8 fanout107 (.A(net111),
    .X(net107));
 sg13g2_buf_8 fanout106 (.A(net111),
    .X(net106));
 sg13g2_buf_8 fanout105 (.A(net111),
    .X(net105));
 sg13g2_nor3_2 _7770_ (.A(net790),
    .B(_0606_),
    .C(net11),
    .Y(_3025_));
 sg13g2_a21o_1 _7771_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_32_ ),
    .B1(_3025_),
    .X(_0483_));
 sg13g2_nor3_2 _7772_ (.A(net790),
    .B(_0655_),
    .C(net11),
    .Y(_3026_));
 sg13g2_a21o_1 _7773_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_33_ ),
    .B1(_3026_),
    .X(_0484_));
 sg13g2_nor3_2 _7774_ (.A(net795),
    .B(_0679_),
    .C(net11),
    .Y(_3027_));
 sg13g2_a21o_1 _7775_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_34_ ),
    .B1(_3027_),
    .X(_0485_));
 sg13g2_nor3_2 _7776_ (.A(net793),
    .B(_0687_),
    .C(net11),
    .Y(_3028_));
 sg13g2_a21o_1 _7777_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_35_ ),
    .B1(_3028_),
    .X(_0486_));
 sg13g2_nor3_2 _7778_ (.A(net794),
    .B(_0690_),
    .C(net10),
    .Y(_3029_));
 sg13g2_a21o_1 _7779_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_36_ ),
    .B1(_3029_),
    .X(_0487_));
 sg13g2_nor3_2 _7780_ (.A(net794),
    .B(_0693_),
    .C(net10),
    .Y(_3030_));
 sg13g2_a21o_1 _7781_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_37_ ),
    .B1(_3030_),
    .X(_0488_));
 sg13g2_nor3_2 _7782_ (.A(net794),
    .B(_0696_),
    .C(net10),
    .Y(_3031_));
 sg13g2_a21o_1 _7783_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_38_ ),
    .B1(_3031_),
    .X(_0489_));
 sg13g2_nor3_2 _7784_ (.A(net793),
    .B(_0699_),
    .C(net10),
    .Y(_3032_));
 sg13g2_a21o_1 _7785_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_39_ ),
    .B1(_3032_),
    .X(_0490_));
 sg13g2_buf_8 fanout104 (.A(net111),
    .X(net104));
 sg13g2_nor3_2 _7787_ (.A(net794),
    .B(_0701_),
    .C(net12),
    .Y(_3034_));
 sg13g2_a21o_1 _7788_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_40_ ),
    .B1(_3034_),
    .X(_0491_));
 sg13g2_nor3_2 _7789_ (.A(net794),
    .B(_0703_),
    .C(net12),
    .Y(_3035_));
 sg13g2_a21o_1 _7790_ (.A2(net14),
    .A1(\i_dm_csrs.sbdata_q_41_ ),
    .B1(_3035_),
    .X(_0492_));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net111));
 sg13g2_buf_4 fanout102 (.X(net102),
    .A(net111));
 sg13g2_nor3_2 _7793_ (.A(net794),
    .B(_0631_),
    .C(net12),
    .Y(_3038_));
 sg13g2_a21o_1 _7794_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_42_ ),
    .B1(_3038_),
    .X(_0493_));
 sg13g2_nor3_2 _7795_ (.A(net794),
    .B(_0633_),
    .C(net12),
    .Y(_3039_));
 sg13g2_a21o_1 _7796_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_43_ ),
    .B1(_3039_),
    .X(_0494_));
 sg13g2_nor3_2 _7797_ (.A(net795),
    .B(_0635_),
    .C(net12),
    .Y(_3040_));
 sg13g2_a21o_1 _7798_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_44_ ),
    .B1(_3040_),
    .X(_0495_));
 sg13g2_nor3_2 _7799_ (.A(net795),
    .B(_2742_),
    .C(net12),
    .Y(_3041_));
 sg13g2_a21o_1 _7800_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_45_ ),
    .B1(_3041_),
    .X(_0496_));
 sg13g2_nor3_2 _7801_ (.A(net794),
    .B(_0638_),
    .C(net11),
    .Y(_3042_));
 sg13g2_a21o_1 _7802_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_46_ ),
    .B1(_3042_),
    .X(_0497_));
 sg13g2_nor3_2 _7803_ (.A(net795),
    .B(_0640_),
    .C(net11),
    .Y(_3043_));
 sg13g2_a21o_1 _7804_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_47_ ),
    .B1(_3043_),
    .X(_0498_));
 sg13g2_nor3_2 _7805_ (.A(net790),
    .B(_0643_),
    .C(net11),
    .Y(_3044_));
 sg13g2_a21o_1 _7806_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_48_ ),
    .B1(_3044_),
    .X(_0499_));
 sg13g2_nor3_2 _7807_ (.A(net790),
    .B(_0646_),
    .C(net11),
    .Y(_3045_));
 sg13g2_a21o_1 _7808_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_49_ ),
    .B1(_3045_),
    .X(_0500_));
 sg13g2_buf_1 fanout101 (.A(slave_addr_i_5_),
    .X(net101));
 sg13g2_nor3_2 _7810_ (.A(net790),
    .B(_0648_),
    .C(net13),
    .Y(_3047_));
 sg13g2_a21o_1 _7811_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_50_ ),
    .B1(_3047_),
    .X(_0501_));
 sg13g2_nor3_2 _7812_ (.A(net790),
    .B(_0650_),
    .C(net13),
    .Y(_3048_));
 sg13g2_a21o_1 _7813_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_51_ ),
    .B1(_3048_),
    .X(_0502_));
 sg13g2_buf_2 fanout100 (.A(slave_addr_i_5_),
    .X(net100));
 sg13g2_buf_2 fanout99 (.A(cmd_12_),
    .X(net99));
 sg13g2_nor3_2 _7816_ (.A(net791),
    .B(_0658_),
    .C(net13),
    .Y(_3051_));
 sg13g2_a21o_1 _7817_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_52_ ),
    .B1(_3051_),
    .X(_0503_));
 sg13g2_nor3_2 _7818_ (.A(net791),
    .B(_0660_),
    .C(net13),
    .Y(_3052_));
 sg13g2_a21o_1 _7819_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_53_ ),
    .B1(_3052_),
    .X(_0504_));
 sg13g2_nor3_2 _7820_ (.A(net791),
    .B(_0662_),
    .C(net13),
    .Y(_3053_));
 sg13g2_a21o_1 _7821_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_54_ ),
    .B1(_3053_),
    .X(_0505_));
 sg13g2_nor3_2 _7822_ (.A(net792),
    .B(_1163_),
    .C(net13),
    .Y(_3054_));
 sg13g2_a21o_1 _7823_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_55_ ),
    .B1(_3054_),
    .X(_0506_));
 sg13g2_nor3_2 _7824_ (.A(net791),
    .B(_0665_),
    .C(net13),
    .Y(_3055_));
 sg13g2_a21o_1 _7825_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_56_ ),
    .B1(_3055_),
    .X(_0507_));
 sg13g2_nor3_2 _7826_ (.A(net791),
    .B(_0667_),
    .C(net13),
    .Y(_3056_));
 sg13g2_a21o_1 _7827_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_57_ ),
    .B1(_3056_),
    .X(_0508_));
 sg13g2_nor3_2 _7828_ (.A(net792),
    .B(_0669_),
    .C(net12),
    .Y(_3057_));
 sg13g2_a21o_1 _7829_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_58_ ),
    .B1(_3057_),
    .X(_0509_));
 sg13g2_nor3_2 _7830_ (.A(net792),
    .B(_0671_),
    .C(net12),
    .Y(_3058_));
 sg13g2_a21o_1 _7831_ (.A2(net17),
    .A1(\i_dm_csrs.sbdata_q_59_ ),
    .B1(_3058_),
    .X(_0510_));
 sg13g2_nor3_2 _7832_ (.A(net796),
    .B(_0673_),
    .C(net10),
    .Y(_3059_));
 sg13g2_a21o_1 _7833_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_60_ ),
    .B1(_3059_),
    .X(_0511_));
 sg13g2_nor3_2 _7834_ (.A(net795),
    .B(_0675_),
    .C(net10),
    .Y(_3060_));
 sg13g2_a21o_1 _7835_ (.A2(net16),
    .A1(\i_dm_csrs.sbdata_q_61_ ),
    .B1(_3060_),
    .X(_0512_));
 sg13g2_nor3_2 _7836_ (.A(net790),
    .B(_0682_),
    .C(net10),
    .Y(_3061_));
 sg13g2_a21o_1 _7837_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_62_ ),
    .B1(_3061_),
    .X(_0513_));
 sg13g2_nor3_2 _7838_ (.A(net790),
    .B(_0684_),
    .C(net10),
    .Y(_3062_));
 sg13g2_a21o_1 _7839_ (.A2(net15),
    .A1(\i_dm_csrs.sbdata_q_63_ ),
    .B1(_3062_),
    .X(_0514_));
 sg13g2_a22oi_1 _7840_ (.Y(_3063_),
    .B1(_2546_),
    .B2(net223),
    .A2(net428),
    .A1(\i_dm_csrs.sbcs_q_20_ ));
 sg13g2_inv_1 _7841_ (.Y(_0515_),
    .A(_3063_));
 sg13g2_a22oi_1 _7842_ (.Y(_3064_),
    .B1(_2546_),
    .B2(net235),
    .A2(net428),
    .A1(\i_dm_csrs.sbcs_q_15_ ));
 sg13g2_inv_1 _7843_ (.Y(_0516_),
    .A(_3064_));
 sg13g2_buf_8 fanout98 (.A(dmactive_o),
    .X(net98));
 sg13g2_inv_1 _7845_ (.Y(_3066_),
    .A(net613));
 sg13g2_buf_16 fanout97 (.X(net97),
    .A(net98));
 sg13g2_buf_2 fanout96 (.A(net98),
    .X(net96));
 sg13g2_nand2_1 _7848_ (.Y(_3069_),
    .A(net643),
    .B(net103));
 sg13g2_o21ai_1 _7849_ (.B1(_3069_),
    .Y(_0517_),
    .A1(net643),
    .A2(net579));
 sg13g2_inv_1 _7850_ (.Y(_3070_),
    .A(net70));
 sg13g2_buf_4 fanout95 (.X(net95),
    .A(net96));
 sg13g2_nand2_1 _7852_ (.Y(_3072_),
    .A(net643),
    .B(net661));
 sg13g2_o21ai_1 _7853_ (.B1(_3072_),
    .Y(_0518_),
    .A1(net643),
    .A2(net578));
 sg13g2_buf_2 fanout94 (.A(net96),
    .X(net94));
 sg13g2_inv_1 _7855_ (.Y(_3074_),
    .A(net67));
 sg13g2_buf_4 fanout93 (.X(net93),
    .A(net96));
 sg13g2_buf_2 fanout92 (.A(net96),
    .X(net92));
 sg13g2_nand2_2 _7858_ (.Y(_3077_),
    .A(net642),
    .B(net100));
 sg13g2_o21ai_1 _7859_ (.B1(_3077_),
    .Y(_0519_),
    .A1(net642),
    .A2(net545));
 sg13g2_inv_1 _7860_ (.Y(_3078_),
    .A(net63));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net96));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net96));
 sg13g2_nand2_2 _7863_ (.Y(_3081_),
    .A(net642),
    .B(net645));
 sg13g2_o21ai_1 _7864_ (.B1(_3081_),
    .Y(_0520_),
    .A1(net642),
    .A2(net576));
 sg13g2_inv_1 _7865_ (.Y(_3082_),
    .A(net59));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net96));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(net96));
 sg13g2_nand2_1 _7868_ (.Y(_3085_),
    .A(net642),
    .B(slave_addr_i_7_));
 sg13g2_o21ai_1 _7869_ (.B1(_3085_),
    .Y(_0521_),
    .A1(net642),
    .A2(net574));
 sg13g2_inv_1 _7870_ (.Y(_3086_),
    .A(\i_dm_mem.rdata_q_0_ ));
 sg13g2_nand2_2 _7871_ (.Y(_3087_),
    .A(slave_addr_i_9_),
    .B(_0706_));
 sg13g2_nor4_2 _7872_ (.A(net102),
    .B(net657),
    .C(net567),
    .Y(_3088_),
    .D(_1136_));
 sg13g2_a21oi_1 _7873_ (.A1(slave_addr_i_9_),
    .A2(net555),
    .Y(_3089_),
    .B1(slave_addr_i_10_));
 sg13g2_nor2_1 _7874_ (.A(slave_addr_i_11_),
    .B(_3089_),
    .Y(_3090_));
 sg13g2_and2_2 _7875_ (.A(net102),
    .B(net656),
    .X(_3091_));
 sg13g2_buf_4 fanout87 (.X(net87),
    .A(net97));
 sg13g2_nand2_1 _7877_ (.Y(_3093_),
    .A(net101),
    .B(_3091_));
 sg13g2_inv_1 _7878_ (.Y(_3094_),
    .A(_3093_));
 sg13g2_and2_2 _7879_ (.A(_0707_),
    .B(_1135_),
    .X(_3095_));
 sg13g2_o21ai_1 _7880_ (.B1(_3095_),
    .Y(_3096_),
    .A1(net644),
    .A2(_3094_));
 sg13g2_nand2b_1 _7881_ (.Y(_3097_),
    .B(_3096_),
    .A_N(_3090_));
 sg13g2_nor2_1 _7882_ (.A(_1745_),
    .B(slave_wdata_i_0_),
    .Y(_3098_));
 sg13g2_or2_1 _7883_ (.X(_3099_),
    .B(\i_dm_mem.state_q_1_ ),
    .A(\i_dm_mem.state_q_0__$_NOT__A_Y ));
 sg13g2_a22oi_1 _7884_ (.Y(_3100_),
    .B1(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .B2(_3099_),
    .A2(\i_dm_mem.state_q_0__$_NOT__A_Y ),
    .A1(\i_dm_mem.state_q_0_ ));
 sg13g2_or2_1 _7885_ (.X(_3101_),
    .B(_3100_),
    .A(_3098_));
 sg13g2_inv_1 _7886_ (.Y(_3102_),
    .A(_3101_));
 sg13g2_nor2b_1 _7887_ (.A(slave_we_i),
    .B_N(net642),
    .Y(_3103_));
 sg13g2_inv_1 _7888_ (.Y(_3104_),
    .A(_3103_));
 sg13g2_a21oi_2 _7889_ (.B1(_3104_),
    .Y(_3105_),
    .A2(_3102_),
    .A1(net543));
 sg13g2_o21ai_1 _7890_ (.B1(_3105_),
    .Y(_3106_),
    .A1(net543),
    .A2(net388));
 sg13g2_buf_4 fanout86 (.X(net86),
    .A(net97));
 sg13g2_buf_2 fanout85 (.A(net97),
    .X(net85));
 sg13g2_and2_1 _7893_ (.A(_3105_),
    .B(net388),
    .X(_3109_));
 sg13g2_inv_1 _7894_ (.Y(_3110_),
    .A(net100));
 sg13g2_nor4_1 _7895_ (.A(cmd_19_),
    .B(net565),
    .C(_1197_),
    .D(_1205_),
    .Y(_3111_));
 sg13g2_nand2_1 _7896_ (.Y(_3112_),
    .A(net565),
    .B(net644));
 sg13g2_nor2_1 _7897_ (.A(net565),
    .B(net645),
    .Y(_3113_));
 sg13g2_nand2_1 _7898_ (.Y(_3114_),
    .A(_3091_),
    .B(_3113_));
 sg13g2_nand2_2 _7899_ (.Y(_3115_),
    .A(_0707_),
    .B(_1135_));
 sg13g2_a21oi_1 _7900_ (.A1(_3112_),
    .A2(_3114_),
    .Y(_3116_),
    .B1(_3115_));
 sg13g2_nand2b_1 _7901_ (.Y(_3117_),
    .B(net441),
    .A_N(_3111_));
 sg13g2_and2_1 _7902_ (.A(net1),
    .B(_3117_),
    .X(_3118_));
 sg13g2_buf_4 fanout84 (.X(net84),
    .A(net97));
 sg13g2_and3_1 _7904_ (.X(_3120_),
    .A(net100),
    .B(net644),
    .C(_1135_));
 sg13g2_buf_16 fanout83 (.X(net83),
    .A(net97));
 sg13g2_and2_1 _7906_ (.A(_0707_),
    .B(net564),
    .X(_3122_));
 sg13g2_buf_2 fanout82 (.A(net97),
    .X(net82));
 sg13g2_buf_2 fanout81 (.A(net97),
    .X(net81));
 sg13g2_buf_2 fanout80 (.A(net97),
    .X(net80));
 sg13g2_buf_2 fanout79 (.A(\i_dm_sba.sbaccess_mask_3__$_AND__B_A_$_AND__Y_A ),
    .X(net79));
 sg13g2_buf_1 fanout78 (.A(net79),
    .X(net78));
 sg13g2_buf_2 fanout77 (.A(net79),
    .X(net77));
 sg13g2_mux4_1 _7913_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_0_ ),
    .A1(\i_dm_csrs.progbuf_o_64_ ),
    .A2(\i_dm_csrs.progbuf_o_128_ ),
    .A3(\i_dm_csrs.progbuf_o_192_ ),
    .S1(net662),
    .X(_3129_));
 sg13g2_nand2b_1 _7914_ (.Y(_3130_),
    .B(slave_addr_i_10_),
    .A_N(slave_addr_i_8_));
 sg13g2_nor4_2 _7915_ (.A(ndmreset_o),
    .B(slave_addr_i_7_),
    .C(_1132_),
    .Y(_3131_),
    .D(_3130_));
 sg13g2_nand2_1 _7916_ (.Y(_3132_),
    .A(_0709_),
    .B(_3131_));
 sg13g2_nor2_1 _7917_ (.A(_3099_),
    .B(_3132_),
    .Y(_3133_));
 sg13g2_a221oi_1 _7918_ (.B2(_3129_),
    .C1(_3133_),
    .B1(net501),
    .A1(data_csrs_mem_0_),
    .Y(_3134_),
    .A2(net35));
 sg13g2_a22oi_1 _7919_ (.Y(_0522_),
    .B1(_3118_),
    .B2(_3134_),
    .A2(net7),
    .A1(_3086_));
 sg13g2_nand2_1 _7920_ (.Y(_3135_),
    .A(_3105_),
    .B(net388));
 sg13g2_nor2b_2 _7921_ (.A(net109),
    .B_N(net657),
    .Y(_3136_));
 sg13g2_nor2b_2 _7922_ (.A(net101),
    .B_N(net645),
    .Y(_3137_));
 sg13g2_nand2_2 _7923_ (.Y(_3138_),
    .A(_3095_),
    .B(_3137_));
 sg13g2_nor3_1 _7924_ (.A(net277),
    .B(_3136_),
    .C(_3138_),
    .Y(_3139_));
 sg13g2_nand4_1 _7925_ (.B(cmd_17_),
    .C(_1199_),
    .A(cmd_16_),
    .Y(_3140_),
    .D(_1204_));
 sg13g2_nor2_2 _7926_ (.A(_1195_),
    .B(_3140_),
    .Y(_3141_));
 sg13g2_nand2_2 _7927_ (.Y(_3142_),
    .A(net549),
    .B(_3141_));
 sg13g2_nor4_1 _7928_ (.A(cmd_0_),
    .B(\cmd_0__$_OR__A_B ),
    .C(cmd_4_),
    .D(cmd_2_),
    .Y(_3143_));
 sg13g2_nand3b_1 _7929_ (.B(\cmd_5__$_NOT__A_Y ),
    .C(_3143_),
    .Y(_3144_),
    .A_N(\cmd_3__$_NOT__A_Y ));
 sg13g2_and2_2 _7930_ (.A(net99),
    .B(_3144_),
    .X(_3145_));
 sg13g2_nand2_1 _7931_ (.Y(_3146_),
    .A(cmd_3_),
    .B(_3145_));
 sg13g2_inv_1 _7932_ (.Y(_3147_),
    .A(net102));
 sg13g2_nor2_2 _7933_ (.A(net558),
    .B(net658),
    .Y(_3148_));
 sg13g2_o21ai_1 _7934_ (.B1(_3148_),
    .Y(_3149_),
    .A1(_3142_),
    .A2(_3146_));
 sg13g2_buf_2 fanout76 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_1_ ),
    .X(net76));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(net76));
 sg13g2_mux4_1 _7938_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_10_ ),
    .A1(\i_dm_csrs.progbuf_o_74_ ),
    .A2(\i_dm_csrs.progbuf_o_138_ ),
    .A3(\i_dm_csrs.progbuf_o_202_ ),
    .S1(net652),
    .X(_3153_));
 sg13g2_a22oi_1 _7939_ (.Y(_3154_),
    .B1(net562),
    .B2(_3153_),
    .A2(net553),
    .A1(data_csrs_mem_10_));
 sg13g2_nand3_1 _7940_ (.B(_3105_),
    .C(net388),
    .A(_0707_),
    .Y(_3155_));
 sg13g2_nor2_1 _7941_ (.A(_3154_),
    .B(_3155_),
    .Y(_3156_));
 sg13g2_a221oi_1 _7942_ (.B2(_3149_),
    .C1(_3156_),
    .B1(_3139_),
    .A1(\i_dm_mem.rdata_q_10_ ),
    .Y(_3157_),
    .A2(net6));
 sg13g2_inv_1 _7943_ (.Y(_0523_),
    .A(_3157_));
 sg13g2_inv_1 _7944_ (.Y(_3158_),
    .A(net99));
 sg13g2_buf_2 fanout73 (.A(net76),
    .X(net73));
 sg13g2_nand2b_2 _7946_ (.Y(_3160_),
    .B(net102),
    .A_N(net656));
 sg13g2_nor4_2 _7947_ (.A(net39),
    .B(_3138_),
    .C(_3160_),
    .Y(_3161_),
    .D(_3142_));
 sg13g2_nand2_1 _7948_ (.Y(_3162_),
    .A(cmd_4_),
    .B(_3161_));
 sg13g2_buf_2 fanout72 (.A(net76),
    .X(net72));
 sg13g2_mux4_1 _7950_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_11_ ),
    .A1(\i_dm_csrs.progbuf_o_75_ ),
    .A2(\i_dm_csrs.progbuf_o_139_ ),
    .A3(\i_dm_csrs.progbuf_o_203_ ),
    .S1(net651),
    .X(_3164_));
 sg13g2_a22oi_1 _7951_ (.Y(_3165_),
    .B1(net500),
    .B2(_3164_),
    .A2(net36),
    .A1(data_csrs_mem_11_));
 sg13g2_a21oi_1 _7952_ (.A1(_3162_),
    .A2(_3165_),
    .Y(_3166_),
    .B1(net275));
 sg13g2_a21o_1 _7953_ (.A2(net7),
    .A1(\i_dm_mem.rdata_q_11_ ),
    .B1(_3166_),
    .X(_0524_));
 sg13g2_nand2_2 _7954_ (.Y(_3167_),
    .A(_1200_),
    .B(_1201_));
 sg13g2_or2_2 _7955_ (.X(_3168_),
    .B(_3140_),
    .A(_1195_));
 sg13g2_nor2_2 _7956_ (.A(_3167_),
    .B(_3168_),
    .Y(_3169_));
 sg13g2_nor2_2 _7957_ (.A(net39),
    .B(_3144_),
    .Y(_3170_));
 sg13g2_or2_2 _7958_ (.X(_3171_),
    .B(net497),
    .A(\i_dm_mem.abstract_cmd_132__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ));
 sg13g2_buf_2 fanout71 (.A(net76),
    .X(net71));
 sg13g2_inv_1 _7960_ (.Y(_3173_),
    .A(\cmd_16__$_NOT__A_Y ));
 sg13g2_nor2_1 _7961_ (.A(cmd_14_),
    .B(cmd_15_),
    .Y(_3174_));
 sg13g2_nand4_1 _7962_ (.B(_1199_),
    .C(_3174_),
    .A(cmd_17_),
    .Y(_3175_),
    .D(_1204_));
 sg13g2_nor3_2 _7963_ (.A(cmd_16_),
    .B(_3173_),
    .C(_3175_),
    .Y(_3176_));
 sg13g2_nand2_2 _7964_ (.Y(_3177_),
    .A(net549),
    .B(_3176_));
 sg13g2_nor2_1 _7965_ (.A(_3145_),
    .B(_3177_),
    .Y(_3178_));
 sg13g2_nand2_1 _7966_ (.Y(_3179_),
    .A(net558),
    .B(net658));
 sg13g2_a221oi_1 _7967_ (.B2(cmd_20_),
    .C1(_3179_),
    .B1(_3178_),
    .A1(_3169_),
    .Y(_3180_),
    .A2(_3171_));
 sg13g2_nor2_2 _7968_ (.A(_1196_),
    .B(_3175_),
    .Y(_3181_));
 sg13g2_nand2_2 _7969_ (.Y(_3182_),
    .A(net549),
    .B(_3181_));
 sg13g2_buf_2 fanout70 (.A(net76),
    .X(net70));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2_ ));
 sg13g2_nand2_2 _7972_ (.Y(_3185_),
    .A(cmd_12_),
    .B(_3144_));
 sg13g2_nor3_1 _7973_ (.A(cmd_20_),
    .B(net658),
    .C(_3185_),
    .Y(_3186_));
 sg13g2_o21ai_1 _7974_ (.B1(net110),
    .Y(_3187_),
    .A1(_3182_),
    .A2(_3186_));
 sg13g2_o21ai_1 _7975_ (.B1(_3114_),
    .Y(_3188_),
    .A1(_3091_),
    .A2(_3112_));
 sg13g2_and2_2 _7976_ (.A(_3095_),
    .B(_3188_),
    .X(_3189_));
 sg13g2_nand3_1 _7977_ (.B(_3187_),
    .C(_3189_),
    .A(net2),
    .Y(_3190_));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2_ ));
 sg13g2_buf_2 fanout67 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2_ ),
    .X(net67));
 sg13g2_mux4_1 _7980_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_12_ ),
    .A1(\i_dm_csrs.progbuf_o_76_ ),
    .A2(\i_dm_csrs.progbuf_o_140_ ),
    .A3(\i_dm_csrs.progbuf_o_204_ ),
    .S1(net647),
    .X(_3193_));
 sg13g2_a22oi_1 _7981_ (.Y(_3194_),
    .B1(net559),
    .B2(_3193_),
    .A2(net550),
    .A1(data_csrs_mem_12_));
 sg13g2_nor2_1 _7982_ (.A(net568),
    .B(_3194_),
    .Y(_3195_));
 sg13g2_a22oi_1 _7983_ (.Y(_3196_),
    .B1(net2),
    .B2(_3195_),
    .A2(net6),
    .A1(\i_dm_mem.rdata_q_12_ ));
 sg13g2_o21ai_1 _7984_ (.B1(_3196_),
    .Y(_0525_),
    .A1(_3180_),
    .A2(_3190_));
 sg13g2_nand2_1 _7985_ (.Y(_3197_),
    .A(net543),
    .B(_3105_));
 sg13g2_a21oi_1 _7986_ (.A1(\i_dm_mem.rdata_q_13_ ),
    .A2(_3197_),
    .Y(_3198_),
    .B1(net2));
 sg13g2_buf_2 fanout66 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3_ ),
    .X(net66));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65));
 sg13g2_mux4_1 _7989_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_13_ ),
    .A1(\i_dm_csrs.progbuf_o_77_ ),
    .A2(\i_dm_csrs.progbuf_o_141_ ),
    .A3(\i_dm_csrs.progbuf_o_205_ ),
    .S1(net646),
    .X(_3201_));
 sg13g2_a22oi_1 _7990_ (.Y(_3202_),
    .B1(net561),
    .B2(_3201_),
    .A2(net552),
    .A1(data_csrs_mem_13_));
 sg13g2_nor2_1 _7991_ (.A(net568),
    .B(_3202_),
    .Y(_3203_));
 sg13g2_buf_2 fanout64 (.A(net66),
    .X(net64));
 sg13g2_and2_1 _7993_ (.A(cmd_21_),
    .B(net658),
    .X(_3205_));
 sg13g2_a21oi_1 _7994_ (.A1(_3178_),
    .A2(_3205_),
    .Y(_3206_),
    .B1(net103));
 sg13g2_nor2_1 _7995_ (.A(_3185_),
    .B(_3182_),
    .Y(_3207_));
 sg13g2_a21oi_1 _7996_ (.A1(cmd_21_),
    .A2(_3207_),
    .Y(_3208_),
    .B1(net658));
 sg13g2_nor3_1 _7997_ (.A(_3138_),
    .B(_3206_),
    .C(_3208_),
    .Y(_3209_));
 sg13g2_nor3_1 _7998_ (.A(net3),
    .B(_3203_),
    .C(_3209_),
    .Y(_3210_));
 sg13g2_nor2_1 _7999_ (.A(_3198_),
    .B(_3210_),
    .Y(_0526_));
 sg13g2_buf_2 fanout63 (.A(net66),
    .X(net63));
 sg13g2_nor3_1 _8001_ (.A(net660),
    .B(_3185_),
    .C(_3182_),
    .Y(_3212_));
 sg13g2_nor3_1 _8002_ (.A(net102),
    .B(_3145_),
    .C(_3177_),
    .Y(_3213_));
 sg13g2_o21ai_1 _8003_ (.B1(cmd_22_),
    .Y(_3214_),
    .A1(_3212_),
    .A2(_3213_));
 sg13g2_o21ai_1 _8004_ (.B1(_3214_),
    .Y(_3215_),
    .A1(net103),
    .A2(net656));
 sg13g2_buf_2 fanout62 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ),
    .X(net62));
 sg13g2_buf_4 fanout61 (.X(net61),
    .A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ));
 sg13g2_mux4_1 _8007_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_14_ ),
    .A1(\i_dm_csrs.progbuf_o_78_ ),
    .A2(\i_dm_csrs.progbuf_o_142_ ),
    .A3(\i_dm_csrs.progbuf_o_206_ ),
    .S1(net653),
    .X(_3218_));
 sg13g2_a22oi_1 _8008_ (.Y(_3219_),
    .B1(net564),
    .B2(_3218_),
    .A2(net555),
    .A1(data_csrs_mem_14_));
 sg13g2_nor2_1 _8009_ (.A(net566),
    .B(_3219_),
    .Y(_3220_));
 sg13g2_a21oi_2 _8010_ (.B1(_3220_),
    .Y(_3221_),
    .A2(_3215_),
    .A1(_3189_));
 sg13g2_buf_2 fanout60 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ),
    .X(net60));
 sg13g2_nand2_1 _8012_ (.Y(_3223_),
    .A(\i_dm_mem.rdata_q_14_ ),
    .B(net4));
 sg13g2_o21ai_1 _8013_ (.B1(_3223_),
    .Y(_0527_),
    .A1(net275),
    .A2(_3221_));
 sg13g2_nor2_1 _8014_ (.A(net543),
    .B(net388),
    .Y(_3224_));
 sg13g2_nor2b_2 _8015_ (.A(_3224_),
    .B_N(_3105_),
    .Y(_3225_));
 sg13g2_buf_2 fanout59 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ),
    .X(net59));
 sg13g2_buf_2 fanout58 (.A(\i_dm_mem.word_enable32_q ),
    .X(net58));
 sg13g2_buf_4 fanout57 (.X(net57),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_mux4_1 _8019_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_15_ ),
    .A1(\i_dm_csrs.progbuf_o_79_ ),
    .A2(\i_dm_csrs.progbuf_o_143_ ),
    .A3(\i_dm_csrs.progbuf_o_207_ ),
    .S1(net648),
    .X(_3229_));
 sg13g2_a22oi_1 _8020_ (.Y(_3230_),
    .B1(net501),
    .B2(_3229_),
    .A2(net37),
    .A1(data_csrs_mem_15_));
 sg13g2_buf_4 fanout56 (.X(net56),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_nor2_1 _8022_ (.A(\i_dm_mem.rdata_q_15_ ),
    .B(net247),
    .Y(_3232_));
 sg13g2_a21oi_1 _8023_ (.A1(net247),
    .A2(_3230_),
    .Y(_0528_),
    .B1(_3232_));
 sg13g2_buf_4 fanout55 (.X(net55),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_nor2_2 _8025_ (.A(\i_dm_mem.abstract_cmd_132__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ),
    .B(_3170_),
    .Y(_3234_));
 sg13g2_o21ai_1 _8026_ (.B1(net659),
    .Y(_3235_),
    .A1(_3234_),
    .A2(_3177_));
 sg13g2_nand2_1 _8027_ (.Y(_3236_),
    .A(_3095_),
    .B(_3188_));
 sg13g2_nor2_1 _8028_ (.A(net103),
    .B(_3236_),
    .Y(_3237_));
 sg13g2_buf_4 fanout54 (.X(net54),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_buf_4 fanout53 (.X(net53),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_mux4_1 _8031_ (.S0(net108),
    .A0(\i_dm_csrs.progbuf_o_16_ ),
    .A1(\i_dm_csrs.progbuf_o_80_ ),
    .A2(\i_dm_csrs.progbuf_o_144_ ),
    .A3(\i_dm_csrs.progbuf_o_208_ ),
    .S1(net652),
    .X(_3240_));
 sg13g2_a22oi_1 _8032_ (.Y(_3241_),
    .B1(net562),
    .B2(_3240_),
    .A2(net553),
    .A1(data_csrs_mem_16_));
 sg13g2_buf_4 fanout52 (.X(net52),
    .A(\i_dm_mem.word_enable32_q ));
 sg13g2_or2_1 _8034_ (.X(_3243_),
    .B(_3175_),
    .A(_1196_));
 sg13g2_nand3_1 _8035_ (.B(net645),
    .C(_1193_),
    .A(_3110_),
    .Y(_3244_));
 sg13g2_o21ai_1 _8036_ (.B1(_3244_),
    .Y(_3245_),
    .A1(net644),
    .A2(_3093_));
 sg13g2_nand3_1 _8037_ (.B(_3095_),
    .C(_3245_),
    .A(net549),
    .Y(_3246_));
 sg13g2_nor3_1 _8038_ (.A(net558),
    .B(_3243_),
    .C(_3246_),
    .Y(_3247_));
 sg13g2_o21ai_1 _8039_ (.B1(_3247_),
    .Y(_3248_),
    .A1(net659),
    .A2(_3145_));
 sg13g2_o21ai_1 _8040_ (.B1(_3248_),
    .Y(_3249_),
    .A1(net567),
    .A2(_3241_));
 sg13g2_a21oi_1 _8041_ (.A1(_3235_),
    .A2(_3237_),
    .Y(_3250_),
    .B1(_3249_));
 sg13g2_nand2_1 _8042_ (.Y(_3251_),
    .A(\i_dm_mem.rdata_q_16_ ),
    .B(net4));
 sg13g2_o21ai_1 _8043_ (.B1(_3251_),
    .Y(_0529_),
    .A1(net273),
    .A2(_3250_));
 sg13g2_mux4_1 _8044_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_17_ ),
    .A1(\i_dm_csrs.progbuf_o_81_ ),
    .A2(\i_dm_csrs.progbuf_o_145_ ),
    .A3(\i_dm_csrs.progbuf_o_209_ ),
    .S1(net650),
    .X(_3252_));
 sg13g2_a22oi_1 _8045_ (.Y(_3253_),
    .B1(net501),
    .B2(_3252_),
    .A2(net37),
    .A1(data_csrs_mem_17_));
 sg13g2_nor2_1 _8046_ (.A(\i_dm_mem.rdata_q_17_ ),
    .B(net248),
    .Y(_3254_));
 sg13g2_a21oi_1 _8047_ (.A1(net247),
    .A2(_3253_),
    .Y(_0530_),
    .B1(_3254_));
 sg13g2_nor2_1 _8048_ (.A(_3167_),
    .B(_3243_),
    .Y(_3255_));
 sg13g2_o21ai_1 _8049_ (.B1(_3255_),
    .Y(_3256_),
    .A1(net102),
    .A2(_3171_));
 sg13g2_o21ai_1 _8050_ (.B1(_3256_),
    .Y(_3257_),
    .A1(net103),
    .A2(net658));
 sg13g2_nand3_1 _8051_ (.B(_3189_),
    .C(_3257_),
    .A(net2),
    .Y(_3258_));
 sg13g2_mux4_1 _8052_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_18_ ),
    .A1(\i_dm_csrs.progbuf_o_82_ ),
    .A2(\i_dm_csrs.progbuf_o_146_ ),
    .A3(\i_dm_csrs.progbuf_o_210_ ),
    .S1(net650),
    .X(_3259_));
 sg13g2_a22oi_1 _8053_ (.Y(_3260_),
    .B1(net562),
    .B2(_3259_),
    .A2(net553),
    .A1(data_csrs_mem_18_));
 sg13g2_nor2_1 _8054_ (.A(_3155_),
    .B(_3260_),
    .Y(_3261_));
 sg13g2_a21oi_1 _8055_ (.A1(\i_dm_mem.rdata_q_18_ ),
    .A2(net6),
    .Y(_3262_),
    .B1(_3261_));
 sg13g2_nand2_1 _8056_ (.Y(_0531_),
    .A(_3258_),
    .B(_3262_));
 sg13g2_mux4_1 _8057_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_19_ ),
    .A1(\i_dm_csrs.progbuf_o_83_ ),
    .A2(\i_dm_csrs.progbuf_o_147_ ),
    .A3(\i_dm_csrs.progbuf_o_211_ ),
    .S1(net650),
    .X(_3263_));
 sg13g2_a22oi_1 _8058_ (.Y(_3264_),
    .B1(net501),
    .B2(_3263_),
    .A2(net37),
    .A1(data_csrs_mem_19_));
 sg13g2_nor2_1 _8059_ (.A(\i_dm_mem.rdata_q_19_ ),
    .B(net248),
    .Y(_3265_));
 sg13g2_a21oi_1 _8060_ (.A1(net247),
    .A2(_3264_),
    .Y(_0532_),
    .B1(_3265_));
 sg13g2_inv_1 _8061_ (.Y(_3266_),
    .A(\i_dm_mem.rdata_q_1_ ));
 sg13g2_mux4_1 _8062_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_1_ ),
    .A1(\i_dm_csrs.progbuf_o_65_ ),
    .A2(\i_dm_csrs.progbuf_o_129_ ),
    .A3(\i_dm_csrs.progbuf_o_193_ ),
    .S1(net653),
    .X(_3267_));
 sg13g2_nor3_1 _8063_ (.A(\i_dm_mem.state_q_0_ ),
    .B(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .C(_3132_),
    .Y(_3268_));
 sg13g2_a221oi_1 _8064_ (.B2(_3267_),
    .C1(_3268_),
    .B1(net499),
    .A1(data_csrs_mem_1_),
    .Y(_3269_),
    .A2(net35));
 sg13g2_a22oi_1 _8065_ (.Y(_0533_),
    .B1(_3118_),
    .B2(_3269_),
    .A2(net7),
    .A1(_3266_));
 sg13g2_mux4_1 _8066_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_20_ ),
    .A1(\i_dm_csrs.progbuf_o_84_ ),
    .A2(\i_dm_csrs.progbuf_o_148_ ),
    .A3(\i_dm_csrs.progbuf_o_212_ ),
    .S1(net646),
    .X(_3270_));
 sg13g2_a22oi_1 _8067_ (.Y(_3271_),
    .B1(net560),
    .B2(_3270_),
    .A2(net551),
    .A1(data_csrs_mem_20_));
 sg13g2_nand2b_1 _8068_ (.Y(_3272_),
    .B(_3091_),
    .A_N(_3111_));
 sg13g2_inv_1 _8069_ (.Y(_3273_),
    .A(_3272_));
 sg13g2_a21o_1 _8070_ (.A2(net40),
    .A1(cmd_0_),
    .B1(net497),
    .X(_3274_));
 sg13g2_nand3_1 _8071_ (.B(_3141_),
    .C(_3274_),
    .A(_3136_),
    .Y(_3275_));
 sg13g2_nand4_1 _8072_ (.B(net99),
    .C(_3148_),
    .A(cmd_0_),
    .Y(_3276_),
    .D(_3176_));
 sg13g2_a21oi_1 _8073_ (.A1(_3275_),
    .A2(_3276_),
    .Y(_3277_),
    .B1(_3167_));
 sg13g2_o21ai_1 _8074_ (.B1(net441),
    .Y(_3278_),
    .A1(_3273_),
    .A2(_3277_));
 sg13g2_o21ai_1 _8075_ (.B1(_3278_),
    .Y(_3279_),
    .A1(net569),
    .A2(_3271_));
 sg13g2_a22oi_1 _8076_ (.Y(_3280_),
    .B1(net2),
    .B2(_3279_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_20_ ));
 sg13g2_inv_1 _8077_ (.Y(_0534_),
    .A(_3280_));
 sg13g2_nand2_1 _8078_ (.Y(_3281_),
    .A(_3091_),
    .B(net441));
 sg13g2_a21oi_1 _8079_ (.A1(net101),
    .A2(_3182_),
    .Y(_3282_),
    .B1(_3281_));
 sg13g2_mux4_1 _8080_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_21_ ),
    .A1(\i_dm_csrs.progbuf_o_85_ ),
    .A2(\i_dm_csrs.progbuf_o_149_ ),
    .A3(\i_dm_csrs.progbuf_o_213_ ),
    .S1(net646),
    .X(_3283_));
 sg13g2_a22oi_1 _8081_ (.Y(_3284_),
    .B1(net560),
    .B2(_3283_),
    .A2(net551),
    .A1(data_csrs_mem_21_));
 sg13g2_nor2_1 _8082_ (.A(net566),
    .B(_3284_),
    .Y(_3285_));
 sg13g2_nand2b_1 _8083_ (.Y(_3286_),
    .B(_3145_),
    .A_N(cmd_1_));
 sg13g2_a22oi_1 _8084_ (.Y(_3287_),
    .B1(_3176_),
    .B2(_3286_),
    .A2(_3171_),
    .A1(_3141_));
 sg13g2_nor4_1 _8085_ (.A(_3167_),
    .B(_3160_),
    .C(_3236_),
    .D(_3287_),
    .Y(_3288_));
 sg13g2_nand3_1 _8086_ (.B(net441),
    .C(_3136_),
    .A(net549),
    .Y(_3289_));
 sg13g2_a21oi_1 _8087_ (.A1(net40),
    .A2(cmd_1_),
    .Y(_3290_),
    .B1(net497));
 sg13g2_nor2_1 _8088_ (.A(_3110_),
    .B(_3091_),
    .Y(_3291_));
 sg13g2_nor4_1 _8089_ (.A(_3168_),
    .B(_3289_),
    .C(_3290_),
    .D(_3291_),
    .Y(_3292_));
 sg13g2_nor4_2 _8090_ (.A(_3282_),
    .B(_3285_),
    .C(_3288_),
    .Y(_3293_),
    .D(_3292_));
 sg13g2_nand2_1 _8091_ (.Y(_3294_),
    .A(\i_dm_mem.rdata_q_21_ ),
    .B(net4));
 sg13g2_o21ai_1 _8092_ (.B1(_3294_),
    .Y(_0535_),
    .A1(net273),
    .A2(_3293_));
 sg13g2_buf_8 fanout51 (.A(master_add_o_0_),
    .X(net51));
 sg13g2_buf_8 fanout50 (.A(master_add_o_2_),
    .X(net50));
 sg13g2_nand2_1 _8095_ (.Y(_3297_),
    .A(net654),
    .B(\i_dm_csrs.progbuf_o_214_ ));
 sg13g2_o21ai_1 _8096_ (.B1(_3297_),
    .Y(_3298_),
    .A1(net654),
    .A2(_2507_));
 sg13g2_nor3_1 _8097_ (.A(net104),
    .B(net654),
    .C(_2280_),
    .Y(_3299_));
 sg13g2_a21o_1 _8098_ (.A2(_3298_),
    .A1(net109),
    .B1(_3299_),
    .X(_3300_));
 sg13g2_a22oi_1 _8099_ (.Y(_3301_),
    .B1(net564),
    .B2(_3300_),
    .A2(net555),
    .A1(data_csrs_mem_22_));
 sg13g2_nor2_1 _8100_ (.A(net567),
    .B(_3301_),
    .Y(_3302_));
 sg13g2_nor2_2 _8101_ (.A(_3115_),
    .B(_3112_),
    .Y(_3303_));
 sg13g2_nand2b_1 _8102_ (.Y(_3304_),
    .B(_3303_),
    .A_N(net657));
 sg13g2_nand2_1 _8103_ (.Y(_3305_),
    .A(net109),
    .B(\i_dm_csrs.progbuf_o_86_ ));
 sg13g2_o21ai_1 _8104_ (.B1(_3305_),
    .Y(_3306_),
    .A1(net107),
    .A2(_2280_));
 sg13g2_or2_1 _8105_ (.X(_3307_),
    .B(_3306_),
    .A(net661));
 sg13g2_nand3_1 _8106_ (.B(net498),
    .C(_3307_),
    .A(\i_dm_csrs.progbuf_o_150_ ),
    .Y(_3308_));
 sg13g2_a21oi_1 _8107_ (.A1(_3304_),
    .A2(_3308_),
    .Y(_3309_),
    .B1(net103));
 sg13g2_nor2_1 _8108_ (.A(net660),
    .B(net101),
    .Y(_3310_));
 sg13g2_nand4_1 _8109_ (.B(cmd_2_),
    .C(net441),
    .A(net99),
    .Y(_3311_),
    .D(_3310_));
 sg13g2_nor3_2 _8110_ (.A(net107),
    .B(_3167_),
    .C(_3168_),
    .Y(_3312_));
 sg13g2_nor2_1 _8111_ (.A(net99),
    .B(_3138_),
    .Y(_3313_));
 sg13g2_nand3_1 _8112_ (.B(_3312_),
    .C(_3313_),
    .A(cmd_2_),
    .Y(_3314_));
 sg13g2_o21ai_1 _8113_ (.B1(_3314_),
    .Y(_3315_),
    .A1(_3177_),
    .A2(_3311_));
 sg13g2_nor3_1 _8114_ (.A(_3302_),
    .B(_3309_),
    .C(_3315_),
    .Y(_3316_));
 sg13g2_nand2_1 _8115_ (.Y(_3317_),
    .A(\i_dm_mem.rdata_q_22_ ),
    .B(net4));
 sg13g2_o21ai_1 _8116_ (.B1(_3317_),
    .Y(_0536_),
    .A1(net273),
    .A2(_3316_));
 sg13g2_inv_1 _8117_ (.Y(_3318_),
    .A(\i_dm_mem.rdata_q_23_ ));
 sg13g2_nand4_1 _8118_ (.B(net549),
    .C(_3171_),
    .A(net557),
    .Y(_3319_),
    .D(_3176_));
 sg13g2_nor2_1 _8119_ (.A(net99),
    .B(_3168_),
    .Y(_3320_));
 sg13g2_nand4_1 _8120_ (.B(net557),
    .C(net549),
    .A(cmd_3_),
    .Y(_3321_),
    .D(_3320_));
 sg13g2_nand3_1 _8121_ (.B(_3319_),
    .C(_3321_),
    .A(net658),
    .Y(_3322_));
 sg13g2_o21ai_1 _8122_ (.B1(net110),
    .Y(_3323_),
    .A1(_3146_),
    .A2(_3177_));
 sg13g2_nand3_1 _8123_ (.B(_3322_),
    .C(_3323_),
    .A(_3189_),
    .Y(_3324_));
 sg13g2_mux4_1 _8124_ (.S0(net102),
    .A0(\i_dm_csrs.progbuf_o_23_ ),
    .A1(\i_dm_csrs.progbuf_o_87_ ),
    .A2(\i_dm_csrs.progbuf_o_151_ ),
    .A3(\i_dm_csrs.progbuf_o_215_ ),
    .S1(net654),
    .X(_3325_));
 sg13g2_a221oi_1 _8125_ (.B2(_3325_),
    .C1(net278),
    .B1(net499),
    .A1(data_csrs_mem_23_),
    .Y(_3326_),
    .A2(net36));
 sg13g2_nand3_1 _8126_ (.B(cmd_18_),
    .C(net549),
    .A(\cmd_17__$_NOT__A_Y ),
    .Y(_3327_));
 sg13g2_nor4_1 _8127_ (.A(net556),
    .B(net388),
    .C(_3197_),
    .D(_3327_),
    .Y(_3328_));
 sg13g2_a221oi_1 _8128_ (.B2(_3326_),
    .C1(_3328_),
    .B1(_3324_),
    .A1(_3318_),
    .Y(_0537_),
    .A2(net7));
 sg13g2_nor2b_2 _8129_ (.A(_3090_),
    .B_N(_3096_),
    .Y(_3329_));
 sg13g2_nand2_1 _8130_ (.Y(_3330_),
    .A(_0900_),
    .B(_3327_));
 sg13g2_nand3_1 _8131_ (.B(_3105_),
    .C(_3330_),
    .A(_3088_),
    .Y(_3331_));
 sg13g2_o21ai_1 _8132_ (.B1(_3331_),
    .Y(_3332_),
    .A1(\i_dm_mem.rdata_q_24_ ),
    .A2(_3088_));
 sg13g2_nand2_1 _8133_ (.Y(_3333_),
    .A(_3148_),
    .B(_3176_));
 sg13g2_a21oi_1 _8134_ (.A1(net40),
    .A2(_3333_),
    .Y(_3334_),
    .B1(_3145_));
 sg13g2_nand3_1 _8135_ (.B(_3141_),
    .C(_3185_),
    .A(_3136_),
    .Y(_3335_));
 sg13g2_a21oi_1 _8136_ (.A1(_3333_),
    .A2(_3335_),
    .Y(_3336_),
    .B1(_3246_));
 sg13g2_o21ai_1 _8137_ (.B1(_3336_),
    .Y(_3337_),
    .A1(cmd_4_),
    .A2(_3334_));
 sg13g2_nor3_1 _8138_ (.A(net659),
    .B(_3168_),
    .C(_3234_),
    .Y(_3338_));
 sg13g2_a21oi_1 _8139_ (.A1(net659),
    .A2(_3181_),
    .Y(_3339_),
    .B1(_3338_));
 sg13g2_nor3_1 _8140_ (.A(net557),
    .B(_3246_),
    .C(_3339_),
    .Y(_3340_));
 sg13g2_mux4_1 _8141_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_24_ ),
    .A1(\i_dm_csrs.progbuf_o_88_ ),
    .A2(\i_dm_csrs.progbuf_o_152_ ),
    .A3(\i_dm_csrs.progbuf_o_216_ ),
    .S1(net647),
    .X(_3341_));
 sg13g2_a22oi_1 _8142_ (.Y(_3342_),
    .B1(net560),
    .B2(_3341_),
    .A2(net551),
    .A1(data_csrs_mem_24_));
 sg13g2_nand2_1 _8143_ (.Y(_3343_),
    .A(_3091_),
    .B(_3303_));
 sg13g2_and2_1 _8144_ (.A(net1),
    .B(_3343_),
    .X(_3344_));
 sg13g2_o21ai_1 _8145_ (.B1(_3344_),
    .Y(_3345_),
    .A1(net567),
    .A2(_3342_));
 sg13g2_nor2_1 _8146_ (.A(_3340_),
    .B(_3345_),
    .Y(_3346_));
 sg13g2_nor2_1 _8147_ (.A(\i_dm_mem.rdata_q_24_ ),
    .B(_3105_),
    .Y(_3347_));
 sg13g2_a221oi_1 _8148_ (.B2(_3346_),
    .C1(_3347_),
    .B1(_3337_),
    .A1(_3329_),
    .Y(_0538_),
    .A2(_3332_));
 sg13g2_nand4_1 _8149_ (.B(_3103_),
    .C(net543),
    .A(net556),
    .Y(_3348_),
    .D(_3098_));
 sg13g2_nor2_1 _8150_ (.A(net388),
    .B(_3348_),
    .Y(_3349_));
 sg13g2_nand2_2 _8151_ (.Y(_3350_),
    .A(_3179_),
    .B(_3160_));
 sg13g2_nor2_2 _8152_ (.A(net558),
    .B(net565),
    .Y(_3351_));
 sg13g2_nor2b_1 _8153_ (.A(net644),
    .B_N(net657),
    .Y(_3352_));
 sg13g2_a22oi_1 _8154_ (.Y(_3353_),
    .B1(_3351_),
    .B2(_3352_),
    .A2(_3350_),
    .A1(_3137_));
 sg13g2_nor2_1 _8155_ (.A(_3115_),
    .B(_3353_),
    .Y(_3354_));
 sg13g2_a21oi_1 _8156_ (.A1(net39),
    .A2(cmd_5_),
    .Y(_3355_),
    .B1(net497));
 sg13g2_nand2b_1 _8157_ (.Y(_3356_),
    .B(_3312_),
    .A_N(_3355_));
 sg13g2_nand2_1 _8158_ (.Y(_3357_),
    .A(_3303_),
    .B(_3350_));
 sg13g2_o21ai_1 _8159_ (.B1(net109),
    .Y(_3358_),
    .A1(net658),
    .A2(_3171_));
 sg13g2_a21o_1 _8160_ (.A2(_3356_),
    .A1(_3358_),
    .B1(_3182_),
    .X(_3359_));
 sg13g2_o21ai_1 _8161_ (.B1(_3359_),
    .Y(_3360_),
    .A1(_3356_),
    .A2(_3357_));
 sg13g2_mux4_1 _8162_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_25_ ),
    .A1(\i_dm_csrs.progbuf_o_89_ ),
    .A2(\i_dm_csrs.progbuf_o_153_ ),
    .A3(\i_dm_csrs.progbuf_o_217_ ),
    .S1(net651),
    .X(_3361_));
 sg13g2_a22oi_1 _8163_ (.Y(_3362_),
    .B1(net560),
    .B2(_3361_),
    .A2(net551),
    .A1(data_csrs_mem_25_));
 sg13g2_o21ai_1 _8164_ (.B1(_3344_),
    .Y(_3363_),
    .A1(net567),
    .A2(_3362_));
 sg13g2_a21oi_1 _8165_ (.A1(_3354_),
    .A2(_3360_),
    .Y(_3364_),
    .B1(_3363_));
 sg13g2_buf_16 fanout49 (.X(master_add_o_4_),
    .A(net49));
 sg13g2_nor2_1 _8167_ (.A(\i_dm_mem.rdata_q_25_ ),
    .B(net251),
    .Y(_3366_));
 sg13g2_nor3_1 _8168_ (.A(_3349_),
    .B(_3364_),
    .C(_3366_),
    .Y(_0539_));
 sg13g2_buf_2 fanout48 (.A(master_add_o_4_),
    .X(net48));
 sg13g2_mux4_1 _8170_ (.S0(net108),
    .A0(\i_dm_csrs.progbuf_o_26_ ),
    .A1(\i_dm_csrs.progbuf_o_90_ ),
    .A2(\i_dm_csrs.progbuf_o_154_ ),
    .A3(\i_dm_csrs.progbuf_o_218_ ),
    .S1(net646),
    .X(_3368_));
 sg13g2_and4_1 _8171_ (.A(cmd_6_),
    .B(_3136_),
    .C(_3169_),
    .D(_3313_),
    .X(_3369_));
 sg13g2_a221oi_1 _8172_ (.B2(_3368_),
    .C1(_3369_),
    .B1(net499),
    .A1(data_csrs_mem_26_),
    .Y(_3370_),
    .A2(net34));
 sg13g2_a21oi_1 _8173_ (.A1(\i_dm_mem.rdata_q_26_ ),
    .A2(net6),
    .Y(_3371_),
    .B1(_3328_));
 sg13g2_o21ai_1 _8174_ (.B1(_3371_),
    .Y(_0540_),
    .A1(net277),
    .A2(_3370_));
 sg13g2_mux4_1 _8175_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_27_ ),
    .A1(\i_dm_csrs.progbuf_o_91_ ),
    .A2(\i_dm_csrs.progbuf_o_155_ ),
    .A3(\i_dm_csrs.progbuf_o_219_ ),
    .S1(net651),
    .X(_3372_));
 sg13g2_a22oi_1 _8176_ (.Y(_3373_),
    .B1(net562),
    .B2(_3372_),
    .A2(net553),
    .A1(data_csrs_mem_27_));
 sg13g2_nor2_1 _8177_ (.A(net566),
    .B(_3373_),
    .Y(_3374_));
 sg13g2_nor2b_1 _8178_ (.A(cmd_16_),
    .B_N(\i_dm_mem.abstract_cmd_132__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ),
    .Y(_3375_));
 sg13g2_o21ai_1 _8179_ (.B1(_3181_),
    .Y(_3376_),
    .A1(_3170_),
    .A2(_3375_));
 sg13g2_nand2_1 _8180_ (.Y(_3377_),
    .A(cmd_7_),
    .B(_3320_));
 sg13g2_a21oi_1 _8181_ (.A1(_3376_),
    .A2(_3377_),
    .Y(_3378_),
    .B1(_3289_));
 sg13g2_a21oi_1 _8182_ (.A1(net656),
    .A2(_3113_),
    .Y(_3379_),
    .B1(_3137_));
 sg13g2_nor2_1 _8183_ (.A(_1196_),
    .B(_3379_),
    .Y(_3380_));
 sg13g2_a21oi_1 _8184_ (.A1(net656),
    .A2(_3137_),
    .Y(_3381_),
    .B1(_3380_));
 sg13g2_nor2_1 _8185_ (.A(_3167_),
    .B(_3175_),
    .Y(_3382_));
 sg13g2_a21oi_1 _8186_ (.A1(net656),
    .A2(_3137_),
    .Y(_3383_),
    .B1(_3382_));
 sg13g2_nor4_2 _8187_ (.A(net557),
    .B(_3115_),
    .C(_3381_),
    .Y(_3384_),
    .D(_3383_));
 sg13g2_nor3_2 _8188_ (.A(_3374_),
    .B(_3378_),
    .C(_3384_),
    .Y(_3385_));
 sg13g2_nand2_1 _8189_ (.Y(_3386_),
    .A(\i_dm_mem.rdata_q_27_ ),
    .B(net3));
 sg13g2_o21ai_1 _8190_ (.B1(_3386_),
    .Y(_0541_),
    .A1(net275),
    .A2(_3385_));
 sg13g2_nand3_1 _8191_ (.B(_3103_),
    .C(_3329_),
    .A(_0900_),
    .Y(_3387_));
 sg13g2_o21ai_1 _8192_ (.B1(_3387_),
    .Y(_3388_),
    .A1(\i_dm_mem.rdata_q_28_ ),
    .A2(_3101_));
 sg13g2_mux4_1 _8193_ (.S0(net107),
    .A0(\i_dm_csrs.progbuf_o_28_ ),
    .A1(\i_dm_csrs.progbuf_o_92_ ),
    .A2(\i_dm_csrs.progbuf_o_156_ ),
    .A3(\i_dm_csrs.progbuf_o_220_ ),
    .S1(net650),
    .X(_3389_));
 sg13g2_a22oi_1 _8194_ (.Y(_3390_),
    .B1(net562),
    .B2(_3389_),
    .A2(net553),
    .A1(data_csrs_mem_28_));
 sg13g2_nor2_1 _8195_ (.A(net566),
    .B(_3390_),
    .Y(_3391_));
 sg13g2_nor2b_1 _8196_ (.A(net99),
    .B_N(cmd_8_),
    .Y(_3392_));
 sg13g2_inv_1 _8197_ (.Y(_3393_),
    .A(_3376_));
 sg13g2_a21oi_1 _8198_ (.A1(_3141_),
    .A2(_3392_),
    .Y(_3394_),
    .B1(_3393_));
 sg13g2_nor3_1 _8199_ (.A(_3179_),
    .B(_3246_),
    .C(_3394_),
    .Y(_3395_));
 sg13g2_nor3_1 _8200_ (.A(_3247_),
    .B(_3391_),
    .C(_3395_),
    .Y(_3396_));
 sg13g2_o21ai_1 _8201_ (.B1(_3103_),
    .Y(_3397_),
    .A1(net543),
    .A2(net388));
 sg13g2_nor2b_1 _8202_ (.A(\i_dm_mem.rdata_q_28_ ),
    .B_N(_3397_),
    .Y(_3398_));
 sg13g2_a221oi_1 _8203_ (.B2(_3344_),
    .C1(_3398_),
    .B1(_3396_),
    .A1(net543),
    .Y(_0542_),
    .A2(_3388_));
 sg13g2_mux4_1 _8204_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_29_ ),
    .A1(\i_dm_csrs.progbuf_o_93_ ),
    .A2(\i_dm_csrs.progbuf_o_157_ ),
    .A3(\i_dm_csrs.progbuf_o_221_ ),
    .S1(net647),
    .X(_3399_));
 sg13g2_a22oi_1 _8205_ (.Y(_3400_),
    .B1(net559),
    .B2(_3399_),
    .A2(net550),
    .A1(data_csrs_mem_29_));
 sg13g2_nor2_1 _8206_ (.A(net566),
    .B(_3400_),
    .Y(_3401_));
 sg13g2_nand2_1 _8207_ (.Y(_3402_),
    .A(cmd_9_),
    .B(_3320_));
 sg13g2_a21oi_1 _8208_ (.A1(_3376_),
    .A2(_3402_),
    .Y(_3403_),
    .B1(_3289_));
 sg13g2_nor3_2 _8209_ (.A(_3384_),
    .B(_3401_),
    .C(_3403_),
    .Y(_3404_));
 sg13g2_nand2_1 _8210_ (.Y(_3405_),
    .A(\i_dm_mem.rdata_q_29_ ),
    .B(net3));
 sg13g2_o21ai_1 _8211_ (.B1(_3405_),
    .Y(_0543_),
    .A1(net275),
    .A2(_3404_));
 sg13g2_inv_1 _8212_ (.Y(_3406_),
    .A(\i_dm_mem.rdata_q_2_ ));
 sg13g2_and4_1 _8213_ (.A(cmd_5_),
    .B(_3303_),
    .C(_3148_),
    .D(_3207_),
    .X(_3407_));
 sg13g2_mux4_1 _8214_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_2_ ),
    .A1(\i_dm_csrs.progbuf_o_66_ ),
    .A2(\i_dm_csrs.progbuf_o_130_ ),
    .A3(\i_dm_csrs.progbuf_o_194_ ),
    .S1(net648),
    .X(_3408_));
 sg13g2_a22oi_1 _8215_ (.Y(_3409_),
    .B1(net561),
    .B2(_3408_),
    .A2(net552),
    .A1(data_csrs_mem_2_));
 sg13g2_o21ai_1 _8216_ (.B1(_3097_),
    .Y(_3410_),
    .A1(net568),
    .A2(_3409_));
 sg13g2_nor3_1 _8217_ (.A(net3),
    .B(_3407_),
    .C(_3410_),
    .Y(_3411_));
 sg13g2_a21oi_1 _8218_ (.A1(_3406_),
    .A2(net6),
    .Y(_0544_),
    .B1(_3411_));
 sg13g2_inv_1 _8219_ (.Y(_3412_),
    .A(\i_dm_mem.rdata_q_30_ ));
 sg13g2_o21ai_1 _8220_ (.B1(_3387_),
    .Y(_3413_),
    .A1(\i_dm_mem.rdata_q_30_ ),
    .A2(_3101_));
 sg13g2_mux4_1 _8221_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_30_ ),
    .A1(\i_dm_csrs.progbuf_o_94_ ),
    .A2(\i_dm_csrs.progbuf_o_158_ ),
    .A3(\i_dm_csrs.progbuf_o_222_ ),
    .S1(net647),
    .X(_3414_));
 sg13g2_a22oi_1 _8222_ (.Y(_3415_),
    .B1(net559),
    .B2(_3414_),
    .A2(net550),
    .A1(data_csrs_mem_30_));
 sg13g2_o21ai_1 _8223_ (.B1(_3344_),
    .Y(_3416_),
    .A1(net567),
    .A2(_3415_));
 sg13g2_a21oi_1 _8224_ (.A1(net39),
    .A2(cmd_10_),
    .Y(_3417_),
    .B1(_3170_));
 sg13g2_nand2b_1 _8225_ (.Y(_3418_),
    .B(_3312_),
    .A_N(_3417_));
 sg13g2_o21ai_1 _8226_ (.B1(_3182_),
    .Y(_3419_),
    .A1(_3357_),
    .A2(_3418_));
 sg13g2_nand2_1 _8227_ (.Y(_3420_),
    .A(_3358_),
    .B(_3418_));
 sg13g2_nand3_1 _8228_ (.B(_3419_),
    .C(_3420_),
    .A(_3354_),
    .Y(_3421_));
 sg13g2_nor2b_1 _8229_ (.A(_3416_),
    .B_N(_3421_),
    .Y(_3422_));
 sg13g2_a221oi_1 _8230_ (.B2(net543),
    .C1(_3422_),
    .B1(_3413_),
    .A1(_3412_),
    .Y(_0545_),
    .A2(_3397_));
 sg13g2_nand4_1 _8231_ (.B(_3136_),
    .C(_3169_),
    .A(cmd_11_),
    .Y(_3423_),
    .D(_3313_));
 sg13g2_mux4_1 _8232_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_31_ ),
    .A1(\i_dm_csrs.progbuf_o_95_ ),
    .A2(\i_dm_csrs.progbuf_o_159_ ),
    .A3(\i_dm_csrs.progbuf_o_223_ ),
    .S1(net654),
    .X(_3424_));
 sg13g2_a22oi_1 _8233_ (.Y(_3425_),
    .B1(net498),
    .B2(_3424_),
    .A2(net35),
    .A1(data_csrs_mem_31_));
 sg13g2_a21oi_1 _8234_ (.A1(_3423_),
    .A2(_3425_),
    .Y(_3426_),
    .B1(_3329_));
 sg13g2_mux2_1 _8235_ (.A0(\i_dm_mem.rdata_q_31_ ),
    .A1(_3426_),
    .S(net251),
    .X(_0546_));
 sg13g2_mux4_1 _8236_ (.S0(net662),
    .A0(\i_dm_csrs.progbuf_o_32_ ),
    .A1(\i_dm_csrs.progbuf_o_160_ ),
    .A2(\i_dm_csrs.progbuf_o_96_ ),
    .A3(\i_dm_csrs.progbuf_o_224_ ),
    .S1(net113),
    .X(_3427_));
 sg13g2_a221oi_1 _8237_ (.B2(_3427_),
    .C1(net441),
    .B1(net501),
    .A1(data_csrs_mem_32_),
    .Y(_3428_),
    .A2(net34));
 sg13g2_nor2_1 _8238_ (.A(\i_dm_mem.rdata_q_32_ ),
    .B(net250),
    .Y(_3429_));
 sg13g2_a21oi_1 _8239_ (.A1(net250),
    .A2(_3428_),
    .Y(_0547_),
    .B1(_3429_));
 sg13g2_mux4_1 _8240_ (.S0(net108),
    .A0(\i_dm_csrs.progbuf_o_33_ ),
    .A1(\i_dm_csrs.progbuf_o_97_ ),
    .A2(\i_dm_csrs.progbuf_o_161_ ),
    .A3(\i_dm_csrs.progbuf_o_225_ ),
    .S1(net655),
    .X(_3430_));
 sg13g2_a221oi_1 _8241_ (.B2(_3430_),
    .C1(net441),
    .B1(net498),
    .A1(data_csrs_mem_33_),
    .Y(_3431_),
    .A2(net34));
 sg13g2_nor2_1 _8242_ (.A(\i_dm_mem.rdata_q_33_ ),
    .B(net250),
    .Y(_3432_));
 sg13g2_a21oi_1 _8243_ (.A1(net250),
    .A2(_3431_),
    .Y(_0548_),
    .B1(_3432_));
 sg13g2_mux4_1 _8244_ (.S0(net104),
    .A0(\i_dm_csrs.progbuf_o_34_ ),
    .A1(\i_dm_csrs.progbuf_o_98_ ),
    .A2(\i_dm_csrs.progbuf_o_162_ ),
    .A3(\i_dm_csrs.progbuf_o_226_ ),
    .S1(net653),
    .X(_3433_));
 sg13g2_nor2_1 _8245_ (.A(_1193_),
    .B(_3236_),
    .Y(_3434_));
 sg13g2_a221oi_1 _8246_ (.B2(_3433_),
    .C1(_3434_),
    .B1(net498),
    .A1(data_csrs_mem_34_),
    .Y(_3435_),
    .A2(net35));
 sg13g2_nor3_1 _8247_ (.A(_3329_),
    .B(net5),
    .C(_3435_),
    .Y(_3436_));
 sg13g2_a21o_1 _8248_ (.A2(net7),
    .A1(\i_dm_mem.rdata_q_34_ ),
    .B1(_3436_),
    .X(_0549_));
 sg13g2_mux4_1 _8249_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_35_ ),
    .A1(\i_dm_csrs.progbuf_o_99_ ),
    .A2(\i_dm_csrs.progbuf_o_163_ ),
    .A3(\i_dm_csrs.progbuf_o_227_ ),
    .S1(net653),
    .X(_3437_));
 sg13g2_a22oi_1 _8250_ (.Y(_3438_),
    .B1(net499),
    .B2(_3437_),
    .A2(net37),
    .A1(data_csrs_mem_35_));
 sg13g2_nor2_1 _8251_ (.A(\i_dm_mem.rdata_q_35_ ),
    .B(net251),
    .Y(_3439_));
 sg13g2_a21oi_1 _8252_ (.A1(net251),
    .A2(_3438_),
    .Y(_0550_),
    .B1(_3439_));
 sg13g2_mux4_1 _8253_ (.S0(net648),
    .A0(\i_dm_csrs.progbuf_o_36_ ),
    .A1(\i_dm_csrs.progbuf_o_164_ ),
    .A2(\i_dm_csrs.progbuf_o_100_ ),
    .A3(\i_dm_csrs.progbuf_o_228_ ),
    .S1(net113),
    .X(_3440_));
 sg13g2_nand3_1 _8254_ (.B(_0707_),
    .C(_1135_),
    .A(net644),
    .Y(_3441_));
 sg13g2_nor2_1 _8255_ (.A(net565),
    .B(_3441_),
    .Y(_3442_));
 sg13g2_nand3_1 _8256_ (.B(_3169_),
    .C(_3185_),
    .A(net109),
    .Y(_3443_));
 sg13g2_o21ai_1 _8257_ (.B1(_3091_),
    .Y(_3444_),
    .A1(_3137_),
    .A2(_3113_));
 sg13g2_nand2_1 _8258_ (.Y(_3445_),
    .A(data_csrs_mem_36_),
    .B(net38));
 sg13g2_o21ai_1 _8259_ (.B1(_3445_),
    .Y(_3446_),
    .A1(_3115_),
    .A2(_3444_));
 sg13g2_a221oi_1 _8260_ (.B2(_3303_),
    .C1(_3446_),
    .B1(_3443_),
    .A1(_3440_),
    .Y(_3447_),
    .A2(_3442_));
 sg13g2_nand2_1 _8261_ (.Y(_3448_),
    .A(\i_dm_mem.rdata_q_36_ ),
    .B(net3));
 sg13g2_o21ai_1 _8262_ (.B1(_3448_),
    .Y(_0551_),
    .A1(net274),
    .A2(_3447_));
 sg13g2_mux4_1 _8263_ (.S0(net651),
    .A0(\i_dm_csrs.progbuf_o_37_ ),
    .A1(\i_dm_csrs.progbuf_o_165_ ),
    .A2(\i_dm_csrs.progbuf_o_101_ ),
    .A3(\i_dm_csrs.progbuf_o_229_ ),
    .S1(net114),
    .X(_3449_));
 sg13g2_a22oi_1 _8264_ (.Y(_3450_),
    .B1(net562),
    .B2(_3449_),
    .A2(net553),
    .A1(data_csrs_mem_37_));
 sg13g2_nor2_1 _8265_ (.A(_3167_),
    .B(_3357_),
    .Y(_3451_));
 sg13g2_and2_1 _8266_ (.A(cmd_16_),
    .B(net103),
    .X(_3452_));
 sg13g2_nor3_1 _8267_ (.A(_3243_),
    .B(_3234_),
    .C(_3452_),
    .Y(_3453_));
 sg13g2_a21oi_1 _8268_ (.A1(cmd_18_),
    .A2(_1206_),
    .Y(_3454_),
    .B1(_3343_));
 sg13g2_a21oi_1 _8269_ (.A1(net424),
    .A2(_3453_),
    .Y(_3455_),
    .B1(_3454_));
 sg13g2_o21ai_1 _8270_ (.B1(_3455_),
    .Y(_3456_),
    .A1(net569),
    .A2(_3450_));
 sg13g2_a22oi_1 _8271_ (.Y(_3457_),
    .B1(net1),
    .B2(_3456_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_37_ ));
 sg13g2_inv_1 _8272_ (.Y(_0552_),
    .A(_3457_));
 sg13g2_mux4_1 _8273_ (.S0(net648),
    .A0(\i_dm_csrs.progbuf_o_38_ ),
    .A1(\i_dm_csrs.progbuf_o_166_ ),
    .A2(\i_dm_csrs.progbuf_o_102_ ),
    .A3(\i_dm_csrs.progbuf_o_230_ ),
    .S1(net113),
    .X(_3458_));
 sg13g2_a22oi_1 _8274_ (.Y(_3459_),
    .B1(net564),
    .B2(_3458_),
    .A2(net552),
    .A1(data_csrs_mem_38_));
 sg13g2_o21ai_1 _8275_ (.B1(_3455_),
    .Y(_3460_),
    .A1(net569),
    .A2(_3459_));
 sg13g2_a22oi_1 _8276_ (.Y(_3461_),
    .B1(net1),
    .B2(_3460_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_38_ ));
 sg13g2_inv_1 _8277_ (.Y(_0553_),
    .A(_3461_));
 sg13g2_mux4_1 _8278_ (.S0(net653),
    .A0(\i_dm_csrs.progbuf_o_39_ ),
    .A1(\i_dm_csrs.progbuf_o_167_ ),
    .A2(\i_dm_csrs.progbuf_o_103_ ),
    .A3(\i_dm_csrs.progbuf_o_231_ ),
    .S1(net113),
    .X(_3462_));
 sg13g2_a22oi_1 _8279_ (.Y(_3463_),
    .B1(net498),
    .B2(_3462_),
    .A2(net36),
    .A1(data_csrs_mem_39_));
 sg13g2_nor2_1 _8280_ (.A(\i_dm_mem.rdata_q_39_ ),
    .B(net251),
    .Y(_3464_));
 sg13g2_a21oi_1 _8281_ (.A1(net251),
    .A2(_3463_),
    .Y(_0554_),
    .B1(_3464_));
 sg13g2_mux4_1 _8282_ (.S0(net108),
    .A0(\i_dm_csrs.progbuf_o_3_ ),
    .A1(\i_dm_csrs.progbuf_o_67_ ),
    .A2(\i_dm_csrs.progbuf_o_131_ ),
    .A3(\i_dm_csrs.progbuf_o_195_ ),
    .S1(net653),
    .X(_3465_));
 sg13g2_a221oi_1 _8283_ (.B2(_3465_),
    .C1(_3329_),
    .B1(net498),
    .A1(data_csrs_mem_3_),
    .Y(_3466_),
    .A2(net35));
 sg13g2_nor2_1 _8284_ (.A(\i_dm_mem.rdata_q_3_ ),
    .B(net251),
    .Y(_3467_));
 sg13g2_a21oi_1 _8285_ (.A1(net251),
    .A2(_3466_),
    .Y(_0555_),
    .B1(_3467_));
 sg13g2_nand2_1 _8286_ (.Y(_3468_),
    .A(\i_dm_csrs.progbuf_o_168_ ),
    .B(net100));
 sg13g2_nor3_1 _8287_ (.A(net655),
    .B(\i_dm_csrs.progbuf_o_40_ ),
    .C(net565),
    .Y(_3469_));
 sg13g2_a21oi_1 _8288_ (.A1(net655),
    .A2(_3468_),
    .Y(_3470_),
    .B1(_3469_));
 sg13g2_nand2_1 _8289_ (.Y(_3471_),
    .A(net645),
    .B(_3470_));
 sg13g2_nor2b_1 _8290_ (.A(\i_dm_csrs.progbuf_o_232_ ),
    .B_N(net645),
    .Y(_3472_));
 sg13g2_a21oi_1 _8291_ (.A1(\i_dm_csrs.progbuf_o_104_ ),
    .A2(net645),
    .Y(_3473_),
    .B1(net655));
 sg13g2_a21oi_1 _8292_ (.A1(net655),
    .A2(_3472_),
    .Y(_3474_),
    .B1(_3473_));
 sg13g2_nand3_1 _8293_ (.B(net100),
    .C(_3474_),
    .A(net110),
    .Y(_3475_));
 sg13g2_o21ai_1 _8294_ (.B1(_3475_),
    .Y(_3476_),
    .A1(net105),
    .A2(_3471_));
 sg13g2_a22oi_1 _8295_ (.Y(_3477_),
    .B1(_3095_),
    .B2(_3476_),
    .A2(net35),
    .A1(data_csrs_mem_40_));
 sg13g2_nor3_1 _8296_ (.A(_3329_),
    .B(net5),
    .C(_3477_),
    .Y(_3478_));
 sg13g2_a21o_1 _8297_ (.A2(net7),
    .A1(\i_dm_mem.rdata_q_40_ ),
    .B1(_3478_),
    .X(_0556_));
 sg13g2_mux4_1 _8298_ (.S0(net652),
    .A0(\i_dm_csrs.progbuf_o_41_ ),
    .A1(\i_dm_csrs.progbuf_o_169_ ),
    .A2(\i_dm_csrs.progbuf_o_105_ ),
    .A3(\i_dm_csrs.progbuf_o_233_ ),
    .S1(net113),
    .X(_3479_));
 sg13g2_a22oi_1 _8299_ (.Y(_3480_),
    .B1(net500),
    .B2(_3479_),
    .A2(net36),
    .A1(data_csrs_mem_41_));
 sg13g2_nor2_1 _8300_ (.A(\i_dm_mem.rdata_q_41_ ),
    .B(net247),
    .Y(_3481_));
 sg13g2_a21oi_1 _8301_ (.A1(net249),
    .A2(_3480_),
    .Y(_0557_),
    .B1(_3481_));
 sg13g2_o21ai_1 _8302_ (.B1(_3350_),
    .Y(_3482_),
    .A1(_3182_),
    .A2(_3234_));
 sg13g2_buf_2 fanout47 (.A(_0728_),
    .X(net47));
 sg13g2_buf_2 fanout46 (.A(_0728_),
    .X(net46));
 sg13g2_buf_4 fanout45 (.X(net45),
    .A(_0728_));
 sg13g2_mux4_1 _8306_ (.S0(net652),
    .A0(\i_dm_csrs.progbuf_o_42_ ),
    .A1(\i_dm_csrs.progbuf_o_170_ ),
    .A2(\i_dm_csrs.progbuf_o_106_ ),
    .A3(\i_dm_csrs.progbuf_o_234_ ),
    .S1(net115),
    .X(_3486_));
 sg13g2_a22oi_1 _8307_ (.Y(_3487_),
    .B1(net563),
    .B2(_3486_),
    .A2(net554),
    .A1(data_csrs_mem_42_));
 sg13g2_nor2_1 _8308_ (.A(net566),
    .B(_3487_),
    .Y(_3488_));
 sg13g2_a21oi_1 _8309_ (.A1(_3189_),
    .A2(_3482_),
    .Y(_3489_),
    .B1(_3488_));
 sg13g2_nand2_1 _8310_ (.Y(_3490_),
    .A(\i_dm_mem.rdata_q_42_ ),
    .B(net3));
 sg13g2_o21ai_1 _8311_ (.B1(_3490_),
    .Y(_0558_),
    .A1(net275),
    .A2(_3489_));
 sg13g2_mux4_1 _8312_ (.S0(net651),
    .A0(\i_dm_csrs.progbuf_o_43_ ),
    .A1(\i_dm_csrs.progbuf_o_171_ ),
    .A2(\i_dm_csrs.progbuf_o_107_ ),
    .A3(\i_dm_csrs.progbuf_o_235_ ),
    .S1(net112),
    .X(_3491_));
 sg13g2_a22oi_1 _8313_ (.Y(_3492_),
    .B1(net500),
    .B2(_3491_),
    .A2(net36),
    .A1(data_csrs_mem_43_));
 sg13g2_nor2_1 _8314_ (.A(\i_dm_mem.rdata_q_43_ ),
    .B(net249),
    .Y(_3493_));
 sg13g2_a21oi_1 _8315_ (.A1(_3225_),
    .A2(_3492_),
    .Y(_0559_),
    .B1(_3493_));
 sg13g2_mux4_1 _8316_ (.S0(net647),
    .A0(\i_dm_csrs.progbuf_o_44_ ),
    .A1(\i_dm_csrs.progbuf_o_172_ ),
    .A2(\i_dm_csrs.progbuf_o_108_ ),
    .A3(\i_dm_csrs.progbuf_o_236_ ),
    .S1(net113),
    .X(_3494_));
 sg13g2_a22oi_1 _8317_ (.Y(_3495_),
    .B1(net559),
    .B2(_3494_),
    .A2(net550),
    .A1(data_csrs_mem_44_));
 sg13g2_nand3_1 _8318_ (.B(_3169_),
    .C(_3185_),
    .A(cmd_20_),
    .Y(_3496_));
 sg13g2_a21o_1 _8319_ (.A2(_3496_),
    .A1(net109),
    .B1(_3304_),
    .X(_3497_));
 sg13g2_o21ai_1 _8320_ (.B1(_3497_),
    .Y(_3498_),
    .A1(net567),
    .A2(_3495_));
 sg13g2_a22oi_1 _8321_ (.Y(_3499_),
    .B1(net1),
    .B2(_3498_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_44_ ));
 sg13g2_inv_1 _8322_ (.Y(_0560_),
    .A(_3499_));
 sg13g2_mux4_1 _8323_ (.S0(net646),
    .A0(\i_dm_csrs.progbuf_o_45_ ),
    .A1(\i_dm_csrs.progbuf_o_173_ ),
    .A2(\i_dm_csrs.progbuf_o_109_ ),
    .A3(\i_dm_csrs.progbuf_o_237_ ),
    .S1(net113),
    .X(_3500_));
 sg13g2_a22oi_1 _8324_ (.Y(_3501_),
    .B1(net561),
    .B2(_3500_),
    .A2(net552),
    .A1(data_csrs_mem_45_));
 sg13g2_and4_1 _8325_ (.A(cmd_21_),
    .B(net109),
    .C(_3141_),
    .D(_3185_),
    .X(_3502_));
 sg13g2_o21ai_1 _8326_ (.B1(net424),
    .Y(_3503_),
    .A1(_3453_),
    .A2(_3502_));
 sg13g2_o21ai_1 _8327_ (.B1(_3503_),
    .Y(_3504_),
    .A1(net568),
    .A2(_3501_));
 sg13g2_a22oi_1 _8328_ (.Y(_3505_),
    .B1(net1),
    .B2(_3504_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_45_ ));
 sg13g2_inv_1 _8329_ (.Y(_0561_),
    .A(_3505_));
 sg13g2_mux4_1 _8330_ (.S0(net653),
    .A0(\i_dm_csrs.progbuf_o_46_ ),
    .A1(\i_dm_csrs.progbuf_o_174_ ),
    .A2(\i_dm_csrs.progbuf_o_110_ ),
    .A3(\i_dm_csrs.progbuf_o_238_ ),
    .S1(net112),
    .X(_3506_));
 sg13g2_a22oi_1 _8331_ (.Y(_3507_),
    .B1(net501),
    .B2(_3506_),
    .A2(net36),
    .A1(data_csrs_mem_46_));
 sg13g2_nor2_1 _8332_ (.A(\i_dm_mem.rdata_q_46_ ),
    .B(net250),
    .Y(_3508_));
 sg13g2_a21oi_1 _8333_ (.A1(net250),
    .A2(_3507_),
    .Y(_0562_),
    .B1(_3508_));
 sg13g2_mux4_1 _8334_ (.S0(net648),
    .A0(\i_dm_csrs.progbuf_o_47_ ),
    .A1(\i_dm_csrs.progbuf_o_175_ ),
    .A2(\i_dm_csrs.progbuf_o_111_ ),
    .A3(\i_dm_csrs.progbuf_o_239_ ),
    .S1(net112),
    .X(_3509_));
 sg13g2_a22oi_1 _8335_ (.Y(_3510_),
    .B1(net500),
    .B2(_3509_),
    .A2(net36),
    .A1(data_csrs_mem_47_));
 sg13g2_nor2_1 _8336_ (.A(\i_dm_mem.rdata_q_47_ ),
    .B(net247),
    .Y(_3511_));
 sg13g2_a21oi_1 _8337_ (.A1(net247),
    .A2(_3510_),
    .Y(_0563_),
    .B1(_3511_));
 sg13g2_mux4_1 _8338_ (.S0(net650),
    .A0(\i_dm_csrs.progbuf_o_48_ ),
    .A1(\i_dm_csrs.progbuf_o_176_ ),
    .A2(\i_dm_csrs.progbuf_o_112_ ),
    .A3(\i_dm_csrs.progbuf_o_240_ ),
    .S1(net113),
    .X(_3512_));
 sg13g2_a22oi_1 _8339_ (.Y(_3513_),
    .B1(net562),
    .B2(_3512_),
    .A2(net553),
    .A1(data_csrs_mem_48_));
 sg13g2_o21ai_1 _8340_ (.B1(net110),
    .Y(_3514_),
    .A1(_3142_),
    .A2(_3234_));
 sg13g2_nand2b_1 _8341_ (.Y(_3515_),
    .B(_3514_),
    .A_N(_3304_));
 sg13g2_o21ai_1 _8342_ (.B1(_3515_),
    .Y(_3516_),
    .A1(net566),
    .A2(_3513_));
 sg13g2_a22oi_1 _8343_ (.Y(_3517_),
    .B1(net1),
    .B2(_3516_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_48_ ));
 sg13g2_inv_1 _8344_ (.Y(_0564_),
    .A(_3517_));
 sg13g2_mux4_1 _8345_ (.S0(net650),
    .A0(\i_dm_csrs.progbuf_o_49_ ),
    .A1(\i_dm_csrs.progbuf_o_177_ ),
    .A2(\i_dm_csrs.progbuf_o_113_ ),
    .A3(\i_dm_csrs.progbuf_o_241_ ),
    .S1(net112),
    .X(_3518_));
 sg13g2_a22oi_1 _8346_ (.Y(_3519_),
    .B1(net500),
    .B2(_3518_),
    .A2(net36),
    .A1(data_csrs_mem_49_));
 sg13g2_nor2_1 _8347_ (.A(\i_dm_mem.rdata_q_49_ ),
    .B(net248),
    .Y(_3520_));
 sg13g2_a21oi_1 _8348_ (.A1(net248),
    .A2(_3519_),
    .Y(_0565_),
    .B1(_3520_));
 sg13g2_nor2_1 _8349_ (.A(_3160_),
    .B(_3171_),
    .Y(_3521_));
 sg13g2_a221oi_1 _8350_ (.B2(_3255_),
    .C1(_3117_),
    .B1(_3521_),
    .A1(_3136_),
    .Y(_3522_),
    .A2(_3178_));
 sg13g2_mux4_1 _8351_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_4_ ),
    .A1(\i_dm_csrs.progbuf_o_68_ ),
    .A2(\i_dm_csrs.progbuf_o_132_ ),
    .A3(\i_dm_csrs.progbuf_o_196_ ),
    .S1(net648),
    .X(_3523_));
 sg13g2_a22oi_1 _8352_ (.Y(_3524_),
    .B1(net564),
    .B2(_3523_),
    .A2(net555),
    .A1(data_csrs_mem_4_));
 sg13g2_nor2_1 _8353_ (.A(_3155_),
    .B(_3524_),
    .Y(_3525_));
 sg13g2_a221oi_1 _8354_ (.B2(_3522_),
    .C1(_3525_),
    .B1(net2),
    .A1(\i_dm_mem.rdata_q_4_ ),
    .Y(_3526_),
    .A2(net6));
 sg13g2_inv_1 _8355_ (.Y(_0566_),
    .A(_3526_));
 sg13g2_mux4_1 _8356_ (.S0(net650),
    .A0(\i_dm_csrs.progbuf_o_50_ ),
    .A1(\i_dm_csrs.progbuf_o_178_ ),
    .A2(\i_dm_csrs.progbuf_o_114_ ),
    .A3(\i_dm_csrs.progbuf_o_242_ ),
    .S1(net115),
    .X(_3527_));
 sg13g2_a22oi_1 _8357_ (.Y(_3528_),
    .B1(net563),
    .B2(_3527_),
    .A2(net554),
    .A1(data_csrs_mem_50_));
 sg13g2_o21ai_1 _8358_ (.B1(_3515_),
    .Y(_3529_),
    .A1(net566),
    .A2(_3528_));
 sg13g2_a22oi_1 _8359_ (.Y(_3530_),
    .B1(net1),
    .B2(_3529_),
    .A2(net8),
    .A1(\i_dm_mem.rdata_q_50_ ));
 sg13g2_inv_1 _8360_ (.Y(_0567_),
    .A(_3530_));
 sg13g2_mux4_1 _8361_ (.S0(net652),
    .A0(\i_dm_csrs.progbuf_o_51_ ),
    .A1(\i_dm_csrs.progbuf_o_179_ ),
    .A2(\i_dm_csrs.progbuf_o_115_ ),
    .A3(\i_dm_csrs.progbuf_o_243_ ),
    .S1(net112),
    .X(_3531_));
 sg13g2_a22oi_1 _8362_ (.Y(_3532_),
    .B1(net500),
    .B2(_3531_),
    .A2(net34),
    .A1(data_csrs_mem_51_));
 sg13g2_nor2_1 _8363_ (.A(\i_dm_mem.rdata_q_51_ ),
    .B(net248),
    .Y(_3533_));
 sg13g2_a21oi_1 _8364_ (.A1(net247),
    .A2(_3532_),
    .Y(_0568_),
    .B1(_3533_));
 sg13g2_mux4_1 _8365_ (.S0(net646),
    .A0(\i_dm_csrs.progbuf_o_52_ ),
    .A1(\i_dm_csrs.progbuf_o_180_ ),
    .A2(\i_dm_csrs.progbuf_o_116_ ),
    .A3(\i_dm_csrs.progbuf_o_244_ ),
    .S1(net112),
    .X(_3534_));
 sg13g2_a22oi_1 _8366_ (.Y(_3535_),
    .B1(net560),
    .B2(_3534_),
    .A2(net551),
    .A1(data_csrs_mem_52_));
 sg13g2_inv_1 _8367_ (.Y(_3536_),
    .A(_3535_));
 sg13g2_nor3_1 _8368_ (.A(_3138_),
    .B(_3160_),
    .C(_3177_),
    .Y(_3537_));
 sg13g2_a221oi_1 _8369_ (.B2(_3274_),
    .C1(_3454_),
    .B1(_3537_),
    .A1(_0707_),
    .Y(_3538_),
    .A2(_3536_));
 sg13g2_nand2_1 _8370_ (.Y(_3539_),
    .A(\i_dm_mem.rdata_q_52_ ),
    .B(net3));
 sg13g2_o21ai_1 _8371_ (.B1(_3539_),
    .Y(_0569_),
    .A1(net275),
    .A2(_3538_));
 sg13g2_buf_8 fanout44 (.A(_0612_),
    .X(net44));
 sg13g2_nand2_2 _8373_ (.Y(_3541_),
    .A(net110),
    .B(_3176_));
 sg13g2_nand3_1 _8374_ (.B(_3181_),
    .C(_3171_),
    .A(net557),
    .Y(_3542_));
 sg13g2_o21ai_1 _8375_ (.B1(_3542_),
    .Y(_3543_),
    .A1(_3290_),
    .A2(_3541_));
 sg13g2_mux4_1 _8376_ (.S0(net646),
    .A0(\i_dm_csrs.progbuf_o_53_ ),
    .A1(\i_dm_csrs.progbuf_o_181_ ),
    .A2(\i_dm_csrs.progbuf_o_117_ ),
    .A3(\i_dm_csrs.progbuf_o_245_ ),
    .S1(net114),
    .X(_3544_));
 sg13g2_a22oi_1 _8377_ (.Y(_3545_),
    .B1(net559),
    .B2(_3544_),
    .A2(net550),
    .A1(data_csrs_mem_53_));
 sg13g2_nor2_1 _8378_ (.A(net569),
    .B(_3545_),
    .Y(_3546_));
 sg13g2_a21oi_1 _8379_ (.A1(net424),
    .A2(_3543_),
    .Y(_3547_),
    .B1(_3546_));
 sg13g2_buf_1 fanout43 (.A(_1249_),
    .X(net43));
 sg13g2_nand2_1 _8381_ (.Y(_3549_),
    .A(\i_dm_mem.rdata_q_53_ ),
    .B(net5));
 sg13g2_o21ai_1 _8382_ (.B1(_3549_),
    .Y(_0570_),
    .A1(net274),
    .A2(_3547_));
 sg13g2_nor3_1 _8383_ (.A(net99),
    .B(_3177_),
    .C(_3304_),
    .Y(_3550_));
 sg13g2_nor2_1 _8384_ (.A(\i_dm_csrs.progbuf_o_54_ ),
    .B(net565),
    .Y(_3551_));
 sg13g2_nand3_1 _8385_ (.B(\i_dm_csrs.progbuf_o_182_ ),
    .C(net100),
    .A(net657),
    .Y(_3552_));
 sg13g2_o21ai_1 _8386_ (.B1(_3552_),
    .Y(_3553_),
    .A1(net657),
    .A2(_3551_));
 sg13g2_mux2_1 _8387_ (.A0(\i_dm_csrs.progbuf_o_118_ ),
    .A1(\i_dm_csrs.progbuf_o_246_ ),
    .S(net657),
    .X(_3554_));
 sg13g2_a22oi_1 _8388_ (.Y(_3555_),
    .B1(_3554_),
    .B2(_3351_),
    .A2(_3553_),
    .A1(net558));
 sg13g2_nor2_1 _8389_ (.A(_3441_),
    .B(_3555_),
    .Y(_3556_));
 sg13g2_a221oi_1 _8390_ (.B2(cmd_2_),
    .C1(_3556_),
    .B1(_3550_),
    .A1(data_csrs_mem_54_),
    .Y(_3557_),
    .A2(net34));
 sg13g2_nand2_1 _8391_ (.Y(_3558_),
    .A(\i_dm_mem.rdata_q_54_ ),
    .B(net5));
 sg13g2_o21ai_1 _8392_ (.B1(_3558_),
    .Y(_0571_),
    .A1(net273),
    .A2(_3557_));
 sg13g2_nor2_1 _8393_ (.A(\i_dm_csrs.progbuf_o_55_ ),
    .B(net565),
    .Y(_3559_));
 sg13g2_nand3_1 _8394_ (.B(\i_dm_csrs.progbuf_o_183_ ),
    .C(net100),
    .A(net655),
    .Y(_3560_));
 sg13g2_o21ai_1 _8395_ (.B1(_3560_),
    .Y(_3561_),
    .A1(net655),
    .A2(_3559_));
 sg13g2_mux2_1 _8396_ (.A0(\i_dm_csrs.progbuf_o_119_ ),
    .A1(\i_dm_csrs.progbuf_o_247_ ),
    .S(net655),
    .X(_3562_));
 sg13g2_a22oi_1 _8397_ (.Y(_3563_),
    .B1(_3562_),
    .B2(_3351_),
    .A2(_3561_),
    .A1(net558));
 sg13g2_nor2_1 _8398_ (.A(_3441_),
    .B(_3563_),
    .Y(_3564_));
 sg13g2_a221oi_1 _8399_ (.B2(cmd_3_),
    .C1(_3564_),
    .B1(_3550_),
    .A1(data_csrs_mem_55_),
    .Y(_3565_),
    .A2(net34));
 sg13g2_nand2_1 _8400_ (.Y(_3566_),
    .A(\i_dm_mem.rdata_q_55_ ),
    .B(net5));
 sg13g2_o21ai_1 _8401_ (.B1(_3566_),
    .Y(_0572_),
    .A1(net273),
    .A2(_3565_));
 sg13g2_a21oi_1 _8402_ (.A1(net39),
    .A2(cmd_4_),
    .Y(_3567_),
    .B1(net497));
 sg13g2_o21ai_1 _8403_ (.B1(_3542_),
    .Y(_3568_),
    .A1(_3541_),
    .A2(_3567_));
 sg13g2_mux4_1 _8404_ (.S0(net647),
    .A0(\i_dm_csrs.progbuf_o_56_ ),
    .A1(\i_dm_csrs.progbuf_o_184_ ),
    .A2(\i_dm_csrs.progbuf_o_120_ ),
    .A3(\i_dm_csrs.progbuf_o_248_ ),
    .S1(net114),
    .X(_3569_));
 sg13g2_a22oi_1 _8405_ (.Y(_3570_),
    .B1(net560),
    .B2(_3569_),
    .A2(net551),
    .A1(data_csrs_mem_56_));
 sg13g2_nor2_1 _8406_ (.A(_3087_),
    .B(_3570_),
    .Y(_3571_));
 sg13g2_a21oi_1 _8407_ (.A1(net424),
    .A2(_3568_),
    .Y(_3572_),
    .B1(_3571_));
 sg13g2_nand2_1 _8408_ (.Y(_3573_),
    .A(\i_dm_mem.rdata_q_56_ ),
    .B(net5));
 sg13g2_o21ai_1 _8409_ (.B1(_3573_),
    .Y(_0573_),
    .A1(net274),
    .A2(_3572_));
 sg13g2_o21ai_1 _8410_ (.B1(_3542_),
    .Y(_3574_),
    .A1(_3355_),
    .A2(_3541_));
 sg13g2_mux4_1 _8411_ (.S0(net651),
    .A0(\i_dm_csrs.progbuf_o_57_ ),
    .A1(\i_dm_csrs.progbuf_o_185_ ),
    .A2(\i_dm_csrs.progbuf_o_121_ ),
    .A3(\i_dm_csrs.progbuf_o_249_ ),
    .S1(net114),
    .X(_3575_));
 sg13g2_a22oi_1 _8412_ (.Y(_3576_),
    .B1(net560),
    .B2(_3575_),
    .A2(net551),
    .A1(data_csrs_mem_57_));
 sg13g2_nor2_1 _8413_ (.A(net568),
    .B(_3576_),
    .Y(_3577_));
 sg13g2_a21oi_1 _8414_ (.A1(net424),
    .A2(_3574_),
    .Y(_3578_),
    .B1(_3577_));
 sg13g2_nand2_1 _8415_ (.Y(_3579_),
    .A(\i_dm_mem.rdata_q_57_ ),
    .B(net5));
 sg13g2_o21ai_1 _8416_ (.B1(_3579_),
    .Y(_0574_),
    .A1(net273),
    .A2(_3578_));
 sg13g2_and2_1 _8417_ (.A(net39),
    .B(_3537_),
    .X(_3580_));
 sg13g2_mux4_1 _8418_ (.S0(net646),
    .A0(\i_dm_csrs.progbuf_o_58_ ),
    .A1(\i_dm_csrs.progbuf_o_186_ ),
    .A2(\i_dm_csrs.progbuf_o_122_ ),
    .A3(\i_dm_csrs.progbuf_o_250_ ),
    .S1(net114),
    .X(_3581_));
 sg13g2_a22oi_1 _8419_ (.Y(_3582_),
    .B1(net559),
    .B2(_3581_),
    .A2(net550),
    .A1(data_csrs_mem_58_));
 sg13g2_nor2_1 _8420_ (.A(net568),
    .B(_3582_),
    .Y(_3583_));
 sg13g2_a21oi_1 _8421_ (.A1(cmd_6_),
    .A2(_3580_),
    .Y(_3584_),
    .B1(_3583_));
 sg13g2_nand2_1 _8422_ (.Y(_3585_),
    .A(\i_dm_mem.rdata_q_58_ ),
    .B(net5));
 sg13g2_o21ai_1 _8423_ (.B1(_3585_),
    .Y(_0575_),
    .A1(net273),
    .A2(_3584_));
 sg13g2_a21oi_1 _8424_ (.A1(net39),
    .A2(cmd_7_),
    .Y(_3586_),
    .B1(net497));
 sg13g2_a21oi_1 _8425_ (.A1(\cmd_16__$_NOT__A_Y ),
    .A2(net557),
    .Y(_3587_),
    .B1(cmd_16_));
 sg13g2_or3_1 _8426_ (.A(_3175_),
    .B(_3234_),
    .C(_3587_),
    .X(_3588_));
 sg13g2_o21ai_1 _8427_ (.B1(_3588_),
    .Y(_3589_),
    .A1(_3541_),
    .A2(_3586_));
 sg13g2_mux4_1 _8428_ (.S0(net651),
    .A0(\i_dm_csrs.progbuf_o_59_ ),
    .A1(\i_dm_csrs.progbuf_o_187_ ),
    .A2(\i_dm_csrs.progbuf_o_123_ ),
    .A3(\i_dm_csrs.progbuf_o_251_ ),
    .S1(net114),
    .X(_3590_));
 sg13g2_a22oi_1 _8429_ (.Y(_3591_),
    .B1(net563),
    .B2(_3590_),
    .A2(net554),
    .A1(data_csrs_mem_59_));
 sg13g2_nor2_1 _8430_ (.A(net569),
    .B(_3591_),
    .Y(_3592_));
 sg13g2_a21oi_1 _8431_ (.A1(net424),
    .A2(_3589_),
    .Y(_3593_),
    .B1(_3592_));
 sg13g2_nand2_1 _8432_ (.Y(_3594_),
    .A(\i_dm_mem.rdata_q_59_ ),
    .B(net4));
 sg13g2_o21ai_1 _8433_ (.B1(_3594_),
    .Y(_0576_),
    .A1(net275),
    .A2(_3593_));
 sg13g2_inv_1 _8434_ (.Y(_3595_),
    .A(\i_dm_mem.rdata_q_5_ ));
 sg13g2_a22oi_1 _8435_ (.Y(_3596_),
    .B1(_3171_),
    .B2(_3350_),
    .A2(_3140_),
    .A1(_3148_));
 sg13g2_o21ai_1 _8436_ (.B1(_3272_),
    .Y(_3597_),
    .A1(_3182_),
    .A2(_3596_));
 sg13g2_nand2_1 _8437_ (.Y(_3598_),
    .A(net441),
    .B(_3597_));
 sg13g2_mux4_1 _8438_ (.S0(net105),
    .A0(\i_dm_csrs.progbuf_o_5_ ),
    .A1(\i_dm_csrs.progbuf_o_69_ ),
    .A2(\i_dm_csrs.progbuf_o_133_ ),
    .A3(\i_dm_csrs.progbuf_o_197_ ),
    .S1(net651),
    .X(_3599_));
 sg13g2_a221oi_1 _8439_ (.B2(_3599_),
    .C1(net278),
    .B1(net500),
    .A1(data_csrs_mem_5_),
    .Y(_3600_),
    .A2(net34));
 sg13g2_a22oi_1 _8440_ (.Y(_0577_),
    .B1(_3598_),
    .B2(_3600_),
    .A2(net7),
    .A1(_3595_));
 sg13g2_nor2_1 _8441_ (.A(net497),
    .B(_3392_),
    .Y(_3601_));
 sg13g2_o21ai_1 _8442_ (.B1(_3588_),
    .Y(_3602_),
    .A1(_3541_),
    .A2(_3601_));
 sg13g2_mux4_1 _8443_ (.S0(net650),
    .A0(\i_dm_csrs.progbuf_o_60_ ),
    .A1(\i_dm_csrs.progbuf_o_188_ ),
    .A2(\i_dm_csrs.progbuf_o_124_ ),
    .A3(\i_dm_csrs.progbuf_o_252_ ),
    .S1(net114),
    .X(_3603_));
 sg13g2_a22oi_1 _8444_ (.Y(_3604_),
    .B1(net562),
    .B2(_3603_),
    .A2(net553),
    .A1(data_csrs_mem_60_));
 sg13g2_nor2_1 _8445_ (.A(net569),
    .B(_3604_),
    .Y(_3605_));
 sg13g2_a21oi_1 _8446_ (.A1(net424),
    .A2(_3602_),
    .Y(_3606_),
    .B1(_3605_));
 sg13g2_nand2_1 _8447_ (.Y(_3607_),
    .A(\i_dm_mem.rdata_q_60_ ),
    .B(net4));
 sg13g2_o21ai_1 _8448_ (.B1(_3607_),
    .Y(_0578_),
    .A1(net276),
    .A2(_3606_));
 sg13g2_a21oi_1 _8449_ (.A1(net39),
    .A2(cmd_9_),
    .Y(_3608_),
    .B1(net497));
 sg13g2_o21ai_1 _8450_ (.B1(_3588_),
    .Y(_3609_),
    .A1(_3541_),
    .A2(_3608_));
 sg13g2_mux4_1 _8451_ (.S0(net647),
    .A0(\i_dm_csrs.progbuf_o_61_ ),
    .A1(\i_dm_csrs.progbuf_o_189_ ),
    .A2(\i_dm_csrs.progbuf_o_125_ ),
    .A3(\i_dm_csrs.progbuf_o_253_ ),
    .S1(net114),
    .X(_3610_));
 sg13g2_a22oi_1 _8452_ (.Y(_3611_),
    .B1(net559),
    .B2(_3610_),
    .A2(net550),
    .A1(data_csrs_mem_61_));
 sg13g2_nor2_1 _8453_ (.A(net569),
    .B(_3611_),
    .Y(_3612_));
 sg13g2_a21oi_1 _8454_ (.A1(_3451_),
    .A2(_3609_),
    .Y(_3613_),
    .B1(_3612_));
 sg13g2_nand2_1 _8455_ (.Y(_3614_),
    .A(\i_dm_mem.rdata_q_61_ ),
    .B(net4));
 sg13g2_o21ai_1 _8456_ (.B1(_3614_),
    .Y(_0579_),
    .A1(net276),
    .A2(_3613_));
 sg13g2_o21ai_1 _8457_ (.B1(_3542_),
    .Y(_3615_),
    .A1(_3417_),
    .A2(_3541_));
 sg13g2_mux4_1 _8458_ (.S0(net649),
    .A0(\i_dm_csrs.progbuf_o_62_ ),
    .A1(\i_dm_csrs.progbuf_o_190_ ),
    .A2(\i_dm_csrs.progbuf_o_126_ ),
    .A3(\i_dm_csrs.progbuf_o_254_ ),
    .S1(net112),
    .X(_3616_));
 sg13g2_a22oi_1 _8459_ (.Y(_3617_),
    .B1(net559),
    .B2(_3616_),
    .A2(net550),
    .A1(data_csrs_mem_62_));
 sg13g2_nor2_1 _8460_ (.A(net568),
    .B(_3617_),
    .Y(_3618_));
 sg13g2_a21oi_1 _8461_ (.A1(net424),
    .A2(_3615_),
    .Y(_3619_),
    .B1(_3618_));
 sg13g2_nand2_1 _8462_ (.Y(_3620_),
    .A(\i_dm_mem.rdata_q_62_ ),
    .B(net4));
 sg13g2_o21ai_1 _8463_ (.B1(_3620_),
    .Y(_0580_),
    .A1(net273),
    .A2(_3619_));
 sg13g2_mux4_1 _8464_ (.S0(net654),
    .A0(\i_dm_csrs.progbuf_o_63_ ),
    .A1(\i_dm_csrs.progbuf_o_191_ ),
    .A2(\i_dm_csrs.progbuf_o_127_ ),
    .A3(\i_dm_csrs.progbuf_o_255_ ),
    .S1(net112),
    .X(_3621_));
 sg13g2_a22oi_1 _8465_ (.Y(_3622_),
    .B1(net564),
    .B2(_3621_),
    .A2(net555),
    .A1(data_csrs_mem_63_));
 sg13g2_nor2_1 _8466_ (.A(net568),
    .B(_3622_),
    .Y(_3623_));
 sg13g2_a21oi_1 _8467_ (.A1(cmd_11_),
    .A2(_3580_),
    .Y(_3624_),
    .B1(_3623_));
 sg13g2_nand2_1 _8468_ (.Y(_3625_),
    .A(\i_dm_mem.rdata_q_63_ ),
    .B(net3));
 sg13g2_o21ai_1 _8469_ (.B1(_3625_),
    .Y(_0581_),
    .A1(net274),
    .A2(_3624_));
 sg13g2_inv_1 _8470_ (.Y(_3626_),
    .A(\i_dm_mem.rdata_q_6_ ));
 sg13g2_nor3_1 _8471_ (.A(net557),
    .B(net659),
    .C(_1196_),
    .Y(_3627_));
 sg13g2_and3_1 _8472_ (.X(_3628_),
    .A(cmd_16_),
    .B(net557),
    .C(net659));
 sg13g2_o21ai_1 _8473_ (.B1(_3382_),
    .Y(_3629_),
    .A1(_3627_),
    .A2(_3628_));
 sg13g2_o21ai_1 _8474_ (.B1(_3272_),
    .Y(_3630_),
    .A1(_3234_),
    .A2(_3629_));
 sg13g2_nand2_1 _8475_ (.Y(_3631_),
    .A(_3116_),
    .B(_3630_));
 sg13g2_mux4_1 _8476_ (.S0(net108),
    .A0(\i_dm_csrs.progbuf_o_6_ ),
    .A1(\i_dm_csrs.progbuf_o_70_ ),
    .A2(\i_dm_csrs.progbuf_o_134_ ),
    .A3(\i_dm_csrs.progbuf_o_198_ ),
    .S1(net648),
    .X(_3632_));
 sg13g2_a221oi_1 _8477_ (.B2(_3632_),
    .C1(net278),
    .B1(net498),
    .A1(data_csrs_mem_6_),
    .Y(_3633_),
    .A2(net34));
 sg13g2_a22oi_1 _8478_ (.Y(_0582_),
    .B1(_3631_),
    .B2(_3633_),
    .A2(net7),
    .A1(_3626_));
 sg13g2_nand2_1 _8479_ (.Y(_3634_),
    .A(cmd_0_),
    .B(_3161_));
 sg13g2_mux4_1 _8480_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_7_ ),
    .A1(\i_dm_csrs.progbuf_o_71_ ),
    .A2(\i_dm_csrs.progbuf_o_135_ ),
    .A3(\i_dm_csrs.progbuf_o_199_ ),
    .S1(net648),
    .X(_3635_));
 sg13g2_a22oi_1 _8481_ (.Y(_3636_),
    .B1(net498),
    .B2(_3635_),
    .A2(net35),
    .A1(data_csrs_mem_7_));
 sg13g2_a21oi_1 _8482_ (.A1(_3634_),
    .A2(_3636_),
    .Y(_3637_),
    .B1(net277));
 sg13g2_a21o_1 _8483_ (.A2(net6),
    .A1(\i_dm_mem.rdata_q_7_ ),
    .B1(_3637_),
    .X(_0583_));
 sg13g2_nand2_1 _8484_ (.Y(_3638_),
    .A(cmd_1_),
    .B(_3145_));
 sg13g2_o21ai_1 _8485_ (.B1(_3148_),
    .Y(_3639_),
    .A1(_3142_),
    .A2(_3638_));
 sg13g2_mux4_1 _8486_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_8_ ),
    .A1(\i_dm_csrs.progbuf_o_72_ ),
    .A2(\i_dm_csrs.progbuf_o_136_ ),
    .A3(\i_dm_csrs.progbuf_o_200_ ),
    .S1(net653),
    .X(_3640_));
 sg13g2_a22oi_1 _8487_ (.Y(_3641_),
    .B1(net564),
    .B2(_3640_),
    .A2(net555),
    .A1(data_csrs_mem_8_));
 sg13g2_nor2_1 _8488_ (.A(_3155_),
    .B(_3641_),
    .Y(_3642_));
 sg13g2_a221oi_1 _8489_ (.B2(_3639_),
    .C1(_3642_),
    .B1(_3139_),
    .A1(\i_dm_mem.rdata_q_8_ ),
    .Y(_3643_),
    .A2(net6));
 sg13g2_inv_1 _8490_ (.Y(_0584_),
    .A(_3643_));
 sg13g2_nand2_1 _8491_ (.Y(_3644_),
    .A(cmd_2_),
    .B(_3161_));
 sg13g2_mux4_1 _8492_ (.S0(net106),
    .A0(\i_dm_csrs.progbuf_o_9_ ),
    .A1(\i_dm_csrs.progbuf_o_73_ ),
    .A2(\i_dm_csrs.progbuf_o_137_ ),
    .A3(\i_dm_csrs.progbuf_o_201_ ),
    .S1(net652),
    .X(_3645_));
 sg13g2_a22oi_1 _8493_ (.Y(_3646_),
    .B1(net500),
    .B2(_3645_),
    .A2(net35),
    .A1(data_csrs_mem_9_));
 sg13g2_a21oi_1 _8494_ (.A1(_3644_),
    .A2(_3646_),
    .Y(_3647_),
    .B1(net275));
 sg13g2_a21o_1 _8495_ (.A2(net8),
    .A1(\i_dm_mem.rdata_q_9_ ),
    .B1(_3647_),
    .X(_0585_));
 sg13g2_nor2_1 _8496_ (.A(slave_wdata_i_0_),
    .B(_1137_),
    .Y(_3648_));
 sg13g2_nand2_2 _8497_ (.Y(_3649_),
    .A(\clear_resumeack_$_AND__Y_A ),
    .B(_1244_));
 sg13g2_a22oi_1 _8498_ (.Y(_3650_),
    .B1(_3649_),
    .B2(\i_dm_csrs.dmstatus_16_ ),
    .A2(_3136_),
    .A1(_3648_));
 sg13g2_nor2_1 _8499_ (.A(ndmreset_o),
    .B(_3650_),
    .Y(\i_dm_mem.resuming_d ));
 sg13g2_nor2_1 _8500_ (.A(\i_dm_csrs.dmstatus_16_ ),
    .B(\i_dm_mem.state_q_0_ ),
    .Y(_3651_));
 sg13g2_or4_1 _8501_ (.A(slave_wdata_i_0_),
    .B(net110),
    .C(net656),
    .D(_3651_),
    .X(_3652_));
 sg13g2_o21ai_1 _8502_ (.B1(\i_dm_mem.state_q_0__$_NOT__A_Y ),
    .Y(_3653_),
    .A1(\i_dm_csrs.dmstatus_16_ ),
    .A2(\i_dm_mem.state_q_0_ ));
 sg13g2_nor2b_1 _8503_ (.A(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .B_N(_3653_),
    .Y(_3654_));
 sg13g2_o21ai_1 _8504_ (.B1(_3654_),
    .Y(_3655_),
    .A1(_1137_),
    .A2(_3652_));
 sg13g2_or4_1 _8505_ (.A(_1745_),
    .B(\i_dm_csrs.dmstatus_16_ ),
    .C(_1703_),
    .D(debug_req_o),
    .X(_3656_));
 sg13g2_nor2_1 _8506_ (.A(\i_dm_mem.state_q_0__$_NOT__A_Y ),
    .B(\i_dm_mem.state_q_1_ ),
    .Y(_3657_));
 sg13g2_a21oi_1 _8507_ (.A1(net556),
    .A2(_3656_),
    .Y(_3658_),
    .B1(_3657_));
 sg13g2_nand2_1 _8508_ (.Y(_3659_),
    .A(net556),
    .B(_3656_));
 sg13g2_and3_1 _8509_ (.X(_3660_),
    .A(cmd_valid),
    .B(halted),
    .C(_1206_));
 sg13g2_o21ai_1 _8510_ (.B1(_3655_),
    .Y(_3661_),
    .A1(_3659_),
    .A2(_3660_));
 sg13g2_o21ai_1 _8511_ (.B1(_3657_),
    .Y(_3662_),
    .A1(_1137_),
    .A2(_3160_));
 sg13g2_nand2b_1 _8512_ (.Y(_3663_),
    .B(_3662_),
    .A_N(_3661_));
 sg13g2_inv_1 _8513_ (.Y(_3664_),
    .A(\i_dm_mem.state_q_0_ ));
 sg13g2_a221oi_1 _8514_ (.B2(_3664_),
    .C1(ndmreset_o),
    .B1(_3663_),
    .A1(_3655_),
    .Y(_0586_),
    .A2(_3658_));
 sg13g2_nor2b_1 _8515_ (.A(\i_dm_mem.state_q_1_ ),
    .B_N(_3661_),
    .Y(_3665_));
 sg13g2_nor3_1 _8516_ (.A(_1137_),
    .B(_3099_),
    .C(_3160_),
    .Y(_3666_));
 sg13g2_nor3_1 _8517_ (.A(_0900_),
    .B(_3657_),
    .C(_3656_),
    .Y(_3667_));
 sg13g2_nor3_1 _8518_ (.A(_3661_),
    .B(_3666_),
    .C(_3667_),
    .Y(_3668_));
 sg13g2_nor3_1 _8519_ (.A(ndmreset_o),
    .B(_3665_),
    .C(_3668_),
    .Y(_0587_));
 sg13g2_inv_1 _8520_ (.Y(_3669_),
    .A(\i_dm_sba.state_q_0_ ));
 sg13g2_or2_1 _8521_ (.X(_3670_),
    .B(\i_dm_sba.state_q_1__$_NOT__A_Y ),
    .A(\i_dm_sba.state_q_0_ ));
 sg13g2_o21ai_1 _8522_ (.B1(_3670_),
    .Y(_3671_),
    .A1(\i_dm_sba.state_q_0__$_NOT__A_Y ),
    .A2(\i_dm_sba.state_q_1_ ));
 sg13g2_nand2b_2 _8523_ (.Y(_3672_),
    .B(_3671_),
    .A_N(\i_dm_sba.state_q_2_ ));
 sg13g2_or2_1 _8524_ (.X(_3673_),
    .B(_2561_),
    .A(net795));
 sg13g2_o21ai_1 _8525_ (.B1(_3673_),
    .Y(_3674_),
    .A1(master_gnt_i),
    .A2(_3672_));
 sg13g2_and2_1 _8526_ (.A(_3669_),
    .B(_3674_),
    .X(_3675_));
 sg13g2_nor3_2 _8527_ (.A(\i_dm_csrs.sbcs_q_12_ ),
    .B(\i_dm_csrs.sbcs_q_13_ ),
    .C(\i_dm_csrs.sbcs_q_14_ ),
    .Y(_3676_));
 sg13g2_nand4_1 _8528_ (.B(_0602_),
    .C(net803),
    .A(net141),
    .Y(_3677_),
    .D(_3676_));
 sg13g2_nand2_1 _8529_ (.Y(_3678_),
    .A(_3669_),
    .B(_3677_));
 sg13g2_nand2_1 _8530_ (.Y(_3679_),
    .A(\i_dm_sba.state_q_0__$_NOT__A_Y ),
    .B(_3678_));
 sg13g2_nor2_1 _8531_ (.A(_3679_),
    .B(_3674_),
    .Y(_3680_));
 sg13g2_nand3_1 _8532_ (.B(_0602_),
    .C(_3676_),
    .A(net142),
    .Y(_3681_));
 sg13g2_a21oi_1 _8533_ (.A1(\i_dm_csrs.sbcs_q_15_ ),
    .A2(_1169_),
    .Y(_3682_),
    .B1(_0611_));
 sg13g2_nor3_1 _8534_ (.A(\i_dm_csrs.sbcs_q_22_ ),
    .B(_3681_),
    .C(_3682_),
    .Y(_3683_));
 sg13g2_nand3_1 _8535_ (.B(net42),
    .C(_3683_),
    .A(net44),
    .Y(_3684_));
 sg13g2_nand4_1 _8536_ (.B(_2364_),
    .C(_2553_),
    .A(\i_dm_csrs.sbcs_q_20_ ),
    .Y(_3685_),
    .D(_3676_));
 sg13g2_and3_1 _8537_ (.X(_3686_),
    .A(_1255_),
    .B(_3684_),
    .C(_3685_));
 sg13g2_nor3_1 _8538_ (.A(\i_dm_sba.state_q_2_ ),
    .B(\i_dm_sba.state_q_1_ ),
    .C(_3686_),
    .Y(_3687_));
 sg13g2_nor2_1 _8539_ (.A(_3674_),
    .B(_3687_),
    .Y(_3688_));
 sg13g2_nor4_1 _8540_ (.A(_2811_),
    .B(_3675_),
    .C(_3680_),
    .D(_3688_),
    .Y(_0588_));
 sg13g2_nor2b_1 _8541_ (.A(\i_dm_sba.state_q_1_ ),
    .B_N(_3674_),
    .Y(_3689_));
 sg13g2_o21ai_1 _8542_ (.B1(\i_dm_sba.state_q_0__$_NOT__A_Y ),
    .Y(_3690_),
    .A1(\i_dm_sba.state_q_0_ ),
    .A2(_3677_));
 sg13g2_nor2_1 _8543_ (.A(_3674_),
    .B(_3690_),
    .Y(_3691_));
 sg13g2_nor4_1 _8544_ (.A(_2811_),
    .B(_3688_),
    .C(_3689_),
    .D(_3691_),
    .Y(_0589_));
 sg13g2_nand2_1 _8545_ (.Y(_3692_),
    .A(\i_dm_sba.state_q_2_ ),
    .B(_3674_));
 sg13g2_nor3_2 _8546_ (.A(\i_dm_sba.state_q_2_ ),
    .B(\i_dm_sba.state_q_0_ ),
    .C(\i_dm_sba.state_q_1__$_NOT__A_Y ),
    .Y(master_we_o));
 sg13g2_nor2b_1 _8547_ (.A(_3686_),
    .B_N(master_we_o),
    .Y(_3693_));
 sg13g2_nand2b_1 _8548_ (.Y(_3694_),
    .B(_3693_),
    .A_N(_3674_));
 sg13g2_a21oi_1 _8549_ (.A1(_3692_),
    .A2(_3694_),
    .Y(_0590_),
    .B1(_2811_));
 sg13g2_o21ai_1 _8550_ (.B1(_2717_),
    .Y(_3695_),
    .A1(_1496_),
    .A2(net546));
 sg13g2_nor3_1 _8551_ (.A(net632),
    .B(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_B ),
    .C(_2558_),
    .Y(_3696_));
 sg13g2_nand2b_1 _8552_ (.Y(_3697_),
    .B(_3696_),
    .A_N(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_A ));
 sg13g2_a21oi_2 _8553_ (.B1(_3672_),
    .Y(master_be_o_3_),
    .A2(_3697_),
    .A1(_3695_));
 sg13g2_nand2b_1 _8554_ (.Y(_3698_),
    .B(_3696_),
    .A_N(net51));
 sg13g2_a21oi_2 _8555_ (.B1(_3672_),
    .Y(master_be_o_2_),
    .A2(_3698_),
    .A1(_3695_));
 sg13g2_nand4_1 _8556_ (.B(_2557_),
    .C(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_B ),
    .A(_2833_),
    .Y(_3699_),
    .D(_2589_));
 sg13g2_and2_1 _8557_ (.A(_3695_),
    .B(_3699_),
    .X(_3700_));
 sg13g2_or4_1 _8558_ (.A(net632),
    .B(master_add_o_1_),
    .C(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_A ),
    .D(_2558_),
    .X(_3701_));
 sg13g2_a21oi_1 _8559_ (.A1(net632),
    .A2(net79),
    .Y(_3702_),
    .B1(net628));
 sg13g2_nand2b_1 _8560_ (.Y(_3703_),
    .B(_3702_),
    .A_N(_3672_));
 sg13g2_a21oi_2 _8561_ (.B1(_3703_),
    .Y(master_be_o_1_),
    .A2(_3701_),
    .A1(_3700_));
 sg13g2_nand3b_1 _8562_ (.B(_1496_),
    .C(_2589_),
    .Y(_3704_),
    .A_N(_2797_));
 sg13g2_a21oi_2 _8563_ (.B1(_3703_),
    .Y(master_be_o_0_),
    .A2(_3704_),
    .A1(_3700_));
 sg13g2_nor2_2 _8564_ (.A(_2811_),
    .B(_3672_),
    .Y(master_req_o));
 sg13g2_buf_2 fanout42 (.A(_1249_),
    .X(net42));
 sg13g2_buf_2 fanout41 (.A(_1255_),
    .X(net41));
 sg13g2_and2_1 _8567_ (.A(\i_dm_csrs.sbdata_o_23_ ),
    .B(net513),
    .X(_3707_));
 sg13g2_a21oi_1 _8568_ (.A1(\i_dm_csrs.sbdata_o_7_ ),
    .A2(net452),
    .Y(_3708_),
    .B1(_3707_));
 sg13g2_buf_1 fanout40 (.A(_3158_),
    .X(net40));
 sg13g2_buf_2 fanout39 (.A(net40),
    .X(net39));
 sg13g2_mux2_1 _8571_ (.A0(\i_dm_csrs.sbdata_o_15_ ),
    .A1(\i_dm_csrs.sbdata_o_31_ ),
    .S(net513),
    .X(_3711_));
 sg13g2_nor2_1 _8572_ (.A(net448),
    .B(_3711_),
    .Y(_3712_));
 sg13g2_a21oi_2 _8573_ (.B1(_3712_),
    .Y(master_wdata_o_31_),
    .A2(_3708_),
    .A1(net448));
 sg13g2_and2_1 _8574_ (.A(\i_dm_csrs.sbdata_o_22_ ),
    .B(net512),
    .X(_3713_));
 sg13g2_a21oi_1 _8575_ (.A1(\i_dm_csrs.sbdata_o_6_ ),
    .A2(net453),
    .Y(_3714_),
    .B1(_3713_));
 sg13g2_mux2_1 _8576_ (.A0(\i_dm_csrs.sbdata_o_14_ ),
    .A1(\i_dm_csrs.sbdata_o_30_ ),
    .S(net514),
    .X(_3715_));
 sg13g2_nor2_1 _8577_ (.A(net444),
    .B(_3715_),
    .Y(_3716_));
 sg13g2_a21oi_2 _8578_ (.B1(_3716_),
    .Y(master_wdata_o_30_),
    .A2(_3714_),
    .A1(net444));
 sg13g2_and2_1 _8579_ (.A(\i_dm_csrs.sbdata_o_21_ ),
    .B(net513),
    .X(_3717_));
 sg13g2_a21oi_1 _8580_ (.A1(\i_dm_csrs.sbdata_o_5_ ),
    .A2(net453),
    .Y(_3718_),
    .B1(_3717_));
 sg13g2_buf_1 fanout38 (.A(_0712_),
    .X(net38));
 sg13g2_nand3_1 _8582_ (.B(net511),
    .C(net449),
    .A(\i_dm_csrs.sbdata_o_13_ ),
    .Y(_3720_));
 sg13g2_o21ai_1 _8583_ (.B1(_3720_),
    .Y(master_wdata_o_21_),
    .A1(net444),
    .A2(_3718_));
 sg13g2_and2_1 _8584_ (.A(\i_dm_csrs.sbdata_o_20_ ),
    .B(net512),
    .X(_3721_));
 sg13g2_a21oi_1 _8585_ (.A1(\i_dm_csrs.sbdata_o_4_ ),
    .A2(net452),
    .Y(_3722_),
    .B1(_3721_));
 sg13g2_nand3_1 _8586_ (.B(net512),
    .C(net446),
    .A(\i_dm_csrs.sbdata_o_12_ ),
    .Y(_3723_));
 sg13g2_o21ai_1 _8587_ (.B1(_3723_),
    .Y(master_wdata_o_20_),
    .A1(net446),
    .A2(_3722_));
 sg13g2_and2_1 _8588_ (.A(\i_dm_csrs.sbdata_o_19_ ),
    .B(net512),
    .X(_3724_));
 sg13g2_a21oi_1 _8589_ (.A1(\i_dm_csrs.sbdata_o_3_ ),
    .A2(net452),
    .Y(_3725_),
    .B1(_3724_));
 sg13g2_nand3_1 _8590_ (.B(net512),
    .C(net447),
    .A(\i_dm_csrs.sbdata_o_11_ ),
    .Y(_3726_));
 sg13g2_o21ai_1 _8591_ (.B1(_3726_),
    .Y(master_wdata_o_19_),
    .A1(net446),
    .A2(_3725_));
 sg13g2_and2_1 _8592_ (.A(\i_dm_csrs.sbdata_o_18_ ),
    .B(net511),
    .X(_3727_));
 sg13g2_a21oi_1 _8593_ (.A1(\i_dm_csrs.sbdata_o_2_ ),
    .A2(net453),
    .Y(_3728_),
    .B1(_3727_));
 sg13g2_nand3_1 _8594_ (.B(net511),
    .C(net449),
    .A(\i_dm_csrs.sbdata_o_10_ ),
    .Y(_3729_));
 sg13g2_o21ai_1 _8595_ (.B1(_3729_),
    .Y(master_wdata_o_18_),
    .A1(net444),
    .A2(_3728_));
 sg13g2_and2_1 _8596_ (.A(\i_dm_csrs.sbdata_o_17_ ),
    .B(net513),
    .X(_3730_));
 sg13g2_a21oi_1 _8597_ (.A1(\i_dm_csrs.sbdata_o_1_ ),
    .A2(net452),
    .Y(_3731_),
    .B1(_3730_));
 sg13g2_nand3_1 _8598_ (.B(net513),
    .C(net448),
    .A(\i_dm_csrs.sbdata_o_9_ ),
    .Y(_3732_));
 sg13g2_o21ai_1 _8599_ (.B1(_3732_),
    .Y(master_wdata_o_17_),
    .A1(net448),
    .A2(_3731_));
 sg13g2_and2_1 _8600_ (.A(\i_dm_csrs.sbdata_o_16_ ),
    .B(net511),
    .X(_3733_));
 sg13g2_a21oi_1 _8601_ (.A1(\i_dm_csrs.sbdata_o_0_ ),
    .A2(net453),
    .Y(_3734_),
    .B1(_3733_));
 sg13g2_nand3_1 _8602_ (.B(net511),
    .C(net445),
    .A(\i_dm_csrs.sbdata_o_8_ ),
    .Y(_3735_));
 sg13g2_o21ai_1 _8603_ (.B1(_3735_),
    .Y(master_wdata_o_16_),
    .A1(net445),
    .A2(_3734_));
 sg13g2_nand2_1 _8604_ (.Y(_3736_),
    .A(\i_dm_csrs.sbdata_o_15_ ),
    .B(_2839_));
 sg13g2_buf_2 fanout37 (.A(net38),
    .X(net37));
 sg13g2_nand2_1 _8606_ (.Y(_3738_),
    .A(\i_dm_csrs.sbdata_o_7_ ),
    .B(net447));
 sg13g2_a21oi_2 _8607_ (.B1(net454),
    .Y(master_wdata_o_15_),
    .A2(_3738_),
    .A1(_3736_));
 sg13g2_nand2_1 _8608_ (.Y(_3739_),
    .A(\i_dm_csrs.sbdata_o_14_ ),
    .B(_2839_));
 sg13g2_nand2_1 _8609_ (.Y(_3740_),
    .A(\i_dm_csrs.sbdata_o_6_ ),
    .B(net445));
 sg13g2_a21oi_2 _8610_ (.B1(net453),
    .Y(master_wdata_o_14_),
    .A2(_3740_),
    .A1(_3739_));
 sg13g2_nand2_1 _8611_ (.Y(_3741_),
    .A(\i_dm_csrs.sbdata_o_13_ ),
    .B(_2839_));
 sg13g2_nand2_1 _8612_ (.Y(_3742_),
    .A(\i_dm_csrs.sbdata_o_5_ ),
    .B(net445));
 sg13g2_a21oi_2 _8613_ (.B1(net453),
    .Y(master_wdata_o_13_),
    .A2(_3742_),
    .A1(_3741_));
 sg13g2_nand2_1 _8614_ (.Y(_3743_),
    .A(\i_dm_csrs.sbdata_o_12_ ),
    .B(net505));
 sg13g2_nand2_1 _8615_ (.Y(_3744_),
    .A(\i_dm_csrs.sbdata_o_4_ ),
    .B(net445));
 sg13g2_a21oi_2 _8616_ (.B1(net453),
    .Y(master_wdata_o_12_),
    .A2(_3744_),
    .A1(_3743_));
 sg13g2_mux2_1 _8617_ (.A0(\i_dm_csrs.sbdata_o_13_ ),
    .A1(\i_dm_csrs.sbdata_o_29_ ),
    .S(net511),
    .X(_3745_));
 sg13g2_nor2_1 _8618_ (.A(net444),
    .B(_3745_),
    .Y(_3746_));
 sg13g2_a21oi_2 _8619_ (.B1(_3746_),
    .Y(master_wdata_o_29_),
    .A2(_3718_),
    .A1(net444));
 sg13g2_nand2_1 _8620_ (.Y(_3747_),
    .A(\i_dm_csrs.sbdata_o_11_ ),
    .B(net505));
 sg13g2_nand2_1 _8621_ (.Y(_3748_),
    .A(\i_dm_csrs.sbdata_o_3_ ),
    .B(net447));
 sg13g2_a21oi_2 _8622_ (.B1(net452),
    .Y(master_wdata_o_11_),
    .A2(_3748_),
    .A1(_3747_));
 sg13g2_nand2_1 _8623_ (.Y(_3749_),
    .A(\i_dm_csrs.sbdata_o_10_ ),
    .B(net505));
 sg13g2_nand2_1 _8624_ (.Y(_3750_),
    .A(\i_dm_csrs.sbdata_o_2_ ),
    .B(net447));
 sg13g2_a21oi_2 _8625_ (.B1(net452),
    .Y(master_wdata_o_10_),
    .A2(_3750_),
    .A1(_3749_));
 sg13g2_nand2_1 _8626_ (.Y(_3751_),
    .A(\i_dm_csrs.sbdata_o_1_ ),
    .B(net449));
 sg13g2_nand2_1 _8627_ (.Y(_3752_),
    .A(\i_dm_csrs.sbdata_o_9_ ),
    .B(net505));
 sg13g2_a21oi_2 _8628_ (.B1(net452),
    .Y(master_wdata_o_9_),
    .A2(_3752_),
    .A1(_3751_));
 sg13g2_nand2_1 _8629_ (.Y(_3753_),
    .A(\i_dm_csrs.sbdata_o_0_ ),
    .B(net447));
 sg13g2_nand2_1 _8630_ (.Y(_3754_),
    .A(\i_dm_csrs.sbdata_o_8_ ),
    .B(net505));
 sg13g2_a21oi_2 _8631_ (.B1(net452),
    .Y(master_wdata_o_8_),
    .A2(_3754_),
    .A1(_3753_));
 sg13g2_and2_2 _8632_ (.A(\i_dm_csrs.sbdata_o_7_ ),
    .B(net426),
    .X(master_wdata_o_7_));
 sg13g2_and2_2 _8633_ (.A(\i_dm_csrs.sbdata_o_6_ ),
    .B(net426),
    .X(master_wdata_o_6_));
 sg13g2_and2_2 _8634_ (.A(\i_dm_csrs.sbdata_o_5_ ),
    .B(net426),
    .X(master_wdata_o_5_));
 sg13g2_and2_2 _8635_ (.A(\i_dm_csrs.sbdata_o_4_ ),
    .B(net426),
    .X(master_wdata_o_4_));
 sg13g2_and2_2 _8636_ (.A(\i_dm_csrs.sbdata_o_3_ ),
    .B(net426),
    .X(master_wdata_o_3_));
 sg13g2_and2_2 _8637_ (.A(\i_dm_csrs.sbdata_o_2_ ),
    .B(net426),
    .X(master_wdata_o_2_));
 sg13g2_mux2_1 _8638_ (.A0(\i_dm_csrs.sbdata_o_12_ ),
    .A1(\i_dm_csrs.sbdata_o_28_ ),
    .S(net513),
    .X(_3755_));
 sg13g2_nor2_1 _8639_ (.A(net448),
    .B(_3755_),
    .Y(_3756_));
 sg13g2_a21oi_2 _8640_ (.B1(_3756_),
    .Y(master_wdata_o_28_),
    .A2(_3722_),
    .A1(net447));
 sg13g2_and2_2 _8641_ (.A(\i_dm_csrs.sbdata_o_1_ ),
    .B(net426),
    .X(master_wdata_o_1_));
 sg13g2_and2_2 _8642_ (.A(\i_dm_csrs.sbdata_o_0_ ),
    .B(net426),
    .X(master_wdata_o_0_));
 sg13g2_mux2_1 _8643_ (.A0(\i_dm_csrs.sbdata_o_11_ ),
    .A1(\i_dm_csrs.sbdata_o_27_ ),
    .S(net511),
    .X(_3757_));
 sg13g2_nor2_1 _8644_ (.A(net445),
    .B(_3757_),
    .Y(_3758_));
 sg13g2_a21oi_2 _8645_ (.B1(_3758_),
    .Y(master_wdata_o_27_),
    .A2(_3725_),
    .A1(net444));
 sg13g2_mux2_1 _8646_ (.A0(\i_dm_csrs.sbdata_o_10_ ),
    .A1(\i_dm_csrs.sbdata_o_26_ ),
    .S(net512),
    .X(_3759_));
 sg13g2_nor2_1 _8647_ (.A(net447),
    .B(_3759_),
    .Y(_3760_));
 sg13g2_a21oi_2 _8648_ (.B1(_3760_),
    .Y(master_wdata_o_26_),
    .A2(_3728_),
    .A1(net446));
 sg13g2_mux2_1 _8649_ (.A0(\i_dm_csrs.sbdata_o_9_ ),
    .A1(\i_dm_csrs.sbdata_o_25_ ),
    .S(net514),
    .X(_3761_));
 sg13g2_nor2_1 _8650_ (.A(net448),
    .B(_3761_),
    .Y(_3762_));
 sg13g2_a21oi_2 _8651_ (.B1(_3762_),
    .Y(master_wdata_o_25_),
    .A2(_3731_),
    .A1(net448));
 sg13g2_mux2_1 _8652_ (.A0(\i_dm_csrs.sbdata_o_8_ ),
    .A1(\i_dm_csrs.sbdata_o_24_ ),
    .S(net512),
    .X(_3763_));
 sg13g2_nor2_1 _8653_ (.A(net444),
    .B(_3763_),
    .Y(_3764_));
 sg13g2_a21oi_2 _8654_ (.B1(_3764_),
    .Y(master_wdata_o_24_),
    .A2(_3734_),
    .A1(net445));
 sg13g2_nand3_1 _8655_ (.B(net512),
    .C(net446),
    .A(\i_dm_csrs.sbdata_o_15_ ),
    .Y(_3765_));
 sg13g2_o21ai_1 _8656_ (.B1(_3765_),
    .Y(master_wdata_o_23_),
    .A1(net446),
    .A2(_3708_));
 sg13g2_nand3_1 _8657_ (.B(net511),
    .C(net446),
    .A(\i_dm_csrs.sbdata_o_14_ ),
    .Y(_3766_));
 sg13g2_o21ai_1 _8658_ (.B1(_3766_),
    .Y(master_wdata_o_22_),
    .A1(net446),
    .A2(_3714_));
 sg13g2_nand3_1 _8659_ (.B(_0893_),
    .C(_1120_),
    .A(ndmreset_o),
    .Y(_3767_));
 sg13g2_o21ai_1 _8660_ (.B1(_3767_),
    .Y(_0591_),
    .A1(_1120_),
    .A2(_0655_));
 sg13g2_buf_4 fanout36 (.X(net36),
    .A(net38));
 sg13g2_buf_4 fanout35 (.X(net35),
    .A(net38));
 sg13g2_mux2_2 _8663_ (.A0(\i_dm_mem.rdata_q_31_ ),
    .A1(\i_dm_mem.rdata_q_63_ ),
    .S(net53),
    .X(_3770_));
 sg13g2_nor2_1 _8664_ (.A(net577),
    .B(net545),
    .Y(_3771_));
 sg13g2_buf_4 fanout34 (.X(net34),
    .A(net38));
 sg13g2_buf_2 fanout33 (.A(_0713_),
    .X(net33));
 sg13g2_nor2_2 _8667_ (.A(net64),
    .B(net61),
    .Y(_3774_));
 sg13g2_nor2b_1 _8668_ (.A(net56),
    .B_N(net610),
    .Y(_3775_));
 sg13g2_nand3_1 _8669_ (.B(_3774_),
    .C(_3775_),
    .A(net496),
    .Y(_3776_));
 sg13g2_buf_2 fanout32 (.A(net440),
    .X(net32));
 sg13g2_buf_4 fanout31 (.X(net31),
    .A(net440));
 sg13g2_buf_4 fanout30 (.X(net30),
    .A(net440));
 sg13g2_buf_2 fanout29 (.A(net440),
    .X(net29));
 sg13g2_buf_2 fanout28 (.A(net440),
    .X(net28));
 sg13g2_inv_2 _8675_ (.Y(_3782_),
    .A(net52));
 sg13g2_nor2_2 _8676_ (.A(net67),
    .B(net575),
    .Y(_3783_));
 sg13g2_o21ai_1 _8677_ (.B1(_3783_),
    .Y(_3784_),
    .A1(net71),
    .A2(net542));
 sg13g2_nand2_1 _8678_ (.Y(_3785_),
    .A(net574),
    .B(_3784_));
 sg13g2_buf_4 fanout27 (.X(net27),
    .A(net440));
 sg13g2_nand2_2 _8680_ (.Y(_3787_),
    .A(net74),
    .B(net59));
 sg13g2_nand3_1 _8681_ (.B(_3785_),
    .C(_3787_),
    .A(net615),
    .Y(_3788_));
 sg13g2_a21oi_2 _8682_ (.B1(net64),
    .Y(_3789_),
    .A2(net68),
    .A1(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__$_NOT__A_Y ));
 sg13g2_nor2_1 _8683_ (.A(net573),
    .B(_3789_),
    .Y(_3790_));
 sg13g2_buf_4 fanout26 (.X(net26),
    .A(net440));
 sg13g2_a21oi_1 _8685_ (.A1(_3776_),
    .A2(_3788_),
    .Y(_3792_),
    .B1(net495));
 sg13g2_buf_2 fanout25 (.A(net440),
    .X(net25));
 sg13g2_buf_8 fanout24 (.A(_2829_),
    .X(net24));
 sg13g2_mux2_2 _8688_ (.A0(_3770_),
    .A1(_3792_),
    .S(net626),
    .X(slave_rdata_o_31_));
 sg13g2_buf_4 fanout23 (.X(net23),
    .A(net24));
 sg13g2_nor2_2 _8690_ (.A(net70),
    .B(net69),
    .Y(_3796_));
 sg13g2_nand2_1 _8691_ (.Y(_3797_),
    .A(net572),
    .B(_3796_));
 sg13g2_a21oi_1 _8692_ (.A1(_3787_),
    .A2(_3797_),
    .Y(_3798_),
    .B1(net616));
 sg13g2_nor2_2 _8693_ (.A(net544),
    .B(net575),
    .Y(_3799_));
 sg13g2_buf_16 fanout22 (.X(net22),
    .A(net24));
 sg13g2_nor2_1 _8695_ (.A(net64),
    .B(net609),
    .Y(_3801_));
 sg13g2_o21ai_1 _8696_ (.B1(net577),
    .Y(_3802_),
    .A1(_3799_),
    .A2(_3801_));
 sg13g2_nand2_1 _8697_ (.Y(_3803_),
    .A(net545),
    .B(_3774_));
 sg13g2_nor2b_2 _8698_ (.A(net61),
    .B_N(net610),
    .Y(_3804_));
 sg13g2_nor2_1 _8699_ (.A(net545),
    .B(_3804_),
    .Y(_3805_));
 sg13g2_o21ai_1 _8700_ (.B1(_3805_),
    .Y(_3806_),
    .A1(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__$_NOT__A_Y ),
    .A2(net572));
 sg13g2_buf_16 fanout21 (.X(net21),
    .A(net24));
 sg13g2_buf_16 fanout20 (.X(net20),
    .A(net24));
 sg13g2_buf_16 fanout19 (.X(net19),
    .A(net24));
 sg13g2_nand2_1 _8704_ (.Y(_3810_),
    .A(net621),
    .B(net541));
 sg13g2_a21oi_1 _8705_ (.A1(net66),
    .A2(net62),
    .Y(_3811_),
    .B1(_3810_));
 sg13g2_nand4_1 _8706_ (.B(_3803_),
    .C(_3806_),
    .A(_3802_),
    .Y(_3812_),
    .D(_3811_));
 sg13g2_buf_16 fanout18 (.X(net18),
    .A(net24));
 sg13g2_buf_4 fanout17 (.X(net17),
    .A(_3021_));
 sg13g2_nand2_1 _8709_ (.Y(_3815_),
    .A(net608),
    .B(_3799_));
 sg13g2_o21ai_1 _8710_ (.B1(_3815_),
    .Y(_3816_),
    .A1(net579),
    .A2(_3799_));
 sg13g2_buf_4 fanout16 (.X(net16),
    .A(_3021_));
 sg13g2_a21oi_1 _8712_ (.A1(net74),
    .A2(_3816_),
    .Y(_3818_),
    .B1(net61));
 sg13g2_nor2_1 _8713_ (.A(net493),
    .B(_3818_),
    .Y(_3819_));
 sg13g2_buf_2 fanout15 (.A(_3021_),
    .X(net15));
 sg13g2_mux2_1 _8715_ (.A0(\i_dm_mem.rdata_q_62_ ),
    .A1(_3819_),
    .S(net619),
    .X(_3821_));
 sg13g2_buf_4 fanout14 (.X(net14),
    .A(_3021_));
 sg13g2_nor3_1 _8717_ (.A(_3412_),
    .B(net618),
    .C(net58),
    .Y(_3823_));
 sg13g2_a21oi_1 _8718_ (.A1(net57),
    .A2(_3821_),
    .Y(_3824_),
    .B1(_3823_));
 sg13g2_o21ai_1 _8719_ (.B1(_3824_),
    .Y(slave_rdata_o_30_),
    .A1(_3798_),
    .A2(_3812_));
 sg13g2_buf_8 fanout13 (.A(_3021_),
    .X(net13));
 sg13g2_nand2_1 _8721_ (.Y(_3826_),
    .A(net63),
    .B(net570));
 sg13g2_a22oi_1 _8722_ (.Y(_3827_),
    .B1(_3826_),
    .B2(net613),
    .A2(_3804_),
    .A1(_3799_));
 sg13g2_buf_8 fanout12 (.A(_3021_),
    .X(net12));
 sg13g2_o21ai_1 _8724_ (.B1(net570),
    .Y(_3829_),
    .A1(net545),
    .A2(net63));
 sg13g2_nand2_1 _8725_ (.Y(_3830_),
    .A(net608),
    .B(_3829_));
 sg13g2_mux2_1 _8726_ (.A0(_3827_),
    .A1(_3830_),
    .S(net578),
    .X(_3831_));
 sg13g2_nor2_1 _8727_ (.A(net493),
    .B(_3831_),
    .Y(_3832_));
 sg13g2_nor2_1 _8728_ (.A(net579),
    .B(net69),
    .Y(_3833_));
 sg13g2_nand2_1 _8729_ (.Y(_3834_),
    .A(net73),
    .B(net575));
 sg13g2_o21ai_1 _8730_ (.B1(_3834_),
    .Y(_3835_),
    .A1(net71),
    .A2(_3826_));
 sg13g2_nand2_1 _8731_ (.Y(_3836_),
    .A(net63),
    .B(net608));
 sg13g2_nand2_1 _8732_ (.Y(_3837_),
    .A(net571),
    .B(_3836_));
 sg13g2_buf_8 fanout11 (.A(_3021_),
    .X(net11));
 sg13g2_buf_8 fanout10 (.A(_3021_),
    .X(net10));
 sg13g2_and2_1 _8735_ (.A(net59),
    .B(net609),
    .X(_3840_));
 sg13g2_a221oi_1 _8736_ (.B2(net72),
    .C1(_3840_),
    .B1(_3837_),
    .A1(_3833_),
    .Y(_3841_),
    .A2(_3835_));
 sg13g2_nor2_1 _8737_ (.A(net493),
    .B(_3841_),
    .Y(_3842_));
 sg13g2_buf_1 fanout9 (.A(_3106_),
    .X(net9));
 sg13g2_buf_2 fanout8 (.A(net9),
    .X(net8));
 sg13g2_mux4_1 _8740_ (.S0(net56),
    .A0(\i_dm_mem.rdata_q_21_ ),
    .A1(\i_dm_mem.rdata_q_53_ ),
    .A2(_3832_),
    .A3(_3842_),
    .S1(net620),
    .X(slave_rdata_o_21_));
 sg13g2_buf_2 fanout7 (.A(net9),
    .X(net7));
 sg13g2_nor2b_1 _8742_ (.A(net58),
    .B_N(\i_dm_mem.rdata_q_20_ ),
    .Y(_3846_));
 sg13g2_a21oi_1 _8743_ (.A1(\i_dm_mem.rdata_q_52_ ),
    .A2(net57),
    .Y(_3847_),
    .B1(_3846_));
 sg13g2_nor2b_2 _8744_ (.A(net495),
    .B_N(net624),
    .Y(_3848_));
 sg13g2_nor2_2 _8745_ (.A(net67),
    .B(net63),
    .Y(_3849_));
 sg13g2_a21oi_1 _8746_ (.A1(net613),
    .A2(_3849_),
    .Y(_3850_),
    .B1(_3799_));
 sg13g2_nor2_1 _8747_ (.A(net544),
    .B(net63),
    .Y(_3851_));
 sg13g2_o21ai_1 _8748_ (.B1(net609),
    .Y(_3852_),
    .A1(_3783_),
    .A2(_3851_));
 sg13g2_mux2_1 _8749_ (.A0(_3850_),
    .A1(_3852_),
    .S(net578),
    .X(_3853_));
 sg13g2_buf_2 fanout6 (.A(net9),
    .X(net6));
 sg13g2_nor2_1 _8751_ (.A(net571),
    .B(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ),
    .Y(_3855_));
 sg13g2_a21oi_1 _8752_ (.A1(net574),
    .A2(_3853_),
    .Y(_3856_),
    .B1(_3855_));
 sg13g2_nand2_1 _8753_ (.Y(_3857_),
    .A(_3848_),
    .B(_3856_));
 sg13g2_nand2_1 _8754_ (.Y(_3858_),
    .A(net62),
    .B(net610));
 sg13g2_nand3_1 _8755_ (.B(net574),
    .C(_3783_),
    .A(net614),
    .Y(_3859_));
 sg13g2_a21oi_1 _8756_ (.A1(_3858_),
    .A2(_3859_),
    .Y(_3860_),
    .B1(net578));
 sg13g2_nand2_1 _8757_ (.Y(_3861_),
    .A(_3848_),
    .B(_3860_));
 sg13g2_mux2_1 _8758_ (.A0(_3857_),
    .A1(_3861_),
    .S(net56),
    .X(_3862_));
 sg13g2_o21ai_1 _8759_ (.B1(_3862_),
    .Y(slave_rdata_o_20_),
    .A1(net624),
    .A2(_3847_));
 sg13g2_buf_2 fanout5 (.A(net9),
    .X(net5));
 sg13g2_nor3_2 _8761_ (.A(net579),
    .B(net75),
    .C(net570),
    .Y(_3864_));
 sg13g2_a21oi_2 _8762_ (.B1(net55),
    .Y(_3865_),
    .A2(_3864_),
    .A1(_3848_));
 sg13g2_nand2b_1 _8763_ (.Y(_3866_),
    .B(\i_dm_mem.rdata_q_19_ ),
    .A_N(net623));
 sg13g2_buf_2 fanout4 (.A(net9),
    .X(net4));
 sg13g2_nor2b_1 _8765_ (.A(net61),
    .B_N(net620),
    .Y(_3868_));
 sg13g2_nand4_1 _8766_ (.B(net75),
    .C(_3783_),
    .A(net614),
    .Y(_3869_),
    .D(_3868_));
 sg13g2_and2_1 _8767_ (.A(net55),
    .B(_3869_),
    .X(_3870_));
 sg13g2_nand2b_1 _8768_ (.Y(_3871_),
    .B(\i_dm_mem.rdata_q_51_ ),
    .A_N(net622));
 sg13g2_a22oi_1 _8769_ (.Y(slave_rdata_o_19_),
    .B1(_3870_),
    .B2(_3871_),
    .A2(_3866_),
    .A1(_3865_));
 sg13g2_buf_2 fanout3 (.A(net9),
    .X(net3));
 sg13g2_nor2_1 _8771_ (.A(net615),
    .B(net496),
    .Y(_3873_));
 sg13g2_o21ai_1 _8772_ (.B1(net576),
    .Y(_3874_),
    .A1(_3796_),
    .A2(_3873_));
 sg13g2_nor2_1 _8773_ (.A(net615),
    .B(net576),
    .Y(_3875_));
 sg13g2_nand2_1 _8774_ (.Y(_3876_),
    .A(net572),
    .B(net54));
 sg13g2_a21oi_1 _8775_ (.A1(net496),
    .A2(_3875_),
    .Y(_3877_),
    .B1(_3876_));
 sg13g2_nand2_1 _8776_ (.Y(_3878_),
    .A(net615),
    .B(net576));
 sg13g2_o21ai_1 _8777_ (.B1(net65),
    .Y(_3879_),
    .A1(net71),
    .A2(net611));
 sg13g2_a22oi_1 _8778_ (.Y(_3880_),
    .B1(_3879_),
    .B2(_3074_),
    .A2(_3878_),
    .A1(net496));
 sg13g2_nor2_1 _8779_ (.A(net60),
    .B(_3880_),
    .Y(_3881_));
 sg13g2_nor2_1 _8780_ (.A(net615),
    .B(net73),
    .Y(_3882_));
 sg13g2_o21ai_1 _8781_ (.B1(_3882_),
    .Y(_3883_),
    .A1(net61),
    .A2(_3799_));
 sg13g2_o21ai_1 _8782_ (.B1(_3883_),
    .Y(_3884_),
    .A1(net610),
    .A2(_3787_));
 sg13g2_nor4_1 _8783_ (.A(net53),
    .B(net494),
    .C(_3881_),
    .D(_3884_),
    .Y(_3885_));
 sg13g2_a21oi_1 _8784_ (.A1(_3874_),
    .A2(_3877_),
    .Y(_3886_),
    .B1(_3885_));
 sg13g2_mux2_1 _8785_ (.A0(\i_dm_mem.rdata_q_18_ ),
    .A1(\i_dm_mem.rdata_q_50_ ),
    .S(net53),
    .X(_3887_));
 sg13g2_nor2_1 _8786_ (.A(net626),
    .B(_3887_),
    .Y(_3888_));
 sg13g2_a21oi_2 _8787_ (.B1(_3888_),
    .Y(slave_rdata_o_18_),
    .A2(_3886_),
    .A1(net626));
 sg13g2_nand2b_1 _8788_ (.Y(_3889_),
    .B(\i_dm_mem.rdata_q_17_ ),
    .A_N(net622));
 sg13g2_nand2b_1 _8789_ (.Y(_3890_),
    .B(\i_dm_mem.rdata_q_49_ ),
    .A_N(net622));
 sg13g2_a22oi_1 _8790_ (.Y(slave_rdata_o_17_),
    .B1(_3890_),
    .B2(_3870_),
    .A2(_3889_),
    .A1(_3865_));
 sg13g2_nor2_1 _8791_ (.A(net53),
    .B(net494),
    .Y(_3891_));
 sg13g2_nor2_2 _8792_ (.A(_3066_),
    .B(net74),
    .Y(_3892_));
 sg13g2_nor2_1 _8793_ (.A(_3774_),
    .B(_3892_),
    .Y(_3893_));
 sg13g2_buf_2 fanout2 (.A(_3109_),
    .X(net2));
 sg13g2_o21ai_1 _8795_ (.B1(net69),
    .Y(_3895_),
    .A1(net65),
    .A2(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ));
 sg13g2_and2_1 _8796_ (.A(net70),
    .B(net612),
    .X(_3896_));
 sg13g2_o21ai_1 _8797_ (.B1(net62),
    .Y(_3897_),
    .A1(_3892_),
    .A2(_3896_));
 sg13g2_o21ai_1 _8798_ (.B1(_3897_),
    .Y(_3898_),
    .A1(_3893_),
    .A2(_3895_));
 sg13g2_nor2_2 _8799_ (.A(net70),
    .B(net544),
    .Y(_3899_));
 sg13g2_a21o_1 _8800_ (.A2(net66),
    .A1(net73),
    .B1(_3899_),
    .X(_3900_));
 sg13g2_nor2b_1 _8801_ (.A(net66),
    .B_N(net609),
    .Y(_3901_));
 sg13g2_nor2_1 _8802_ (.A(net71),
    .B(net575),
    .Y(_3902_));
 sg13g2_a21o_1 _8803_ (.A2(_3901_),
    .A1(net73),
    .B1(_3902_),
    .X(_3903_));
 sg13g2_a22oi_1 _8804_ (.Y(_3904_),
    .B1(_3903_),
    .B2(net69),
    .A2(_3900_),
    .A1(net616));
 sg13g2_inv_1 _8805_ (.Y(_3905_),
    .A(_3904_));
 sg13g2_nor2_2 _8806_ (.A(net59),
    .B(net542),
    .Y(_3906_));
 sg13g2_a22oi_1 _8807_ (.Y(_3907_),
    .B1(_3905_),
    .B2(_3906_),
    .A2(_3898_),
    .A1(_3891_));
 sg13g2_mux2_1 _8808_ (.A0(\i_dm_mem.rdata_q_16_ ),
    .A1(\i_dm_mem.rdata_q_48_ ),
    .S(net53),
    .X(_3908_));
 sg13g2_nor2_1 _8809_ (.A(net620),
    .B(_3908_),
    .Y(_3909_));
 sg13g2_a21oi_2 _8810_ (.B1(_3909_),
    .Y(slave_rdata_o_16_),
    .A2(_3907_),
    .A1(net621));
 sg13g2_nand2b_1 _8811_ (.Y(_3910_),
    .B(\i_dm_mem.rdata_q_15_ ),
    .A_N(net623));
 sg13g2_nand2b_1 _8812_ (.Y(_3911_),
    .B(\i_dm_mem.rdata_q_47_ ),
    .A_N(net622));
 sg13g2_a22oi_1 _8813_ (.Y(slave_rdata_o_15_),
    .B1(_3911_),
    .B2(_3870_),
    .A2(_3910_),
    .A1(_3865_));
 sg13g2_mux2_1 _8814_ (.A0(\i_dm_mem.rdata_q_14_ ),
    .A1(\i_dm_mem.rdata_q_46_ ),
    .S(net54),
    .X(_3912_));
 sg13g2_a21oi_1 _8815_ (.A1(net73),
    .A2(net56),
    .Y(_3913_),
    .B1(_3775_));
 sg13g2_o21ai_1 _8816_ (.B1(_3074_),
    .Y(_3914_),
    .A1(net575),
    .A2(_3913_));
 sg13g2_nand2_1 _8817_ (.Y(_3915_),
    .A(net573),
    .B(_3914_));
 sg13g2_nand4_1 _8818_ (.B(net542),
    .C(_3789_),
    .A(net62),
    .Y(_3916_),
    .D(_3892_));
 sg13g2_nand3_1 _8819_ (.B(net52),
    .C(_3899_),
    .A(net611),
    .Y(_3917_));
 sg13g2_o21ai_1 _8820_ (.B1(_3917_),
    .Y(_3918_),
    .A1(net67),
    .A2(_3913_));
 sg13g2_nand2_1 _8821_ (.Y(_3919_),
    .A(net577),
    .B(net542));
 sg13g2_nand3_1 _8822_ (.B(net68),
    .C(net52),
    .A(net73),
    .Y(_3920_));
 sg13g2_a21oi_1 _8823_ (.A1(_3919_),
    .A2(_3920_),
    .Y(_3921_),
    .B1(_3878_));
 sg13g2_a21oi_1 _8824_ (.A1(net65),
    .A2(_3918_),
    .Y(_3922_),
    .B1(_3921_));
 sg13g2_a21oi_1 _8825_ (.A1(_3915_),
    .A2(_3916_),
    .Y(_3923_),
    .B1(_3922_));
 sg13g2_nand2b_1 _8826_ (.Y(_3924_),
    .B(net625),
    .A_N(_3923_));
 sg13g2_o21ai_1 _8827_ (.B1(_3924_),
    .Y(_3925_),
    .A1(net625),
    .A2(_3912_));
 sg13g2_inv_16 _8828_ (.A(_3925_),
    .Y(slave_rdata_o_14_));
 sg13g2_nor2b_1 _8829_ (.A(net58),
    .B_N(\i_dm_mem.rdata_q_13_ ),
    .Y(_3926_));
 sg13g2_a21oi_2 _8830_ (.B1(_3926_),
    .Y(_3927_),
    .A2(net57),
    .A1(\i_dm_mem.rdata_q_45_ ));
 sg13g2_nand3_1 _8831_ (.B(net69),
    .C(net65),
    .A(net614),
    .Y(_3928_));
 sg13g2_a21oi_1 _8832_ (.A1(net574),
    .A2(_3928_),
    .Y(_3929_),
    .B1(net76));
 sg13g2_nor2_1 _8833_ (.A(net576),
    .B(net61),
    .Y(_3930_));
 sg13g2_and2_1 _8834_ (.A(net67),
    .B(net608),
    .X(_3931_));
 sg13g2_o21ai_1 _8835_ (.B1(net75),
    .Y(_3932_),
    .A1(_3930_),
    .A2(_3931_));
 sg13g2_nand3_1 _8836_ (.B(_3858_),
    .C(_3932_),
    .A(net58),
    .Y(_3933_));
 sg13g2_o21ai_1 _8837_ (.B1(net625),
    .Y(_3934_),
    .A1(net573),
    .A2(_3789_));
 sg13g2_nand2_1 _8838_ (.Y(_3935_),
    .A(net64),
    .B(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ));
 sg13g2_nand2_1 _8839_ (.Y(_3936_),
    .A(net69),
    .B(_3896_));
 sg13g2_o21ai_1 _8840_ (.B1(_3936_),
    .Y(_3937_),
    .A1(net68),
    .A2(_3935_));
 sg13g2_nor3_1 _8841_ (.A(net60),
    .B(net57),
    .C(_3937_),
    .Y(_3938_));
 sg13g2_nor2_1 _8842_ (.A(_3934_),
    .B(_3938_),
    .Y(_3939_));
 sg13g2_o21ai_1 _8843_ (.B1(_3939_),
    .Y(_3940_),
    .A1(_3929_),
    .A2(_3933_));
 sg13g2_o21ai_1 _8844_ (.B1(_3940_),
    .Y(slave_rdata_o_13_),
    .A1(net625),
    .A2(_3927_));
 sg13g2_buf_4 fanout1 (.X(net1),
    .A(_3109_));
 sg13g2_nand2_1 _8846_ (.Y(_3942_),
    .A(_3789_),
    .B(_3892_));
 sg13g2_nor2_2 _8847_ (.A(net577),
    .B(net68),
    .Y(_3943_));
 sg13g2_nor2_1 _8848_ (.A(_3899_),
    .B(_3943_),
    .Y(_3944_));
 sg13g2_nand2_1 _8849_ (.Y(_3945_),
    .A(net612),
    .B(_3796_));
 sg13g2_o21ai_1 _8850_ (.B1(_3945_),
    .Y(_3946_),
    .A1(_3066_),
    .A2(_3944_));
 sg13g2_a221oi_1 _8851_ (.B2(net65),
    .C1(net60),
    .B1(_3946_),
    .A1(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ),
    .Y(_3947_),
    .A2(_3851_));
 sg13g2_a21oi_1 _8852_ (.A1(net62),
    .A2(_3942_),
    .Y(_3948_),
    .B1(_3947_));
 sg13g2_inv_1 _8853_ (.Y(_3949_),
    .A(_3849_));
 sg13g2_nand2b_1 _8854_ (.Y(_3950_),
    .B(net63),
    .A_N(net609));
 sg13g2_a21oi_1 _8855_ (.A1(_3949_),
    .A2(_3950_),
    .Y(_3951_),
    .B1(net72));
 sg13g2_nor2_1 _8856_ (.A(net616),
    .B(net64),
    .Y(_3952_));
 sg13g2_nor4_1 _8857_ (.A(net496),
    .B(_3876_),
    .C(_3951_),
    .D(_3952_),
    .Y(_3953_));
 sg13g2_a21oi_1 _8858_ (.A1(net542),
    .A2(_3948_),
    .Y(_3954_),
    .B1(_3953_));
 sg13g2_mux2_1 _8859_ (.A0(\i_dm_mem.rdata_q_12_ ),
    .A1(\i_dm_mem.rdata_q_44_ ),
    .S(net54),
    .X(_3955_));
 sg13g2_nor2_1 _8860_ (.A(net619),
    .B(_3955_),
    .Y(_3956_));
 sg13g2_a21oi_2 _8861_ (.B1(_3956_),
    .Y(slave_rdata_o_12_),
    .A2(_3954_),
    .A1(net621));
 sg13g2_nand2_1 _8862_ (.Y(_3957_),
    .A(net575),
    .B(net611));
 sg13g2_o21ai_1 _8863_ (.B1(net573),
    .Y(_3958_),
    .A1(net544),
    .A2(_3957_));
 sg13g2_nand2_1 _8864_ (.Y(_3959_),
    .A(_3070_),
    .B(_3958_));
 sg13g2_o21ai_1 _8865_ (.B1(net573),
    .Y(_3960_),
    .A1(net67),
    .A2(net575));
 sg13g2_a22oi_1 _8866_ (.Y(_3961_),
    .B1(_3960_),
    .B2(net615),
    .A2(_3804_),
    .A1(net496));
 sg13g2_a21oi_1 _8867_ (.A1(_3959_),
    .A2(_3961_),
    .Y(_3962_),
    .B1(_3790_));
 sg13g2_nand3_1 _8868_ (.B(net63),
    .C(net608),
    .A(net68),
    .Y(_3963_));
 sg13g2_o21ai_1 _8869_ (.B1(_3963_),
    .Y(_3964_),
    .A1(net579),
    .A2(net67));
 sg13g2_nand2_1 _8870_ (.Y(_3965_),
    .A(net73),
    .B(_3964_));
 sg13g2_nand2_1 _8871_ (.Y(_3966_),
    .A(net61),
    .B(_3789_));
 sg13g2_o21ai_1 _8872_ (.B1(_3966_),
    .Y(_3967_),
    .A1(net60),
    .A2(_3965_));
 sg13g2_mux4_1 _8873_ (.S0(net56),
    .A0(\i_dm_mem.rdata_q_29_ ),
    .A1(\i_dm_mem.rdata_q_61_ ),
    .A2(_3962_),
    .A3(_3967_),
    .S1(net625),
    .X(slave_rdata_o_29_));
 sg13g2_nor2b_1 _8874_ (.A(net58),
    .B_N(\i_dm_mem.rdata_q_11_ ),
    .Y(_3968_));
 sg13g2_a21oi_1 _8875_ (.A1(\i_dm_mem.rdata_q_43_ ),
    .A2(net57),
    .Y(_3969_),
    .B1(_3968_));
 sg13g2_mux2_1 _8876_ (.A0(net610),
    .A1(net614),
    .S(net68),
    .X(_3970_));
 sg13g2_nand4_1 _8877_ (.B(_3868_),
    .C(_3902_),
    .A(net56),
    .Y(_3971_),
    .D(_3970_));
 sg13g2_o21ai_1 _8878_ (.B1(_3971_),
    .Y(_3972_),
    .A1(net55),
    .A2(_3861_));
 sg13g2_inv_1 _8879_ (.Y(_3973_),
    .A(_3972_));
 sg13g2_o21ai_1 _8880_ (.B1(_3973_),
    .Y(slave_rdata_o_11_),
    .A1(net624),
    .A2(_3969_));
 sg13g2_nand2_1 _8881_ (.Y(_3974_),
    .A(net577),
    .B(_3774_));
 sg13g2_a21oi_1 _8882_ (.A1(_3787_),
    .A2(_3974_),
    .Y(_3975_),
    .B1(net616));
 sg13g2_nor2_1 _8883_ (.A(net577),
    .B(net609),
    .Y(_3976_));
 sg13g2_o21ai_1 _8884_ (.B1(net65),
    .Y(_3977_),
    .A1(net60),
    .A2(_3976_));
 sg13g2_nand2_1 _8885_ (.Y(_3978_),
    .A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__$_NOT__A_Y ),
    .B(net67));
 sg13g2_o21ai_1 _8886_ (.B1(_3978_),
    .Y(_3979_),
    .A1(net71),
    .A2(net609));
 sg13g2_nand2_1 _8887_ (.Y(_3980_),
    .A(net62),
    .B(_3979_));
 sg13g2_nand3_1 _8888_ (.B(_3977_),
    .C(_3980_),
    .A(_3803_),
    .Y(_3981_));
 sg13g2_nor2_1 _8889_ (.A(_3975_),
    .B(_3981_),
    .Y(_3982_));
 sg13g2_nor2_2 _8890_ (.A(net544),
    .B(net61),
    .Y(_3983_));
 sg13g2_nand2_1 _8891_ (.Y(_3984_),
    .A(net570),
    .B(_3952_));
 sg13g2_o21ai_1 _8892_ (.B1(_3984_),
    .Y(_3985_),
    .A1(net608),
    .A2(_3983_));
 sg13g2_a221oi_1 _8893_ (.B2(net72),
    .C1(net494),
    .B1(_3985_),
    .A1(net571),
    .Y(_3986_),
    .A2(_3849_));
 sg13g2_mux4_1 _8894_ (.S0(net56),
    .A0(\i_dm_mem.rdata_q_10_ ),
    .A1(\i_dm_mem.rdata_q_42_ ),
    .A2(_3982_),
    .A3(_3986_),
    .S1(net620),
    .X(slave_rdata_o_10_));
 sg13g2_nand2_1 _8895_ (.Y(_3987_),
    .A(\i_dm_mem.rdata_q_41_ ),
    .B(net55));
 sg13g2_nand2_1 _8896_ (.Y(_3988_),
    .A(\i_dm_mem.rdata_q_9_ ),
    .B(_3782_));
 sg13g2_a21oi_2 _8897_ (.B1(net623),
    .Y(slave_rdata_o_9_),
    .A2(_3988_),
    .A1(_3987_));
 sg13g2_inv_1 _8898_ (.Y(_3989_),
    .A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ));
 sg13g2_nand2b_1 _8899_ (.Y(_3990_),
    .B(net578),
    .A_N(_3836_));
 sg13g2_o21ai_1 _8900_ (.B1(_3990_),
    .Y(_3991_),
    .A1(net65),
    .A2(_3989_));
 sg13g2_a22oi_1 _8901_ (.Y(_3992_),
    .B1(_3983_),
    .B2(_3991_),
    .A2(_3840_),
    .A1(net70));
 sg13g2_nor2_1 _8902_ (.A(net493),
    .B(_3992_),
    .Y(_3993_));
 sg13g2_o21ai_1 _8903_ (.B1(_3836_),
    .Y(_3994_),
    .A1(net71),
    .A2(_3952_));
 sg13g2_a22oi_1 _8904_ (.Y(_3995_),
    .B1(_3983_),
    .B2(_3994_),
    .A2(_3840_),
    .A1(net578));
 sg13g2_nor2_1 _8905_ (.A(net493),
    .B(_3995_),
    .Y(_3996_));
 sg13g2_mux4_1 _8906_ (.S0(net541),
    .A0(\i_dm_mem.rdata_q_40_ ),
    .A1(\i_dm_mem.rdata_q_8_ ),
    .A2(_3993_),
    .A3(_3996_),
    .S1(net620),
    .X(slave_rdata_o_8_));
 sg13g2_mux2_1 _8907_ (.A0(\i_dm_mem.rdata_q_7_ ),
    .A1(\i_dm_mem.rdata_q_39_ ),
    .S(net54),
    .X(_3997_));
 sg13g2_nand2b_1 _8908_ (.Y(_3998_),
    .B(_3997_),
    .A_N(net619));
 sg13g2_o21ai_1 _8909_ (.B1(_3998_),
    .Y(slave_rdata_o_7_),
    .A1(net54),
    .A2(_3869_));
 sg13g2_and2_1 _8910_ (.A(\i_dm_mem.rdata_q_38_ ),
    .B(net52),
    .X(_3999_));
 sg13g2_a21oi_1 _8911_ (.A1(\i_dm_mem.rdata_q_6_ ),
    .A2(_3782_),
    .Y(_4000_),
    .B1(_3999_));
 sg13g2_a21oi_1 _8912_ (.A1(net69),
    .A2(_3957_),
    .Y(_4001_),
    .B1(_3875_));
 sg13g2_nand2_1 _8913_ (.Y(_4002_),
    .A(net73),
    .B(_3801_));
 sg13g2_o21ai_1 _8914_ (.B1(_4002_),
    .Y(_4003_),
    .A1(net72),
    .A2(_4001_));
 sg13g2_nor2_1 _8915_ (.A(net615),
    .B(net577),
    .Y(_4004_));
 sg13g2_a22oi_1 _8916_ (.Y(_4005_),
    .B1(_4004_),
    .B2(_3960_),
    .A2(_4003_),
    .A1(net573));
 sg13g2_nor2b_1 _8917_ (.A(net74),
    .B_N(net610),
    .Y(_4006_));
 sg13g2_nand2_1 _8918_ (.Y(_4007_),
    .A(_3906_),
    .B(_3965_));
 sg13g2_a21oi_1 _8919_ (.A1(_3783_),
    .A2(_4006_),
    .Y(_4008_),
    .B1(_4007_));
 sg13g2_nor2_1 _8920_ (.A(_3934_),
    .B(_4008_),
    .Y(_4009_));
 sg13g2_o21ai_1 _8921_ (.B1(_4009_),
    .Y(_4010_),
    .A1(net54),
    .A2(_4005_));
 sg13g2_o21ai_1 _8922_ (.B1(_4010_),
    .Y(slave_rdata_o_6_),
    .A1(net625),
    .A2(_4000_));
 sg13g2_o21ai_1 _8923_ (.B1(net74),
    .Y(_4011_),
    .A1(net544),
    .A2(net611));
 sg13g2_nand2_1 _8924_ (.Y(_4012_),
    .A(net575),
    .B(_4011_));
 sg13g2_o21ai_1 _8925_ (.B1(_4012_),
    .Y(_4013_),
    .A1(net617),
    .A2(_3944_));
 sg13g2_a21oi_1 _8926_ (.A1(net573),
    .A2(_4013_),
    .Y(_4014_),
    .B1(net495));
 sg13g2_nor2b_1 _8927_ (.A(_3875_),
    .B_N(_4002_),
    .Y(_4015_));
 sg13g2_nand2_1 _8928_ (.Y(_4016_),
    .A(_3899_),
    .B(_3957_));
 sg13g2_o21ai_1 _8929_ (.B1(_4016_),
    .Y(_4017_),
    .A1(net68),
    .A2(_4015_));
 sg13g2_a21oi_1 _8930_ (.A1(net573),
    .A2(_4017_),
    .Y(_4018_),
    .B1(net495));
 sg13g2_mux4_1 _8931_ (.S0(_3782_),
    .A0(\i_dm_mem.rdata_q_37_ ),
    .A1(\i_dm_mem.rdata_q_5_ ),
    .A2(_4014_),
    .A3(_4018_),
    .S1(net626),
    .X(slave_rdata_o_5_));
 sg13g2_a21oi_1 _8932_ (.A1(net65),
    .A2(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ),
    .Y(_4019_),
    .B1(net68));
 sg13g2_o21ai_1 _8933_ (.B1(_3950_),
    .Y(_4020_),
    .A1(net64),
    .A2(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ));
 sg13g2_a21o_1 _8934_ (.A2(_3796_),
    .A1(_3066_),
    .B1(_3976_),
    .X(_4021_));
 sg13g2_a22oi_1 _8935_ (.Y(_4022_),
    .B1(_4021_),
    .B2(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3_ ),
    .A2(_4020_),
    .A1(net69));
 sg13g2_nor2_1 _8936_ (.A(net541),
    .B(_4022_),
    .Y(_4023_));
 sg13g2_a21oi_1 _8937_ (.A1(net542),
    .A2(_4019_),
    .Y(_4024_),
    .B1(_4023_));
 sg13g2_nand2_1 _8938_ (.Y(_4025_),
    .A(net615),
    .B(net72));
 sg13g2_nor2_1 _8939_ (.A(net54),
    .B(_4006_),
    .Y(_4026_));
 sg13g2_a21oi_1 _8940_ (.A1(_4025_),
    .A2(_4026_),
    .Y(_4027_),
    .B1(_3966_));
 sg13g2_a21oi_1 _8941_ (.A1(net572),
    .A2(_4024_),
    .Y(_4028_),
    .B1(_4027_));
 sg13g2_mux2_1 _8942_ (.A0(\i_dm_mem.rdata_q_4_ ),
    .A1(\i_dm_mem.rdata_q_36_ ),
    .S(net53),
    .X(_4029_));
 sg13g2_nor2_1 _8943_ (.A(net621),
    .B(_4029_),
    .Y(_4030_));
 sg13g2_a21oi_2 _8944_ (.B1(_4030_),
    .Y(slave_rdata_o_4_),
    .A2(_4028_),
    .A1(net621));
 sg13g2_or2_1 _8945_ (.X(_4031_),
    .B(_3810_),
    .A(net494));
 sg13g2_a21oi_1 _8946_ (.A1(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_2__$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ),
    .A2(_3774_),
    .Y(_4032_),
    .B1(_3864_));
 sg13g2_nor2b_1 _8947_ (.A(net618),
    .B_N(\i_dm_mem.rdata_q_3_ ),
    .Y(_4033_));
 sg13g2_nand2b_1 _8948_ (.Y(_4034_),
    .B(\i_dm_mem.rdata_q_35_ ),
    .A_N(net618));
 sg13g2_a21oi_1 _8949_ (.A1(_3869_),
    .A2(_4034_),
    .Y(_4035_),
    .B1(net541));
 sg13g2_a21oi_1 _8950_ (.A1(net541),
    .A2(_4033_),
    .Y(_4036_),
    .B1(_4035_));
 sg13g2_o21ai_1 _8951_ (.B1(_4036_),
    .Y(slave_rdata_o_3_),
    .A1(_4031_),
    .A2(_4032_));
 sg13g2_nand3_1 _8952_ (.B(net570),
    .C(_3931_),
    .A(net66),
    .Y(_4037_));
 sg13g2_o21ai_1 _8953_ (.B1(_4037_),
    .Y(_4038_),
    .A1(net579),
    .A2(net570));
 sg13g2_a22oi_1 _8954_ (.Y(_4039_),
    .B1(_4038_),
    .B2(net577),
    .A2(_3774_),
    .A1(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_2__$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ));
 sg13g2_nand3_1 _8955_ (.B(net70),
    .C(_3783_),
    .A(net616),
    .Y(_4040_));
 sg13g2_nand2_1 _8956_ (.Y(_4041_),
    .A(_3899_),
    .B(_3901_));
 sg13g2_a21oi_1 _8957_ (.A1(_4040_),
    .A2(_4041_),
    .Y(_4042_),
    .B1(net60));
 sg13g2_mux2_1 _8958_ (.A0(\i_dm_mem.rdata_q_34_ ),
    .A1(_4042_),
    .S(net618),
    .X(_4043_));
 sg13g2_nor3_1 _8959_ (.A(_3406_),
    .B(net618),
    .C(net58),
    .Y(_4044_));
 sg13g2_a21oi_1 _8960_ (.A1(net57),
    .A2(_4043_),
    .Y(_4045_),
    .B1(_4044_));
 sg13g2_o21ai_1 _8961_ (.B1(_4045_),
    .Y(slave_rdata_o_2_),
    .A1(_4031_),
    .A2(_4039_));
 sg13g2_or2_1 _8962_ (.X(_4046_),
    .B(_3931_),
    .A(net59));
 sg13g2_a22oi_1 _8963_ (.Y(_4047_),
    .B1(_4046_),
    .B2(net74),
    .A2(_3833_),
    .A1(_3930_));
 sg13g2_a21oi_1 _8964_ (.A1(_3830_),
    .A2(_4047_),
    .Y(_4048_),
    .B1(net493));
 sg13g2_o21ai_1 _8965_ (.B1(net614),
    .Y(_4049_),
    .A1(_3799_),
    .A2(_3943_));
 sg13g2_or2_1 _8966_ (.X(_4050_),
    .B(net611),
    .A(net64));
 sg13g2_a21oi_1 _8967_ (.A1(_3771_),
    .A2(_4050_),
    .Y(_4051_),
    .B1(net60));
 sg13g2_a21oi_1 _8968_ (.A1(_4049_),
    .A2(_4051_),
    .Y(_4052_),
    .B1(net494));
 sg13g2_mux4_1 _8969_ (.S0(net56),
    .A0(\i_dm_mem.rdata_q_28_ ),
    .A1(\i_dm_mem.rdata_q_60_ ),
    .A2(_4048_),
    .A3(_4052_),
    .S1(net620),
    .X(slave_rdata_o_28_));
 sg13g2_nand2_1 _8970_ (.Y(_4053_),
    .A(\i_dm_mem.rdata_q_33_ ),
    .B(net52));
 sg13g2_o21ai_1 _8971_ (.B1(_4053_),
    .Y(_4054_),
    .A1(_3266_),
    .A2(net55));
 sg13g2_nor2_1 _8972_ (.A(net622),
    .B(_4054_),
    .Y(_4055_));
 sg13g2_a21oi_2 _8973_ (.B1(_4055_),
    .Y(slave_rdata_o_1_),
    .A2(net495),
    .A1(net622));
 sg13g2_nand2_1 _8974_ (.Y(_4056_),
    .A(\i_dm_mem.rdata_q_32_ ),
    .B(net52));
 sg13g2_o21ai_1 _8975_ (.B1(_4056_),
    .Y(_4057_),
    .A1(_3086_),
    .A2(net55));
 sg13g2_nor2_1 _8976_ (.A(net622),
    .B(_4057_),
    .Y(_4058_));
 sg13g2_a21oi_2 _8977_ (.B1(_4058_),
    .Y(slave_rdata_o_0_),
    .A2(net495),
    .A1(net622));
 sg13g2_o21ai_1 _8978_ (.B1(_3826_),
    .Y(_4059_),
    .A1(net571),
    .A2(net608));
 sg13g2_nand2_1 _8979_ (.Y(_4060_),
    .A(net608),
    .B(_3834_));
 sg13g2_nand2_1 _8980_ (.Y(_4061_),
    .A(net545),
    .B(net570));
 sg13g2_a21oi_1 _8981_ (.A1(_3787_),
    .A2(_4061_),
    .Y(_4062_),
    .B1(net613));
 sg13g2_a221oi_1 _8982_ (.B2(_3983_),
    .C1(_4062_),
    .B1(_4060_),
    .A1(net578),
    .Y(_4063_),
    .A2(_4059_));
 sg13g2_o21ai_1 _8983_ (.B1(net62),
    .Y(_4064_),
    .A1(net71),
    .A2(net610));
 sg13g2_and2_1 _8984_ (.A(net52),
    .B(_4064_),
    .X(_4065_));
 sg13g2_a21oi_1 _8985_ (.A1(_3965_),
    .A2(_4065_),
    .Y(_4066_),
    .B1(net495));
 sg13g2_o21ai_1 _8986_ (.B1(_4066_),
    .Y(_4067_),
    .A1(net54),
    .A2(_4063_));
 sg13g2_mux2_1 _8987_ (.A0(\i_dm_mem.rdata_q_27_ ),
    .A1(\i_dm_mem.rdata_q_59_ ),
    .S(net53),
    .X(_4068_));
 sg13g2_nor2_1 _8988_ (.A(net624),
    .B(_4068_),
    .Y(_4069_));
 sg13g2_a21oi_2 _8989_ (.B1(_4069_),
    .Y(slave_rdata_o_27_),
    .A2(_4067_),
    .A1(net625));
 sg13g2_nor2_1 _8990_ (.A(net60),
    .B(_3949_),
    .Y(_4070_));
 sg13g2_a21oi_1 _8991_ (.A1(net75),
    .A2(_4070_),
    .Y(_4071_),
    .B1(_3864_));
 sg13g2_nor2b_1 _8992_ (.A(net618),
    .B_N(\i_dm_mem.rdata_q_26_ ),
    .Y(_4072_));
 sg13g2_nand2b_1 _8993_ (.Y(_4073_),
    .B(\i_dm_mem.rdata_q_58_ ),
    .A_N(net618));
 sg13g2_a21oi_1 _8994_ (.A1(_3869_),
    .A2(_4073_),
    .Y(_4074_),
    .B1(net541));
 sg13g2_a21oi_1 _8995_ (.A1(net541),
    .A2(_4072_),
    .Y(_4075_),
    .B1(_4074_));
 sg13g2_o21ai_1 _8996_ (.B1(_4075_),
    .Y(slave_rdata_o_26_),
    .A1(_4031_),
    .A2(_4071_));
 sg13g2_o21ai_1 _8997_ (.B1(net614),
    .Y(_4076_),
    .A1(net59),
    .A2(_3943_));
 sg13g2_nand3_1 _8998_ (.B(_3771_),
    .C(_3804_),
    .A(net66),
    .Y(_4077_));
 sg13g2_and2_1 _8999_ (.A(_4076_),
    .B(_4077_),
    .X(_4078_));
 sg13g2_a21oi_1 _9000_ (.A1(_3959_),
    .A2(_4078_),
    .Y(_4079_),
    .B1(net494));
 sg13g2_o21ai_1 _9001_ (.B1(_3990_),
    .Y(_4080_),
    .A1(net579),
    .A2(_3834_));
 sg13g2_nand2_1 _9002_ (.Y(_4081_),
    .A(net570),
    .B(_3963_));
 sg13g2_a221oi_1 _9003_ (.B2(net72),
    .C1(_3840_),
    .B1(_4081_),
    .A1(net544),
    .Y(_4082_),
    .A2(_4080_));
 sg13g2_nor2_1 _9004_ (.A(net493),
    .B(_4082_),
    .Y(_4083_));
 sg13g2_mux4_1 _9005_ (.S0(net55),
    .A0(\i_dm_mem.rdata_q_25_ ),
    .A1(\i_dm_mem.rdata_q_57_ ),
    .A2(_4079_),
    .A3(_4083_),
    .S1(net619),
    .X(slave_rdata_o_25_));
 sg13g2_nor2b_1 _9006_ (.A(net57),
    .B_N(\i_dm_mem.rdata_q_24_ ),
    .Y(_4084_));
 sg13g2_a21oi_1 _9007_ (.A1(\i_dm_mem.rdata_q_56_ ),
    .A2(net57),
    .Y(_4085_),
    .B1(_4084_));
 sg13g2_a21oi_1 _9008_ (.A1(net544),
    .A2(_3902_),
    .Y(_4086_),
    .B1(net59));
 sg13g2_nand2_1 _9009_ (.Y(_4087_),
    .A(net74),
    .B(_3983_));
 sg13g2_o21ai_1 _9010_ (.B1(_4087_),
    .Y(_4088_),
    .A1(net70),
    .A2(net64));
 sg13g2_o21ai_1 _9011_ (.B1(net542),
    .Y(_4089_),
    .A1(net70),
    .A2(net574));
 sg13g2_a221oi_1 _9012_ (.B2(net610),
    .C1(_4089_),
    .B1(_4088_),
    .A1(_3774_),
    .Y(_4090_),
    .A2(_3943_));
 sg13g2_o21ai_1 _9013_ (.B1(_4090_),
    .Y(_4091_),
    .A1(net579),
    .A2(_4086_));
 sg13g2_nand3_1 _9014_ (.B(_4007_),
    .C(_4091_),
    .A(_3848_),
    .Y(_4092_));
 sg13g2_o21ai_1 _9015_ (.B1(_4092_),
    .Y(slave_rdata_o_24_),
    .A1(net625),
    .A2(_4085_));
 sg13g2_a21oi_1 _9016_ (.A1(net613),
    .A2(_3774_),
    .Y(_4093_),
    .B1(_3840_));
 sg13g2_a221oi_1 _9017_ (.B2(net613),
    .C1(net72),
    .B1(_4061_),
    .A1(_3804_),
    .Y(_4094_),
    .A2(_3849_));
 sg13g2_a21oi_1 _9018_ (.A1(net75),
    .A2(_4093_),
    .Y(_4095_),
    .B1(_4094_));
 sg13g2_o21ai_1 _9019_ (.B1(net616),
    .Y(_4096_),
    .A1(_3783_),
    .A2(_3851_));
 sg13g2_a21oi_1 _9020_ (.A1(_3963_),
    .A2(_4096_),
    .Y(_4097_),
    .B1(net71));
 sg13g2_a21o_1 _9021_ (.A2(_3901_),
    .A1(net496),
    .B1(_4097_),
    .X(_4098_));
 sg13g2_a22oi_1 _9022_ (.Y(_4099_),
    .B1(_4098_),
    .B2(_3906_),
    .A2(_4095_),
    .A1(_3891_));
 sg13g2_nand2_1 _9023_ (.Y(_4100_),
    .A(\i_dm_mem.rdata_q_55_ ),
    .B(net52));
 sg13g2_o21ai_1 _9024_ (.B1(_4100_),
    .Y(_4101_),
    .A1(_3318_),
    .A2(net55));
 sg13g2_nor2_1 _9025_ (.A(net618),
    .B(_4101_),
    .Y(_4102_));
 sg13g2_a21oi_2 _9026_ (.B1(_4102_),
    .Y(slave_rdata_o_23_),
    .A2(_4099_),
    .A1(net621));
 sg13g2_a22oi_1 _9027_ (.Y(_4103_),
    .B1(_3829_),
    .B2(net613),
    .A2(_3804_),
    .A1(_3799_));
 sg13g2_nand4_1 _9028_ (.B(net75),
    .C(net545),
    .A(net613),
    .Y(_4104_),
    .D(_3930_));
 sg13g2_o21ai_1 _9029_ (.B1(_4104_),
    .Y(_4105_),
    .A1(net72),
    .A2(_4103_));
 sg13g2_nor2_1 _9030_ (.A(net541),
    .B(net493),
    .Y(_4106_));
 sg13g2_nand2_1 _9031_ (.Y(_4107_),
    .A(net74),
    .B(_3949_));
 sg13g2_a22oi_1 _9032_ (.Y(_4108_),
    .B1(_4107_),
    .B2(net616),
    .A2(_3901_),
    .A1(net496));
 sg13g2_nor3_1 _9033_ (.A(net59),
    .B(net58),
    .C(_4108_),
    .Y(_4109_));
 sg13g2_a21oi_1 _9034_ (.A1(_4105_),
    .A2(_4106_),
    .Y(_4110_),
    .B1(_4109_));
 sg13g2_mux2_1 _9035_ (.A0(\i_dm_mem.rdata_q_22_ ),
    .A1(\i_dm_mem.rdata_q_54_ ),
    .S(net53),
    .X(_4111_));
 sg13g2_nor2_1 _9036_ (.A(net619),
    .B(_4111_),
    .Y(_4112_));
 sg13g2_a21oi_2 _9037_ (.B1(_4112_),
    .Y(slave_rdata_o_22_),
    .A2(_4110_),
    .A1(net621));
 sg13g2_dfrbp_2 cmd_0__reg (.RESET_B(net747),
    .D(_0003_),
    .Q(cmd_0_),
    .Q_N(_4678_),
    .CLK(clknet_leaf_72_clk_i));
 sg13g2_dfrbp_1 cmd_10__reg (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net746),
    .D(_0004_),
    .Q_N(_4677_),
    .Q(cmd_10_));
 sg13g2_dfrbp_2 cmd_11__reg (.RESET_B(net746),
    .D(_0005_),
    .Q(cmd_11_),
    .Q_N(_4676_),
    .CLK(clknet_leaf_41_clk_i));
 sg13g2_dfrbp_1 cmd_12__reg (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net733),
    .D(_0006_),
    .Q_N(\i_dm_mem.abstract_cmd_132__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ),
    .Q(cmd_12_));
 sg13g2_dfrbp_1 cmd_14__reg (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net743),
    .D(_0007_),
    .Q_N(_4675_),
    .Q(cmd_14_));
 sg13g2_dfrbp_1 cmd_15__reg (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net743),
    .D(_0008_),
    .Q_N(_4674_),
    .Q(cmd_15_));
 sg13g2_dfrbp_2 cmd_16__reg (.RESET_B(net731),
    .D(_0009_),
    .Q(cmd_16_),
    .Q_N(\cmd_16__$_NOT__A_Y ),
    .CLK(clknet_leaf_73_clk_i));
 sg13g2_dfrbp_1 cmd_17__reg (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net731),
    .D(_0010_),
    .Q_N(\cmd_17__$_NOT__A_Y ),
    .Q(cmd_17_));
 sg13g2_dfrbp_1 cmd_18__reg (.CLK(clknet_leaf_74_clk_i),
    .RESET_B(net731),
    .D(_0011_),
    .Q_N(_4673_),
    .Q(cmd_18_));
 sg13g2_dfrbp_1 cmd_19__reg (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net742),
    .D(_0012_),
    .Q_N(_4672_),
    .Q(cmd_19_));
 sg13g2_dfrbp_1 cmd_1__reg (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net733),
    .D(_0013_),
    .Q_N(\cmd_0__$_OR__A_B ),
    .Q(cmd_1_));
 sg13g2_dfrbp_2 cmd_20__reg (.RESET_B(net746),
    .D(_0014_),
    .Q(cmd_20_),
    .Q_N(_4671_),
    .CLK(clknet_leaf_73_clk_i));
 sg13g2_dfrbp_2 cmd_21__reg (.RESET_B(net746),
    .D(_0015_),
    .Q(cmd_21_),
    .Q_N(_4670_),
    .CLK(clknet_leaf_73_clk_i));
 sg13g2_dfrbp_1 cmd_22__reg (.CLK(clknet_leaf_73_clk_i),
    .RESET_B(net731),
    .D(_0016_),
    .Q_N(\cmd_19__$_OR__B_A_$_OR__Y_B_$_AND__Y_A ),
    .Q(cmd_22_));
 sg13g2_dfrbp_1 cmd_24__reg (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(_0017_),
    .Q_N(_4669_),
    .Q(cmd_24_));
 sg13g2_dfrbp_1 cmd_25__reg (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(_0018_),
    .Q_N(_4668_),
    .Q(cmd_25_));
 sg13g2_dfrbp_1 cmd_26__reg (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(_0019_),
    .Q_N(_4667_),
    .Q(cmd_26_));
 sg13g2_dfrbp_1 cmd_27__reg (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net723),
    .D(_0020_),
    .Q_N(_4666_),
    .Q(cmd_27_));
 sg13g2_dfrbp_1 cmd_28__reg (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net755),
    .D(_0021_),
    .Q_N(_4665_),
    .Q(cmd_28_));
 sg13g2_dfrbp_1 cmd_29__reg (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net755),
    .D(_0022_),
    .Q_N(_4664_),
    .Q(cmd_29_));
 sg13g2_dfrbp_2 cmd_2__reg (.RESET_B(net747),
    .D(_0023_),
    .Q(cmd_2_),
    .Q_N(_4663_),
    .CLK(clknet_leaf_72_clk_i));
 sg13g2_dfrbp_1 cmd_30__reg (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net755),
    .D(_0024_),
    .Q_N(_4662_),
    .Q(cmd_30_));
 sg13g2_dfrbp_1 cmd_31__reg (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net755),
    .D(_0025_),
    .Q_N(_4661_),
    .Q(cmd_31_));
 sg13g2_dfrbp_2 cmd_3__reg (.RESET_B(net733),
    .D(_0026_),
    .Q(cmd_3_),
    .Q_N(\cmd_3__$_NOT__A_Y ),
    .CLK(clknet_leaf_71_clk_i));
 sg13g2_dfrbp_2 cmd_4__reg (.RESET_B(net747),
    .D(_0027_),
    .Q(cmd_4_),
    .Q_N(_4660_),
    .CLK(clknet_leaf_72_clk_i));
 sg13g2_dfrbp_1 cmd_5__reg (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net733),
    .D(_0028_),
    .Q_N(\cmd_5__$_NOT__A_Y ),
    .Q(cmd_5_));
 sg13g2_dfrbp_2 cmd_6__reg (.RESET_B(net743),
    .D(_0029_),
    .Q(cmd_6_),
    .Q_N(_4659_),
    .CLK(clknet_leaf_40_clk_i));
 sg13g2_dfrbp_1 cmd_7__reg (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net742),
    .D(_0030_),
    .Q_N(_4658_),
    .Q(cmd_7_));
 sg13g2_dfrbp_1 cmd_8__reg (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net746),
    .D(_0031_),
    .Q_N(_4657_),
    .Q(cmd_8_));
 sg13g2_dfrbp_1 cmd_9__reg (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net746),
    .D(_0032_),
    .Q_N(_4679_),
    .Q(cmd_9_));
 sg13g2_dfrbp_1 cmd_valid_reg (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net715),
    .D(cmd_valid_reg_D),
    .Q_N(_4656_),
    .Q(cmd_valid));
 sg13g2_dfrbp_1 data_csrs_mem_0__reg (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net693),
    .D(_0033_),
    .Q_N(_4655_),
    .Q(data_csrs_mem_0_));
 sg13g2_dfrbp_1 data_csrs_mem_10__reg (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net713),
    .D(_0034_),
    .Q_N(_4654_),
    .Q(data_csrs_mem_10_));
 sg13g2_dfrbp_1 data_csrs_mem_11__reg (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net713),
    .D(_0035_),
    .Q_N(_4653_),
    .Q(data_csrs_mem_11_));
 sg13g2_dfrbp_1 data_csrs_mem_12__reg (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net678),
    .D(_0036_),
    .Q_N(_4652_),
    .Q(data_csrs_mem_12_));
 sg13g2_dfrbp_1 data_csrs_mem_13__reg (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net690),
    .D(_0037_),
    .Q_N(_4651_),
    .Q(data_csrs_mem_13_));
 sg13g2_dfrbp_1 data_csrs_mem_14__reg (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net693),
    .D(_0038_),
    .Q_N(_4650_),
    .Q(data_csrs_mem_14_));
 sg13g2_dfrbp_1 data_csrs_mem_15__reg (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net715),
    .D(_0039_),
    .Q_N(_4649_),
    .Q(data_csrs_mem_15_));
 sg13g2_dfrbp_1 data_csrs_mem_16__reg (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net702),
    .D(_0040_),
    .Q_N(_4648_),
    .Q(data_csrs_mem_16_));
 sg13g2_dfrbp_1 data_csrs_mem_17__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net702),
    .D(_0041_),
    .Q_N(_4647_),
    .Q(data_csrs_mem_17_));
 sg13g2_dfrbp_1 data_csrs_mem_18__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net703),
    .D(_0042_),
    .Q_N(_4646_),
    .Q(data_csrs_mem_18_));
 sg13g2_dfrbp_1 data_csrs_mem_19__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net703),
    .D(_0043_),
    .Q_N(_4645_),
    .Q(data_csrs_mem_19_));
 sg13g2_dfrbp_1 data_csrs_mem_1__reg (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net693),
    .D(_0044_),
    .Q_N(_4644_),
    .Q(data_csrs_mem_1_));
 sg13g2_dfrbp_1 data_csrs_mem_20__reg (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net702),
    .D(_0045_),
    .Q_N(_4643_),
    .Q(data_csrs_mem_20_));
 sg13g2_dfrbp_1 data_csrs_mem_21__reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net702),
    .D(_0046_),
    .Q_N(_4642_),
    .Q(data_csrs_mem_21_));
 sg13g2_dfrbp_2 data_csrs_mem_22__reg (.RESET_B(net703),
    .D(_0047_),
    .Q(data_csrs_mem_22_),
    .Q_N(_4641_),
    .CLK(clknet_leaf_20_clk_i));
 sg13g2_dfrbp_2 data_csrs_mem_23__reg (.RESET_B(net679),
    .D(_0048_),
    .Q(data_csrs_mem_23_),
    .Q_N(_4640_),
    .CLK(clknet_leaf_12_clk_i));
 sg13g2_dfrbp_1 data_csrs_mem_24__reg (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net679),
    .D(_0049_),
    .Q_N(_4639_),
    .Q(data_csrs_mem_24_));
 sg13g2_dfrbp_1 data_csrs_mem_25__reg (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net679),
    .D(_0050_),
    .Q_N(_4638_),
    .Q(data_csrs_mem_25_));
 sg13g2_dfrbp_2 data_csrs_mem_26__reg (.RESET_B(net678),
    .D(_0051_),
    .Q(data_csrs_mem_26_),
    .Q_N(_4637_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_1 data_csrs_mem_27__reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net679),
    .D(_0052_),
    .Q_N(_4636_),
    .Q(data_csrs_mem_27_));
 sg13g2_dfrbp_1 data_csrs_mem_28__reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net679),
    .D(_0053_),
    .Q_N(_4635_),
    .Q(data_csrs_mem_28_));
 sg13g2_dfrbp_1 data_csrs_mem_29__reg (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net678),
    .D(_0054_),
    .Q_N(_4634_),
    .Q(data_csrs_mem_29_));
 sg13g2_dfrbp_1 data_csrs_mem_2__reg (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net690),
    .D(_0055_),
    .Q_N(_4633_),
    .Q(data_csrs_mem_2_));
 sg13g2_dfrbp_1 data_csrs_mem_30__reg (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net678),
    .D(_0056_),
    .Q_N(_4632_),
    .Q(data_csrs_mem_30_));
 sg13g2_dfrbp_2 data_csrs_mem_31__reg (.RESET_B(net690),
    .D(_0057_),
    .Q(data_csrs_mem_31_),
    .Q_N(_4631_),
    .CLK(clknet_leaf_92_clk_i));
 sg13g2_dfrbp_1 data_csrs_mem_32__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net693),
    .D(_0058_),
    .Q_N(_4630_),
    .Q(data_csrs_mem_32_));
 sg13g2_dfrbp_1 data_csrs_mem_33__reg (.CLK(clknet_leaf_88_clk_i),
    .RESET_B(net693),
    .D(_0059_),
    .Q_N(_4629_),
    .Q(data_csrs_mem_33_));
 sg13g2_dfrbp_1 data_csrs_mem_34__reg (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net690),
    .D(_0060_),
    .Q_N(_4628_),
    .Q(data_csrs_mem_34_));
 sg13g2_dfrbp_1 data_csrs_mem_35__reg (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net692),
    .D(_0061_),
    .Q_N(_4627_),
    .Q(data_csrs_mem_35_));
 sg13g2_dfrbp_1 data_csrs_mem_36__reg (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net692),
    .D(_0062_),
    .Q_N(_4626_),
    .Q(data_csrs_mem_36_));
 sg13g2_dfrbp_1 data_csrs_mem_37__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net691),
    .D(_0063_),
    .Q_N(_4625_),
    .Q(data_csrs_mem_37_));
 sg13g2_dfrbp_1 data_csrs_mem_38__reg (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net691),
    .D(_0064_),
    .Q_N(_4624_),
    .Q(data_csrs_mem_38_));
 sg13g2_dfrbp_1 data_csrs_mem_39__reg (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net690),
    .D(_0065_),
    .Q_N(_4623_),
    .Q(data_csrs_mem_39_));
 sg13g2_dfrbp_1 data_csrs_mem_3__reg (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net692),
    .D(_0066_),
    .Q_N(_4622_),
    .Q(data_csrs_mem_3_));
 sg13g2_dfrbp_1 data_csrs_mem_40__reg (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net692),
    .D(_0067_),
    .Q_N(_4621_),
    .Q(data_csrs_mem_40_));
 sg13g2_dfrbp_1 data_csrs_mem_41__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net691),
    .D(_0068_),
    .Q_N(_4620_),
    .Q(data_csrs_mem_41_));
 sg13g2_dfrbp_1 data_csrs_mem_42__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net713),
    .D(_0069_),
    .Q_N(_4619_),
    .Q(data_csrs_mem_42_));
 sg13g2_dfrbp_1 data_csrs_mem_43__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net713),
    .D(_0070_),
    .Q_N(_4618_),
    .Q(data_csrs_mem_43_));
 sg13g2_dfrbp_1 data_csrs_mem_44__reg (.CLK(clknet_leaf_11_clk_i),
    .RESET_B(net680),
    .D(_0071_),
    .Q_N(_4617_),
    .Q(data_csrs_mem_44_));
 sg13g2_dfrbp_1 data_csrs_mem_45__reg (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net690),
    .D(_0072_),
    .Q_N(_4616_),
    .Q(data_csrs_mem_45_));
 sg13g2_dfrbp_1 data_csrs_mem_46__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net693),
    .D(_0073_),
    .Q_N(_4615_),
    .Q(data_csrs_mem_46_));
 sg13g2_dfrbp_1 data_csrs_mem_47__reg (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net713),
    .D(_0074_),
    .Q_N(_4614_),
    .Q(data_csrs_mem_47_));
 sg13g2_dfrbp_1 data_csrs_mem_48__reg (.CLK(clknet_leaf_13_clk_i),
    .RESET_B(net680),
    .D(_0075_),
    .Q_N(_4613_),
    .Q(data_csrs_mem_48_));
 sg13g2_dfrbp_1 data_csrs_mem_49__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net713),
    .D(_0076_),
    .Q_N(_4612_),
    .Q(data_csrs_mem_49_));
 sg13g2_dfrbp_1 data_csrs_mem_4__reg (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net692),
    .D(_0077_),
    .Q_N(_4611_),
    .Q(data_csrs_mem_4_));
 sg13g2_dfrbp_1 data_csrs_mem_50__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net713),
    .D(_0078_),
    .Q_N(_4610_),
    .Q(data_csrs_mem_50_));
 sg13g2_dfrbp_1 data_csrs_mem_51__reg (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net713),
    .D(_0079_),
    .Q_N(_4609_),
    .Q(data_csrs_mem_51_));
 sg13g2_dfrbp_1 data_csrs_mem_52__reg (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net702),
    .D(_0080_),
    .Q_N(_4608_),
    .Q(data_csrs_mem_52_));
 sg13g2_dfrbp_1 data_csrs_mem_53__reg (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net702),
    .D(_0081_),
    .Q_N(_4607_),
    .Q(data_csrs_mem_53_));
 sg13g2_dfrbp_2 data_csrs_mem_54__reg (.RESET_B(net703),
    .D(_0082_),
    .Q(data_csrs_mem_54_),
    .Q_N(_4606_),
    .CLK(clknet_leaf_20_clk_i));
 sg13g2_dfrbp_2 data_csrs_mem_55__reg (.RESET_B(net691),
    .D(_0083_),
    .Q(data_csrs_mem_55_),
    .Q_N(_4605_),
    .CLK(clknet_leaf_12_clk_i));
 sg13g2_dfrbp_1 data_csrs_mem_56__reg (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net679),
    .D(_0084_),
    .Q_N(_4604_),
    .Q(data_csrs_mem_56_));
 sg13g2_dfrbp_1 data_csrs_mem_57__reg (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net679),
    .D(_0085_),
    .Q_N(_4603_),
    .Q(data_csrs_mem_57_));
 sg13g2_dfrbp_1 data_csrs_mem_58__reg (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net678),
    .D(_0086_),
    .Q_N(_4602_),
    .Q(data_csrs_mem_58_));
 sg13g2_dfrbp_1 data_csrs_mem_59__reg (.CLK(clknet_leaf_12_clk_i),
    .RESET_B(net691),
    .D(_0087_),
    .Q_N(_4601_),
    .Q(data_csrs_mem_59_));
 sg13g2_dfrbp_1 data_csrs_mem_5__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net695),
    .D(_0088_),
    .Q_N(_4600_),
    .Q(data_csrs_mem_5_));
 sg13g2_dfrbp_1 data_csrs_mem_60__reg (.CLK(clknet_leaf_9_clk_i),
    .RESET_B(net679),
    .D(_0089_),
    .Q_N(_4599_),
    .Q(data_csrs_mem_60_));
 sg13g2_dfrbp_1 data_csrs_mem_61__reg (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net678),
    .D(_0090_),
    .Q_N(_4598_),
    .Q(data_csrs_mem_61_));
 sg13g2_dfrbp_1 data_csrs_mem_62__reg (.CLK(clknet_leaf_10_clk_i),
    .RESET_B(net680),
    .D(_0091_),
    .Q_N(_4597_),
    .Q(data_csrs_mem_62_));
 sg13g2_dfrbp_2 data_csrs_mem_63__reg (.RESET_B(net690),
    .D(_0092_),
    .Q(data_csrs_mem_63_),
    .Q_N(_4596_),
    .CLK(clknet_leaf_11_clk_i));
 sg13g2_dfrbp_1 data_csrs_mem_6__reg (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net695),
    .D(_0093_),
    .Q_N(_4595_),
    .Q(data_csrs_mem_6_));
 sg13g2_dfrbp_1 data_csrs_mem_7__reg (.CLK(clknet_leaf_91_clk_i),
    .RESET_B(net691),
    .D(_0094_),
    .Q_N(_4594_),
    .Q(data_csrs_mem_7_));
 sg13g2_dfrbp_1 data_csrs_mem_8__reg (.CLK(clknet_leaf_89_clk_i),
    .RESET_B(net692),
    .D(_0095_),
    .Q_N(_4593_),
    .Q(data_csrs_mem_8_));
 sg13g2_dfrbp_1 data_csrs_mem_9__reg (.CLK(clknet_leaf_14_clk_i),
    .RESET_B(net695),
    .D(_0096_),
    .Q_N(_4592_),
    .Q(data_csrs_mem_9_));
 sg13g2_dfrbp_2 debug_req_o_reg (.RESET_B(net742),
    .D(_0097_),
    .Q(debug_req_o),
    .Q_N(_4591_),
    .CLK(clknet_leaf_40_clk_i));
 sg13g2_dfrbp_2 dmactive_o_reg (.RESET_B(net748),
    .D(_0098_),
    .Q(dmactive_o),
    .Q_N(\ndmreset_o_reg_E_$_AND__Y_B_$_OR__Y_A ),
    .CLK(clknet_leaf_44_clk_i));
 sg13g2_dfrbp_2 halted_reg (.RESET_B(net715),
    .D(_0099_),
    .Q(halted),
    .Q_N(\i_dm_csrs.dmstatus_11__$_AND__Y_A ),
    .CLK(clknet_leaf_39_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_0__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net722),
    .D(_0100_),
    .Q_N(_4590_),
    .Q(\i_dm_csrs.abstractauto_q_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_16__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net714),
    .D(_0101_),
    .Q_N(_4589_),
    .Q(\i_dm_csrs.abstractauto_q_16_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_17__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net714),
    .D(_0102_),
    .Q_N(_4588_),
    .Q(\i_dm_csrs.abstractauto_q_17_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_18__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net721),
    .D(_0103_),
    .Q_N(_4587_),
    .Q(\i_dm_csrs.abstractauto_q_18_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_19__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net716),
    .D(_0104_),
    .Q_N(_4586_),
    .Q(\i_dm_csrs.abstractauto_q_19_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_1__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net722),
    .D(_0105_),
    .Q_N(_4585_),
    .Q(\i_dm_csrs.abstractauto_q_1_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_20__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net717),
    .D(_0106_),
    .Q_N(_4584_),
    .Q(\i_dm_csrs.abstractauto_q_20_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_21__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net717),
    .D(_0107_),
    .Q_N(_4583_),
    .Q(\i_dm_csrs.abstractauto_q_21_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_22__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net721),
    .D(_0108_),
    .Q_N(_4582_),
    .Q(\i_dm_csrs.abstractauto_q_22_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.abstractauto_q_23__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net721),
    .D(_0109_),
    .Q_N(_4680_),
    .Q(\i_dm_csrs.abstractauto_q_23_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.cmderr_q_0__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net742),
    .D(\i_dm_csrs.cmderr_q_0__reg_D ),
    .Q_N(_4681_),
    .Q(\i_dm_csrs.cmderr_q_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.cmderr_q_1__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net715),
    .D(\i_dm_csrs.cmderr_q_1__reg_D ),
    .Q_N(_4682_),
    .Q(\i_dm_csrs.cmderr_q_1_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.cmderr_q_2__reg  (.RESET_B(net715),
    .D(\i_dm_csrs.cmderr_q_2__reg_D ),
    .Q(\i_dm_csrs.cmderr_q_2_ ),
    .Q_N(_4581_),
    .CLK(clknet_leaf_39_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.havereset_q_reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net714),
    .D(_0002_),
    .Q_N(\i_dm_csrs.dmstatus_18_ ),
    .Q(_0000_));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_0__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net768),
    .D(_0110_),
    .Q_N(_4580_),
    .Q(\i_dm_csrs.i_fifo.mem_q_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_10__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net767),
    .D(_0111_),
    .Q_N(_4579_),
    .Q(\i_dm_csrs.i_fifo.mem_q_10_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_11__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net768),
    .D(_0112_),
    .Q_N(_4578_),
    .Q(\i_dm_csrs.i_fifo.mem_q_11_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_12__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net774),
    .D(_0113_),
    .Q_N(_4577_),
    .Q(\i_dm_csrs.i_fifo.mem_q_12_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_13__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net765),
    .D(_0114_),
    .Q_N(_4576_),
    .Q(\i_dm_csrs.i_fifo.mem_q_13_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_14__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net772),
    .D(_0115_),
    .Q_N(_4575_),
    .Q(\i_dm_csrs.i_fifo.mem_q_14_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_15__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net767),
    .D(_0116_),
    .Q_N(_4574_),
    .Q(\i_dm_csrs.i_fifo.mem_q_15_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_16__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0117_),
    .Q_N(_4573_),
    .Q(\i_dm_csrs.i_fifo.mem_q_16_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_17__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net772),
    .D(_0118_),
    .Q_N(_4572_),
    .Q(\i_dm_csrs.i_fifo.mem_q_17_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_18__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net768),
    .D(_0119_),
    .Q_N(_4571_),
    .Q(\i_dm_csrs.i_fifo.mem_q_18_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_19__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0120_),
    .Q_N(_4570_),
    .Q(\i_dm_csrs.i_fifo.mem_q_19_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_1__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net768),
    .D(_0121_),
    .Q_N(_4569_),
    .Q(\i_dm_csrs.i_fifo.mem_q_1_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_20__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net767),
    .D(_0122_),
    .Q_N(_4568_),
    .Q(\i_dm_csrs.i_fifo.mem_q_20_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_21__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0123_),
    .Q_N(_4567_),
    .Q(\i_dm_csrs.i_fifo.mem_q_21_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_22__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net772),
    .D(_0124_),
    .Q_N(_4566_),
    .Q(\i_dm_csrs.i_fifo.mem_q_22_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_23__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net774),
    .D(_0125_),
    .Q_N(_4565_),
    .Q(\i_dm_csrs.i_fifo.mem_q_23_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_24__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0126_),
    .Q_N(_4564_),
    .Q(\i_dm_csrs.i_fifo.mem_q_24_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_25__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net772),
    .D(_0127_),
    .Q_N(_4563_),
    .Q(\i_dm_csrs.i_fifo.mem_q_25_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_26__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net774),
    .D(_0128_),
    .Q_N(_4562_),
    .Q(\i_dm_csrs.i_fifo.mem_q_26_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_27__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0129_),
    .Q_N(_4561_),
    .Q(\i_dm_csrs.i_fifo.mem_q_27_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_28__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net764),
    .D(_0130_),
    .Q_N(_4560_),
    .Q(\i_dm_csrs.i_fifo.mem_q_28_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_29__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net765),
    .D(_0131_),
    .Q_N(_4559_),
    .Q(\i_dm_csrs.i_fifo.mem_q_29_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_2__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net772),
    .D(_0132_),
    .Q_N(_4558_),
    .Q(\i_dm_csrs.i_fifo.mem_q_2_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_30__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net774),
    .D(_0133_),
    .Q_N(_4557_),
    .Q(\i_dm_csrs.i_fifo.mem_q_30_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_31__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net764),
    .D(_0134_),
    .Q_N(_4556_),
    .Q(\i_dm_csrs.i_fifo.mem_q_31_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_32__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0135_),
    .Q_N(_4555_),
    .Q(\i_dm_csrs.i_fifo.mem_q_32_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_33__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net768),
    .D(_0136_),
    .Q_N(_4554_),
    .Q(\i_dm_csrs.i_fifo.mem_q_33_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_34__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net768),
    .D(_0137_),
    .Q_N(_4553_),
    .Q(\i_dm_csrs.i_fifo.mem_q_34_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_35__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net768),
    .D(_0138_),
    .Q_N(_4552_),
    .Q(\i_dm_csrs.i_fifo.mem_q_35_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_36__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net772),
    .D(_0139_),
    .Q_N(_4551_),
    .Q(\i_dm_csrs.i_fifo.mem_q_36_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_37__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net773),
    .D(_0140_),
    .Q_N(_4550_),
    .Q(\i_dm_csrs.i_fifo.mem_q_37_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_38__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net774),
    .D(_0141_),
    .Q_N(_4549_),
    .Q(\i_dm_csrs.i_fifo.mem_q_38_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_39__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net766),
    .D(_0142_),
    .Q_N(_4548_),
    .Q(\i_dm_csrs.i_fifo.mem_q_39_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_3__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net773),
    .D(_0143_),
    .Q_N(_4547_),
    .Q(\i_dm_csrs.i_fifo.mem_q_3_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_40__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net767),
    .D(_0144_),
    .Q_N(_4546_),
    .Q(\i_dm_csrs.i_fifo.mem_q_40_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_41__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net764),
    .D(_0145_),
    .Q_N(_4545_),
    .Q(\i_dm_csrs.i_fifo.mem_q_41_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_42__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net764),
    .D(_0146_),
    .Q_N(_4544_),
    .Q(\i_dm_csrs.i_fifo.mem_q_42_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_43__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net775),
    .D(_0147_),
    .Q_N(_4543_),
    .Q(\i_dm_csrs.i_fifo.mem_q_43_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_44__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net767),
    .D(_0148_),
    .Q_N(_4542_),
    .Q(\i_dm_csrs.i_fifo.mem_q_44_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_45__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net769),
    .D(_0149_),
    .Q_N(_4541_),
    .Q(\i_dm_csrs.i_fifo.mem_q_45_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_46__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net775),
    .D(_0150_),
    .Q_N(_4540_),
    .Q(\i_dm_csrs.i_fifo.mem_q_46_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_47__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net765),
    .D(_0151_),
    .Q_N(_4539_),
    .Q(\i_dm_csrs.i_fifo.mem_q_47_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_48__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net772),
    .D(_0152_),
    .Q_N(_4538_),
    .Q(\i_dm_csrs.i_fifo.mem_q_48_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_49__reg  (.CLK(clknet_leaf_64_clk_i),
    .RESET_B(net767),
    .D(_0153_),
    .Q_N(_4537_),
    .Q(\i_dm_csrs.i_fifo.mem_q_49_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_4__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net774),
    .D(_0154_),
    .Q_N(_4536_),
    .Q(\i_dm_csrs.i_fifo.mem_q_4_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_50__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0155_),
    .Q_N(_4535_),
    .Q(\i_dm_csrs.i_fifo.mem_q_50_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_51__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net772),
    .D(_0156_),
    .Q_N(_4534_),
    .Q(\i_dm_csrs.i_fifo.mem_q_51_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_52__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net768),
    .D(_0157_),
    .Q_N(_4533_),
    .Q(\i_dm_csrs.i_fifo.mem_q_52_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_53__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0158_),
    .Q_N(_4532_),
    .Q(\i_dm_csrs.i_fifo.mem_q_53_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_54__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net767),
    .D(_0159_),
    .Q_N(_4531_),
    .Q(\i_dm_csrs.i_fifo.mem_q_54_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_55__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0160_),
    .Q_N(_4530_),
    .Q(\i_dm_csrs.i_fifo.mem_q_55_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_56__reg  (.CLK(clknet_leaf_59_clk_i),
    .RESET_B(net773),
    .D(_0161_),
    .Q_N(_4529_),
    .Q(\i_dm_csrs.i_fifo.mem_q_56_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_57__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net774),
    .D(_0162_),
    .Q_N(_4528_),
    .Q(\i_dm_csrs.i_fifo.mem_q_57_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_58__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0163_),
    .Q_N(_4527_),
    .Q(\i_dm_csrs.i_fifo.mem_q_58_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_59__reg  (.CLK(clknet_leaf_58_clk_i),
    .RESET_B(net773),
    .D(_0164_),
    .Q_N(_4526_),
    .Q(\i_dm_csrs.i_fifo.mem_q_59_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_5__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net766),
    .D(_0165_),
    .Q_N(_4525_),
    .Q(\i_dm_csrs.i_fifo.mem_q_5_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_60__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net775),
    .D(_0166_),
    .Q_N(_4524_),
    .Q(\i_dm_csrs.i_fifo.mem_q_60_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_61__reg  (.CLK(clknet_leaf_56_clk_i),
    .RESET_B(net776),
    .D(_0167_),
    .Q_N(_4523_),
    .Q(\i_dm_csrs.i_fifo.mem_q_61_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_62__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net764),
    .D(_0168_),
    .Q_N(_4522_),
    .Q(\i_dm_csrs.i_fifo.mem_q_62_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_63__reg  (.CLK(clknet_leaf_63_clk_i),
    .RESET_B(net765),
    .D(_0169_),
    .Q_N(_4521_),
    .Q(\i_dm_csrs.i_fifo.mem_q_63_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_64__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net774),
    .D(_0170_),
    .Q_N(_4520_),
    .Q(\i_dm_csrs.i_fifo.mem_q_64_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_65__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net764),
    .D(_0171_),
    .Q_N(_4519_),
    .Q(\i_dm_csrs.i_fifo.mem_q_65_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_66__reg  (.CLK(clknet_leaf_65_clk_i),
    .RESET_B(net766),
    .D(_0172_),
    .Q_N(_4518_),
    .Q(\i_dm_csrs.i_fifo.mem_q_66_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_67__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net769),
    .D(_0173_),
    .Q_N(_4517_),
    .Q(\i_dm_csrs.i_fifo.mem_q_67_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_6__reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net767),
    .D(_0174_),
    .Q_N(_4516_),
    .Q(\i_dm_csrs.i_fifo.mem_q_6_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_7__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net764),
    .D(_0175_),
    .Q_N(_4515_),
    .Q(\i_dm_csrs.i_fifo.mem_q_7_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_8__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net764),
    .D(_0176_),
    .Q_N(_4514_),
    .Q(\i_dm_csrs.i_fifo.mem_q_8_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.mem_q_9__reg  (.CLK(clknet_leaf_57_clk_i),
    .RESET_B(net775),
    .D(_0177_),
    .Q_N(_4513_),
    .Q(\i_dm_csrs.i_fifo.mem_q_9_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.i_fifo.read_pointer_q_reg  (.RESET_B(net773),
    .D(_0178_),
    .Q(\i_dm_csrs.i_fifo.read_pointer_q ),
    .Q_N(\i_dm_csrs.i_fifo.read_pointer_n ),
    .CLK(clknet_leaf_60_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.status_cnt_q_1__reg  (.CLK(clknet_leaf_61_clk_i),
    .RESET_B(net773),
    .D(_0179_),
    .Q_N(\i_dm_csrs.i_fifo.full_o_$_NOT__Y_A_$_OR__Y_B ),
    .Q(\i_dm_csrs.i_fifo.status_cnt_q_1_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.usage_o_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net773),
    .D(_0180_),
    .Q_N(\i_dm_csrs.i_fifo.status_cnt_n_0_ ),
    .Q(\i_dm_csrs.i_fifo.status_cnt_q_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.i_fifo.write_pointer_q_reg  (.CLK(clknet_leaf_60_clk_i),
    .RESET_B(net769),
    .D(_0181_),
    .Q_N(\i_dm_csrs.i_fifo.write_pointer_n ),
    .Q(\i_dm_csrs.i_fifo.write_pointer_q ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_0__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net693),
    .D(_0182_),
    .Q_N(_4512_),
    .Q(\i_dm_csrs.progbuf_o_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_100__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net683),
    .D(_0183_),
    .Q_N(_4511_),
    .Q(\i_dm_csrs.progbuf_o_100_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_101__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net698),
    .D(_0184_),
    .Q_N(_4510_),
    .Q(\i_dm_csrs.progbuf_o_101_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_102__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net691),
    .D(_0185_),
    .Q_N(_4509_),
    .Q(\i_dm_csrs.progbuf_o_102_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_103__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net682),
    .D(_0186_),
    .Q_N(_4508_),
    .Q(\i_dm_csrs.progbuf_o_103_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_104__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0187_),
    .Q_N(_4507_),
    .Q(\i_dm_csrs.progbuf_o_104_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_105__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net717),
    .D(_0188_),
    .Q_N(_4506_),
    .Q(\i_dm_csrs.progbuf_o_105_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_106__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net705),
    .D(_0189_),
    .Q_N(_4505_),
    .Q(\i_dm_csrs.progbuf_o_106_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_107__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net675),
    .D(_0190_),
    .Q_N(_4504_),
    .Q(\i_dm_csrs.progbuf_o_107_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_108__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net674),
    .D(_0191_),
    .Q_N(_4503_),
    .Q(\i_dm_csrs.progbuf_o_108_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_109__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net669),
    .D(_0192_),
    .Q_N(_4502_),
    .Q(\i_dm_csrs.progbuf_o_109_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_10__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net705),
    .D(_0193_),
    .Q_N(_4501_),
    .Q(\i_dm_csrs.progbuf_o_10_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_110__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net685),
    .D(_0194_),
    .Q_N(_4500_),
    .Q(\i_dm_csrs.progbuf_o_110_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_111__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net681),
    .D(_0195_),
    .Q_N(_4499_),
    .Q(\i_dm_csrs.progbuf_o_111_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_112__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net704),
    .D(_0196_),
    .Q_N(_4498_),
    .Q(\i_dm_csrs.progbuf_o_112_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_113__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0197_),
    .Q_N(_4497_),
    .Q(\i_dm_csrs.progbuf_o_113_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_114__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net700),
    .D(_0198_),
    .Q_N(_4496_),
    .Q(\i_dm_csrs.progbuf_o_114_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_115__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net708),
    .D(_0199_),
    .Q_N(_4495_),
    .Q(\i_dm_csrs.progbuf_o_115_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_116__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net666),
    .D(_0200_),
    .Q_N(_4494_),
    .Q(\i_dm_csrs.progbuf_o_116_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_117__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net665),
    .D(_0201_),
    .Q_N(_4493_),
    .Q(\i_dm_csrs.progbuf_o_117_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_118__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net731),
    .D(_0202_),
    .Q_N(_4492_),
    .Q(\i_dm_csrs.progbuf_o_118_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_119__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net727),
    .D(_0203_),
    .Q_N(_4491_),
    .Q(\i_dm_csrs.progbuf_o_119_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_11__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net675),
    .D(_0204_),
    .Q_N(_4490_),
    .Q(\i_dm_csrs.progbuf_o_11_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_120__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net675),
    .D(_0205_),
    .Q_N(_4489_),
    .Q(\i_dm_csrs.progbuf_o_120_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_121__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net697),
    .D(_0206_),
    .Q_N(_4488_),
    .Q(\i_dm_csrs.progbuf_o_121_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_122__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net663),
    .D(_0207_),
    .Q_N(_4487_),
    .Q(\i_dm_csrs.progbuf_o_122_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_123__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net704),
    .D(_0208_),
    .Q_N(_4486_),
    .Q(\i_dm_csrs.progbuf_o_123_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_124__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net699),
    .D(_0209_),
    .Q_N(_4485_),
    .Q(\i_dm_csrs.progbuf_o_124_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_125__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net663),
    .D(_0210_),
    .Q_N(_4484_),
    .Q(\i_dm_csrs.progbuf_o_125_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_126__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net669),
    .D(_0211_),
    .Q_N(_4483_),
    .Q(\i_dm_csrs.progbuf_o_126_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_127__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0212_),
    .Q_N(_4482_),
    .Q(\i_dm_csrs.progbuf_o_127_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_128__reg  (.CLK(clknet_leaf_16_clk_i),
    .RESET_B(net693),
    .D(_0213_),
    .Q_N(_4481_),
    .Q(\i_dm_csrs.progbuf_o_128_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_129__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0214_),
    .Q_N(_4480_),
    .Q(\i_dm_csrs.progbuf_o_129_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_12__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net674),
    .D(_0215_),
    .Q_N(_4479_),
    .Q(\i_dm_csrs.progbuf_o_12_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_130__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net681),
    .D(_0216_),
    .Q_N(_4478_),
    .Q(\i_dm_csrs.progbuf_o_130_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_131__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net687),
    .D(_0217_),
    .Q_N(_4477_),
    .Q(\i_dm_csrs.progbuf_o_131_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_132__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net667),
    .D(_0218_),
    .Q_N(_4476_),
    .Q(\i_dm_csrs.progbuf_o_132_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_133__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net698),
    .D(_0219_),
    .Q_N(_4475_),
    .Q(\i_dm_csrs.progbuf_o_133_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_134__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net683),
    .D(_0220_),
    .Q_N(_4474_),
    .Q(\i_dm_csrs.progbuf_o_134_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_135__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net681),
    .D(_0221_),
    .Q_N(_4473_),
    .Q(\i_dm_csrs.progbuf_o_135_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_136__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net687),
    .D(_0222_),
    .Q_N(_4472_),
    .Q(\i_dm_csrs.progbuf_o_136_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_137__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net716),
    .D(_0223_),
    .Q_N(_4471_),
    .Q(\i_dm_csrs.progbuf_o_137_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_138__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net705),
    .D(_0224_),
    .Q_N(_4470_),
    .Q(\i_dm_csrs.progbuf_o_138_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_139__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net675),
    .D(_0225_),
    .Q_N(_4469_),
    .Q(\i_dm_csrs.progbuf_o_139_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_13__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0226_),
    .Q_N(_4468_),
    .Q(\i_dm_csrs.progbuf_o_13_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_140__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net674),
    .D(_0227_),
    .Q_N(_4467_),
    .Q(\i_dm_csrs.progbuf_o_140_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_141__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0228_),
    .Q_N(_4466_),
    .Q(\i_dm_csrs.progbuf_o_141_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_142__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net685),
    .D(_0229_),
    .Q_N(_4465_),
    .Q(\i_dm_csrs.progbuf_o_142_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_143__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net667),
    .D(_0230_),
    .Q_N(_4464_),
    .Q(\i_dm_csrs.progbuf_o_143_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_144__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net704),
    .D(_0231_),
    .Q_N(_4463_),
    .Q(\i_dm_csrs.progbuf_o_144_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_145__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0232_),
    .Q_N(_4462_),
    .Q(\i_dm_csrs.progbuf_o_145_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_146__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net700),
    .D(_0233_),
    .Q_N(_4461_),
    .Q(\i_dm_csrs.progbuf_o_146_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_147__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net708),
    .D(_0234_),
    .Q_N(_4460_),
    .Q(\i_dm_csrs.progbuf_o_147_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_148__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net666),
    .D(_0235_),
    .Q_N(_4459_),
    .Q(\i_dm_csrs.progbuf_o_148_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_149__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net665),
    .D(_0236_),
    .Q_N(_4458_),
    .Q(\i_dm_csrs.progbuf_o_149_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_14__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net682),
    .D(_0237_),
    .Q_N(_4457_),
    .Q(\i_dm_csrs.progbuf_o_14_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_150__reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net692),
    .D(_0238_),
    .Q_N(_4456_),
    .Q(\i_dm_csrs.progbuf_o_150_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_151__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net687),
    .D(_0239_),
    .Q_N(_4455_),
    .Q(\i_dm_csrs.progbuf_o_151_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_152__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0240_),
    .Q_N(_4454_),
    .Q(\i_dm_csrs.progbuf_o_152_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_153__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net699),
    .D(_0241_),
    .Q_N(_4453_),
    .Q(\i_dm_csrs.progbuf_o_153_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_154__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net663),
    .D(_0242_),
    .Q_N(_4452_),
    .Q(\i_dm_csrs.progbuf_o_154_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_155__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net698),
    .D(_0243_),
    .Q_N(_4451_),
    .Q(\i_dm_csrs.progbuf_o_155_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_156__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net699),
    .D(_0244_),
    .Q_N(_4450_),
    .Q(\i_dm_csrs.progbuf_o_156_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_157__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0245_),
    .Q_N(_4449_),
    .Q(\i_dm_csrs.progbuf_o_157_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_158__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net669),
    .D(_0246_),
    .Q_N(_4448_),
    .Q(\i_dm_csrs.progbuf_o_158_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_159__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0247_),
    .Q_N(_4447_),
    .Q(\i_dm_csrs.progbuf_o_159_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_15__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net668),
    .D(_0248_),
    .Q_N(_4446_),
    .Q(\i_dm_csrs.progbuf_o_15_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_160__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net731),
    .D(_0249_),
    .Q_N(_4445_),
    .Q(\i_dm_csrs.progbuf_o_160_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_161__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0250_),
    .Q_N(_4444_),
    .Q(\i_dm_csrs.progbuf_o_161_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_162__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net682),
    .D(_0251_),
    .Q_N(_4443_),
    .Q(\i_dm_csrs.progbuf_o_162_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_163__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net687),
    .D(_0252_),
    .Q_N(_4442_),
    .Q(\i_dm_csrs.progbuf_o_163_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_164__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net681),
    .D(_0253_),
    .Q_N(_4441_),
    .Q(\i_dm_csrs.progbuf_o_164_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_165__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net698),
    .D(_0254_),
    .Q_N(_4440_),
    .Q(\i_dm_csrs.progbuf_o_165_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_166__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net683),
    .D(_0255_),
    .Q_N(_4439_),
    .Q(\i_dm_csrs.progbuf_o_166_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_167__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net682),
    .D(_0256_),
    .Q_N(_4438_),
    .Q(\i_dm_csrs.progbuf_o_167_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_168__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0257_),
    .Q_N(_4437_),
    .Q(\i_dm_csrs.progbuf_o_168_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_169__reg  (.CLK(clknet_leaf_32_clk_i),
    .RESET_B(net719),
    .D(_0258_),
    .Q_N(_4436_),
    .Q(\i_dm_csrs.progbuf_o_169_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_16__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net704),
    .D(_0259_),
    .Q_N(_4435_),
    .Q(\i_dm_csrs.progbuf_o_16_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_170__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net714),
    .D(_0260_),
    .Q_N(_4434_),
    .Q(\i_dm_csrs.progbuf_o_170_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_171__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net675),
    .D(_0261_),
    .Q_N(_4433_),
    .Q(\i_dm_csrs.progbuf_o_171_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_172__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net674),
    .D(_0262_),
    .Q_N(_4432_),
    .Q(\i_dm_csrs.progbuf_o_172_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_173__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0263_),
    .Q_N(_4431_),
    .Q(\i_dm_csrs.progbuf_o_173_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_174__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net685),
    .D(_0264_),
    .Q_N(_4430_),
    .Q(\i_dm_csrs.progbuf_o_174_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_175__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net681),
    .D(_0265_),
    .Q_N(_4429_),
    .Q(\i_dm_csrs.progbuf_o_175_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_176__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net704),
    .D(_0266_),
    .Q_N(_4428_),
    .Q(\i_dm_csrs.progbuf_o_176_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_177__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net712),
    .D(_0267_),
    .Q_N(_4427_),
    .Q(\i_dm_csrs.progbuf_o_177_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_178__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0268_),
    .Q_N(_4426_),
    .Q(\i_dm_csrs.progbuf_o_178_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_179__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net710),
    .D(_0269_),
    .Q_N(_4425_),
    .Q(\i_dm_csrs.progbuf_o_179_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_17__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0270_),
    .Q_N(_4424_),
    .Q(\i_dm_csrs.progbuf_o_17_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_180__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net666),
    .D(_0271_),
    .Q_N(_4423_),
    .Q(\i_dm_csrs.progbuf_o_180_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_181__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net665),
    .D(_0272_),
    .Q_N(_4422_),
    .Q(\i_dm_csrs.progbuf_o_181_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_182__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net727),
    .D(_0273_),
    .Q_N(_4421_),
    .Q(\i_dm_csrs.progbuf_o_182_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_183__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0274_),
    .Q_N(_4420_),
    .Q(\i_dm_csrs.progbuf_o_183_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_184__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0275_),
    .Q_N(_4419_),
    .Q(\i_dm_csrs.progbuf_o_184_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_185__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net697),
    .D(_0276_),
    .Q_N(_4418_),
    .Q(\i_dm_csrs.progbuf_o_185_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_186__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net663),
    .D(_0277_),
    .Q_N(_4417_),
    .Q(\i_dm_csrs.progbuf_o_186_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_187__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net698),
    .D(_0278_),
    .Q_N(_4416_),
    .Q(\i_dm_csrs.progbuf_o_187_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_188__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net707),
    .D(_0279_),
    .Q_N(_4415_),
    .Q(\i_dm_csrs.progbuf_o_188_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_189__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net663),
    .D(_0280_),
    .Q_N(_4414_),
    .Q(\i_dm_csrs.progbuf_o_189_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_18__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net700),
    .D(_0281_),
    .Q_N(_4413_),
    .Q(\i_dm_csrs.progbuf_o_18_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_190__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net669),
    .D(_0282_),
    .Q_N(_4412_),
    .Q(\i_dm_csrs.progbuf_o_190_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_191__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net686),
    .D(_0283_),
    .Q_N(_4411_),
    .Q(\i_dm_csrs.progbuf_o_191_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_192__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net694),
    .D(_0284_),
    .Q_N(_4410_),
    .Q(\i_dm_csrs.progbuf_o_192_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_193__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0285_),
    .Q_N(_4409_),
    .Q(\i_dm_csrs.progbuf_o_193_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_194__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net681),
    .D(_0286_),
    .Q_N(_4408_),
    .Q(\i_dm_csrs.progbuf_o_194_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_195__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net687),
    .D(_0287_),
    .Q_N(_4407_),
    .Q(\i_dm_csrs.progbuf_o_195_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_196__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net668),
    .D(_0288_),
    .Q_N(_4406_),
    .Q(\i_dm_csrs.progbuf_o_196_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_197__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net698),
    .D(_0289_),
    .Q_N(_4405_),
    .Q(\i_dm_csrs.progbuf_o_197_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_198__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net683),
    .D(_0290_),
    .Q_N(_4404_),
    .Q(\i_dm_csrs.progbuf_o_198_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_199__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net683),
    .D(_0291_),
    .Q_N(_4403_),
    .Q(\i_dm_csrs.progbuf_o_199_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_19__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net708),
    .D(_0292_),
    .Q_N(_4402_),
    .Q(\i_dm_csrs.progbuf_o_19_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_1__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0293_),
    .Q_N(_4401_),
    .Q(\i_dm_csrs.progbuf_o_1_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_200__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net688),
    .D(_0294_),
    .Q_N(_4400_),
    .Q(\i_dm_csrs.progbuf_o_200_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_201__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net719),
    .D(_0295_),
    .Q_N(_4399_),
    .Q(\i_dm_csrs.progbuf_o_201_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_202__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net705),
    .D(_0296_),
    .Q_N(_4398_),
    .Q(\i_dm_csrs.progbuf_o_202_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_203__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net676),
    .D(_0297_),
    .Q_N(_4397_),
    .Q(\i_dm_csrs.progbuf_o_203_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_204__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net674),
    .D(_0298_),
    .Q_N(_4396_),
    .Q(\i_dm_csrs.progbuf_o_204_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_205__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0299_),
    .Q_N(_4395_),
    .Q(\i_dm_csrs.progbuf_o_205_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_206__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net685),
    .D(_0300_),
    .Q_N(_4394_),
    .Q(\i_dm_csrs.progbuf_o_206_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_207__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net668),
    .D(_0301_),
    .Q_N(_4393_),
    .Q(\i_dm_csrs.progbuf_o_207_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_208__reg  (.CLK(clknet_leaf_25_clk_i),
    .RESET_B(net704),
    .D(_0302_),
    .Q_N(_4392_),
    .Q(\i_dm_csrs.progbuf_o_208_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_209__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net712),
    .D(_0303_),
    .Q_N(_4391_),
    .Q(\i_dm_csrs.progbuf_o_209_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_20__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net666),
    .D(_0304_),
    .Q_N(_4390_),
    .Q(\i_dm_csrs.progbuf_o_20_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_210__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0305_),
    .Q_N(_4389_),
    .Q(\i_dm_csrs.progbuf_o_210_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_211__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net710),
    .D(_0306_),
    .Q_N(_4388_),
    .Q(\i_dm_csrs.progbuf_o_211_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_212__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net666),
    .D(_0307_),
    .Q_N(_4387_),
    .Q(\i_dm_csrs.progbuf_o_212_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_213__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net665),
    .D(_0308_),
    .Q_N(_4386_),
    .Q(\i_dm_csrs.progbuf_o_213_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_214__reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net694),
    .D(_0309_),
    .Q_N(_4385_),
    .Q(\i_dm_csrs.progbuf_o_214_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_215__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net688),
    .D(_0310_),
    .Q_N(_4384_),
    .Q(\i_dm_csrs.progbuf_o_215_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_216__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0311_),
    .Q_N(_4383_),
    .Q(\i_dm_csrs.progbuf_o_216_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_217__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net697),
    .D(_0312_),
    .Q_N(_4382_),
    .Q(\i_dm_csrs.progbuf_o_217_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_218__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net663),
    .D(_0313_),
    .Q_N(_4381_),
    .Q(\i_dm_csrs.progbuf_o_218_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_219__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net698),
    .D(_0314_),
    .Q_N(_4380_),
    .Q(\i_dm_csrs.progbuf_o_219_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_21__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net665),
    .D(_0315_),
    .Q_N(_4379_),
    .Q(\i_dm_csrs.progbuf_o_21_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_220__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net699),
    .D(_0316_),
    .Q_N(_4378_),
    .Q(\i_dm_csrs.progbuf_o_220_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_221__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net663),
    .D(_0317_),
    .Q_N(_4377_),
    .Q(\i_dm_csrs.progbuf_o_221_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_222__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net669),
    .D(_0318_),
    .Q_N(_4376_),
    .Q(\i_dm_csrs.progbuf_o_222_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_223__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net686),
    .D(_0319_),
    .Q_N(_4375_),
    .Q(\i_dm_csrs.progbuf_o_223_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_224__reg  (.CLK(clknet_leaf_39_clk_i),
    .RESET_B(net735),
    .D(_0320_),
    .Q_N(_4374_),
    .Q(\i_dm_csrs.progbuf_o_224_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_225__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0321_),
    .Q_N(_4373_),
    .Q(\i_dm_csrs.progbuf_o_225_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_226__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net682),
    .D(_0322_),
    .Q_N(_4372_),
    .Q(\i_dm_csrs.progbuf_o_226_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_227__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net687),
    .D(_0323_),
    .Q_N(_4371_),
    .Q(\i_dm_csrs.progbuf_o_227_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_228__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net682),
    .D(_0324_),
    .Q_N(_4370_),
    .Q(\i_dm_csrs.progbuf_o_228_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_229__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net702),
    .D(_0325_),
    .Q_N(_4369_),
    .Q(\i_dm_csrs.progbuf_o_229_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_22__reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net694),
    .D(_0326_),
    .Q_N(_4368_),
    .Q(\i_dm_csrs.progbuf_o_22_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_230__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net683),
    .D(_0327_),
    .Q_N(_4367_),
    .Q(\i_dm_csrs.progbuf_o_230_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_231__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net684),
    .D(_0328_),
    .Q_N(_4366_),
    .Q(\i_dm_csrs.progbuf_o_231_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_232__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0329_),
    .Q_N(_4365_),
    .Q(\i_dm_csrs.progbuf_o_232_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_233__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net719),
    .D(_0330_),
    .Q_N(_4364_),
    .Q(\i_dm_csrs.progbuf_o_233_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_234__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net716),
    .D(_0331_),
    .Q_N(_4363_),
    .Q(\i_dm_csrs.progbuf_o_234_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_235__reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net676),
    .D(_0332_),
    .Q_N(_4362_),
    .Q(\i_dm_csrs.progbuf_o_235_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_236__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net674),
    .D(_0333_),
    .Q_N(_4361_),
    .Q(\i_dm_csrs.progbuf_o_236_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_237__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0334_),
    .Q_N(_4360_),
    .Q(\i_dm_csrs.progbuf_o_237_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_238__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net685),
    .D(_0335_),
    .Q_N(_4359_),
    .Q(\i_dm_csrs.progbuf_o_238_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_239__reg  (.CLK(clknet_leaf_102_clk_i),
    .RESET_B(net681),
    .D(_0336_),
    .Q_N(_4358_),
    .Q(\i_dm_csrs.progbuf_o_239_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_23__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net688),
    .D(_0337_),
    .Q_N(_4357_),
    .Q(\i_dm_csrs.progbuf_o_23_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_240__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net704),
    .D(_0338_),
    .Q_N(_4356_),
    .Q(\i_dm_csrs.progbuf_o_240_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_241__reg  (.CLK(clknet_leaf_29_clk_i),
    .RESET_B(net712),
    .D(_0339_),
    .Q_N(_4355_),
    .Q(\i_dm_csrs.progbuf_o_241_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_242__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net705),
    .D(_0340_),
    .Q_N(_4354_),
    .Q(\i_dm_csrs.progbuf_o_242_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_243__reg  (.CLK(clknet_leaf_31_clk_i),
    .RESET_B(net710),
    .D(_0341_),
    .Q_N(_4353_),
    .Q(\i_dm_csrs.progbuf_o_243_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_244__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net666),
    .D(_0342_),
    .Q_N(_4352_),
    .Q(\i_dm_csrs.progbuf_o_244_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_245__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net669),
    .D(_0343_),
    .Q_N(_4351_),
    .Q(\i_dm_csrs.progbuf_o_245_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_246__reg  (.CLK(clknet_leaf_87_clk_i),
    .RESET_B(net731),
    .D(_0344_),
    .Q_N(_4350_),
    .Q(\i_dm_csrs.progbuf_o_246_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_247__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0345_),
    .Q_N(_4349_),
    .Q(\i_dm_csrs.progbuf_o_247_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_248__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0346_),
    .Q_N(_4348_),
    .Q(\i_dm_csrs.progbuf_o_248_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_249__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net697),
    .D(_0347_),
    .Q_N(_4347_),
    .Q(\i_dm_csrs.progbuf_o_249_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_24__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net675),
    .D(_0348_),
    .Q_N(_4346_),
    .Q(\i_dm_csrs.progbuf_o_24_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_250__reg  (.CLK(clknet_leaf_0_clk_i),
    .RESET_B(net663),
    .D(_0349_),
    .Q_N(_4345_),
    .Q(\i_dm_csrs.progbuf_o_250_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_251__reg  (.CLK(clknet_leaf_20_clk_i),
    .RESET_B(net702),
    .D(_0350_),
    .Q_N(_4344_),
    .Q(\i_dm_csrs.progbuf_o_251_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_252__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net699),
    .D(_0351_),
    .Q_N(_4343_),
    .Q(\i_dm_csrs.progbuf_o_252_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_253__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net664),
    .D(_0352_),
    .Q_N(_4342_),
    .Q(\i_dm_csrs.progbuf_o_253_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_254__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net670),
    .D(_0353_),
    .Q_N(_4341_),
    .Q(\i_dm_csrs.progbuf_o_254_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_255__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0354_),
    .Q_N(_4340_),
    .Q(\i_dm_csrs.progbuf_o_255_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_25__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net697),
    .D(_0355_),
    .Q_N(_4339_),
    .Q(\i_dm_csrs.progbuf_o_25_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_26__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net664),
    .D(_0356_),
    .Q_N(_4338_),
    .Q(\i_dm_csrs.progbuf_o_26_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_27__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net700),
    .D(_0357_),
    .Q_N(_4337_),
    .Q(\i_dm_csrs.progbuf_o_27_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_28__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net699),
    .D(_0358_),
    .Q_N(_4336_),
    .Q(\i_dm_csrs.progbuf_o_28_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_29__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net673),
    .D(_0359_),
    .Q_N(_4335_),
    .Q(\i_dm_csrs.progbuf_o_29_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_2__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net681),
    .D(_0360_),
    .Q_N(_4334_),
    .Q(\i_dm_csrs.progbuf_o_2_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_30__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net669),
    .D(_0361_),
    .Q_N(_4333_),
    .Q(\i_dm_csrs.progbuf_o_30_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_31__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0362_),
    .Q_N(_4332_),
    .Q(\i_dm_csrs.progbuf_o_31_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_32__reg  (.CLK(clknet_4_6_0_clk_i),
    .RESET_B(net715),
    .D(_0363_),
    .Q_N(_4331_),
    .Q(\i_dm_csrs.progbuf_o_32_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_33__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0364_),
    .Q_N(_4330_),
    .Q(\i_dm_csrs.progbuf_o_33_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_34__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net684),
    .D(_0365_),
    .Q_N(_4329_),
    .Q(\i_dm_csrs.progbuf_o_34_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_35__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net687),
    .D(_0366_),
    .Q_N(_4328_),
    .Q(\i_dm_csrs.progbuf_o_35_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_36__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net670),
    .D(_0367_),
    .Q_N(_4327_),
    .Q(\i_dm_csrs.progbuf_o_36_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_37__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net697),
    .D(_0368_),
    .Q_N(_4326_),
    .Q(\i_dm_csrs.progbuf_o_37_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_38__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net690),
    .D(_0369_),
    .Q_N(_4325_),
    .Q(\i_dm_csrs.progbuf_o_38_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_39__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net683),
    .D(_0370_),
    .Q_N(_4324_),
    .Q(\i_dm_csrs.progbuf_o_39_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_3__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net687),
    .D(_0371_),
    .Q_N(_4323_),
    .Q(\i_dm_csrs.progbuf_o_3_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_40__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net727),
    .D(_0372_),
    .Q_N(_4322_),
    .Q(\i_dm_csrs.progbuf_o_40_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_41__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net717),
    .D(_0373_),
    .Q_N(_4321_),
    .Q(\i_dm_csrs.progbuf_o_41_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_42__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net708),
    .D(_0374_),
    .Q_N(_4320_),
    .Q(\i_dm_csrs.progbuf_o_42_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_43__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net676),
    .D(_0375_),
    .Q_N(_4319_),
    .Q(\i_dm_csrs.progbuf_o_43_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_44__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net676),
    .D(_0376_),
    .Q_N(_4318_),
    .Q(\i_dm_csrs.progbuf_o_44_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_45__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net669),
    .D(_0377_),
    .Q_N(_4317_),
    .Q(\i_dm_csrs.progbuf_o_45_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_46__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net685),
    .D(_0378_),
    .Q_N(_4316_),
    .Q(\i_dm_csrs.progbuf_o_46_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_47__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net668),
    .D(_0379_),
    .Q_N(_4315_),
    .Q(\i_dm_csrs.progbuf_o_47_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_48__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net708),
    .D(_0380_),
    .Q_N(_4314_),
    .Q(\i_dm_csrs.progbuf_o_48_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_49__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0381_),
    .Q_N(_4313_),
    .Q(\i_dm_csrs.progbuf_o_49_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_4__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net670),
    .D(_0382_),
    .Q_N(_4312_),
    .Q(\i_dm_csrs.progbuf_o_4_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_50__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net700),
    .D(_0383_),
    .Q_N(_4311_),
    .Q(\i_dm_csrs.progbuf_o_50_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_51__reg  (.CLK(clknet_leaf_27_clk_i),
    .RESET_B(net708),
    .D(_0384_),
    .Q_N(_4310_),
    .Q(\i_dm_csrs.progbuf_o_51_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_52__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net666),
    .D(_0385_),
    .Q_N(_4309_),
    .Q(\i_dm_csrs.progbuf_o_52_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_53__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net665),
    .D(_0386_),
    .Q_N(_4308_),
    .Q(\i_dm_csrs.progbuf_o_53_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_54__reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net731),
    .D(_0387_),
    .Q_N(_4307_),
    .Q(\i_dm_csrs.progbuf_o_54_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_55__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net730),
    .D(_0388_),
    .Q_N(_4306_),
    .Q(\i_dm_csrs.progbuf_o_55_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_56__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net675),
    .D(_0389_),
    .Q_N(_4305_),
    .Q(\i_dm_csrs.progbuf_o_56_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_57__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net697),
    .D(_0390_),
    .Q_N(_4304_),
    .Q(\i_dm_csrs.progbuf_o_57_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_58__reg  (.CLK(clknet_leaf_2_clk_i),
    .RESET_B(net664),
    .D(_0391_),
    .Q_N(_4303_),
    .Q(\i_dm_csrs.progbuf_o_58_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_59__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net700),
    .D(_0392_),
    .Q_N(_4302_),
    .Q(\i_dm_csrs.progbuf_o_59_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_5__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net676),
    .D(_0393_),
    .Q_N(_4301_),
    .Q(\i_dm_csrs.progbuf_o_5_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_60__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net699),
    .D(_0394_),
    .Q_N(_4300_),
    .Q(\i_dm_csrs.progbuf_o_60_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_61__reg  (.CLK(clknet_leaf_8_clk_i),
    .RESET_B(net673),
    .D(_0395_),
    .Q_N(_4299_),
    .Q(\i_dm_csrs.progbuf_o_61_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_62__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net678),
    .D(_0396_),
    .Q_N(_4298_),
    .Q(\i_dm_csrs.progbuf_o_62_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_63__reg  (.CLK(clknet_leaf_83_clk_i),
    .RESET_B(net728),
    .D(_0397_),
    .Q_N(_4297_),
    .Q(\i_dm_csrs.progbuf_o_63_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_64__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net694),
    .D(_0398_),
    .Q_N(_4296_),
    .Q(\i_dm_csrs.progbuf_o_64_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_65__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net685),
    .D(_0399_),
    .Q_N(_4295_),
    .Q(\i_dm_csrs.progbuf_o_65_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_66__reg  (.CLK(clknet_leaf_97_clk_i),
    .RESET_B(net682),
    .D(_0400_),
    .Q_N(_4294_),
    .Q(\i_dm_csrs.progbuf_o_66_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_67__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net692),
    .D(_0401_),
    .Q_N(_4293_),
    .Q(\i_dm_csrs.progbuf_o_67_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_68__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net670),
    .D(_0402_),
    .Q_N(_4292_),
    .Q(\i_dm_csrs.progbuf_o_68_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_69__reg  (.CLK(clknet_leaf_7_clk_i),
    .RESET_B(net676),
    .D(_0403_),
    .Q_N(_4291_),
    .Q(\i_dm_csrs.progbuf_o_69_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_6__reg  (.CLK(clknet_leaf_100_clk_i),
    .RESET_B(net670),
    .D(_0404_),
    .Q_N(_4290_),
    .Q(\i_dm_csrs.progbuf_o_6_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_70__reg  (.CLK(clknet_leaf_92_clk_i),
    .RESET_B(net670),
    .D(_0405_),
    .Q_N(_4289_),
    .Q(\i_dm_csrs.progbuf_o_70_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_71__reg  (.CLK(clknet_leaf_99_clk_i),
    .RESET_B(net684),
    .D(_0406_),
    .Q_N(_4288_),
    .Q(\i_dm_csrs.progbuf_o_71_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_72__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net688),
    .D(_0407_),
    .Q_N(_4287_),
    .Q(\i_dm_csrs.progbuf_o_72_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_73__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net716),
    .D(_0408_),
    .Q_N(_4286_),
    .Q(\i_dm_csrs.progbuf_o_73_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_74__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net708),
    .D(_0409_),
    .Q_N(_4285_),
    .Q(\i_dm_csrs.progbuf_o_74_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_75__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net676),
    .D(_0410_),
    .Q_N(_4284_),
    .Q(\i_dm_csrs.progbuf_o_75_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_76__reg  (.CLK(clknet_leaf_4_clk_i),
    .RESET_B(net677),
    .D(_0411_),
    .Q_N(_4283_),
    .Q(\i_dm_csrs.progbuf_o_76_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_77__reg  (.CLK(clknet_leaf_103_clk_i),
    .RESET_B(net667),
    .D(_0412_),
    .Q_N(_4282_),
    .Q(\i_dm_csrs.progbuf_o_77_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_78__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net685),
    .D(_0413_),
    .Q_N(_4281_),
    .Q(\i_dm_csrs.progbuf_o_78_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_79__reg  (.CLK(clknet_leaf_101_clk_i),
    .RESET_B(net668),
    .D(_0414_),
    .Q_N(_4280_),
    .Q(\i_dm_csrs.progbuf_o_79_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_7__reg  (.CLK(clknet_leaf_98_clk_i),
    .RESET_B(net683),
    .D(_0415_),
    .Q_N(_4279_),
    .Q(\i_dm_csrs.progbuf_o_7_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_80__reg  (.CLK(clknet_leaf_19_clk_i),
    .RESET_B(net704),
    .D(_0416_),
    .Q_N(_4278_),
    .Q(\i_dm_csrs.progbuf_o_80_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_81__reg  (.CLK(clknet_leaf_28_clk_i),
    .RESET_B(net707),
    .D(_0417_),
    .Q_N(_4277_),
    .Q(\i_dm_csrs.progbuf_o_81_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_82__reg  (.CLK(clknet_leaf_24_clk_i),
    .RESET_B(net700),
    .D(_0418_),
    .Q_N(_4276_),
    .Q(\i_dm_csrs.progbuf_o_82_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_83__reg  (.CLK(clknet_leaf_26_clk_i),
    .RESET_B(net708),
    .D(_0419_),
    .Q_N(_4275_),
    .Q(\i_dm_csrs.progbuf_o_83_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_84__reg  (.CLK(clknet_leaf_104_clk_i),
    .RESET_B(net666),
    .D(_0420_),
    .Q_N(_4274_),
    .Q(\i_dm_csrs.progbuf_o_84_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_85__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net672),
    .D(_0421_),
    .Q_N(_4273_),
    .Q(\i_dm_csrs.progbuf_o_85_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_86__reg  (.CLK(clknet_leaf_90_clk_i),
    .RESET_B(net694),
    .D(_0422_),
    .Q_N(_4272_),
    .Q(\i_dm_csrs.progbuf_o_86_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_87__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net688),
    .D(_0423_),
    .Q_N(_4271_),
    .Q(\i_dm_csrs.progbuf_o_87_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_88__reg  (.CLK(clknet_leaf_6_clk_i),
    .RESET_B(net675),
    .D(_0424_),
    .Q_N(_4270_),
    .Q(\i_dm_csrs.progbuf_o_88_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_89__reg  (.CLK(clknet_leaf_21_clk_i),
    .RESET_B(net697),
    .D(_0425_),
    .Q_N(_4269_),
    .Q(\i_dm_csrs.progbuf_o_89_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_8__reg  (.CLK(clknet_leaf_94_clk_i),
    .RESET_B(net688),
    .D(_0426_),
    .Q_N(_4268_),
    .Q(\i_dm_csrs.progbuf_o_8_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_90__reg  (.CLK(clknet_leaf_1_clk_i),
    .RESET_B(net664),
    .D(_0427_),
    .Q_N(_4267_),
    .Q(\i_dm_csrs.progbuf_o_90_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_91__reg  (.CLK(clknet_leaf_22_clk_i),
    .RESET_B(net700),
    .D(_0428_),
    .Q_N(_4266_),
    .Q(\i_dm_csrs.progbuf_o_91_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_92__reg  (.CLK(clknet_leaf_23_clk_i),
    .RESET_B(net699),
    .D(_0429_),
    .Q_N(_4265_),
    .Q(\i_dm_csrs.progbuf_o_92_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_93__reg  (.CLK(clknet_leaf_5_clk_i),
    .RESET_B(net673),
    .D(_0430_),
    .Q_N(_4264_),
    .Q(\i_dm_csrs.progbuf_o_93_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_94__reg  (.CLK(clknet_leaf_3_clk_i),
    .RESET_B(net678),
    .D(_0431_),
    .Q_N(_4263_),
    .Q(\i_dm_csrs.progbuf_o_94_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_95__reg  (.CLK(clknet_leaf_95_clk_i),
    .RESET_B(net686),
    .D(_0432_),
    .Q_N(_4262_),
    .Q(\i_dm_csrs.progbuf_o_95_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_96__reg  (.CLK(clknet_leaf_17_clk_i),
    .RESET_B(net726),
    .D(_0433_),
    .Q_N(_4261_),
    .Q(\i_dm_csrs.progbuf_o_96_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_97__reg  (.CLK(clknet_leaf_82_clk_i),
    .RESET_B(net728),
    .D(_0434_),
    .Q_N(_4260_),
    .Q(\i_dm_csrs.progbuf_o_97_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_98__reg  (.CLK(clknet_leaf_96_clk_i),
    .RESET_B(net684),
    .D(_0435_),
    .Q_N(_4259_),
    .Q(\i_dm_csrs.progbuf_o_98_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_99__reg  (.CLK(clknet_leaf_93_clk_i),
    .RESET_B(net684),
    .D(_0436_),
    .Q_N(_4258_),
    .Q(\i_dm_csrs.progbuf_o_99_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.progbuf_o_9__reg  (.CLK(clknet_leaf_18_clk_i),
    .RESET_B(net716),
    .D(_0437_),
    .Q_N(_4683_),
    .Q(\i_dm_csrs.progbuf_o_9_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.resumeack_i_reg  (.RESET_B(net735),
    .D(\i_dm_mem.resuming_d ),
    .Q(\i_dm_csrs.dmstatus_16_ ),
    .Q_N(_4684_),
    .CLK(clknet_leaf_88_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.resumereq_o_reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net742),
    .D(\i_dm_csrs.resumereq_o_reg_D ),
    .Q_N(\clear_resumeack_$_AND__Y_A ),
    .Q(\i_dm_csrs.resumereq_o ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaccess_o_0__reg  (.CLK(clknet_leaf_69_clk_i),
    .RESET_B(net763),
    .D(_0438_),
    .Q_N(\i_dm_sba.sbaccess_mask_3__$_AND__B_A_$_AND__Y_A ),
    .Q(\i_dm_csrs.sbaccess_o_0_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaccess_o_1__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net748),
    .D(_0439_),
    .Q_N(\i_dm_csrs.sbaccess_o_1_ ),
    .Q(_0001_));
 sg13g2_dfrbp_2 \i_dm_csrs.sbaccess_o_2__reg  (.RESET_B(net763),
    .D(_0440_),
    .Q(\i_dm_csrs.sbaccess_o_2_ ),
    .Q_N(\i_dm_sba.sbaccess_mask_3_ ),
    .CLK(clknet_leaf_69_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_32__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_32__reg_D ),
    .Q_N(_4685_),
    .Q(\i_dm_csrs.sbaddr_q_32_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_33__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_33__reg_D ),
    .Q_N(_4686_),
    .Q(\i_dm_csrs.sbaddr_q_33_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_34__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_34__reg_D ),
    .Q_N(_4687_),
    .Q(\i_dm_csrs.sbaddr_q_34_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_35__reg  (.CLK(clknet_leaf_70_clk_i),
    .RESET_B(net747),
    .D(\i_dm_csrs.sbaddr_q_35__reg_D ),
    .Q_N(_4688_),
    .Q(\i_dm_csrs.sbaddr_q_35_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_36__reg  (.CLK(clknet_leaf_72_clk_i),
    .RESET_B(net747),
    .D(\i_dm_csrs.sbaddr_q_36__reg_D ),
    .Q_N(_4689_),
    .Q(\i_dm_csrs.sbaddr_q_36_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_37__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net746),
    .D(\i_dm_csrs.sbaddr_q_37__reg_D ),
    .Q_N(_4690_),
    .Q(\i_dm_csrs.sbaddr_q_37_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_38__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net746),
    .D(\i_dm_csrs.sbaddr_q_38__reg_D ),
    .Q_N(_4691_),
    .Q(\i_dm_csrs.sbaddr_q_38_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_39__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net742),
    .D(\i_dm_csrs.sbaddr_q_39__reg_D ),
    .Q_N(_4692_),
    .Q(\i_dm_csrs.sbaddr_q_39_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_40__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_40__reg_D ),
    .Q_N(_4693_),
    .Q(\i_dm_csrs.sbaddr_q_40_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_41__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_41__reg_D ),
    .Q_N(_4694_),
    .Q(\i_dm_csrs.sbaddr_q_41_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_42__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net748),
    .D(\i_dm_csrs.sbaddr_q_42__reg_D ),
    .Q_N(_4695_),
    .Q(\i_dm_csrs.sbaddr_q_42_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_43__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net747),
    .D(\i_dm_csrs.sbaddr_q_43__reg_D ),
    .Q_N(_4696_),
    .Q(\i_dm_csrs.sbaddr_q_43_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_44__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net757),
    .D(\i_dm_csrs.sbaddr_q_44__reg_D ),
    .Q_N(_4697_),
    .Q(\i_dm_csrs.sbaddr_q_44_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_45__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net752),
    .D(\i_dm_csrs.sbaddr_q_45__reg_D ),
    .Q_N(_4698_),
    .Q(\i_dm_csrs.sbaddr_q_45_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_46__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_46__reg_D ),
    .Q_N(_4699_),
    .Q(\i_dm_csrs.sbaddr_q_46_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_47__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_47__reg_D ),
    .Q_N(_4700_),
    .Q(\i_dm_csrs.sbaddr_q_47_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_48__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net752),
    .D(\i_dm_csrs.sbaddr_q_48__reg_D ),
    .Q_N(_4701_),
    .Q(\i_dm_csrs.sbaddr_q_48_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_49__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_49__reg_D ),
    .Q_N(_4702_),
    .Q(\i_dm_csrs.sbaddr_q_49_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_50__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_50__reg_D ),
    .Q_N(_4703_),
    .Q(\i_dm_csrs.sbaddr_q_50_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_51__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_51__reg_D ),
    .Q_N(_4704_),
    .Q(\i_dm_csrs.sbaddr_q_51_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_52__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net752),
    .D(\i_dm_csrs.sbaddr_q_52__reg_D ),
    .Q_N(_4705_),
    .Q(\i_dm_csrs.sbaddr_q_52_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_53__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net755),
    .D(\i_dm_csrs.sbaddr_q_53__reg_D ),
    .Q_N(_4706_),
    .Q(\i_dm_csrs.sbaddr_q_53_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_54__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net744),
    .D(\i_dm_csrs.sbaddr_q_54__reg_D ),
    .Q_N(_4707_),
    .Q(\i_dm_csrs.sbaddr_q_54_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_55__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net755),
    .D(\i_dm_csrs.sbaddr_q_55__reg_D ),
    .Q_N(_4708_),
    .Q(\i_dm_csrs.sbaddr_q_55_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_56__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(\i_dm_csrs.sbaddr_q_56__reg_D ),
    .Q_N(_4709_),
    .Q(\i_dm_csrs.sbaddr_q_56_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_57__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net754),
    .D(\i_dm_csrs.sbaddr_q_57__reg_D ),
    .Q_N(_4710_),
    .Q(\i_dm_csrs.sbaddr_q_57_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_58__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(\i_dm_csrs.sbaddr_q_58__reg_D ),
    .Q_N(_4711_),
    .Q(\i_dm_csrs.sbaddr_q_58_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_59__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net723),
    .D(\i_dm_csrs.sbaddr_q_59__reg_D ),
    .Q_N(_4712_),
    .Q(\i_dm_csrs.sbaddr_q_59_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_60__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net755),
    .D(\i_dm_csrs.sbaddr_q_60__reg_D ),
    .Q_N(_4713_),
    .Q(\i_dm_csrs.sbaddr_q_60_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_61__reg  (.CLK(clknet_leaf_45_clk_i),
    .RESET_B(net757),
    .D(\i_dm_csrs.sbaddr_q_61__reg_D ),
    .Q_N(_4714_),
    .Q(\i_dm_csrs.sbaddr_q_61_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_62__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net752),
    .D(\i_dm_csrs.sbaddr_q_62__reg_D ),
    .Q_N(_4715_),
    .Q(\i_dm_csrs.sbaddr_q_62_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbaddr_q_63__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net752),
    .D(\i_dm_csrs.sbaddr_q_63__reg_D ),
    .Q_N(_4257_),
    .Q(\i_dm_csrs.sbaddr_q_63_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.sbautoincrement_o_reg  (.RESET_B(net757),
    .D(_0441_),
    .Q(\i_dm_csrs.sbautoincrement_o ),
    .Q_N(_4256_),
    .CLK(clknet_leaf_52_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_12__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net757),
    .D(_0442_),
    .Q_N(_4255_),
    .Q(\i_dm_csrs.sbcs_q_12_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_13__reg  (.CLK(clknet_leaf_44_clk_i),
    .RESET_B(net757),
    .D(_0443_),
    .Q_N(_4254_),
    .Q(\i_dm_csrs.sbcs_q_13_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_14__reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net757),
    .D(_0444_),
    .Q_N(_4716_),
    .Q(\i_dm_csrs.sbcs_q_14_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_21__reg  (.CLK(clknet_leaf_51_clk_i),
    .RESET_B(net758),
    .D(\i_dm_csrs.sbcs_q_21__reg_D ),
    .Q_N(_4717_),
    .Q(\i_dm_csrs.sbcs_q_21_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.sbcs_q_22__reg  (.RESET_B(net722),
    .D(\i_dm_csrs.sbcs_q_22__reg_D ),
    .Q(\i_dm_csrs.sbcs_q_22_ ),
    .Q_N(_4253_),
    .CLK(clknet_leaf_37_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_23__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net758),
    .D(_0445_),
    .Q_N(_4252_),
    .Q(\i_dm_csrs.sbcs_q_23_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_24__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net756),
    .D(_0446_),
    .Q_N(_4251_),
    .Q(\i_dm_csrs.sbcs_q_24_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_25__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net756),
    .D(_0447_),
    .Q_N(_4250_),
    .Q(\i_dm_csrs.sbcs_q_25_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_26__reg  (.CLK(clknet_leaf_49_clk_i),
    .RESET_B(net756),
    .D(_0448_),
    .Q_N(_4249_),
    .Q(\i_dm_csrs.sbcs_q_26_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_27__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net756),
    .D(_0449_),
    .Q_N(_4248_),
    .Q(\i_dm_csrs.sbcs_q_27_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_28__reg  (.CLK(clknet_leaf_50_clk_i),
    .RESET_B(net758),
    .D(_0450_),
    .Q_N(_4718_),
    .Q(\i_dm_csrs.sbcs_q_28_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbcs_q_29__reg  (.CLK(clknet_leaf_43_clk_i),
    .RESET_B(net749),
    .D(net83),
    .Q_N(_4247_),
    .Q(\i_dm_csrs.sbcs_q_0_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_0__reg  (.RESET_B(net722),
    .D(_0451_),
    .Q(\i_dm_csrs.sbdata_o_0_ ),
    .Q_N(_4246_),
    .CLK(clknet_leaf_35_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_10__reg  (.RESET_B(net722),
    .D(_0452_),
    .Q(\i_dm_csrs.sbdata_o_10_ ),
    .Q_N(_4245_),
    .CLK(clknet_leaf_37_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_11__reg  (.RESET_B(net724),
    .D(_0453_),
    .Q(\i_dm_csrs.sbdata_o_11_ ),
    .Q_N(_4244_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_12__reg  (.RESET_B(net710),
    .D(_0454_),
    .Q(\i_dm_csrs.sbdata_o_12_ ),
    .Q_N(_4243_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_13__reg  (.RESET_B(net716),
    .D(_0455_),
    .Q(\i_dm_csrs.sbdata_o_13_ ),
    .Q_N(_4242_),
    .CLK(clknet_leaf_31_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_14__reg  (.RESET_B(net716),
    .D(_0456_),
    .Q(\i_dm_csrs.sbdata_o_14_ ),
    .Q_N(_4241_),
    .CLK(clknet_leaf_32_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_15__reg  (.RESET_B(net718),
    .D(_0457_),
    .Q(\i_dm_csrs.sbdata_o_15_ ),
    .Q_N(_4240_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_16__reg  (.RESET_B(net709),
    .D(_0458_),
    .Q(\i_dm_csrs.sbdata_o_16_ ),
    .Q_N(_4239_),
    .CLK(clknet_leaf_31_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_17__reg  (.RESET_B(net710),
    .D(_0459_),
    .Q(\i_dm_csrs.sbdata_o_17_ ),
    .Q_N(_4238_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_18__reg  (.RESET_B(net709),
    .D(_0460_),
    .Q(\i_dm_csrs.sbdata_o_18_ ),
    .Q_N(_4237_),
    .CLK(clknet_leaf_31_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_19__reg  (.RESET_B(net710),
    .D(_0461_),
    .Q(\i_dm_csrs.sbdata_o_19_ ),
    .Q_N(_4236_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_1__reg  (.RESET_B(net718),
    .D(_0462_),
    .Q(\i_dm_csrs.sbdata_o_1_ ),
    .Q_N(_4235_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_20__reg  (.RESET_B(net718),
    .D(_0463_),
    .Q(\i_dm_csrs.sbdata_o_20_ ),
    .Q_N(_4234_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_21__reg  (.RESET_B(net718),
    .D(_0464_),
    .Q(\i_dm_csrs.sbdata_o_21_ ),
    .Q_N(_4233_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_22__reg  (.RESET_B(net718),
    .D(_0465_),
    .Q(\i_dm_csrs.sbdata_o_22_ ),
    .Q_N(_4232_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_23__reg  (.RESET_B(net718),
    .D(_0466_),
    .Q(\i_dm_csrs.sbdata_o_23_ ),
    .Q_N(_4231_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_24__reg  (.RESET_B(net710),
    .D(_0467_),
    .Q(\i_dm_csrs.sbdata_o_24_ ),
    .Q_N(_4230_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_25__reg  (.RESET_B(net718),
    .D(_0468_),
    .Q(\i_dm_csrs.sbdata_o_25_ ),
    .Q_N(_4229_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_26__reg  (.RESET_B(net710),
    .D(_0469_),
    .Q(\i_dm_csrs.sbdata_o_26_ ),
    .Q_N(_4228_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_27__reg  (.RESET_B(net709),
    .D(_0470_),
    .Q(\i_dm_csrs.sbdata_o_27_ ),
    .Q_N(_4227_),
    .CLK(clknet_leaf_31_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_28__reg  (.RESET_B(net711),
    .D(_0471_),
    .Q(\i_dm_csrs.sbdata_o_28_ ),
    .Q_N(_4226_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_29__reg  (.RESET_B(net709),
    .D(_0472_),
    .Q(\i_dm_csrs.sbdata_o_29_ ),
    .Q_N(_4225_),
    .CLK(clknet_leaf_30_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_2__reg  (.RESET_B(net721),
    .D(_0473_),
    .Q(\i_dm_csrs.sbdata_o_2_ ),
    .Q_N(_4224_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_30__reg  (.RESET_B(net716),
    .D(_0474_),
    .Q(\i_dm_csrs.sbdata_o_30_ ),
    .Q_N(_4223_),
    .CLK(clknet_leaf_31_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_31__reg  (.RESET_B(net718),
    .D(_0475_),
    .Q(\i_dm_csrs.sbdata_o_31_ ),
    .Q_N(_4222_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_3__reg  (.RESET_B(net724),
    .D(_0476_),
    .Q(\i_dm_csrs.sbdata_o_3_ ),
    .Q_N(_4221_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_4__reg  (.RESET_B(net724),
    .D(_0477_),
    .Q(\i_dm_csrs.sbdata_o_4_ ),
    .Q_N(_4220_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_5__reg  (.RESET_B(net721),
    .D(_0478_),
    .Q(\i_dm_csrs.sbdata_o_5_ ),
    .Q_N(_4219_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_6__reg  (.RESET_B(net721),
    .D(_0479_),
    .Q(\i_dm_csrs.sbdata_o_6_ ),
    .Q_N(_4218_),
    .CLK(clknet_leaf_33_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_7__reg  (.RESET_B(net723),
    .D(_0480_),
    .Q(\i_dm_csrs.sbdata_o_7_ ),
    .Q_N(_4217_),
    .CLK(clknet_leaf_35_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_8__reg  (.RESET_B(net721),
    .D(_0481_),
    .Q(\i_dm_csrs.sbdata_o_8_ ),
    .Q_N(_4216_),
    .CLK(clknet_leaf_34_clk_i));
 sg13g2_dfrbp_2 \i_dm_csrs.sbdata_o_9__reg  (.RESET_B(net723),
    .D(_0482_),
    .Q(\i_dm_csrs.sbdata_o_9_ ),
    .Q_N(_4215_),
    .CLK(clknet_leaf_35_clk_i));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_32__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net753),
    .D(_0483_),
    .Q_N(_4214_),
    .Q(\i_dm_csrs.sbdata_q_32_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_33__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net753),
    .D(_0484_),
    .Q_N(_4213_),
    .Q(\i_dm_csrs.sbdata_q_33_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_34__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net752),
    .D(_0485_),
    .Q_N(_4212_),
    .Q(\i_dm_csrs.sbdata_q_34_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_35__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net742),
    .D(_0486_),
    .Q_N(_4211_),
    .Q(\i_dm_csrs.sbdata_q_35_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_36__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net743),
    .D(_0487_),
    .Q_N(_4210_),
    .Q(\i_dm_csrs.sbdata_q_36_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_37__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net743),
    .D(_0488_),
    .Q_N(_4209_),
    .Q(\i_dm_csrs.sbdata_q_37_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_38__reg  (.CLK(clknet_leaf_40_clk_i),
    .RESET_B(net743),
    .D(_0489_),
    .Q_N(_4208_),
    .Q(\i_dm_csrs.sbdata_q_38_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_39__reg  (.CLK(clknet_leaf_41_clk_i),
    .RESET_B(net743),
    .D(_0490_),
    .Q_N(_4207_),
    .Q(\i_dm_csrs.sbdata_q_39_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_40__reg  (.CLK(clknet_leaf_42_clk_i),
    .RESET_B(net744),
    .D(_0491_),
    .Q_N(_4206_),
    .Q(\i_dm_csrs.sbdata_q_40_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_41__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net744),
    .D(_0492_),
    .Q_N(_4205_),
    .Q(\i_dm_csrs.sbdata_q_41_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_42__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net745),
    .D(_0493_),
    .Q_N(_4204_),
    .Q(\i_dm_csrs.sbdata_q_42_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_43__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net745),
    .D(_0494_),
    .Q_N(_4203_),
    .Q(\i_dm_csrs.sbdata_q_43_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_44__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net752),
    .D(_0495_),
    .Q_N(_4202_),
    .Q(\i_dm_csrs.sbdata_q_44_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_45__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net752),
    .D(_0496_),
    .Q_N(_4201_),
    .Q(\i_dm_csrs.sbdata_q_45_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_46__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net745),
    .D(_0497_),
    .Q_N(_4200_),
    .Q(\i_dm_csrs.sbdata_q_46_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_47__reg  (.CLK(clknet_leaf_46_clk_i),
    .RESET_B(net745),
    .D(_0498_),
    .Q_N(_4199_),
    .Q(\i_dm_csrs.sbdata_q_47_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_48__reg  (.CLK(clknet_leaf_37_clk_i),
    .RESET_B(net722),
    .D(_0499_),
    .Q_N(_4198_),
    .Q(\i_dm_csrs.sbdata_q_48_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_49__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net754),
    .D(_0500_),
    .Q_N(_4197_),
    .Q(\i_dm_csrs.sbdata_q_49_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_50__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net722),
    .D(_0501_),
    .Q_N(_4196_),
    .Q(\i_dm_csrs.sbdata_q_50_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_51__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net723),
    .D(_0502_),
    .Q_N(_4195_),
    .Q(\i_dm_csrs.sbdata_q_51_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_52__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net721),
    .D(_0503_),
    .Q_N(_4194_),
    .Q(\i_dm_csrs.sbdata_q_52_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_53__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net719),
    .D(_0504_),
    .Q_N(_4193_),
    .Q(\i_dm_csrs.sbdata_q_53_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_54__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net723),
    .D(_0505_),
    .Q_N(_4192_),
    .Q(\i_dm_csrs.sbdata_q_54_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_55__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net723),
    .D(_0506_),
    .Q_N(_4191_),
    .Q(\i_dm_csrs.sbdata_q_55_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_56__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net724),
    .D(_0507_),
    .Q_N(_4190_),
    .Q(\i_dm_csrs.sbdata_q_56_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_57__reg  (.CLK(clknet_leaf_35_clk_i),
    .RESET_B(net724),
    .D(_0508_),
    .Q_N(_4189_),
    .Q(\i_dm_csrs.sbdata_q_57_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_58__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net723),
    .D(_0509_),
    .Q_N(_4188_),
    .Q(\i_dm_csrs.sbdata_q_58_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_59__reg  (.CLK(clknet_leaf_36_clk_i),
    .RESET_B(net724),
    .D(_0510_),
    .Q_N(_4187_),
    .Q(\i_dm_csrs.sbdata_q_59_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_60__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net755),
    .D(_0511_),
    .Q_N(_4186_),
    .Q(\i_dm_csrs.sbdata_q_60_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_61__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net753),
    .D(_0512_),
    .Q_N(_4185_),
    .Q(\i_dm_csrs.sbdata_q_61_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_62__reg  (.CLK(clknet_leaf_47_clk_i),
    .RESET_B(net753),
    .D(_0513_),
    .Q_N(_4184_),
    .Q(\i_dm_csrs.sbdata_q_62_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbdata_q_63__reg  (.CLK(clknet_leaf_48_clk_i),
    .RESET_B(net754),
    .D(_0514_),
    .Q_N(_4183_),
    .Q(\i_dm_csrs.sbdata_q_63_ ));
 sg13g2_dfrbp_1 \i_dm_csrs.sbreadonaddr_o_reg  (.CLK(clknet_leaf_52_clk_i),
    .RESET_B(net757),
    .D(_0515_),
    .Q_N(_4182_),
    .Q(\i_dm_csrs.sbcs_q_20_ ));
 sg13g2_dfrbp_2 \i_dm_csrs.sbreadondata_o_reg  (.RESET_B(net749),
    .D(_0516_),
    .Q(\i_dm_csrs.sbcs_q_15_ ),
    .Q_N(_4719_),
    .CLK(clknet_leaf_44_clk_i));
 sg13g2_dfrbp_1 \i_dm_mem.fwd_rom_q_reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net761),
    .D(slave_addr_i_11_),
    .Q_N(_4181_),
    .Q(\i_dm_mem.fwd_rom_q ));
 sg13g2_dfrbp_1 \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_0__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net739),
    .D(_0517_),
    .Q_N(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_42__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ),
    .Q(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_0_ ));
 sg13g2_dfrbp_2 \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_1__reg  (.RESET_B(net740),
    .D(_0518_),
    .Q(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_1_ ),
    .Q_N(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_20__$_MUX__Y_A_$_MUX__Y_B ),
    .CLK(clknet_leaf_81_clk_i));
 sg13g2_dfrbp_1 \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net740),
    .D(_0519_),
    .Q_N(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_2__$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ),
    .Q(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_2_ ));
 sg13g2_dfrbp_1 \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__reg  (.CLK(clknet_leaf_81_clk_i),
    .RESET_B(net740),
    .D(_0520_),
    .Q_N(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3__$_NOT__A_Y ),
    .Q(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_3_ ));
 sg13g2_dfrbp_1 \i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net741),
    .D(_0521_),
    .Q_N(_4180_),
    .Q(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_4_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_0__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net732),
    .D(_0522_),
    .Q_N(_4179_),
    .Q(\i_dm_mem.rdata_q_0_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_10__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net734),
    .D(_0523_),
    .Q_N(_4178_),
    .Q(\i_dm_mem.rdata_q_10_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_11__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net732),
    .D(_0524_),
    .Q_N(_4177_),
    .Q(\i_dm_mem.rdata_q_11_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_12__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net734),
    .D(_0525_),
    .Q_N(_4176_),
    .Q(\i_dm_mem.rdata_q_12_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_13__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net729),
    .D(_0526_),
    .Q_N(_4175_),
    .Q(\i_dm_mem.rdata_q_13_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_14__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net738),
    .D(_0527_),
    .Q_N(_4174_),
    .Q(\i_dm_mem.rdata_q_14_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_15__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net762),
    .D(_0528_),
    .Q_N(_4173_),
    .Q(\i_dm_mem.rdata_q_15_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_16__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net736),
    .D(_0529_),
    .Q_N(_4172_),
    .Q(\i_dm_mem.rdata_q_16_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_17__reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net762),
    .D(_0530_),
    .Q_N(_4171_),
    .Q(\i_dm_mem.rdata_q_17_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_18__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net732),
    .D(_0531_),
    .Q_N(_4170_),
    .Q(\i_dm_mem.rdata_q_18_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_19__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net762),
    .D(_0532_),
    .Q_N(_4169_),
    .Q(\i_dm_mem.rdata_q_19_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_1__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net732),
    .D(_0533_),
    .Q_N(_4168_),
    .Q(\i_dm_mem.rdata_q_1_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_20__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net732),
    .D(_0534_),
    .Q_N(_4167_),
    .Q(\i_dm_mem.rdata_q_20_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_21__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net736),
    .D(_0535_),
    .Q_N(_4166_),
    .Q(\i_dm_mem.rdata_q_21_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_22__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net736),
    .D(_0536_),
    .Q_N(_4165_),
    .Q(\i_dm_mem.rdata_q_22_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_23__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net734),
    .D(_0537_),
    .Q_N(_4164_),
    .Q(\i_dm_mem.rdata_q_23_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_24__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net734),
    .D(_0538_),
    .Q_N(_4163_),
    .Q(\i_dm_mem.rdata_q_24_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_25__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0539_),
    .Q_N(_4162_),
    .Q(\i_dm_mem.rdata_q_25_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_26__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net729),
    .D(_0540_),
    .Q_N(_4161_),
    .Q(\i_dm_mem.rdata_q_26_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_27__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net737),
    .D(_0541_),
    .Q_N(_4160_),
    .Q(\i_dm_mem.rdata_q_27_ ));
 sg13g2_dfrbp_2 \i_dm_mem.rdata_q_28__reg  (.RESET_B(net730),
    .D(_0542_),
    .Q(\i_dm_mem.rdata_q_28_ ),
    .Q_N(_4159_),
    .CLK(clknet_leaf_84_clk_i));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_29__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net737),
    .D(_0543_),
    .Q_N(_4158_),
    .Q(\i_dm_mem.rdata_q_29_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_2__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0544_),
    .Q_N(_4157_),
    .Q(\i_dm_mem.rdata_q_2_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_30__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net730),
    .D(_0545_),
    .Q_N(_4156_),
    .Q(\i_dm_mem.rdata_q_30_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_31__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0546_),
    .Q_N(_4155_),
    .Q(\i_dm_mem.rdata_q_31_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_32__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net738),
    .D(_0547_),
    .Q_N(_4154_),
    .Q(\i_dm_mem.rdata_q_32_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_33__reg  (.CLK(clknet_4_11_0_clk_i),
    .RESET_B(net738),
    .D(_0548_),
    .Q_N(_4153_),
    .Q(\i_dm_mem.rdata_q_33_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_34__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net734),
    .D(_0549_),
    .Q_N(_4152_),
    .Q(\i_dm_mem.rdata_q_34_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_35__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net740),
    .D(_0550_),
    .Q_N(_4151_),
    .Q(\i_dm_mem.rdata_q_35_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_36__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0551_),
    .Q_N(_4150_),
    .Q(\i_dm_mem.rdata_q_36_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_37__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net737),
    .D(_0552_),
    .Q_N(_4149_),
    .Q(\i_dm_mem.rdata_q_37_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_38__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net737),
    .D(_0553_),
    .Q_N(_4148_),
    .Q(\i_dm_mem.rdata_q_38_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_39__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net740),
    .D(_0554_),
    .Q_N(_4147_),
    .Q(\i_dm_mem.rdata_q_39_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_3__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net740),
    .D(_0555_),
    .Q_N(_4146_),
    .Q(\i_dm_mem.rdata_q_3_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_40__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net734),
    .D(_0556_),
    .Q_N(_4145_),
    .Q(\i_dm_mem.rdata_q_40_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_41__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net761),
    .D(_0557_),
    .Q_N(_4144_),
    .Q(\i_dm_mem.rdata_q_41_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_42__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net737),
    .D(_0558_),
    .Q_N(_4143_),
    .Q(\i_dm_mem.rdata_q_42_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_43__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net761),
    .D(_0559_),
    .Q_N(_4142_),
    .Q(\i_dm_mem.rdata_q_43_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_44__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net736),
    .D(_0560_),
    .Q_N(_4141_),
    .Q(\i_dm_mem.rdata_q_44_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_45__reg  (.CLK(clknet_leaf_86_clk_i),
    .RESET_B(net734),
    .D(_0561_),
    .Q_N(_4140_),
    .Q(\i_dm_mem.rdata_q_45_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_46__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net738),
    .D(_0562_),
    .Q_N(_4139_),
    .Q(\i_dm_mem.rdata_q_46_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_47__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net762),
    .D(_0563_),
    .Q_N(_4138_),
    .Q(\i_dm_mem.rdata_q_47_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_48__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net737),
    .D(_0564_),
    .Q_N(_4137_),
    .Q(\i_dm_mem.rdata_q_48_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_49__reg  (.CLK(clknet_leaf_67_clk_i),
    .RESET_B(net762),
    .D(_0565_),
    .Q_N(_4136_),
    .Q(\i_dm_mem.rdata_q_49_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_4__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0566_),
    .Q_N(_4135_),
    .Q(\i_dm_mem.rdata_q_4_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_50__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net732),
    .D(_0567_),
    .Q_N(_4134_),
    .Q(\i_dm_mem.rdata_q_50_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_51__reg  (.CLK(clknet_leaf_66_clk_i),
    .RESET_B(net762),
    .D(_0568_),
    .Q_N(_4133_),
    .Q(\i_dm_mem.rdata_q_51_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_52__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net732),
    .D(_0569_),
    .Q_N(_4132_),
    .Q(\i_dm_mem.rdata_q_52_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_53__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net736),
    .D(_0570_),
    .Q_N(_4131_),
    .Q(\i_dm_mem.rdata_q_53_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_54__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net736),
    .D(_0571_),
    .Q_N(_4130_),
    .Q(\i_dm_mem.rdata_q_54_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_55__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net736),
    .D(_0572_),
    .Q_N(_4129_),
    .Q(\i_dm_mem.rdata_q_55_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_56__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net739),
    .D(_0573_),
    .Q_N(_4128_),
    .Q(\i_dm_mem.rdata_q_56_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_57__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net740),
    .D(_0574_),
    .Q_N(_4127_),
    .Q(\i_dm_mem.rdata_q_57_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_58__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net740),
    .D(_0575_),
    .Q_N(_4126_),
    .Q(\i_dm_mem.rdata_q_58_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_59__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net737),
    .D(_0576_),
    .Q_N(_4125_),
    .Q(\i_dm_mem.rdata_q_59_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_5__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net733),
    .D(_0577_),
    .Q_N(_4124_),
    .Q(\i_dm_mem.rdata_q_5_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_60__reg  (.CLK(clknet_leaf_79_clk_i),
    .RESET_B(net738),
    .D(_0578_),
    .Q_N(_4123_),
    .Q(\i_dm_mem.rdata_q_60_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_61__reg  (.CLK(clknet_leaf_76_clk_i),
    .RESET_B(net738),
    .D(_0579_),
    .Q_N(_4122_),
    .Q(\i_dm_mem.rdata_q_61_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_62__reg  (.CLK(clknet_leaf_78_clk_i),
    .RESET_B(net736),
    .D(_0580_),
    .Q_N(_4121_),
    .Q(\i_dm_mem.rdata_q_62_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_63__reg  (.CLK(clknet_leaf_85_clk_i),
    .RESET_B(net729),
    .D(_0581_),
    .Q_N(_4120_),
    .Q(\i_dm_mem.rdata_q_63_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_6__reg  (.CLK(clknet_leaf_75_clk_i),
    .RESET_B(net732),
    .D(_0582_),
    .Q_N(_4119_),
    .Q(\i_dm_mem.rdata_q_6_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_7__reg  (.CLK(clknet_leaf_84_clk_i),
    .RESET_B(net730),
    .D(_0583_),
    .Q_N(_4118_),
    .Q(\i_dm_mem.rdata_q_7_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_8__reg  (.CLK(clknet_leaf_77_clk_i),
    .RESET_B(net734),
    .D(_0584_),
    .Q_N(_4117_),
    .Q(\i_dm_mem.rdata_q_8_ ));
 sg13g2_dfrbp_1 \i_dm_mem.rdata_q_9__reg  (.CLK(clknet_leaf_71_clk_i),
    .RESET_B(net738),
    .D(_0585_),
    .Q_N(_4116_),
    .Q(\i_dm_mem.rdata_q_9_ ));
 sg13g2_dfrbp_2 \i_dm_mem.state_q_0__reg  (.RESET_B(net735),
    .D(_0586_),
    .Q(\i_dm_mem.state_q_0_ ),
    .Q_N(\i_dm_mem.state_q_0__$_NOT__A_Y ),
    .CLK(clknet_leaf_74_clk_i));
 sg13g2_dfrbp_1 \i_dm_mem.state_q_1__reg  (.CLK(clknet_leaf_15_clk_i),
    .RESET_B(net694),
    .D(_0587_),
    .Q_N(\i_dm_mem.state_q_1__$_NOT__A_Y ),
    .Q(\i_dm_mem.state_q_1_ ));
 sg13g2_dfrbp_2 \i_dm_mem.word_enable32_q_reg  (.RESET_B(net737),
    .D(slave_addr_i_2_),
    .Q(\i_dm_mem.word_enable32_q ),
    .Q_N(_4115_),
    .CLK(clknet_leaf_79_clk_i));
 sg13g2_dfrbp_2 \i_dm_sba.state_q_0__reg  (.RESET_B(net771),
    .D(_0588_),
    .Q(\i_dm_sba.state_q_0_ ),
    .Q_N(\i_dm_sba.state_q_0__$_NOT__A_Y ),
    .CLK(clknet_leaf_61_clk_i));
 sg13g2_dfrbp_2 \i_dm_sba.state_q_1__reg  (.RESET_B(net771),
    .D(_0589_),
    .Q(\i_dm_sba.state_q_1_ ),
    .Q_N(\i_dm_sba.state_q_1__$_NOT__A_Y ),
    .CLK(clknet_leaf_61_clk_i));
 sg13g2_dfrbp_2 \i_dm_sba.state_q_2__reg  (.RESET_B(net759),
    .D(_0590_),
    .Q(\i_dm_sba.state_q_2_ ),
    .Q_N(\i_dm_csrs.sbbusy_i_$_OR__Y_A_$_OR__A_B ),
    .CLK(clknet_leaf_61_clk_i));
 sg13g2_dfrbp_2 \master_add_o[0]_reg  (.RESET_B(net771),
    .D(\master_add_o[0]_reg_D ),
    .Q(master_add_o_0_),
    .Q_N(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_A ),
    .CLK(clknet_leaf_62_clk_i));
 sg13g2_dfrbp_2 \master_add_o[10]_reg  (.RESET_B(net761),
    .D(\master_add_o[10]_reg_D ),
    .Q(master_add_o_10_),
    .Q_N(_4720_),
    .CLK(clknet_leaf_70_clk_i));
 sg13g2_dfrbp_2 \master_add_o[11]_reg  (.RESET_B(net747),
    .D(\master_add_o[11]_reg_D ),
    .Q(master_add_o_11_),
    .Q_N(_4721_),
    .CLK(clknet_leaf_70_clk_i));
 sg13g2_dfrbp_2 \master_add_o[12]_reg  (.RESET_B(net761),
    .D(\master_add_o[12]_reg_D ),
    .Q(master_add_o_12_),
    .Q_N(_4722_),
    .CLK(clknet_leaf_70_clk_i));
 sg13g2_dfrbp_2 \master_add_o[13]_reg  (.RESET_B(net761),
    .D(\master_add_o[13]_reg_D ),
    .Q(master_add_o_13_),
    .Q_N(_4723_),
    .CLK(clknet_leaf_70_clk_i));
 sg13g2_dfrbp_2 \master_add_o[14]_reg  (.RESET_B(net761),
    .D(\master_add_o[14]_reg_D ),
    .Q(master_add_o_14_),
    .Q_N(_4724_),
    .CLK(clknet_leaf_70_clk_i));
 sg13g2_dfrbp_2 \master_add_o[15]_reg  (.RESET_B(net750),
    .D(\master_add_o[15]_reg_D ),
    .Q(master_add_o_15_),
    .Q_N(_4725_),
    .CLK(clknet_leaf_69_clk_i));
 sg13g2_dfrbp_2 \master_add_o[16]_reg  (.RESET_B(net749),
    .D(\master_add_o[16]_reg_D ),
    .Q(master_add_o_16_),
    .Q_N(_4726_),
    .CLK(clknet_leaf_69_clk_i));
 sg13g2_dfrbp_2 \master_add_o[17]_reg  (.RESET_B(net763),
    .D(\master_add_o[17]_reg_D ),
    .Q(master_add_o_17_),
    .Q_N(_4727_),
    .CLK(clknet_leaf_69_clk_i));
 sg13g2_dfrbp_2 \master_add_o[18]_reg  (.RESET_B(net749),
    .D(\master_add_o[18]_reg_D ),
    .Q(master_add_o_18_),
    .Q_N(_4728_),
    .CLK(clknet_leaf_44_clk_i));
 sg13g2_dfrbp_2 \master_add_o[19]_reg  (.RESET_B(net758),
    .D(\master_add_o[19]_reg_D ),
    .Q(master_add_o_19_),
    .Q_N(_4729_),
    .CLK(clknet_leaf_51_clk_i));
 sg13g2_dfrbp_2 \master_add_o[1]_reg  (.RESET_B(net771),
    .D(\master_add_o[1]_reg_D ),
    .Q(master_add_o_1_),
    .Q_N(\i_dm_sba.be_mask_3__$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_NOT__Y_A_$_OR__Y_B ),
    .CLK(clknet_leaf_53_clk_i));
 sg13g2_dfrbp_2 \master_add_o[20]_reg  (.RESET_B(net758),
    .D(\master_add_o[20]_reg_D ),
    .Q(master_add_o_20_),
    .Q_N(_4730_),
    .CLK(clknet_leaf_51_clk_i));
 sg13g2_dfrbp_2 \master_add_o[21]_reg  (.RESET_B(net758),
    .D(\master_add_o[21]_reg_D ),
    .Q(master_add_o_21_),
    .Q_N(_4731_),
    .CLK(clknet_leaf_51_clk_i));
 sg13g2_dfrbp_2 \master_add_o[22]_reg  (.RESET_B(net757),
    .D(\master_add_o[22]_reg_D ),
    .Q(master_add_o_22_),
    .Q_N(_4732_),
    .CLK(clknet_leaf_52_clk_i));
 sg13g2_dfrbp_2 \master_add_o[23]_reg  (.RESET_B(net758),
    .D(\master_add_o[23]_reg_D ),
    .Q(master_add_o_23_),
    .Q_N(_4733_),
    .CLK(clknet_leaf_50_clk_i));
 sg13g2_dfrbp_2 \master_add_o[24]_reg  (.RESET_B(net759),
    .D(\master_add_o[24]_reg_D ),
    .Q(master_add_o_24_),
    .Q_N(_4734_),
    .CLK(clknet_leaf_51_clk_i));
 sg13g2_dfrbp_2 \master_add_o[25]_reg  (.RESET_B(net759),
    .D(\master_add_o[25]_reg_D ),
    .Q(master_add_o_25_),
    .Q_N(_4735_),
    .CLK(clknet_4_12_0_clk_i));
 sg13g2_dfrbp_2 \master_add_o[26]_reg  (.RESET_B(net771),
    .D(\master_add_o[26]_reg_D ),
    .Q(master_add_o_26_),
    .Q_N(_4736_),
    .CLK(clknet_leaf_54_clk_i));
 sg13g2_dfrbp_2 \master_add_o[27]_reg  (.RESET_B(net777),
    .D(\master_add_o[27]_reg_D ),
    .Q(master_add_o_27_),
    .Q_N(_4737_),
    .CLK(clknet_leaf_54_clk_i));
 sg13g2_dfrbp_2 \master_add_o[28]_reg  (.RESET_B(net759),
    .D(\master_add_o[28]_reg_D ),
    .Q(master_add_o_28_),
    .Q_N(_4738_),
    .CLK(clknet_leaf_54_clk_i));
 sg13g2_dfrbp_2 \master_add_o[29]_reg  (.RESET_B(net759),
    .D(\master_add_o[29]_reg_D ),
    .Q(master_add_o_29_),
    .Q_N(_4739_),
    .CLK(clknet_leaf_52_clk_i));
 sg13g2_dfrbp_2 \master_add_o[2]_reg  (.RESET_B(net763),
    .D(\master_add_o[2]_reg_D ),
    .Q(master_add_o_2_),
    .Q_N(_4740_),
    .CLK(clknet_leaf_67_clk_i));
 sg13g2_dfrbp_2 \master_add_o[30]_reg  (.RESET_B(net771),
    .D(\master_add_o[30]_reg_D ),
    .Q(master_add_o_30_),
    .Q_N(_4741_),
    .CLK(clknet_leaf_53_clk_i));
 sg13g2_dfrbp_2 \master_add_o[31]_reg  (.RESET_B(net771),
    .D(\master_add_o[31]_reg_D ),
    .Q(master_add_o_31_),
    .Q_N(_4742_),
    .CLK(clknet_leaf_53_clk_i));
 sg13g2_dfrbp_2 \master_add_o[3]_reg  (.RESET_B(net771),
    .D(\master_add_o[3]_reg_D ),
    .Q(master_add_o_3_),
    .Q_N(_4743_),
    .CLK(clknet_leaf_53_clk_i));
 sg13g2_dfrbp_1 \master_add_o[4]_reg  (.CLK(clknet_leaf_68_clk_i),
    .RESET_B(net763),
    .D(\master_add_o[4]_reg_D ),
    .Q_N(_4744_),
    .Q(net49));
 sg13g2_dfrbp_2 \master_add_o[5]_reg  (.RESET_B(net761),
    .D(\master_add_o[5]_reg_D ),
    .Q(master_add_o_5_),
    .Q_N(_4745_),
    .CLK(clknet_leaf_67_clk_i));
 sg13g2_dfrbp_2 \master_add_o[6]_reg  (.RESET_B(net763),
    .D(\master_add_o[6]_reg_D ),
    .Q(master_add_o_6_),
    .Q_N(_4746_),
    .CLK(clknet_leaf_62_clk_i));
 sg13g2_dfrbp_2 \master_add_o[7]_reg  (.RESET_B(net762),
    .D(\master_add_o[7]_reg_D ),
    .Q(master_add_o_7_),
    .Q_N(_4747_),
    .CLK(clknet_leaf_67_clk_i));
 sg13g2_dfrbp_2 \master_add_o[8]_reg  (.RESET_B(net758),
    .D(\master_add_o[8]_reg_D ),
    .Q(master_add_o_8_),
    .Q_N(_4748_),
    .CLK(clknet_leaf_50_clk_i));
 sg13g2_dfrbp_2 \master_add_o[9]_reg  (.RESET_B(net777),
    .D(\master_add_o[9]_reg_D ),
    .Q(master_add_o_9_),
    .Q_N(_4114_),
    .CLK(clknet_leaf_54_clk_i));
 sg13g2_dfrbp_2 ndmreset_o_reg (.RESET_B(net742),
    .D(_0591_),
    .Q(ndmreset_o),
    .Q_N(_4113_),
    .CLK(clknet_leaf_40_clk_i));
 sg13g2_buf_2 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(net449),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(net449),
    .X(net448));
 sg13g2_buf_1 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(_2856_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(net454),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(net453));
 sg13g2_buf_2 fanout453 (.A(net454),
    .X(net453));
 sg13g2_buf_4 fanout454 (.X(net454),
    .A(_2834_));
 sg13g2_buf_8 fanout455 (.A(_2657_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_2657_),
    .X(net456));
 sg13g2_buf_4 fanout457 (.X(net457),
    .A(net460));
 sg13g2_buf_1 fanout458 (.A(net460),
    .X(net458));
 sg13g2_buf_4 fanout459 (.X(net459),
    .A(net460));
 sg13g2_buf_2 fanout460 (.A(_2368_),
    .X(net460));
 sg13g2_buf_4 fanout461 (.X(net461),
    .A(net462));
 sg13g2_buf_4 fanout462 (.X(net462),
    .A(_2368_));
 sg13g2_buf_4 fanout463 (.X(net463),
    .A(net465));
 sg13g2_buf_4 fanout464 (.X(net464),
    .A(net465));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_2266_));
 sg13g2_buf_4 fanout466 (.X(net466),
    .A(net467));
 sg13g2_buf_4 fanout467 (.X(net467),
    .A(_2266_));
 sg13g2_buf_4 fanout468 (.X(net468),
    .A(net470));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(net470));
 sg13g2_buf_4 fanout470 (.X(net470),
    .A(_2176_));
 sg13g2_buf_4 fanout471 (.X(net471),
    .A(net472));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_2176_));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(net475));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(net475));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(_2092_));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(net477));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_2092_));
 sg13g2_buf_4 fanout478 (.X(net478),
    .A(net480));
 sg13g2_buf_4 fanout479 (.X(net479),
    .A(net480));
 sg13g2_buf_2 fanout480 (.A(_1772_),
    .X(net480));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(net482));
 sg13g2_buf_4 fanout482 (.X(net482),
    .A(_1772_));
 sg13g2_buf_2 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net487),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(net487),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(net487),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_1317_),
    .X(net487));
 sg13g2_buf_4 fanout488 (.X(net488),
    .A(net490));
 sg13g2_buf_4 fanout489 (.X(net489),
    .A(net490));
 sg13g2_buf_2 fanout490 (.A(_1292_),
    .X(net490));
 sg13g2_buf_4 fanout491 (.X(net491),
    .A(net492));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_1292_));
 sg13g2_buf_2 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(net495),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_3790_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_3771_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_3170_),
    .X(net497));
 sg13g2_buf_4 fanout498 (.X(net498),
    .A(_3122_));
 sg13g2_buf_1 fanout499 (.A(_3122_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_3122_),
    .X(net501));
 sg13g2_buf_16 fanout502 (.X(net502),
    .A(net505));
 sg13g2_buf_16 fanout503 (.X(net503),
    .A(net504));
 sg13g2_buf_16 fanout504 (.X(net504),
    .A(net505));
 sg13g2_buf_8 fanout505 (.A(_2839_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(net509),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(net509),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(net515),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(net514),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(net513),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_4 fanout515 (.X(net515),
    .A(_2835_));
 sg13g2_buf_4 fanout516 (.X(net516),
    .A(net518));
 sg13g2_buf_4 fanout517 (.X(net517),
    .A(net518));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(_2012_));
 sg13g2_buf_4 fanout519 (.X(net519),
    .A(net520));
 sg13g2_buf_4 fanout520 (.X(net520),
    .A(_2012_));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(net523));
 sg13g2_buf_4 fanout522 (.X(net522),
    .A(net523));
 sg13g2_buf_4 fanout523 (.X(net523),
    .A(_1906_));
 sg13g2_buf_4 fanout524 (.X(net524),
    .A(net525));
 sg13g2_buf_4 fanout525 (.X(net525),
    .A(_1906_));
 sg13g2_buf_2 fanout526 (.A(_1480_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_2 fanout529 (.A(_1364_),
    .X(net529));
 sg13g2_buf_4 fanout530 (.X(net530),
    .A(net531));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(net532));
 sg13g2_buf_4 fanout532 (.X(net532),
    .A(_1355_));
 sg13g2_buf_2 fanout533 (.A(net534),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(net535),
    .X(net534));
 sg13g2_buf_4 fanout535 (.X(net535),
    .A(_1327_));
 sg13g2_buf_4 fanout536 (.X(net536),
    .A(net537));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(net540));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(net540));
 sg13g2_buf_2 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_0898_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_3782_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_3088_),
    .X(net543));
 sg13g2_buf_4 fanout544 (.X(net544),
    .A(net545));
 sg13g2_buf_2 fanout545 (.A(_3074_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_2557_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_1210_),
    .X(net547));
 sg13g2_buf_1 fanout548 (.A(_1210_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_1202_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(net552),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(net552),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(net554),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(net554),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(net555),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_0710_),
    .X(net555));
 sg13g2_buf_4 fanout556 (.X(net556),
    .A(_0609_));
 sg13g2_buf_2 fanout557 (.A(net558),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_3147_),
    .X(net558));
 sg13g2_buf_4 fanout559 (.X(net559),
    .A(net561));
 sg13g2_buf_2 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(net563),
    .X(net561));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(net563));
 sg13g2_buf_2 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_3120_));
 sg13g2_buf_2 fanout565 (.A(_3110_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(net567),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_3087_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_3087_),
    .X(net569));
 sg13g2_buf_2 fanout570 (.A(net572),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(net572),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_3082_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_3082_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_3078_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_3070_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_3066_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_1322_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(net585),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(net585),
    .X(net583));
 sg13g2_buf_1 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_1179_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_1179_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_1179_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(net589),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_4 fanout590 (.X(net590),
    .A(net591));
 sg13g2_buf_4 fanout591 (.X(net591),
    .A(_1172_));
 sg13g2_buf_2 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(net595),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net595),
    .X(net594));
 sg13g2_buf_1 fanout595 (.A(net599),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(net599),
    .X(net597));
 sg13g2_buf_16 fanout598 (.X(net598),
    .A(net599));
 sg13g2_buf_16 fanout599 (.X(net599),
    .A(_1165_));
 sg13g2_buf_2 fanout600 (.A(net607),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net603),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_1 fanout603 (.A(net607),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(net606),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(net606),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(net607),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_0895_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(net612),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net612),
    .X(net610));
 sg13g2_buf_1 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_1 fanout612 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.rdata_o_42__$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(net617),
    .X(net613));
 sg13g2_buf_2 fanout614 (.A(net617),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net616),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_1 fanout617 (.A(\i_dm_mem.gen_rom_snd_scratch.i_debug_rom.addr_q_0_ ),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(net621),
    .X(net620));
 sg13g2_buf_4 fanout621 (.X(net621),
    .A(net627));
 sg13g2_buf_2 fanout622 (.A(net623),
    .X(net622));
 sg13g2_buf_1 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(net627),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(net627),
    .X(net625));
 sg13g2_buf_1 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(\i_dm_mem.fwd_rom_q ),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(\i_dm_csrs.sbaccess_o_2_ ),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(\i_dm_csrs.sbaccess_o_1_ ),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(net633),
    .X(net631));
 sg13g2_buf_1 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_1 fanout633 (.A(\i_dm_csrs.sbaccess_o_0_ ),
    .X(net633));
 sg13g2_buf_4 fanout634 (.X(net634),
    .A(net636));
 sg13g2_buf_4 fanout635 (.X(net635),
    .A(net636));
 sg13g2_buf_2 fanout636 (.A(\i_dm_csrs.i_fifo.read_pointer_q ),
    .X(net636));
 sg13g2_buf_4 fanout637 (.X(net637),
    .A(net638));
 sg13g2_buf_4 fanout638 (.X(net638),
    .A(\i_dm_csrs.i_fifo.read_pointer_q ));
 sg13g2_buf_2 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_1 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(\ndmreset_o_reg_E_$_AND__Y_B_$_OR__Y_A ),
    .X(net641));
 sg13g2_buf_4 fanout642 (.X(net642),
    .A(slave_req_i));
 sg13g2_buf_2 fanout643 (.A(slave_req_i),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(slave_addr_i_6_),
    .X(net645));
 sg13g2_buf_4 fanout646 (.X(net646),
    .A(net649));
 sg13g2_buf_4 fanout647 (.X(net647),
    .A(net649));
 sg13g2_buf_4 fanout648 (.X(net648),
    .A(net649));
 sg13g2_buf_2 fanout649 (.A(slave_addr_i_4_),
    .X(net649));
 sg13g2_buf_4 fanout650 (.X(net650),
    .A(net652));
 sg13g2_buf_4 fanout651 (.X(net651),
    .A(net652));
 sg13g2_buf_8 fanout652 (.A(slave_addr_i_4_),
    .X(net652));
 sg13g2_buf_4 fanout653 (.X(net653),
    .A(net654));
 sg13g2_buf_4 fanout654 (.X(net654),
    .A(net661));
 sg13g2_buf_2 fanout655 (.A(net661),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net660),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(net660),
    .X(net658));
 sg13g2_buf_1 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(slave_addr_i_4_),
    .X(net662));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(net665));
 sg13g2_buf_2 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_4 fanout665 (.X(net665),
    .A(net672));
 sg13g2_buf_4 fanout666 (.X(net666),
    .A(net672));
 sg13g2_buf_4 fanout667 (.X(net667),
    .A(net671));
 sg13g2_buf_2 fanout668 (.A(net671),
    .X(net668));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(net671));
 sg13g2_buf_4 fanout670 (.X(net670),
    .A(net671));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net696),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(net677));
 sg13g2_buf_4 fanout674 (.X(net674),
    .A(net677));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(net676));
 sg13g2_buf_4 fanout676 (.X(net676),
    .A(net677));
 sg13g2_buf_2 fanout677 (.A(net696),
    .X(net677));
 sg13g2_buf_4 fanout678 (.X(net678),
    .A(net680));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(net680));
 sg13g2_buf_4 fanout680 (.X(net680),
    .A(net696));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(net682));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(net684));
 sg13g2_buf_4 fanout683 (.X(net683),
    .A(net684));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(net696));
 sg13g2_buf_4 fanout685 (.X(net685),
    .A(net689));
 sg13g2_buf_4 fanout686 (.X(net686),
    .A(net689));
 sg13g2_buf_4 fanout687 (.X(net687),
    .A(net689));
 sg13g2_buf_4 fanout688 (.X(net688),
    .A(net689));
 sg13g2_buf_2 fanout689 (.A(net696),
    .X(net689));
 sg13g2_buf_4 fanout690 (.X(net690),
    .A(net691));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(net695));
 sg13g2_buf_4 fanout692 (.X(net692),
    .A(net694));
 sg13g2_buf_4 fanout693 (.X(net693),
    .A(net694));
 sg13g2_buf_4 fanout694 (.X(net694),
    .A(net695));
 sg13g2_buf_2 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_4 fanout696 (.X(net696),
    .A(net779));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(net701));
 sg13g2_buf_4 fanout698 (.X(net698),
    .A(net701));
 sg13g2_buf_4 fanout699 (.X(net699),
    .A(net701));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(net701));
 sg13g2_buf_2 fanout701 (.A(net706),
    .X(net701));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(net706));
 sg13g2_buf_2 fanout703 (.A(net706),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(net705));
 sg13g2_buf_4 fanout705 (.X(net705),
    .A(net706));
 sg13g2_buf_2 fanout706 (.A(net726),
    .X(net706));
 sg13g2_buf_4 fanout707 (.X(net707),
    .A(net712));
 sg13g2_buf_4 fanout708 (.X(net708),
    .A(net711));
 sg13g2_buf_2 fanout709 (.A(net711),
    .X(net709));
 sg13g2_buf_4 fanout710 (.X(net710),
    .A(net711));
 sg13g2_buf_2 fanout711 (.A(net712),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(net726),
    .X(net712));
 sg13g2_buf_4 fanout713 (.X(net713),
    .A(net715));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_4 fanout715 (.X(net715),
    .A(net726));
 sg13g2_buf_4 fanout716 (.X(net716),
    .A(net720));
 sg13g2_buf_2 fanout717 (.A(net720),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(net720));
 sg13g2_buf_2 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(net725),
    .X(net720));
 sg13g2_buf_4 fanout721 (.X(net721),
    .A(net725));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(net725));
 sg13g2_buf_4 fanout723 (.X(net723),
    .A(net724));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(net725));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_4 fanout726 (.X(net726),
    .A(net779));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(net728));
 sg13g2_buf_4 fanout728 (.X(net728),
    .A(net730));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(net730));
 sg13g2_buf_4 fanout730 (.X(net730),
    .A(net741));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(net735));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(net733));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(net735));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(net735));
 sg13g2_buf_4 fanout735 (.X(net735),
    .A(net741));
 sg13g2_buf_4 fanout736 (.X(net736),
    .A(net739));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(net738));
 sg13g2_buf_4 fanout738 (.X(net738),
    .A(net739));
 sg13g2_buf_2 fanout739 (.A(net741),
    .X(net739));
 sg13g2_buf_4 fanout740 (.X(net740),
    .A(net741));
 sg13g2_buf_4 fanout741 (.X(net741),
    .A(net779));
 sg13g2_buf_4 fanout742 (.X(net742),
    .A(net743));
 sg13g2_buf_4 fanout743 (.X(net743),
    .A(net751));
 sg13g2_buf_4 fanout744 (.X(net744),
    .A(net751));
 sg13g2_buf_2 fanout745 (.A(net751),
    .X(net745));
 sg13g2_buf_4 fanout746 (.X(net746),
    .A(net747));
 sg13g2_buf_4 fanout747 (.X(net747),
    .A(net750));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(net750));
 sg13g2_buf_2 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net751),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(net760),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(net753));
 sg13g2_buf_2 fanout753 (.A(net760),
    .X(net753));
 sg13g2_buf_4 fanout754 (.X(net754),
    .A(net756));
 sg13g2_buf_4 fanout755 (.X(net755),
    .A(net756));
 sg13g2_buf_2 fanout756 (.A(net760),
    .X(net756));
 sg13g2_buf_4 fanout757 (.X(net757),
    .A(net759));
 sg13g2_buf_4 fanout758 (.X(net758),
    .A(net759));
 sg13g2_buf_4 fanout759 (.X(net759),
    .A(net760));
 sg13g2_buf_2 fanout760 (.A(net778),
    .X(net760));
 sg13g2_buf_4 fanout761 (.X(net761),
    .A(net762));
 sg13g2_buf_4 fanout762 (.X(net762),
    .A(net763));
 sg13g2_buf_4 fanout763 (.X(net763),
    .A(net778));
 sg13g2_buf_4 fanout764 (.X(net764),
    .A(net770));
 sg13g2_buf_2 fanout765 (.A(net770),
    .X(net765));
 sg13g2_buf_4 fanout766 (.X(net766),
    .A(net770));
 sg13g2_buf_4 fanout767 (.X(net767),
    .A(net769));
 sg13g2_buf_4 fanout768 (.X(net768),
    .A(net769));
 sg13g2_buf_2 fanout769 (.A(net770),
    .X(net769));
 sg13g2_buf_1 fanout770 (.A(net778),
    .X(net770));
 sg13g2_buf_4 fanout771 (.X(net771),
    .A(net777));
 sg13g2_buf_4 fanout772 (.X(net772),
    .A(net773));
 sg13g2_buf_4 fanout773 (.X(net773),
    .A(net777));
 sg13g2_buf_4 fanout774 (.X(net774),
    .A(net776));
 sg13g2_buf_2 fanout775 (.A(net776),
    .X(net775));
 sg13g2_buf_4 fanout776 (.X(net776),
    .A(net777));
 sg13g2_buf_2 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_4 fanout779 (.X(net779),
    .A(rst_ni));
 sg13g2_buf_2 fanout780 (.A(net789),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(net789),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(net784),
    .X(net782));
 sg13g2_buf_1 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_1 fanout784 (.A(net789),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(net789),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(net796),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(net792),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net793),
    .X(net791));
 sg13g2_buf_1 fanout792 (.A(net793),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(net796),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net796),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(master_r_valid_i),
    .X(net796));
 sg13g2_buf_4 fanout797 (.X(net797),
    .A(dmi_req_i_36_));
 sg13g2_buf_4 fanout798 (.X(net798),
    .A(net799));
 sg13g2_buf_8 fanout799 (.A(dmi_req_i_23_),
    .X(net799));
 sg13g2_buf_2 fanout800 (.A(net801),
    .X(net800));
 sg13g2_buf_4 fanout801 (.X(net801),
    .A(net802));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(dmi_req_i_13_));
 sg13g2_buf_2 rebuffer803 (.A(_2553_),
    .X(net803));
 sg13g2_buf_16 clkbuf_leaf_0_clk_i (.X(clknet_leaf_0_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_1_clk_i (.X(clknet_leaf_1_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_2_clk_i (.X(clknet_leaf_2_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_3_clk_i (.X(clknet_leaf_3_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_4_clk_i (.X(clknet_leaf_4_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_5_clk_i (.X(clknet_leaf_5_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_6_clk_i (.X(clknet_leaf_6_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_7_clk_i (.X(clknet_leaf_7_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_8_clk_i (.X(clknet_leaf_8_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_9_clk_i (.X(clknet_leaf_9_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_10_clk_i (.X(clknet_leaf_10_clk_i),
    .A(clknet_4_1_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_11_clk_i (.X(clknet_leaf_11_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_12_clk_i (.X(clknet_leaf_12_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_13_clk_i (.X(clknet_leaf_13_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_14_clk_i (.X(clknet_leaf_14_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_15_clk_i (.X(clknet_leaf_15_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_16_clk_i (.X(clknet_leaf_16_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_17_clk_i (.X(clknet_leaf_17_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_18_clk_i (.X(clknet_leaf_18_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_19_clk_i (.X(clknet_leaf_19_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_20_clk_i (.X(clknet_leaf_20_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_21_clk_i (.X(clknet_leaf_21_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_22_clk_i (.X(clknet_leaf_22_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_23_clk_i (.X(clknet_leaf_23_clk_i),
    .A(clknet_4_4_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_24_clk_i (.X(clknet_leaf_24_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_25_clk_i (.X(clknet_leaf_25_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_26_clk_i (.X(clknet_leaf_26_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_27_clk_i (.X(clknet_leaf_27_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_28_clk_i (.X(clknet_leaf_28_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_29_clk_i (.X(clknet_leaf_29_clk_i),
    .A(clknet_4_5_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_30_clk_i (.X(clknet_leaf_30_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_31_clk_i (.X(clknet_leaf_31_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_32_clk_i (.X(clknet_leaf_32_clk_i),
    .A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_33_clk_i (.X(clknet_leaf_33_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_34_clk_i (.X(clknet_leaf_34_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_35_clk_i (.X(clknet_leaf_35_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_36_clk_i (.X(clknet_leaf_36_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_37_clk_i (.X(clknet_leaf_37_clk_i),
    .A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_39_clk_i (.X(clknet_leaf_39_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_40_clk_i (.X(clknet_leaf_40_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_41_clk_i (.X(clknet_leaf_41_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_42_clk_i (.X(clknet_leaf_42_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_43_clk_i (.X(clknet_leaf_43_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_44_clk_i (.X(clknet_leaf_44_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_45_clk_i (.X(clknet_leaf_45_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_46_clk_i (.X(clknet_leaf_46_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_47_clk_i (.X(clknet_leaf_47_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_48_clk_i (.X(clknet_leaf_48_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_49_clk_i (.X(clknet_leaf_49_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_50_clk_i (.X(clknet_leaf_50_clk_i),
    .A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_51_clk_i (.X(clknet_leaf_51_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_52_clk_i (.X(clknet_leaf_52_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_53_clk_i (.X(clknet_leaf_53_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_54_clk_i (.X(clknet_leaf_54_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_56_clk_i (.X(clknet_leaf_56_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_57_clk_i (.X(clknet_leaf_57_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_58_clk_i (.X(clknet_leaf_58_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_59_clk_i (.X(clknet_leaf_59_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_60_clk_i (.X(clknet_leaf_60_clk_i),
    .A(clknet_4_15_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_61_clk_i (.X(clknet_leaf_61_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_62_clk_i (.X(clknet_leaf_62_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_63_clk_i (.X(clknet_leaf_63_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_64_clk_i (.X(clknet_leaf_64_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_65_clk_i (.X(clknet_leaf_65_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_66_clk_i (.X(clknet_leaf_66_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_67_clk_i (.X(clknet_leaf_67_clk_i),
    .A(clknet_4_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_68_clk_i (.X(clknet_leaf_68_clk_i),
    .A(clknet_4_14_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_69_clk_i (.X(clknet_leaf_69_clk_i),
    .A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_70_clk_i (.X(clknet_leaf_70_clk_i),
    .A(clknet_4_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_71_clk_i (.X(clknet_leaf_71_clk_i),
    .A(clknet_4_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_72_clk_i (.X(clknet_leaf_72_clk_i),
    .A(clknet_4_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_73_clk_i (.X(clknet_leaf_73_clk_i),
    .A(clknet_4_9_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_74_clk_i (.X(clknet_leaf_74_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_75_clk_i (.X(clknet_leaf_75_clk_i),
    .A(clknet_4_11_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_76_clk_i (.X(clknet_leaf_76_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_77_clk_i (.X(clknet_leaf_77_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_78_clk_i (.X(clknet_leaf_78_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_79_clk_i (.X(clknet_leaf_79_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_81_clk_i (.X(clknet_leaf_81_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_82_clk_i (.X(clknet_leaf_82_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_83_clk_i (.X(clknet_leaf_83_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_84_clk_i (.X(clknet_leaf_84_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_85_clk_i (.X(clknet_leaf_85_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_86_clk_i (.X(clknet_leaf_86_clk_i),
    .A(clknet_4_10_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_87_clk_i (.X(clknet_leaf_87_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_88_clk_i (.X(clknet_leaf_88_clk_i),
    .A(clknet_4_8_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_89_clk_i (.X(clknet_leaf_89_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_90_clk_i (.X(clknet_leaf_90_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_91_clk_i (.X(clknet_leaf_91_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_92_clk_i (.X(clknet_leaf_92_clk_i),
    .A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_93_clk_i (.X(clknet_leaf_93_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_94_clk_i (.X(clknet_leaf_94_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_95_clk_i (.X(clknet_leaf_95_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_96_clk_i (.X(clknet_leaf_96_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_97_clk_i (.X(clknet_leaf_97_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_98_clk_i (.X(clknet_leaf_98_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_99_clk_i (.X(clknet_leaf_99_clk_i),
    .A(clknet_4_2_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_100_clk_i (.X(clknet_leaf_100_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_101_clk_i (.X(clknet_leaf_101_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_102_clk_i (.X(clknet_leaf_102_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_103_clk_i (.X(clknet_leaf_103_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_16 clkbuf_leaf_104_clk_i (.X(clknet_leaf_104_clk_i),
    .A(clknet_4_0_0_clk_i));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_0_0_clk_i (.X(clknet_4_0_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_1_0_clk_i (.X(clknet_4_1_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_2_0_clk_i (.X(clknet_4_2_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_3_0_clk_i (.X(clknet_4_3_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_4_0_clk_i (.X(clknet_4_4_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_5_0_clk_i (.X(clknet_4_5_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_6_0_clk_i (.X(clknet_4_6_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_7_0_clk_i (.X(clknet_4_7_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_8_0_clk_i (.X(clknet_4_8_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_9_0_clk_i (.X(clknet_4_9_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_10_0_clk_i (.X(clknet_4_10_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_11_0_clk_i (.X(clknet_4_11_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_12_0_clk_i (.X(clknet_4_12_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_13_0_clk_i (.X(clknet_4_13_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_14_0_clk_i (.X(clknet_4_14_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_15_0_clk_i (.X(clknet_4_15_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkload0 (.A(clknet_4_3_0_clk_i));
 sg13g2_buf_16 clkload1 (.A(clknet_4_5_0_clk_i));
 sg13g2_inv_4 clkload2 (.A(clknet_4_6_0_clk_i));
 sg13g2_buf_16 clkload3 (.A(clknet_4_7_0_clk_i));
 sg13g2_buf_16 clkload4 (.A(clknet_4_9_0_clk_i));
 sg13g2_inv_8 clkload5 (.A(clknet_4_11_0_clk_i));
 sg13g2_inv_4 clkload6 (.A(clknet_4_12_0_clk_i));
 sg13g2_buf_16 clkload7 (.A(clknet_4_13_0_clk_i));
 sg13g2_buf_16 clkload8 (.A(clknet_4_15_0_clk_i));
 sg13g2_inv_2 clkload9 (.A(clknet_leaf_2_clk_i));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_100_clk_i));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_101_clk_i));
 sg13g2_inv_4 clkload12 (.A(clknet_leaf_104_clk_i));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_3_clk_i));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_8_clk_i));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_10_clk_i));
 sg13g2_inv_1 clkload16 (.A(clknet_leaf_97_clk_i));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_99_clk_i));
 sg13g2_buf_2 clkload18 (.A(clknet_leaf_11_clk_i));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_12_clk_i));
 sg13g2_inv_2 clkload20 (.A(clknet_leaf_89_clk_i));
 sg13g2_inv_2 clkload21 (.A(clknet_leaf_91_clk_i));
 sg13g2_buf_2 clkload22 (.A(clknet_leaf_92_clk_i));
 sg13g2_inv_1 clkload23 (.A(clknet_leaf_7_clk_i));
 sg13g2_inv_4 clkload24 (.A(clknet_leaf_9_clk_i));
 sg13g2_buf_16 clkload25 (.A(clknet_leaf_19_clk_i));
 sg13g2_buf_2 clkload26 (.A(clknet_leaf_21_clk_i));
 sg13g2_inv_1 clkload27 (.A(clknet_leaf_22_clk_i));
 sg13g2_inv_2 clkload28 (.A(clknet_leaf_23_clk_i));
 sg13g2_inv_1 clkload29 (.A(clknet_leaf_24_clk_i));
 sg13g2_inv_1 clkload30 (.A(clknet_leaf_25_clk_i));
 sg13g2_buf_8 clkload31 (.A(clknet_leaf_26_clk_i));
 sg13g2_inv_1 clkload32 (.A(clknet_leaf_27_clk_i));
 sg13g2_buf_16 clkload33 (.A(clknet_leaf_29_clk_i));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_13_clk_i));
 sg13g2_buf_2 clkload35 (.A(clknet_leaf_14_clk_i));
 sg13g2_buf_2 clkload36 (.A(clknet_leaf_16_clk_i));
 sg13g2_inv_4 clkload37 (.A(clknet_leaf_17_clk_i));
 sg13g2_buf_2 clkload38 (.A(clknet_leaf_18_clk_i));
 sg13g2_buf_4 clkload39 (.A(clknet_leaf_31_clk_i));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_33_clk_i));
 sg13g2_buf_2 clkload41 (.A(clknet_leaf_35_clk_i));
 sg13g2_buf_2 clkload42 (.A(clknet_leaf_37_clk_i));
 sg13g2_buf_16 clkload43 (.A(clknet_leaf_74_clk_i));
 sg13g2_buf_4 clkload44 (.A(clknet_leaf_82_clk_i));
 sg13g2_buf_4 clkload45 (.A(clknet_leaf_83_clk_i));
 sg13g2_buf_2 clkload46 (.A(clknet_leaf_84_clk_i));
 sg13g2_buf_16 clkload47 (.A(clknet_leaf_87_clk_i));
 sg13g2_buf_16 clkload48 (.A(clknet_leaf_88_clk_i));
 sg13g2_buf_8 clkload49 (.A(clknet_leaf_15_clk_i));
 sg13g2_buf_8 clkload50 (.A(clknet_leaf_39_clk_i));
 sg13g2_inv_1 clkload51 (.A(clknet_leaf_42_clk_i));
 sg13g2_inv_2 clkload52 (.A(clknet_leaf_43_clk_i));
 sg13g2_buf_8 clkload53 (.A(clknet_leaf_73_clk_i));
 sg13g2_inv_1 clkload54 (.A(clknet_leaf_77_clk_i));
 sg13g2_buf_2 clkload55 (.A(clknet_leaf_79_clk_i));
 sg13g2_inv_4 clkload56 (.A(clknet_leaf_81_clk_i));
 sg13g2_inv_4 clkload57 (.A(clknet_leaf_86_clk_i));
 sg13g2_inv_2 clkload58 (.A(clknet_leaf_70_clk_i));
 sg13g2_buf_2 clkload59 (.A(clknet_leaf_71_clk_i));
 sg13g2_buf_2 clkload60 (.A(clknet_leaf_75_clk_i));
 sg13g2_buf_2 clkload61 (.A(clknet_leaf_45_clk_i));
 sg13g2_buf_2 clkload62 (.A(clknet_leaf_51_clk_i));
 sg13g2_inv_2 clkload63 (.A(clknet_leaf_53_clk_i));
 sg13g2_buf_2 clkload64 (.A(clknet_leaf_69_clk_i));
 sg13g2_inv_2 clkload65 (.A(clknet_leaf_50_clk_i));
 sg13g2_inv_4 clkload66 (.A(clknet_leaf_61_clk_i));
 sg13g2_buf_16 clkload67 (.A(clknet_leaf_62_clk_i));
 sg13g2_inv_4 clkload68 (.A(clknet_leaf_68_clk_i));
 sg13g2_inv_4 clkload69 (.A(clknet_leaf_54_clk_i));
 sg13g2_inv_2 clkload70 (.A(clknet_leaf_60_clk_i));
 sg13g2_antennanp ANTENNA_1 (.A(_1134_));
 sg13g2_antennanp ANTENNA_2 (.A(_1408_));
 sg13g2_antennanp ANTENNA_3 (.A(_1419_));
 sg13g2_antennanp ANTENNA_4 (.A(_1455_));
 sg13g2_antennanp ANTENNA_5 (.A(_1553_));
 sg13g2_antennanp ANTENNA_6 (.A(_1573_));
 sg13g2_antennanp ANTENNA_7 (.A(_1573_));
 sg13g2_antennanp ANTENNA_8 (.A(_1637_));
 sg13g2_antennanp ANTENNA_9 (.A(_1659_));
 sg13g2_antennanp ANTENNA_10 (.A(_1714_));
 sg13g2_antennanp ANTENNA_11 (.A(_1744_));
 sg13g2_antennanp ANTENNA_12 (.A(_1798_));
 sg13g2_antennanp ANTENNA_13 (.A(net221));
 sg13g2_antennanp ANTENNA_14 (.A(net221));
 sg13g2_antennanp ANTENNA_15 (.A(net221));
 sg13g2_antennanp ANTENNA_16 (.A(net221));
 sg13g2_antennanp ANTENNA_17 (.A(net221));
 sg13g2_antennanp ANTENNA_18 (.A(net221));
 sg13g2_antennanp ANTENNA_19 (.A(net221));
 sg13g2_antennanp ANTENNA_20 (.A(net221));
 sg13g2_antennanp ANTENNA_21 (.A(net221));
 sg13g2_antennanp ANTENNA_22 (.A(net128));
 sg13g2_antennanp ANTENNA_23 (.A(net128));
 sg13g2_antennanp ANTENNA_24 (.A(net128));
 sg13g2_antennanp ANTENNA_25 (.A(net128));
 sg13g2_antennanp ANTENNA_26 (.A(net128));
 sg13g2_antennanp ANTENNA_27 (.A(net128));
 sg13g2_antennanp ANTENNA_28 (.A(net128));
 sg13g2_antennanp ANTENNA_29 (.A(net128));
 sg13g2_antennanp ANTENNA_30 (.A(net128));
 sg13g2_antennanp ANTENNA_31 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_32 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_33 (.A(hartinfo_i_13_));
 sg13g2_antennanp ANTENNA_34 (.A(hartinfo_i_18_));
 sg13g2_antennanp ANTENNA_35 (.A(hartinfo_i_19_));
 sg13g2_antennanp ANTENNA_36 (.A(hartinfo_i_22_));
 sg13g2_antennanp ANTENNA_37 (.A(hartinfo_i_26_));
 sg13g2_antennanp ANTENNA_38 (.A(hartinfo_i_30_));
 sg13g2_antennanp ANTENNA_39 (.A(hartinfo_i_3_));
 sg13g2_antennanp ANTENNA_40 (.A(hartinfo_i_5_));
 sg13g2_antennanp ANTENNA_41 (.A(hartinfo_i_9_));
 sg13g2_antennanp ANTENNA_42 (.A(master_r_rdata_i_26_));
 sg13g2_antennanp ANTENNA_43 (.A(master_r_rdata_i_26_));
 sg13g2_antennanp ANTENNA_44 (.A(master_r_rdata_i_26_));
 sg13g2_antennanp ANTENNA_45 (.A(master_r_rdata_i_26_));
 sg13g2_antennanp ANTENNA_46 (.A(next_dm_addr_i_13_));
 sg13g2_antennanp ANTENNA_47 (.A(next_dm_addr_i_14_));
 sg13g2_antennanp ANTENNA_48 (.A(next_dm_addr_i_16_));
 sg13g2_antennanp ANTENNA_49 (.A(next_dm_addr_i_17_));
 sg13g2_antennanp ANTENNA_50 (.A(next_dm_addr_i_19_));
 sg13g2_antennanp ANTENNA_51 (.A(next_dm_addr_i_1_));
 sg13g2_antennanp ANTENNA_52 (.A(next_dm_addr_i_20_));
 sg13g2_antennanp ANTENNA_53 (.A(next_dm_addr_i_26_));
 sg13g2_antennanp ANTENNA_54 (.A(next_dm_addr_i_28_));
 sg13g2_antennanp ANTENNA_55 (.A(next_dm_addr_i_2_));
 sg13g2_antennanp ANTENNA_56 (.A(next_dm_addr_i_30_));
 sg13g2_antennanp ANTENNA_57 (.A(next_dm_addr_i_8_));
 sg13g2_antennanp ANTENNA_58 (.A(slave_addr_i_6_));
 sg13g2_antennanp ANTENNA_59 (.A(slave_addr_i_9_));
 sg13g2_antennanp ANTENNA_60 (.A(slave_addr_i_9_));
 sg13g2_antennanp ANTENNA_61 (.A(slave_addr_i_9_));
 sg13g2_antennanp ANTENNA_62 (.A(slave_addr_i_9_));
 sg13g2_antennanp ANTENNA_63 (.A(slave_addr_i_9_));
 sg13g2_antennanp ANTENNA_64 (.A(net779));
 sg13g2_antennanp ANTENNA_65 (.A(net779));
 sg13g2_antennanp ANTENNA_66 (.A(net779));
 sg13g2_antennanp ANTENNA_67 (.A(net779));
 sg13g2_antennanp ANTENNA_68 (.A(_1134_));
 sg13g2_antennanp ANTENNA_69 (.A(_1408_));
 sg13g2_antennanp ANTENNA_70 (.A(_1419_));
 sg13g2_antennanp ANTENNA_71 (.A(_1455_));
 sg13g2_antennanp ANTENNA_72 (.A(_1553_));
 sg13g2_antennanp ANTENNA_73 (.A(_1553_));
 sg13g2_antennanp ANTENNA_74 (.A(_1573_));
 sg13g2_antennanp ANTENNA_75 (.A(_1637_));
 sg13g2_antennanp ANTENNA_76 (.A(_1659_));
 sg13g2_antennanp ANTENNA_77 (.A(_1714_));
 sg13g2_antennanp ANTENNA_78 (.A(_1744_));
 sg13g2_antennanp ANTENNA_79 (.A(_1798_));
 sg13g2_antennanp ANTENNA_80 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_81 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_82 (.A(hartinfo_i_18_));
 sg13g2_antennanp ANTENNA_83 (.A(hartinfo_i_19_));
 sg13g2_antennanp ANTENNA_84 (.A(hartinfo_i_26_));
 sg13g2_antennanp ANTENNA_85 (.A(hartinfo_i_5_));
 sg13g2_antennanp ANTENNA_86 (.A(next_dm_addr_i_13_));
 sg13g2_antennanp ANTENNA_87 (.A(next_dm_addr_i_14_));
 sg13g2_antennanp ANTENNA_88 (.A(next_dm_addr_i_19_));
 sg13g2_antennanp ANTENNA_89 (.A(next_dm_addr_i_1_));
 sg13g2_antennanp ANTENNA_90 (.A(next_dm_addr_i_20_));
 sg13g2_antennanp ANTENNA_91 (.A(next_dm_addr_i_28_));
 sg13g2_antennanp ANTENNA_92 (.A(next_dm_addr_i_2_));
 sg13g2_antennanp ANTENNA_93 (.A(next_dm_addr_i_30_));
 sg13g2_antennanp ANTENNA_94 (.A(next_dm_addr_i_3_));
 sg13g2_antennanp ANTENNA_95 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_96 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_97 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_98 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_99 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_100 (.A(slave_addr_i_6_));
 sg13g2_antennanp ANTENNA_101 (.A(_1134_));
 sg13g2_antennanp ANTENNA_102 (.A(_1408_));
 sg13g2_antennanp ANTENNA_103 (.A(_1419_));
 sg13g2_antennanp ANTENNA_104 (.A(_1455_));
 sg13g2_antennanp ANTENNA_105 (.A(_1553_));
 sg13g2_antennanp ANTENNA_106 (.A(_1553_));
 sg13g2_antennanp ANTENNA_107 (.A(_1573_));
 sg13g2_antennanp ANTENNA_108 (.A(_1637_));
 sg13g2_antennanp ANTENNA_109 (.A(_1659_));
 sg13g2_antennanp ANTENNA_110 (.A(_1714_));
 sg13g2_antennanp ANTENNA_111 (.A(_1744_));
 sg13g2_antennanp ANTENNA_112 (.A(_1798_));
 sg13g2_antennanp ANTENNA_113 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_114 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_115 (.A(hartinfo_i_18_));
 sg13g2_antennanp ANTENNA_116 (.A(hartinfo_i_19_));
 sg13g2_antennanp ANTENNA_117 (.A(hartinfo_i_26_));
 sg13g2_antennanp ANTENNA_118 (.A(hartinfo_i_28_));
 sg13g2_antennanp ANTENNA_119 (.A(next_dm_addr_i_13_));
 sg13g2_antennanp ANTENNA_120 (.A(next_dm_addr_i_14_));
 sg13g2_antennanp ANTENNA_121 (.A(next_dm_addr_i_1_));
 sg13g2_antennanp ANTENNA_122 (.A(next_dm_addr_i_20_));
 sg13g2_antennanp ANTENNA_123 (.A(next_dm_addr_i_2_));
 sg13g2_antennanp ANTENNA_124 (.A(next_dm_addr_i_30_));
 sg13g2_antennanp ANTENNA_125 (.A(next_dm_addr_i_3_));
 sg13g2_antennanp ANTENNA_126 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_127 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_128 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_129 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_130 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_131 (.A(_1134_));
 sg13g2_antennanp ANTENNA_132 (.A(_1408_));
 sg13g2_antennanp ANTENNA_133 (.A(_1419_));
 sg13g2_antennanp ANTENNA_134 (.A(_1455_));
 sg13g2_antennanp ANTENNA_135 (.A(_1455_));
 sg13g2_antennanp ANTENNA_136 (.A(_1553_));
 sg13g2_antennanp ANTENNA_137 (.A(_1553_));
 sg13g2_antennanp ANTENNA_138 (.A(_1573_));
 sg13g2_antennanp ANTENNA_139 (.A(_1573_));
 sg13g2_antennanp ANTENNA_140 (.A(_1637_));
 sg13g2_antennanp ANTENNA_141 (.A(_1659_));
 sg13g2_antennanp ANTENNA_142 (.A(_1714_));
 sg13g2_antennanp ANTENNA_143 (.A(_1744_));
 sg13g2_antennanp ANTENNA_144 (.A(_1798_));
 sg13g2_antennanp ANTENNA_145 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_146 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_147 (.A(hartinfo_i_18_));
 sg13g2_antennanp ANTENNA_148 (.A(hartinfo_i_19_));
 sg13g2_antennanp ANTENNA_149 (.A(hartinfo_i_26_));
 sg13g2_antennanp ANTENNA_150 (.A(next_dm_addr_i_13_));
 sg13g2_antennanp ANTENNA_151 (.A(next_dm_addr_i_14_));
 sg13g2_antennanp ANTENNA_152 (.A(next_dm_addr_i_20_));
 sg13g2_antennanp ANTENNA_153 (.A(next_dm_addr_i_2_));
 sg13g2_antennanp ANTENNA_154 (.A(next_dm_addr_i_30_));
 sg13g2_antennanp ANTENNA_155 (.A(next_dm_addr_i_3_));
 sg13g2_antennanp ANTENNA_156 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_157 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_158 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_159 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_160 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_161 (.A(_1134_));
 sg13g2_antennanp ANTENNA_162 (.A(_1408_));
 sg13g2_antennanp ANTENNA_163 (.A(_1419_));
 sg13g2_antennanp ANTENNA_164 (.A(_1455_));
 sg13g2_antennanp ANTENNA_165 (.A(_1455_));
 sg13g2_antennanp ANTENNA_166 (.A(_1553_));
 sg13g2_antennanp ANTENNA_167 (.A(_1553_));
 sg13g2_antennanp ANTENNA_168 (.A(_1573_));
 sg13g2_antennanp ANTENNA_169 (.A(_1637_));
 sg13g2_antennanp ANTENNA_170 (.A(_1659_));
 sg13g2_antennanp ANTENNA_171 (.A(_1714_));
 sg13g2_antennanp ANTENNA_172 (.A(_1744_));
 sg13g2_antennanp ANTENNA_173 (.A(_1798_));
 sg13g2_antennanp ANTENNA_174 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_175 (.A(dmi_req_i_8_));
 sg13g2_antennanp ANTENNA_176 (.A(hartinfo_i_18_));
 sg13g2_antennanp ANTENNA_177 (.A(hartinfo_i_19_));
 sg13g2_antennanp ANTENNA_178 (.A(hartinfo_i_26_));
 sg13g2_antennanp ANTENNA_179 (.A(hartinfo_i_28_));
 sg13g2_antennanp ANTENNA_180 (.A(next_dm_addr_i_13_));
 sg13g2_antennanp ANTENNA_181 (.A(next_dm_addr_i_14_));
 sg13g2_antennanp ANTENNA_182 (.A(next_dm_addr_i_20_));
 sg13g2_antennanp ANTENNA_183 (.A(next_dm_addr_i_2_));
 sg13g2_antennanp ANTENNA_184 (.A(next_dm_addr_i_30_));
 sg13g2_antennanp ANTENNA_185 (.A(next_dm_addr_i_3_));
 sg13g2_antennanp ANTENNA_186 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_187 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_188 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_189 (.A(slave_addr_i_11_));
 sg13g2_antennanp ANTENNA_190 (.A(slave_addr_i_11_));
 sg13g2_fill_8 FILLER_0_0 ();
 sg13g2_fill_8 FILLER_0_8 ();
 sg13g2_fill_8 FILLER_0_16 ();
 sg13g2_fill_8 FILLER_0_24 ();
 sg13g2_fill_8 FILLER_0_32 ();
 sg13g2_fill_8 FILLER_0_40 ();
 sg13g2_fill_8 FILLER_0_48 ();
 sg13g2_fill_8 FILLER_0_56 ();
 sg13g2_fill_8 FILLER_0_64 ();
 sg13g2_fill_8 FILLER_0_72 ();
 sg13g2_fill_8 FILLER_0_80 ();
 sg13g2_fill_8 FILLER_0_88 ();
 sg13g2_fill_8 FILLER_0_96 ();
 sg13g2_fill_8 FILLER_0_104 ();
 sg13g2_fill_8 FILLER_0_112 ();
 sg13g2_fill_8 FILLER_0_120 ();
 sg13g2_fill_8 FILLER_0_128 ();
 sg13g2_fill_8 FILLER_0_136 ();
 sg13g2_fill_8 FILLER_0_144 ();
 sg13g2_fill_8 FILLER_0_152 ();
 sg13g2_fill_8 FILLER_0_160 ();
 sg13g2_fill_8 FILLER_0_168 ();
 sg13g2_fill_8 FILLER_0_176 ();
 sg13g2_fill_8 FILLER_0_184 ();
 sg13g2_fill_8 FILLER_0_192 ();
 sg13g2_fill_8 FILLER_0_200 ();
 sg13g2_fill_8 FILLER_0_208 ();
 sg13g2_fill_8 FILLER_0_216 ();
 sg13g2_fill_8 FILLER_0_224 ();
 sg13g2_fill_8 FILLER_0_232 ();
 sg13g2_fill_8 FILLER_0_240 ();
 sg13g2_fill_8 FILLER_0_248 ();
 sg13g2_fill_8 FILLER_0_256 ();
 sg13g2_fill_8 FILLER_0_264 ();
 sg13g2_fill_8 FILLER_0_272 ();
 sg13g2_fill_8 FILLER_0_280 ();
 sg13g2_fill_8 FILLER_0_288 ();
 sg13g2_fill_8 FILLER_0_296 ();
 sg13g2_fill_8 FILLER_0_304 ();
 sg13g2_fill_8 FILLER_0_312 ();
 sg13g2_fill_8 FILLER_0_320 ();
 sg13g2_fill_8 FILLER_0_328 ();
 sg13g2_fill_8 FILLER_0_336 ();
 sg13g2_fill_8 FILLER_0_344 ();
 sg13g2_fill_8 FILLER_0_352 ();
 sg13g2_fill_8 FILLER_0_360 ();
 sg13g2_fill_8 FILLER_0_368 ();
 sg13g2_fill_8 FILLER_0_376 ();
 sg13g2_fill_8 FILLER_0_384 ();
 sg13g2_fill_8 FILLER_0_392 ();
 sg13g2_fill_8 FILLER_0_400 ();
 sg13g2_fill_8 FILLER_0_408 ();
 sg13g2_fill_8 FILLER_0_416 ();
 sg13g2_fill_8 FILLER_0_424 ();
 sg13g2_fill_8 FILLER_0_432 ();
 sg13g2_fill_8 FILLER_0_440 ();
 sg13g2_fill_8 FILLER_0_448 ();
 sg13g2_fill_8 FILLER_0_456 ();
 sg13g2_fill_8 FILLER_0_464 ();
 sg13g2_fill_8 FILLER_0_472 ();
 sg13g2_fill_8 FILLER_0_480 ();
 sg13g2_fill_8 FILLER_0_488 ();
 sg13g2_fill_8 FILLER_0_496 ();
 sg13g2_fill_8 FILLER_0_504 ();
 sg13g2_fill_8 FILLER_0_512 ();
 sg13g2_fill_8 FILLER_0_520 ();
 sg13g2_fill_8 FILLER_0_528 ();
 sg13g2_fill_8 FILLER_0_536 ();
 sg13g2_fill_8 FILLER_0_544 ();
 sg13g2_fill_8 FILLER_0_552 ();
 sg13g2_fill_8 FILLER_0_560 ();
 sg13g2_fill_8 FILLER_0_568 ();
 sg13g2_fill_8 FILLER_0_576 ();
 sg13g2_fill_8 FILLER_0_584 ();
 sg13g2_fill_8 FILLER_0_592 ();
 sg13g2_fill_8 FILLER_0_600 ();
 sg13g2_fill_8 FILLER_0_608 ();
 sg13g2_fill_8 FILLER_0_616 ();
 sg13g2_fill_8 FILLER_0_624 ();
 sg13g2_fill_8 FILLER_0_632 ();
 sg13g2_fill_8 FILLER_0_640 ();
 sg13g2_fill_8 FILLER_0_648 ();
 sg13g2_fill_8 FILLER_0_656 ();
 sg13g2_fill_8 FILLER_0_664 ();
 sg13g2_fill_8 FILLER_0_672 ();
 sg13g2_fill_8 FILLER_0_680 ();
 sg13g2_fill_8 FILLER_0_688 ();
 sg13g2_fill_8 FILLER_0_696 ();
 sg13g2_fill_8 FILLER_0_704 ();
 sg13g2_fill_8 FILLER_0_712 ();
 sg13g2_fill_8 FILLER_0_720 ();
 sg13g2_fill_8 FILLER_0_728 ();
 sg13g2_fill_8 FILLER_0_736 ();
 sg13g2_fill_8 FILLER_0_744 ();
 sg13g2_fill_8 FILLER_0_752 ();
 sg13g2_fill_8 FILLER_0_760 ();
 sg13g2_fill_8 FILLER_0_768 ();
 sg13g2_fill_8 FILLER_0_776 ();
 sg13g2_fill_8 FILLER_0_784 ();
 sg13g2_fill_8 FILLER_0_792 ();
 sg13g2_fill_8 FILLER_0_800 ();
 sg13g2_fill_8 FILLER_0_808 ();
 sg13g2_fill_8 FILLER_0_816 ();
 sg13g2_fill_8 FILLER_0_824 ();
 sg13g2_fill_8 FILLER_0_832 ();
 sg13g2_fill_8 FILLER_0_840 ();
 sg13g2_fill_8 FILLER_0_848 ();
 sg13g2_fill_8 FILLER_0_856 ();
 sg13g2_fill_8 FILLER_0_864 ();
 sg13g2_fill_8 FILLER_0_872 ();
 sg13g2_fill_8 FILLER_0_880 ();
 sg13g2_fill_8 FILLER_0_888 ();
 sg13g2_fill_8 FILLER_0_896 ();
 sg13g2_fill_8 FILLER_0_904 ();
 sg13g2_fill_8 FILLER_0_912 ();
 sg13g2_fill_8 FILLER_0_920 ();
 sg13g2_fill_8 FILLER_0_928 ();
 sg13g2_fill_8 FILLER_0_936 ();
 sg13g2_fill_8 FILLER_0_944 ();
 sg13g2_fill_8 FILLER_0_952 ();
 sg13g2_fill_8 FILLER_0_960 ();
 sg13g2_fill_8 FILLER_0_968 ();
 sg13g2_fill_8 FILLER_0_976 ();
 sg13g2_fill_8 FILLER_0_984 ();
 sg13g2_fill_8 FILLER_0_992 ();
 sg13g2_fill_8 FILLER_0_1000 ();
 sg13g2_fill_8 FILLER_0_1008 ();
 sg13g2_fill_8 FILLER_0_1016 ();
 sg13g2_fill_8 FILLER_0_1024 ();
 sg13g2_fill_8 FILLER_0_1032 ();
 sg13g2_fill_8 FILLER_0_1040 ();
 sg13g2_fill_8 FILLER_0_1048 ();
 sg13g2_fill_8 FILLER_0_1056 ();
 sg13g2_fill_8 FILLER_0_1064 ();
 sg13g2_fill_8 FILLER_0_1072 ();
 sg13g2_fill_8 FILLER_0_1080 ();
 sg13g2_fill_8 FILLER_0_1088 ();
 sg13g2_fill_8 FILLER_0_1096 ();
 sg13g2_fill_8 FILLER_0_1104 ();
 sg13g2_fill_8 FILLER_0_1112 ();
 sg13g2_fill_8 FILLER_0_1120 ();
 sg13g2_fill_8 FILLER_0_1128 ();
 sg13g2_fill_8 FILLER_0_1136 ();
 sg13g2_fill_8 FILLER_0_1144 ();
 sg13g2_fill_8 FILLER_0_1152 ();
 sg13g2_fill_4 FILLER_0_1160 ();
 sg13g2_fill_2 FILLER_0_1164 ();
 sg13g2_fill_8 FILLER_1_0 ();
 sg13g2_fill_8 FILLER_1_8 ();
 sg13g2_fill_8 FILLER_1_16 ();
 sg13g2_fill_8 FILLER_1_24 ();
 sg13g2_fill_8 FILLER_1_32 ();
 sg13g2_fill_8 FILLER_1_40 ();
 sg13g2_fill_8 FILLER_1_48 ();
 sg13g2_fill_8 FILLER_1_56 ();
 sg13g2_fill_8 FILLER_1_64 ();
 sg13g2_fill_8 FILLER_1_72 ();
 sg13g2_fill_8 FILLER_1_80 ();
 sg13g2_fill_8 FILLER_1_88 ();
 sg13g2_fill_8 FILLER_1_96 ();
 sg13g2_fill_8 FILLER_1_104 ();
 sg13g2_fill_8 FILLER_1_112 ();
 sg13g2_fill_8 FILLER_1_120 ();
 sg13g2_fill_8 FILLER_1_128 ();
 sg13g2_fill_8 FILLER_1_136 ();
 sg13g2_fill_8 FILLER_1_144 ();
 sg13g2_fill_8 FILLER_1_152 ();
 sg13g2_fill_8 FILLER_1_160 ();
 sg13g2_fill_8 FILLER_1_168 ();
 sg13g2_fill_8 FILLER_1_176 ();
 sg13g2_fill_8 FILLER_1_184 ();
 sg13g2_fill_8 FILLER_1_192 ();
 sg13g2_fill_8 FILLER_1_200 ();
 sg13g2_fill_8 FILLER_1_208 ();
 sg13g2_fill_8 FILLER_1_216 ();
 sg13g2_fill_8 FILLER_1_224 ();
 sg13g2_fill_8 FILLER_1_232 ();
 sg13g2_fill_8 FILLER_1_240 ();
 sg13g2_fill_8 FILLER_1_248 ();
 sg13g2_fill_8 FILLER_1_256 ();
 sg13g2_fill_8 FILLER_1_264 ();
 sg13g2_fill_8 FILLER_1_272 ();
 sg13g2_fill_8 FILLER_1_280 ();
 sg13g2_fill_8 FILLER_1_288 ();
 sg13g2_fill_8 FILLER_1_296 ();
 sg13g2_fill_8 FILLER_1_304 ();
 sg13g2_fill_8 FILLER_1_312 ();
 sg13g2_fill_8 FILLER_1_320 ();
 sg13g2_fill_8 FILLER_1_328 ();
 sg13g2_fill_8 FILLER_1_336 ();
 sg13g2_fill_8 FILLER_1_344 ();
 sg13g2_fill_8 FILLER_1_352 ();
 sg13g2_fill_8 FILLER_1_360 ();
 sg13g2_fill_8 FILLER_1_368 ();
 sg13g2_fill_8 FILLER_1_376 ();
 sg13g2_fill_8 FILLER_1_384 ();
 sg13g2_fill_8 FILLER_1_392 ();
 sg13g2_fill_8 FILLER_1_400 ();
 sg13g2_fill_8 FILLER_1_408 ();
 sg13g2_fill_8 FILLER_1_416 ();
 sg13g2_fill_8 FILLER_1_424 ();
 sg13g2_fill_8 FILLER_1_432 ();
 sg13g2_fill_8 FILLER_1_440 ();
 sg13g2_fill_8 FILLER_1_448 ();
 sg13g2_fill_8 FILLER_1_456 ();
 sg13g2_fill_8 FILLER_1_464 ();
 sg13g2_fill_8 FILLER_1_472 ();
 sg13g2_fill_8 FILLER_1_480 ();
 sg13g2_fill_8 FILLER_1_488 ();
 sg13g2_fill_8 FILLER_1_496 ();
 sg13g2_fill_8 FILLER_1_504 ();
 sg13g2_fill_8 FILLER_1_512 ();
 sg13g2_fill_8 FILLER_1_520 ();
 sg13g2_fill_8 FILLER_1_528 ();
 sg13g2_fill_8 FILLER_1_536 ();
 sg13g2_fill_8 FILLER_1_544 ();
 sg13g2_fill_8 FILLER_1_552 ();
 sg13g2_fill_8 FILLER_1_560 ();
 sg13g2_fill_8 FILLER_1_568 ();
 sg13g2_fill_8 FILLER_1_576 ();
 sg13g2_fill_8 FILLER_1_584 ();
 sg13g2_fill_8 FILLER_1_592 ();
 sg13g2_fill_8 FILLER_1_600 ();
 sg13g2_fill_8 FILLER_1_608 ();
 sg13g2_fill_8 FILLER_1_616 ();
 sg13g2_fill_8 FILLER_1_624 ();
 sg13g2_fill_8 FILLER_1_632 ();
 sg13g2_fill_8 FILLER_1_640 ();
 sg13g2_fill_8 FILLER_1_648 ();
 sg13g2_fill_8 FILLER_1_656 ();
 sg13g2_fill_8 FILLER_1_664 ();
 sg13g2_fill_8 FILLER_1_672 ();
 sg13g2_fill_8 FILLER_1_680 ();
 sg13g2_fill_8 FILLER_1_688 ();
 sg13g2_fill_8 FILLER_1_696 ();
 sg13g2_fill_8 FILLER_1_704 ();
 sg13g2_fill_8 FILLER_1_712 ();
 sg13g2_fill_8 FILLER_1_720 ();
 sg13g2_fill_8 FILLER_1_728 ();
 sg13g2_fill_8 FILLER_1_736 ();
 sg13g2_fill_8 FILLER_1_744 ();
 sg13g2_fill_8 FILLER_1_752 ();
 sg13g2_fill_8 FILLER_1_760 ();
 sg13g2_fill_8 FILLER_1_768 ();
 sg13g2_fill_8 FILLER_1_776 ();
 sg13g2_fill_8 FILLER_1_784 ();
 sg13g2_fill_8 FILLER_1_792 ();
 sg13g2_fill_8 FILLER_1_800 ();
 sg13g2_fill_8 FILLER_1_808 ();
 sg13g2_fill_8 FILLER_1_816 ();
 sg13g2_fill_8 FILLER_1_824 ();
 sg13g2_fill_8 FILLER_1_832 ();
 sg13g2_fill_8 FILLER_1_840 ();
 sg13g2_fill_8 FILLER_1_848 ();
 sg13g2_fill_8 FILLER_1_856 ();
 sg13g2_fill_8 FILLER_1_864 ();
 sg13g2_fill_8 FILLER_1_872 ();
 sg13g2_fill_8 FILLER_1_880 ();
 sg13g2_fill_8 FILLER_1_888 ();
 sg13g2_fill_8 FILLER_1_896 ();
 sg13g2_fill_8 FILLER_1_904 ();
 sg13g2_fill_8 FILLER_1_912 ();
 sg13g2_fill_8 FILLER_1_920 ();
 sg13g2_fill_8 FILLER_1_928 ();
 sg13g2_fill_8 FILLER_1_936 ();
 sg13g2_fill_8 FILLER_1_944 ();
 sg13g2_fill_8 FILLER_1_952 ();
 sg13g2_fill_8 FILLER_1_960 ();
 sg13g2_fill_8 FILLER_1_968 ();
 sg13g2_fill_8 FILLER_1_976 ();
 sg13g2_fill_8 FILLER_1_984 ();
 sg13g2_fill_8 FILLER_1_992 ();
 sg13g2_fill_8 FILLER_1_1000 ();
 sg13g2_fill_8 FILLER_1_1008 ();
 sg13g2_fill_8 FILLER_1_1016 ();
 sg13g2_fill_8 FILLER_1_1024 ();
 sg13g2_fill_8 FILLER_1_1032 ();
 sg13g2_fill_8 FILLER_1_1040 ();
 sg13g2_fill_8 FILLER_1_1048 ();
 sg13g2_fill_8 FILLER_1_1056 ();
 sg13g2_fill_8 FILLER_1_1064 ();
 sg13g2_fill_8 FILLER_1_1072 ();
 sg13g2_fill_8 FILLER_1_1080 ();
 sg13g2_fill_8 FILLER_1_1088 ();
 sg13g2_fill_8 FILLER_1_1096 ();
 sg13g2_fill_8 FILLER_1_1104 ();
 sg13g2_fill_8 FILLER_1_1112 ();
 sg13g2_fill_8 FILLER_1_1120 ();
 sg13g2_fill_8 FILLER_1_1128 ();
 sg13g2_fill_8 FILLER_1_1136 ();
 sg13g2_fill_8 FILLER_1_1144 ();
 sg13g2_fill_8 FILLER_1_1152 ();
 sg13g2_fill_4 FILLER_1_1160 ();
 sg13g2_fill_2 FILLER_1_1164 ();
 sg13g2_fill_8 FILLER_2_0 ();
 sg13g2_fill_8 FILLER_2_8 ();
 sg13g2_fill_8 FILLER_2_16 ();
 sg13g2_fill_8 FILLER_2_24 ();
 sg13g2_fill_8 FILLER_2_32 ();
 sg13g2_fill_8 FILLER_2_40 ();
 sg13g2_fill_8 FILLER_2_48 ();
 sg13g2_fill_8 FILLER_2_56 ();
 sg13g2_fill_8 FILLER_2_64 ();
 sg13g2_fill_8 FILLER_2_72 ();
 sg13g2_fill_8 FILLER_2_80 ();
 sg13g2_fill_8 FILLER_2_88 ();
 sg13g2_fill_8 FILLER_2_96 ();
 sg13g2_fill_8 FILLER_2_104 ();
 sg13g2_fill_8 FILLER_2_112 ();
 sg13g2_fill_8 FILLER_2_120 ();
 sg13g2_fill_8 FILLER_2_128 ();
 sg13g2_fill_8 FILLER_2_136 ();
 sg13g2_fill_8 FILLER_2_144 ();
 sg13g2_fill_8 FILLER_2_152 ();
 sg13g2_fill_8 FILLER_2_160 ();
 sg13g2_fill_8 FILLER_2_168 ();
 sg13g2_fill_8 FILLER_2_176 ();
 sg13g2_fill_8 FILLER_2_184 ();
 sg13g2_fill_8 FILLER_2_192 ();
 sg13g2_fill_8 FILLER_2_200 ();
 sg13g2_fill_8 FILLER_2_208 ();
 sg13g2_fill_8 FILLER_2_216 ();
 sg13g2_fill_8 FILLER_2_224 ();
 sg13g2_fill_8 FILLER_2_232 ();
 sg13g2_fill_8 FILLER_2_240 ();
 sg13g2_fill_8 FILLER_2_248 ();
 sg13g2_fill_8 FILLER_2_256 ();
 sg13g2_fill_8 FILLER_2_264 ();
 sg13g2_fill_8 FILLER_2_272 ();
 sg13g2_fill_8 FILLER_2_280 ();
 sg13g2_fill_8 FILLER_2_288 ();
 sg13g2_fill_8 FILLER_2_296 ();
 sg13g2_fill_8 FILLER_2_304 ();
 sg13g2_fill_8 FILLER_2_312 ();
 sg13g2_fill_8 FILLER_2_320 ();
 sg13g2_fill_8 FILLER_2_328 ();
 sg13g2_fill_8 FILLER_2_336 ();
 sg13g2_fill_8 FILLER_2_344 ();
 sg13g2_fill_8 FILLER_2_352 ();
 sg13g2_fill_8 FILLER_2_360 ();
 sg13g2_fill_8 FILLER_2_368 ();
 sg13g2_fill_8 FILLER_2_376 ();
 sg13g2_fill_8 FILLER_2_384 ();
 sg13g2_fill_8 FILLER_2_392 ();
 sg13g2_fill_8 FILLER_2_400 ();
 sg13g2_fill_8 FILLER_2_408 ();
 sg13g2_fill_8 FILLER_2_416 ();
 sg13g2_fill_8 FILLER_2_424 ();
 sg13g2_fill_8 FILLER_2_432 ();
 sg13g2_fill_8 FILLER_2_440 ();
 sg13g2_fill_8 FILLER_2_448 ();
 sg13g2_fill_8 FILLER_2_456 ();
 sg13g2_fill_8 FILLER_2_464 ();
 sg13g2_fill_8 FILLER_2_472 ();
 sg13g2_fill_8 FILLER_2_480 ();
 sg13g2_fill_8 FILLER_2_488 ();
 sg13g2_fill_8 FILLER_2_496 ();
 sg13g2_fill_8 FILLER_2_504 ();
 sg13g2_fill_8 FILLER_2_512 ();
 sg13g2_fill_8 FILLER_2_520 ();
 sg13g2_fill_8 FILLER_2_528 ();
 sg13g2_fill_8 FILLER_2_536 ();
 sg13g2_fill_8 FILLER_2_544 ();
 sg13g2_fill_8 FILLER_2_552 ();
 sg13g2_fill_8 FILLER_2_560 ();
 sg13g2_fill_8 FILLER_2_568 ();
 sg13g2_fill_8 FILLER_2_576 ();
 sg13g2_fill_8 FILLER_2_584 ();
 sg13g2_fill_8 FILLER_2_592 ();
 sg13g2_fill_8 FILLER_2_600 ();
 sg13g2_fill_8 FILLER_2_608 ();
 sg13g2_fill_8 FILLER_2_616 ();
 sg13g2_fill_8 FILLER_2_624 ();
 sg13g2_fill_8 FILLER_2_632 ();
 sg13g2_fill_8 FILLER_2_640 ();
 sg13g2_fill_8 FILLER_2_648 ();
 sg13g2_fill_8 FILLER_2_656 ();
 sg13g2_fill_8 FILLER_2_664 ();
 sg13g2_fill_8 FILLER_2_672 ();
 sg13g2_fill_8 FILLER_2_680 ();
 sg13g2_fill_8 FILLER_2_688 ();
 sg13g2_fill_8 FILLER_2_696 ();
 sg13g2_fill_8 FILLER_2_704 ();
 sg13g2_fill_8 FILLER_2_712 ();
 sg13g2_fill_8 FILLER_2_720 ();
 sg13g2_fill_8 FILLER_2_728 ();
 sg13g2_fill_8 FILLER_2_736 ();
 sg13g2_fill_8 FILLER_2_744 ();
 sg13g2_fill_8 FILLER_2_752 ();
 sg13g2_fill_8 FILLER_2_760 ();
 sg13g2_fill_8 FILLER_2_768 ();
 sg13g2_fill_8 FILLER_2_776 ();
 sg13g2_fill_8 FILLER_2_784 ();
 sg13g2_fill_8 FILLER_2_792 ();
 sg13g2_fill_8 FILLER_2_800 ();
 sg13g2_fill_8 FILLER_2_808 ();
 sg13g2_fill_8 FILLER_2_816 ();
 sg13g2_fill_8 FILLER_2_824 ();
 sg13g2_fill_8 FILLER_2_832 ();
 sg13g2_fill_8 FILLER_2_840 ();
 sg13g2_fill_8 FILLER_2_848 ();
 sg13g2_fill_8 FILLER_2_856 ();
 sg13g2_fill_8 FILLER_2_864 ();
 sg13g2_fill_8 FILLER_2_872 ();
 sg13g2_fill_8 FILLER_2_880 ();
 sg13g2_fill_8 FILLER_2_888 ();
 sg13g2_fill_8 FILLER_2_896 ();
 sg13g2_fill_8 FILLER_2_904 ();
 sg13g2_fill_8 FILLER_2_912 ();
 sg13g2_fill_8 FILLER_2_920 ();
 sg13g2_fill_8 FILLER_2_928 ();
 sg13g2_fill_8 FILLER_2_936 ();
 sg13g2_fill_8 FILLER_2_944 ();
 sg13g2_fill_8 FILLER_2_952 ();
 sg13g2_fill_8 FILLER_2_960 ();
 sg13g2_fill_8 FILLER_2_968 ();
 sg13g2_fill_8 FILLER_2_976 ();
 sg13g2_fill_8 FILLER_2_984 ();
 sg13g2_fill_8 FILLER_2_992 ();
 sg13g2_fill_8 FILLER_2_1000 ();
 sg13g2_fill_8 FILLER_2_1008 ();
 sg13g2_fill_8 FILLER_2_1016 ();
 sg13g2_fill_8 FILLER_2_1024 ();
 sg13g2_fill_8 FILLER_2_1032 ();
 sg13g2_fill_8 FILLER_2_1040 ();
 sg13g2_fill_8 FILLER_2_1048 ();
 sg13g2_fill_8 FILLER_2_1056 ();
 sg13g2_fill_8 FILLER_2_1064 ();
 sg13g2_fill_8 FILLER_2_1072 ();
 sg13g2_fill_8 FILLER_2_1080 ();
 sg13g2_fill_8 FILLER_2_1088 ();
 sg13g2_fill_8 FILLER_2_1096 ();
 sg13g2_fill_8 FILLER_2_1104 ();
 sg13g2_fill_8 FILLER_2_1112 ();
 sg13g2_fill_8 FILLER_2_1120 ();
 sg13g2_fill_8 FILLER_2_1128 ();
 sg13g2_fill_8 FILLER_2_1136 ();
 sg13g2_fill_8 FILLER_2_1144 ();
 sg13g2_fill_8 FILLER_2_1152 ();
 sg13g2_fill_4 FILLER_2_1160 ();
 sg13g2_fill_2 FILLER_2_1164 ();
 sg13g2_fill_8 FILLER_3_0 ();
 sg13g2_fill_8 FILLER_3_8 ();
 sg13g2_fill_8 FILLER_3_16 ();
 sg13g2_fill_8 FILLER_3_24 ();
 sg13g2_fill_8 FILLER_3_32 ();
 sg13g2_fill_8 FILLER_3_40 ();
 sg13g2_fill_8 FILLER_3_48 ();
 sg13g2_fill_8 FILLER_3_56 ();
 sg13g2_fill_8 FILLER_3_64 ();
 sg13g2_fill_8 FILLER_3_72 ();
 sg13g2_fill_8 FILLER_3_80 ();
 sg13g2_fill_8 FILLER_3_88 ();
 sg13g2_fill_8 FILLER_3_96 ();
 sg13g2_fill_8 FILLER_3_104 ();
 sg13g2_fill_8 FILLER_3_112 ();
 sg13g2_fill_8 FILLER_3_120 ();
 sg13g2_fill_8 FILLER_3_128 ();
 sg13g2_fill_8 FILLER_3_136 ();
 sg13g2_fill_8 FILLER_3_144 ();
 sg13g2_fill_8 FILLER_3_152 ();
 sg13g2_fill_8 FILLER_3_160 ();
 sg13g2_fill_8 FILLER_3_168 ();
 sg13g2_fill_8 FILLER_3_176 ();
 sg13g2_fill_8 FILLER_3_184 ();
 sg13g2_fill_8 FILLER_3_192 ();
 sg13g2_fill_8 FILLER_3_200 ();
 sg13g2_fill_8 FILLER_3_208 ();
 sg13g2_fill_8 FILLER_3_216 ();
 sg13g2_fill_8 FILLER_3_224 ();
 sg13g2_fill_8 FILLER_3_232 ();
 sg13g2_fill_8 FILLER_3_240 ();
 sg13g2_fill_8 FILLER_3_248 ();
 sg13g2_fill_8 FILLER_3_256 ();
 sg13g2_fill_8 FILLER_3_264 ();
 sg13g2_fill_8 FILLER_3_272 ();
 sg13g2_fill_8 FILLER_3_280 ();
 sg13g2_fill_8 FILLER_3_288 ();
 sg13g2_fill_8 FILLER_3_296 ();
 sg13g2_fill_8 FILLER_3_304 ();
 sg13g2_fill_8 FILLER_3_312 ();
 sg13g2_fill_8 FILLER_3_320 ();
 sg13g2_fill_8 FILLER_3_328 ();
 sg13g2_fill_8 FILLER_3_336 ();
 sg13g2_fill_8 FILLER_3_344 ();
 sg13g2_fill_8 FILLER_3_352 ();
 sg13g2_fill_8 FILLER_3_360 ();
 sg13g2_fill_8 FILLER_3_368 ();
 sg13g2_fill_8 FILLER_3_376 ();
 sg13g2_fill_8 FILLER_3_384 ();
 sg13g2_fill_8 FILLER_3_392 ();
 sg13g2_fill_8 FILLER_3_400 ();
 sg13g2_fill_8 FILLER_3_408 ();
 sg13g2_fill_8 FILLER_3_416 ();
 sg13g2_fill_8 FILLER_3_424 ();
 sg13g2_fill_8 FILLER_3_432 ();
 sg13g2_fill_8 FILLER_3_440 ();
 sg13g2_fill_8 FILLER_3_448 ();
 sg13g2_fill_8 FILLER_3_456 ();
 sg13g2_fill_8 FILLER_3_464 ();
 sg13g2_fill_8 FILLER_3_472 ();
 sg13g2_fill_8 FILLER_3_480 ();
 sg13g2_fill_8 FILLER_3_488 ();
 sg13g2_fill_8 FILLER_3_496 ();
 sg13g2_fill_8 FILLER_3_504 ();
 sg13g2_fill_8 FILLER_3_512 ();
 sg13g2_fill_8 FILLER_3_520 ();
 sg13g2_fill_8 FILLER_3_528 ();
 sg13g2_fill_8 FILLER_3_536 ();
 sg13g2_fill_8 FILLER_3_544 ();
 sg13g2_fill_8 FILLER_3_552 ();
 sg13g2_fill_8 FILLER_3_560 ();
 sg13g2_fill_8 FILLER_3_568 ();
 sg13g2_fill_8 FILLER_3_576 ();
 sg13g2_fill_8 FILLER_3_584 ();
 sg13g2_fill_8 FILLER_3_592 ();
 sg13g2_fill_8 FILLER_3_600 ();
 sg13g2_fill_8 FILLER_3_608 ();
 sg13g2_fill_8 FILLER_3_616 ();
 sg13g2_fill_8 FILLER_3_624 ();
 sg13g2_fill_8 FILLER_3_632 ();
 sg13g2_fill_8 FILLER_3_640 ();
 sg13g2_fill_8 FILLER_3_648 ();
 sg13g2_fill_8 FILLER_3_656 ();
 sg13g2_fill_8 FILLER_3_664 ();
 sg13g2_fill_8 FILLER_3_672 ();
 sg13g2_fill_8 FILLER_3_680 ();
 sg13g2_fill_8 FILLER_3_688 ();
 sg13g2_fill_8 FILLER_3_696 ();
 sg13g2_fill_8 FILLER_3_704 ();
 sg13g2_fill_8 FILLER_3_712 ();
 sg13g2_fill_8 FILLER_3_720 ();
 sg13g2_fill_8 FILLER_3_728 ();
 sg13g2_fill_8 FILLER_3_736 ();
 sg13g2_fill_8 FILLER_3_744 ();
 sg13g2_fill_8 FILLER_3_752 ();
 sg13g2_fill_8 FILLER_3_760 ();
 sg13g2_fill_8 FILLER_3_768 ();
 sg13g2_fill_8 FILLER_3_776 ();
 sg13g2_fill_8 FILLER_3_784 ();
 sg13g2_fill_8 FILLER_3_792 ();
 sg13g2_fill_8 FILLER_3_800 ();
 sg13g2_fill_8 FILLER_3_808 ();
 sg13g2_fill_8 FILLER_3_816 ();
 sg13g2_fill_8 FILLER_3_824 ();
 sg13g2_fill_8 FILLER_3_832 ();
 sg13g2_fill_8 FILLER_3_840 ();
 sg13g2_fill_8 FILLER_3_848 ();
 sg13g2_fill_8 FILLER_3_856 ();
 sg13g2_fill_8 FILLER_3_864 ();
 sg13g2_fill_8 FILLER_3_872 ();
 sg13g2_fill_8 FILLER_3_880 ();
 sg13g2_fill_8 FILLER_3_888 ();
 sg13g2_fill_8 FILLER_3_896 ();
 sg13g2_fill_8 FILLER_3_904 ();
 sg13g2_fill_8 FILLER_3_912 ();
 sg13g2_fill_8 FILLER_3_920 ();
 sg13g2_fill_8 FILLER_3_928 ();
 sg13g2_fill_8 FILLER_3_936 ();
 sg13g2_fill_8 FILLER_3_944 ();
 sg13g2_fill_8 FILLER_3_952 ();
 sg13g2_fill_8 FILLER_3_960 ();
 sg13g2_fill_8 FILLER_3_968 ();
 sg13g2_fill_8 FILLER_3_976 ();
 sg13g2_fill_8 FILLER_3_984 ();
 sg13g2_fill_8 FILLER_3_992 ();
 sg13g2_fill_8 FILLER_3_1000 ();
 sg13g2_fill_8 FILLER_3_1008 ();
 sg13g2_fill_8 FILLER_3_1016 ();
 sg13g2_fill_8 FILLER_3_1024 ();
 sg13g2_fill_8 FILLER_3_1032 ();
 sg13g2_fill_8 FILLER_3_1040 ();
 sg13g2_fill_8 FILLER_3_1048 ();
 sg13g2_fill_8 FILLER_3_1056 ();
 sg13g2_fill_8 FILLER_3_1064 ();
 sg13g2_fill_8 FILLER_3_1072 ();
 sg13g2_fill_8 FILLER_3_1080 ();
 sg13g2_fill_8 FILLER_3_1088 ();
 sg13g2_fill_8 FILLER_3_1096 ();
 sg13g2_fill_8 FILLER_3_1104 ();
 sg13g2_fill_8 FILLER_3_1112 ();
 sg13g2_fill_8 FILLER_3_1120 ();
 sg13g2_fill_8 FILLER_3_1128 ();
 sg13g2_fill_8 FILLER_3_1136 ();
 sg13g2_fill_8 FILLER_3_1144 ();
 sg13g2_fill_8 FILLER_3_1152 ();
 sg13g2_fill_4 FILLER_3_1160 ();
 sg13g2_fill_2 FILLER_3_1164 ();
 sg13g2_fill_8 FILLER_4_0 ();
 sg13g2_fill_8 FILLER_4_8 ();
 sg13g2_fill_8 FILLER_4_16 ();
 sg13g2_fill_8 FILLER_4_24 ();
 sg13g2_fill_8 FILLER_4_32 ();
 sg13g2_fill_8 FILLER_4_40 ();
 sg13g2_fill_8 FILLER_4_48 ();
 sg13g2_fill_8 FILLER_4_56 ();
 sg13g2_fill_8 FILLER_4_64 ();
 sg13g2_fill_8 FILLER_4_72 ();
 sg13g2_fill_8 FILLER_4_80 ();
 sg13g2_fill_8 FILLER_4_88 ();
 sg13g2_fill_8 FILLER_4_96 ();
 sg13g2_fill_8 FILLER_4_104 ();
 sg13g2_fill_8 FILLER_4_112 ();
 sg13g2_fill_8 FILLER_4_120 ();
 sg13g2_fill_8 FILLER_4_128 ();
 sg13g2_fill_8 FILLER_4_136 ();
 sg13g2_fill_8 FILLER_4_144 ();
 sg13g2_fill_8 FILLER_4_152 ();
 sg13g2_fill_8 FILLER_4_160 ();
 sg13g2_fill_8 FILLER_4_168 ();
 sg13g2_fill_8 FILLER_4_176 ();
 sg13g2_fill_8 FILLER_4_184 ();
 sg13g2_fill_8 FILLER_4_192 ();
 sg13g2_fill_8 FILLER_4_200 ();
 sg13g2_fill_8 FILLER_4_208 ();
 sg13g2_fill_8 FILLER_4_216 ();
 sg13g2_fill_8 FILLER_4_224 ();
 sg13g2_fill_8 FILLER_4_232 ();
 sg13g2_fill_8 FILLER_4_240 ();
 sg13g2_fill_8 FILLER_4_248 ();
 sg13g2_fill_8 FILLER_4_256 ();
 sg13g2_fill_8 FILLER_4_264 ();
 sg13g2_fill_8 FILLER_4_272 ();
 sg13g2_fill_8 FILLER_4_280 ();
 sg13g2_fill_8 FILLER_4_288 ();
 sg13g2_fill_8 FILLER_4_296 ();
 sg13g2_fill_8 FILLER_4_304 ();
 sg13g2_fill_8 FILLER_4_312 ();
 sg13g2_fill_8 FILLER_4_320 ();
 sg13g2_fill_8 FILLER_4_328 ();
 sg13g2_fill_8 FILLER_4_336 ();
 sg13g2_fill_8 FILLER_4_344 ();
 sg13g2_fill_8 FILLER_4_352 ();
 sg13g2_fill_8 FILLER_4_360 ();
 sg13g2_fill_8 FILLER_4_368 ();
 sg13g2_fill_8 FILLER_4_376 ();
 sg13g2_fill_8 FILLER_4_384 ();
 sg13g2_fill_8 FILLER_4_392 ();
 sg13g2_fill_8 FILLER_4_400 ();
 sg13g2_fill_8 FILLER_4_408 ();
 sg13g2_fill_8 FILLER_4_416 ();
 sg13g2_fill_8 FILLER_4_424 ();
 sg13g2_fill_8 FILLER_4_432 ();
 sg13g2_fill_8 FILLER_4_440 ();
 sg13g2_fill_8 FILLER_4_448 ();
 sg13g2_fill_8 FILLER_4_456 ();
 sg13g2_fill_8 FILLER_4_464 ();
 sg13g2_fill_8 FILLER_4_472 ();
 sg13g2_fill_8 FILLER_4_480 ();
 sg13g2_fill_8 FILLER_4_488 ();
 sg13g2_fill_8 FILLER_4_496 ();
 sg13g2_fill_8 FILLER_4_504 ();
 sg13g2_fill_8 FILLER_4_512 ();
 sg13g2_fill_8 FILLER_4_520 ();
 sg13g2_fill_8 FILLER_4_528 ();
 sg13g2_fill_8 FILLER_4_536 ();
 sg13g2_fill_8 FILLER_4_544 ();
 sg13g2_fill_8 FILLER_4_552 ();
 sg13g2_fill_8 FILLER_4_560 ();
 sg13g2_fill_8 FILLER_4_568 ();
 sg13g2_fill_8 FILLER_4_576 ();
 sg13g2_fill_8 FILLER_4_584 ();
 sg13g2_fill_8 FILLER_4_592 ();
 sg13g2_fill_8 FILLER_4_600 ();
 sg13g2_fill_8 FILLER_4_608 ();
 sg13g2_fill_8 FILLER_4_616 ();
 sg13g2_fill_8 FILLER_4_624 ();
 sg13g2_fill_8 FILLER_4_632 ();
 sg13g2_fill_8 FILLER_4_640 ();
 sg13g2_fill_8 FILLER_4_648 ();
 sg13g2_fill_8 FILLER_4_656 ();
 sg13g2_fill_8 FILLER_4_664 ();
 sg13g2_fill_8 FILLER_4_672 ();
 sg13g2_fill_8 FILLER_4_680 ();
 sg13g2_fill_8 FILLER_4_688 ();
 sg13g2_fill_8 FILLER_4_696 ();
 sg13g2_fill_8 FILLER_4_704 ();
 sg13g2_fill_8 FILLER_4_712 ();
 sg13g2_fill_8 FILLER_4_720 ();
 sg13g2_fill_8 FILLER_4_728 ();
 sg13g2_fill_8 FILLER_4_736 ();
 sg13g2_fill_8 FILLER_4_744 ();
 sg13g2_fill_8 FILLER_4_752 ();
 sg13g2_fill_8 FILLER_4_760 ();
 sg13g2_fill_8 FILLER_4_768 ();
 sg13g2_fill_8 FILLER_4_776 ();
 sg13g2_fill_8 FILLER_4_784 ();
 sg13g2_fill_8 FILLER_4_792 ();
 sg13g2_fill_8 FILLER_4_800 ();
 sg13g2_fill_8 FILLER_4_808 ();
 sg13g2_fill_8 FILLER_4_816 ();
 sg13g2_fill_8 FILLER_4_824 ();
 sg13g2_fill_8 FILLER_4_832 ();
 sg13g2_fill_8 FILLER_4_840 ();
 sg13g2_fill_8 FILLER_4_848 ();
 sg13g2_fill_8 FILLER_4_856 ();
 sg13g2_fill_8 FILLER_4_864 ();
 sg13g2_fill_8 FILLER_4_872 ();
 sg13g2_fill_8 FILLER_4_880 ();
 sg13g2_fill_8 FILLER_4_888 ();
 sg13g2_fill_8 FILLER_4_896 ();
 sg13g2_fill_8 FILLER_4_904 ();
 sg13g2_fill_8 FILLER_4_912 ();
 sg13g2_fill_8 FILLER_4_920 ();
 sg13g2_fill_8 FILLER_4_928 ();
 sg13g2_fill_8 FILLER_4_936 ();
 sg13g2_fill_8 FILLER_4_944 ();
 sg13g2_fill_8 FILLER_4_952 ();
 sg13g2_fill_8 FILLER_4_960 ();
 sg13g2_fill_8 FILLER_4_968 ();
 sg13g2_fill_8 FILLER_4_976 ();
 sg13g2_fill_8 FILLER_4_984 ();
 sg13g2_fill_8 FILLER_4_992 ();
 sg13g2_fill_8 FILLER_4_1000 ();
 sg13g2_fill_8 FILLER_4_1008 ();
 sg13g2_fill_8 FILLER_4_1016 ();
 sg13g2_fill_8 FILLER_4_1024 ();
 sg13g2_fill_8 FILLER_4_1032 ();
 sg13g2_fill_8 FILLER_4_1040 ();
 sg13g2_fill_8 FILLER_4_1048 ();
 sg13g2_fill_8 FILLER_4_1056 ();
 sg13g2_fill_8 FILLER_4_1064 ();
 sg13g2_fill_8 FILLER_4_1072 ();
 sg13g2_fill_8 FILLER_4_1080 ();
 sg13g2_fill_8 FILLER_4_1088 ();
 sg13g2_fill_8 FILLER_4_1096 ();
 sg13g2_fill_8 FILLER_4_1104 ();
 sg13g2_fill_8 FILLER_4_1112 ();
 sg13g2_fill_8 FILLER_4_1120 ();
 sg13g2_fill_8 FILLER_4_1128 ();
 sg13g2_fill_8 FILLER_4_1136 ();
 sg13g2_fill_8 FILLER_4_1144 ();
 sg13g2_fill_8 FILLER_4_1152 ();
 sg13g2_fill_4 FILLER_4_1160 ();
 sg13g2_fill_2 FILLER_4_1164 ();
 sg13g2_fill_8 FILLER_5_0 ();
 sg13g2_fill_8 FILLER_5_8 ();
 sg13g2_fill_8 FILLER_5_16 ();
 sg13g2_fill_8 FILLER_5_24 ();
 sg13g2_fill_8 FILLER_5_32 ();
 sg13g2_fill_8 FILLER_5_40 ();
 sg13g2_fill_8 FILLER_5_48 ();
 sg13g2_fill_8 FILLER_5_56 ();
 sg13g2_fill_8 FILLER_5_64 ();
 sg13g2_fill_8 FILLER_5_72 ();
 sg13g2_fill_8 FILLER_5_80 ();
 sg13g2_fill_8 FILLER_5_88 ();
 sg13g2_fill_8 FILLER_5_96 ();
 sg13g2_fill_8 FILLER_5_104 ();
 sg13g2_fill_8 FILLER_5_112 ();
 sg13g2_fill_8 FILLER_5_120 ();
 sg13g2_fill_8 FILLER_5_128 ();
 sg13g2_fill_8 FILLER_5_136 ();
 sg13g2_fill_8 FILLER_5_144 ();
 sg13g2_fill_8 FILLER_5_152 ();
 sg13g2_fill_8 FILLER_5_160 ();
 sg13g2_fill_8 FILLER_5_168 ();
 sg13g2_fill_8 FILLER_5_176 ();
 sg13g2_fill_8 FILLER_5_184 ();
 sg13g2_fill_8 FILLER_5_192 ();
 sg13g2_fill_8 FILLER_5_200 ();
 sg13g2_fill_8 FILLER_5_208 ();
 sg13g2_fill_8 FILLER_5_216 ();
 sg13g2_fill_8 FILLER_5_224 ();
 sg13g2_fill_8 FILLER_5_232 ();
 sg13g2_fill_8 FILLER_5_240 ();
 sg13g2_fill_8 FILLER_5_248 ();
 sg13g2_fill_8 FILLER_5_256 ();
 sg13g2_fill_8 FILLER_5_264 ();
 sg13g2_fill_8 FILLER_5_272 ();
 sg13g2_fill_8 FILLER_5_280 ();
 sg13g2_fill_8 FILLER_5_288 ();
 sg13g2_fill_8 FILLER_5_296 ();
 sg13g2_fill_8 FILLER_5_304 ();
 sg13g2_fill_8 FILLER_5_312 ();
 sg13g2_fill_8 FILLER_5_320 ();
 sg13g2_fill_8 FILLER_5_328 ();
 sg13g2_fill_8 FILLER_5_336 ();
 sg13g2_fill_8 FILLER_5_344 ();
 sg13g2_fill_8 FILLER_5_352 ();
 sg13g2_fill_8 FILLER_5_360 ();
 sg13g2_fill_8 FILLER_5_368 ();
 sg13g2_fill_8 FILLER_5_376 ();
 sg13g2_fill_8 FILLER_5_384 ();
 sg13g2_fill_8 FILLER_5_392 ();
 sg13g2_fill_8 FILLER_5_400 ();
 sg13g2_fill_8 FILLER_5_408 ();
 sg13g2_fill_4 FILLER_5_416 ();
 sg13g2_fill_2 FILLER_5_420 ();
 sg13g2_fill_1 FILLER_5_422 ();
 sg13g2_fill_8 FILLER_5_426 ();
 sg13g2_fill_8 FILLER_5_434 ();
 sg13g2_fill_8 FILLER_5_442 ();
 sg13g2_fill_8 FILLER_5_450 ();
 sg13g2_fill_8 FILLER_5_458 ();
 sg13g2_fill_8 FILLER_5_466 ();
 sg13g2_fill_8 FILLER_5_474 ();
 sg13g2_fill_8 FILLER_5_482 ();
 sg13g2_fill_8 FILLER_5_490 ();
 sg13g2_fill_8 FILLER_5_498 ();
 sg13g2_fill_8 FILLER_5_506 ();
 sg13g2_fill_8 FILLER_5_514 ();
 sg13g2_fill_8 FILLER_5_522 ();
 sg13g2_fill_8 FILLER_5_530 ();
 sg13g2_fill_8 FILLER_5_538 ();
 sg13g2_fill_8 FILLER_5_546 ();
 sg13g2_fill_8 FILLER_5_554 ();
 sg13g2_fill_8 FILLER_5_562 ();
 sg13g2_fill_8 FILLER_5_570 ();
 sg13g2_fill_8 FILLER_5_578 ();
 sg13g2_fill_8 FILLER_5_586 ();
 sg13g2_fill_8 FILLER_5_594 ();
 sg13g2_fill_8 FILLER_5_602 ();
 sg13g2_fill_8 FILLER_5_610 ();
 sg13g2_fill_8 FILLER_5_618 ();
 sg13g2_fill_8 FILLER_5_626 ();
 sg13g2_fill_8 FILLER_5_634 ();
 sg13g2_fill_8 FILLER_5_642 ();
 sg13g2_fill_8 FILLER_5_650 ();
 sg13g2_fill_8 FILLER_5_658 ();
 sg13g2_fill_8 FILLER_5_666 ();
 sg13g2_fill_8 FILLER_5_674 ();
 sg13g2_fill_8 FILLER_5_682 ();
 sg13g2_fill_8 FILLER_5_690 ();
 sg13g2_fill_8 FILLER_5_698 ();
 sg13g2_fill_8 FILLER_5_706 ();
 sg13g2_fill_8 FILLER_5_714 ();
 sg13g2_fill_8 FILLER_5_722 ();
 sg13g2_fill_8 FILLER_5_730 ();
 sg13g2_fill_8 FILLER_5_738 ();
 sg13g2_fill_8 FILLER_5_746 ();
 sg13g2_fill_8 FILLER_5_754 ();
 sg13g2_fill_8 FILLER_5_762 ();
 sg13g2_fill_8 FILLER_5_770 ();
 sg13g2_fill_8 FILLER_5_778 ();
 sg13g2_fill_8 FILLER_5_786 ();
 sg13g2_fill_8 FILLER_5_794 ();
 sg13g2_fill_8 FILLER_5_802 ();
 sg13g2_fill_8 FILLER_5_810 ();
 sg13g2_fill_8 FILLER_5_818 ();
 sg13g2_fill_8 FILLER_5_826 ();
 sg13g2_fill_8 FILLER_5_834 ();
 sg13g2_fill_8 FILLER_5_842 ();
 sg13g2_fill_8 FILLER_5_850 ();
 sg13g2_fill_8 FILLER_5_858 ();
 sg13g2_fill_8 FILLER_5_866 ();
 sg13g2_fill_8 FILLER_5_874 ();
 sg13g2_fill_8 FILLER_5_882 ();
 sg13g2_fill_8 FILLER_5_890 ();
 sg13g2_fill_8 FILLER_5_898 ();
 sg13g2_fill_8 FILLER_5_906 ();
 sg13g2_fill_8 FILLER_5_914 ();
 sg13g2_fill_8 FILLER_5_922 ();
 sg13g2_fill_8 FILLER_5_930 ();
 sg13g2_fill_8 FILLER_5_938 ();
 sg13g2_fill_8 FILLER_5_946 ();
 sg13g2_fill_8 FILLER_5_954 ();
 sg13g2_fill_8 FILLER_5_962 ();
 sg13g2_fill_8 FILLER_5_970 ();
 sg13g2_fill_8 FILLER_5_978 ();
 sg13g2_fill_8 FILLER_5_986 ();
 sg13g2_fill_8 FILLER_5_994 ();
 sg13g2_fill_8 FILLER_5_1002 ();
 sg13g2_fill_8 FILLER_5_1010 ();
 sg13g2_fill_8 FILLER_5_1018 ();
 sg13g2_fill_8 FILLER_5_1026 ();
 sg13g2_fill_8 FILLER_5_1034 ();
 sg13g2_fill_8 FILLER_5_1042 ();
 sg13g2_fill_8 FILLER_5_1050 ();
 sg13g2_fill_8 FILLER_5_1058 ();
 sg13g2_fill_8 FILLER_5_1066 ();
 sg13g2_fill_8 FILLER_5_1074 ();
 sg13g2_fill_8 FILLER_5_1082 ();
 sg13g2_fill_8 FILLER_5_1090 ();
 sg13g2_fill_8 FILLER_5_1098 ();
 sg13g2_fill_8 FILLER_5_1106 ();
 sg13g2_fill_8 FILLER_5_1114 ();
 sg13g2_fill_8 FILLER_5_1122 ();
 sg13g2_fill_8 FILLER_5_1130 ();
 sg13g2_fill_8 FILLER_5_1138 ();
 sg13g2_fill_8 FILLER_5_1146 ();
 sg13g2_fill_8 FILLER_5_1154 ();
 sg13g2_fill_4 FILLER_5_1162 ();
 sg13g2_fill_8 FILLER_6_0 ();
 sg13g2_fill_8 FILLER_6_8 ();
 sg13g2_fill_8 FILLER_6_16 ();
 sg13g2_fill_8 FILLER_6_24 ();
 sg13g2_fill_8 FILLER_6_32 ();
 sg13g2_fill_8 FILLER_6_40 ();
 sg13g2_fill_8 FILLER_6_48 ();
 sg13g2_fill_8 FILLER_6_56 ();
 sg13g2_fill_8 FILLER_6_64 ();
 sg13g2_fill_8 FILLER_6_72 ();
 sg13g2_fill_8 FILLER_6_80 ();
 sg13g2_fill_8 FILLER_6_88 ();
 sg13g2_fill_8 FILLER_6_96 ();
 sg13g2_fill_8 FILLER_6_104 ();
 sg13g2_fill_8 FILLER_6_112 ();
 sg13g2_fill_8 FILLER_6_120 ();
 sg13g2_fill_8 FILLER_6_128 ();
 sg13g2_fill_8 FILLER_6_136 ();
 sg13g2_fill_8 FILLER_6_144 ();
 sg13g2_fill_8 FILLER_6_152 ();
 sg13g2_fill_8 FILLER_6_160 ();
 sg13g2_fill_8 FILLER_6_168 ();
 sg13g2_fill_8 FILLER_6_176 ();
 sg13g2_fill_8 FILLER_6_184 ();
 sg13g2_fill_8 FILLER_6_192 ();
 sg13g2_fill_8 FILLER_6_200 ();
 sg13g2_fill_8 FILLER_6_208 ();
 sg13g2_fill_8 FILLER_6_216 ();
 sg13g2_fill_8 FILLER_6_224 ();
 sg13g2_fill_8 FILLER_6_232 ();
 sg13g2_fill_8 FILLER_6_240 ();
 sg13g2_fill_8 FILLER_6_248 ();
 sg13g2_fill_8 FILLER_6_256 ();
 sg13g2_fill_8 FILLER_6_264 ();
 sg13g2_fill_8 FILLER_6_272 ();
 sg13g2_fill_8 FILLER_6_280 ();
 sg13g2_fill_8 FILLER_6_288 ();
 sg13g2_fill_8 FILLER_6_296 ();
 sg13g2_fill_8 FILLER_6_304 ();
 sg13g2_fill_8 FILLER_6_312 ();
 sg13g2_fill_8 FILLER_6_320 ();
 sg13g2_fill_8 FILLER_6_328 ();
 sg13g2_fill_8 FILLER_6_336 ();
 sg13g2_fill_8 FILLER_6_344 ();
 sg13g2_fill_8 FILLER_6_352 ();
 sg13g2_fill_8 FILLER_6_360 ();
 sg13g2_fill_8 FILLER_6_368 ();
 sg13g2_fill_8 FILLER_6_376 ();
 sg13g2_fill_8 FILLER_6_384 ();
 sg13g2_fill_8 FILLER_6_392 ();
 sg13g2_fill_8 FILLER_6_400 ();
 sg13g2_fill_8 FILLER_6_408 ();
 sg13g2_fill_8 FILLER_6_441 ();
 sg13g2_fill_8 FILLER_6_449 ();
 sg13g2_fill_8 FILLER_6_457 ();
 sg13g2_fill_8 FILLER_6_465 ();
 sg13g2_fill_8 FILLER_6_473 ();
 sg13g2_fill_8 FILLER_6_481 ();
 sg13g2_fill_2 FILLER_6_492 ();
 sg13g2_fill_8 FILLER_6_500 ();
 sg13g2_fill_8 FILLER_6_508 ();
 sg13g2_fill_8 FILLER_6_516 ();
 sg13g2_fill_8 FILLER_6_524 ();
 sg13g2_fill_8 FILLER_6_532 ();
 sg13g2_fill_8 FILLER_6_540 ();
 sg13g2_fill_8 FILLER_6_548 ();
 sg13g2_fill_8 FILLER_6_556 ();
 sg13g2_fill_8 FILLER_6_564 ();
 sg13g2_fill_8 FILLER_6_572 ();
 sg13g2_fill_8 FILLER_6_580 ();
 sg13g2_fill_8 FILLER_6_588 ();
 sg13g2_fill_8 FILLER_6_596 ();
 sg13g2_fill_8 FILLER_6_604 ();
 sg13g2_fill_8 FILLER_6_612 ();
 sg13g2_fill_8 FILLER_6_620 ();
 sg13g2_fill_8 FILLER_6_628 ();
 sg13g2_fill_8 FILLER_6_636 ();
 sg13g2_fill_8 FILLER_6_644 ();
 sg13g2_fill_8 FILLER_6_652 ();
 sg13g2_fill_8 FILLER_6_660 ();
 sg13g2_fill_8 FILLER_6_668 ();
 sg13g2_fill_8 FILLER_6_676 ();
 sg13g2_fill_8 FILLER_6_684 ();
 sg13g2_fill_8 FILLER_6_692 ();
 sg13g2_fill_8 FILLER_6_700 ();
 sg13g2_fill_8 FILLER_6_708 ();
 sg13g2_fill_8 FILLER_6_716 ();
 sg13g2_fill_8 FILLER_6_724 ();
 sg13g2_fill_8 FILLER_6_732 ();
 sg13g2_fill_8 FILLER_6_740 ();
 sg13g2_fill_8 FILLER_6_748 ();
 sg13g2_fill_8 FILLER_6_756 ();
 sg13g2_fill_8 FILLER_6_764 ();
 sg13g2_fill_8 FILLER_6_772 ();
 sg13g2_fill_8 FILLER_6_780 ();
 sg13g2_fill_8 FILLER_6_788 ();
 sg13g2_fill_8 FILLER_6_796 ();
 sg13g2_fill_8 FILLER_6_804 ();
 sg13g2_fill_8 FILLER_6_812 ();
 sg13g2_fill_8 FILLER_6_820 ();
 sg13g2_fill_8 FILLER_6_828 ();
 sg13g2_fill_8 FILLER_6_836 ();
 sg13g2_fill_8 FILLER_6_844 ();
 sg13g2_fill_8 FILLER_6_852 ();
 sg13g2_fill_8 FILLER_6_860 ();
 sg13g2_fill_8 FILLER_6_868 ();
 sg13g2_fill_8 FILLER_6_876 ();
 sg13g2_fill_8 FILLER_6_884 ();
 sg13g2_fill_8 FILLER_6_892 ();
 sg13g2_fill_8 FILLER_6_900 ();
 sg13g2_fill_8 FILLER_6_908 ();
 sg13g2_fill_8 FILLER_6_916 ();
 sg13g2_fill_8 FILLER_6_924 ();
 sg13g2_fill_8 FILLER_6_932 ();
 sg13g2_fill_8 FILLER_6_940 ();
 sg13g2_fill_8 FILLER_6_948 ();
 sg13g2_fill_8 FILLER_6_956 ();
 sg13g2_fill_8 FILLER_6_964 ();
 sg13g2_fill_8 FILLER_6_972 ();
 sg13g2_fill_8 FILLER_6_980 ();
 sg13g2_fill_8 FILLER_6_988 ();
 sg13g2_fill_8 FILLER_6_996 ();
 sg13g2_fill_8 FILLER_6_1004 ();
 sg13g2_fill_8 FILLER_6_1012 ();
 sg13g2_fill_8 FILLER_6_1020 ();
 sg13g2_fill_8 FILLER_6_1028 ();
 sg13g2_fill_8 FILLER_6_1036 ();
 sg13g2_fill_8 FILLER_6_1044 ();
 sg13g2_fill_8 FILLER_6_1052 ();
 sg13g2_fill_8 FILLER_6_1060 ();
 sg13g2_fill_8 FILLER_6_1068 ();
 sg13g2_fill_8 FILLER_6_1076 ();
 sg13g2_fill_8 FILLER_6_1084 ();
 sg13g2_fill_8 FILLER_6_1092 ();
 sg13g2_fill_8 FILLER_6_1100 ();
 sg13g2_fill_8 FILLER_6_1108 ();
 sg13g2_fill_8 FILLER_6_1116 ();
 sg13g2_fill_8 FILLER_6_1124 ();
 sg13g2_fill_8 FILLER_6_1132 ();
 sg13g2_fill_8 FILLER_6_1140 ();
 sg13g2_fill_8 FILLER_6_1148 ();
 sg13g2_fill_8 FILLER_6_1156 ();
 sg13g2_fill_2 FILLER_6_1164 ();
 sg13g2_fill_8 FILLER_7_0 ();
 sg13g2_fill_8 FILLER_7_8 ();
 sg13g2_fill_8 FILLER_7_16 ();
 sg13g2_fill_8 FILLER_7_24 ();
 sg13g2_fill_8 FILLER_7_32 ();
 sg13g2_fill_8 FILLER_7_40 ();
 sg13g2_fill_8 FILLER_7_48 ();
 sg13g2_fill_8 FILLER_7_56 ();
 sg13g2_fill_8 FILLER_7_64 ();
 sg13g2_fill_8 FILLER_7_72 ();
 sg13g2_fill_8 FILLER_7_80 ();
 sg13g2_fill_8 FILLER_7_88 ();
 sg13g2_fill_8 FILLER_7_96 ();
 sg13g2_fill_8 FILLER_7_104 ();
 sg13g2_fill_8 FILLER_7_112 ();
 sg13g2_fill_8 FILLER_7_120 ();
 sg13g2_fill_8 FILLER_7_128 ();
 sg13g2_fill_8 FILLER_7_136 ();
 sg13g2_fill_8 FILLER_7_144 ();
 sg13g2_fill_8 FILLER_7_152 ();
 sg13g2_fill_8 FILLER_7_160 ();
 sg13g2_fill_8 FILLER_7_168 ();
 sg13g2_fill_8 FILLER_7_176 ();
 sg13g2_fill_8 FILLER_7_184 ();
 sg13g2_fill_8 FILLER_7_192 ();
 sg13g2_fill_8 FILLER_7_200 ();
 sg13g2_fill_8 FILLER_7_208 ();
 sg13g2_fill_8 FILLER_7_216 ();
 sg13g2_fill_8 FILLER_7_224 ();
 sg13g2_fill_8 FILLER_7_232 ();
 sg13g2_fill_8 FILLER_7_240 ();
 sg13g2_fill_8 FILLER_7_248 ();
 sg13g2_fill_8 FILLER_7_256 ();
 sg13g2_fill_8 FILLER_7_264 ();
 sg13g2_fill_8 FILLER_7_272 ();
 sg13g2_fill_8 FILLER_7_280 ();
 sg13g2_fill_8 FILLER_7_288 ();
 sg13g2_fill_8 FILLER_7_296 ();
 sg13g2_fill_4 FILLER_7_304 ();
 sg13g2_fill_2 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_315 ();
 sg13g2_fill_8 FILLER_7_322 ();
 sg13g2_fill_4 FILLER_7_330 ();
 sg13g2_fill_2 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_336 ();
 sg13g2_fill_8 FILLER_7_363 ();
 sg13g2_fill_8 FILLER_7_371 ();
 sg13g2_fill_8 FILLER_7_379 ();
 sg13g2_fill_8 FILLER_7_387 ();
 sg13g2_fill_8 FILLER_7_395 ();
 sg13g2_fill_2 FILLER_7_403 ();
 sg13g2_fill_1 FILLER_7_405 ();
 sg13g2_fill_2 FILLER_7_437 ();
 sg13g2_fill_8 FILLER_7_465 ();
 sg13g2_fill_8 FILLER_7_473 ();
 sg13g2_fill_8 FILLER_7_507 ();
 sg13g2_fill_8 FILLER_7_515 ();
 sg13g2_fill_8 FILLER_7_523 ();
 sg13g2_fill_8 FILLER_7_531 ();
 sg13g2_fill_8 FILLER_7_539 ();
 sg13g2_fill_8 FILLER_7_547 ();
 sg13g2_fill_8 FILLER_7_555 ();
 sg13g2_fill_8 FILLER_7_563 ();
 sg13g2_fill_8 FILLER_7_571 ();
 sg13g2_fill_8 FILLER_7_579 ();
 sg13g2_fill_8 FILLER_7_587 ();
 sg13g2_fill_8 FILLER_7_595 ();
 sg13g2_fill_8 FILLER_7_603 ();
 sg13g2_fill_8 FILLER_7_611 ();
 sg13g2_fill_8 FILLER_7_619 ();
 sg13g2_fill_8 FILLER_7_627 ();
 sg13g2_fill_8 FILLER_7_635 ();
 sg13g2_fill_8 FILLER_7_643 ();
 sg13g2_fill_8 FILLER_7_651 ();
 sg13g2_fill_8 FILLER_7_659 ();
 sg13g2_fill_8 FILLER_7_667 ();
 sg13g2_fill_8 FILLER_7_675 ();
 sg13g2_fill_8 FILLER_7_683 ();
 sg13g2_fill_8 FILLER_7_691 ();
 sg13g2_fill_8 FILLER_7_699 ();
 sg13g2_fill_8 FILLER_7_707 ();
 sg13g2_fill_8 FILLER_7_715 ();
 sg13g2_fill_8 FILLER_7_723 ();
 sg13g2_fill_8 FILLER_7_731 ();
 sg13g2_fill_8 FILLER_7_739 ();
 sg13g2_fill_8 FILLER_7_747 ();
 sg13g2_fill_8 FILLER_7_755 ();
 sg13g2_fill_8 FILLER_7_763 ();
 sg13g2_fill_8 FILLER_7_771 ();
 sg13g2_fill_8 FILLER_7_779 ();
 sg13g2_fill_8 FILLER_7_787 ();
 sg13g2_fill_8 FILLER_7_795 ();
 sg13g2_fill_8 FILLER_7_803 ();
 sg13g2_fill_8 FILLER_7_811 ();
 sg13g2_fill_8 FILLER_7_819 ();
 sg13g2_fill_8 FILLER_7_827 ();
 sg13g2_fill_8 FILLER_7_835 ();
 sg13g2_fill_8 FILLER_7_843 ();
 sg13g2_fill_8 FILLER_7_851 ();
 sg13g2_fill_8 FILLER_7_859 ();
 sg13g2_fill_8 FILLER_7_867 ();
 sg13g2_fill_8 FILLER_7_875 ();
 sg13g2_fill_8 FILLER_7_883 ();
 sg13g2_fill_8 FILLER_7_891 ();
 sg13g2_fill_8 FILLER_7_899 ();
 sg13g2_fill_8 FILLER_7_907 ();
 sg13g2_fill_8 FILLER_7_915 ();
 sg13g2_fill_8 FILLER_7_923 ();
 sg13g2_fill_8 FILLER_7_931 ();
 sg13g2_fill_8 FILLER_7_939 ();
 sg13g2_fill_8 FILLER_7_947 ();
 sg13g2_fill_8 FILLER_7_955 ();
 sg13g2_fill_8 FILLER_7_963 ();
 sg13g2_fill_8 FILLER_7_971 ();
 sg13g2_fill_8 FILLER_7_979 ();
 sg13g2_fill_8 FILLER_7_987 ();
 sg13g2_fill_8 FILLER_7_995 ();
 sg13g2_fill_8 FILLER_7_1003 ();
 sg13g2_fill_8 FILLER_7_1011 ();
 sg13g2_fill_8 FILLER_7_1019 ();
 sg13g2_fill_8 FILLER_7_1027 ();
 sg13g2_fill_8 FILLER_7_1035 ();
 sg13g2_fill_8 FILLER_7_1043 ();
 sg13g2_fill_8 FILLER_7_1051 ();
 sg13g2_fill_8 FILLER_7_1059 ();
 sg13g2_fill_8 FILLER_7_1067 ();
 sg13g2_fill_8 FILLER_7_1075 ();
 sg13g2_fill_8 FILLER_7_1083 ();
 sg13g2_fill_8 FILLER_7_1091 ();
 sg13g2_fill_8 FILLER_7_1099 ();
 sg13g2_fill_8 FILLER_7_1107 ();
 sg13g2_fill_8 FILLER_7_1115 ();
 sg13g2_fill_8 FILLER_7_1123 ();
 sg13g2_fill_8 FILLER_7_1131 ();
 sg13g2_fill_8 FILLER_7_1139 ();
 sg13g2_fill_8 FILLER_7_1147 ();
 sg13g2_fill_8 FILLER_7_1155 ();
 sg13g2_fill_2 FILLER_7_1163 ();
 sg13g2_fill_1 FILLER_7_1165 ();
 sg13g2_fill_8 FILLER_8_0 ();
 sg13g2_fill_8 FILLER_8_8 ();
 sg13g2_fill_8 FILLER_8_16 ();
 sg13g2_fill_8 FILLER_8_24 ();
 sg13g2_fill_8 FILLER_8_32 ();
 sg13g2_fill_8 FILLER_8_40 ();
 sg13g2_fill_8 FILLER_8_48 ();
 sg13g2_fill_8 FILLER_8_56 ();
 sg13g2_fill_8 FILLER_8_64 ();
 sg13g2_fill_8 FILLER_8_72 ();
 sg13g2_fill_8 FILLER_8_80 ();
 sg13g2_fill_8 FILLER_8_88 ();
 sg13g2_fill_8 FILLER_8_96 ();
 sg13g2_fill_8 FILLER_8_104 ();
 sg13g2_fill_8 FILLER_8_112 ();
 sg13g2_fill_8 FILLER_8_120 ();
 sg13g2_fill_8 FILLER_8_128 ();
 sg13g2_fill_8 FILLER_8_136 ();
 sg13g2_fill_8 FILLER_8_144 ();
 sg13g2_fill_8 FILLER_8_152 ();
 sg13g2_fill_8 FILLER_8_160 ();
 sg13g2_fill_2 FILLER_8_168 ();
 sg13g2_fill_1 FILLER_8_170 ();
 sg13g2_fill_8 FILLER_8_197 ();
 sg13g2_fill_8 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_213 ();
 sg13g2_fill_8 FILLER_8_217 ();
 sg13g2_fill_8 FILLER_8_225 ();
 sg13g2_fill_4 FILLER_8_233 ();
 sg13g2_fill_8 FILLER_8_263 ();
 sg13g2_fill_8 FILLER_8_271 ();
 sg13g2_fill_8 FILLER_8_279 ();
 sg13g2_fill_8 FILLER_8_287 ();
 sg13g2_fill_4 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_299 ();
 sg13g2_fill_1 FILLER_8_301 ();
 sg13g2_fill_4 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_332 ();
 sg13g2_fill_8 FILLER_8_370 ();
 sg13g2_fill_2 FILLER_8_378 ();
 sg13g2_fill_8 FILLER_8_461 ();
 sg13g2_fill_4 FILLER_8_469 ();
 sg13g2_fill_1 FILLER_8_473 ();
 sg13g2_fill_8 FILLER_8_531 ();
 sg13g2_fill_8 FILLER_8_539 ();
 sg13g2_fill_8 FILLER_8_547 ();
 sg13g2_fill_8 FILLER_8_555 ();
 sg13g2_fill_8 FILLER_8_563 ();
 sg13g2_fill_8 FILLER_8_571 ();
 sg13g2_fill_8 FILLER_8_579 ();
 sg13g2_fill_8 FILLER_8_587 ();
 sg13g2_fill_8 FILLER_8_595 ();
 sg13g2_fill_8 FILLER_8_603 ();
 sg13g2_fill_8 FILLER_8_611 ();
 sg13g2_fill_8 FILLER_8_619 ();
 sg13g2_fill_8 FILLER_8_627 ();
 sg13g2_fill_8 FILLER_8_635 ();
 sg13g2_fill_8 FILLER_8_643 ();
 sg13g2_fill_8 FILLER_8_651 ();
 sg13g2_fill_8 FILLER_8_659 ();
 sg13g2_fill_8 FILLER_8_667 ();
 sg13g2_fill_8 FILLER_8_675 ();
 sg13g2_fill_8 FILLER_8_683 ();
 sg13g2_fill_8 FILLER_8_691 ();
 sg13g2_fill_8 FILLER_8_699 ();
 sg13g2_fill_8 FILLER_8_707 ();
 sg13g2_fill_8 FILLER_8_715 ();
 sg13g2_fill_8 FILLER_8_723 ();
 sg13g2_fill_8 FILLER_8_731 ();
 sg13g2_fill_8 FILLER_8_739 ();
 sg13g2_fill_8 FILLER_8_747 ();
 sg13g2_fill_8 FILLER_8_755 ();
 sg13g2_fill_8 FILLER_8_763 ();
 sg13g2_fill_8 FILLER_8_771 ();
 sg13g2_fill_8 FILLER_8_779 ();
 sg13g2_fill_8 FILLER_8_787 ();
 sg13g2_fill_8 FILLER_8_795 ();
 sg13g2_fill_8 FILLER_8_803 ();
 sg13g2_fill_8 FILLER_8_811 ();
 sg13g2_fill_8 FILLER_8_819 ();
 sg13g2_fill_8 FILLER_8_827 ();
 sg13g2_fill_8 FILLER_8_835 ();
 sg13g2_fill_8 FILLER_8_843 ();
 sg13g2_fill_8 FILLER_8_851 ();
 sg13g2_fill_8 FILLER_8_859 ();
 sg13g2_fill_8 FILLER_8_867 ();
 sg13g2_fill_8 FILLER_8_875 ();
 sg13g2_fill_8 FILLER_8_883 ();
 sg13g2_fill_8 FILLER_8_891 ();
 sg13g2_fill_8 FILLER_8_899 ();
 sg13g2_fill_8 FILLER_8_907 ();
 sg13g2_fill_8 FILLER_8_915 ();
 sg13g2_fill_8 FILLER_8_923 ();
 sg13g2_fill_8 FILLER_8_931 ();
 sg13g2_fill_8 FILLER_8_939 ();
 sg13g2_fill_8 FILLER_8_947 ();
 sg13g2_fill_8 FILLER_8_955 ();
 sg13g2_fill_8 FILLER_8_963 ();
 sg13g2_fill_8 FILLER_8_971 ();
 sg13g2_fill_8 FILLER_8_979 ();
 sg13g2_fill_8 FILLER_8_987 ();
 sg13g2_fill_8 FILLER_8_995 ();
 sg13g2_fill_8 FILLER_8_1003 ();
 sg13g2_fill_8 FILLER_8_1011 ();
 sg13g2_fill_8 FILLER_8_1019 ();
 sg13g2_fill_8 FILLER_8_1027 ();
 sg13g2_fill_8 FILLER_8_1035 ();
 sg13g2_fill_8 FILLER_8_1043 ();
 sg13g2_fill_8 FILLER_8_1051 ();
 sg13g2_fill_8 FILLER_8_1059 ();
 sg13g2_fill_8 FILLER_8_1067 ();
 sg13g2_fill_8 FILLER_8_1075 ();
 sg13g2_fill_8 FILLER_8_1083 ();
 sg13g2_fill_8 FILLER_8_1091 ();
 sg13g2_fill_8 FILLER_8_1099 ();
 sg13g2_fill_8 FILLER_8_1107 ();
 sg13g2_fill_8 FILLER_8_1115 ();
 sg13g2_fill_8 FILLER_8_1123 ();
 sg13g2_fill_8 FILLER_8_1131 ();
 sg13g2_fill_8 FILLER_8_1139 ();
 sg13g2_fill_8 FILLER_8_1147 ();
 sg13g2_fill_8 FILLER_8_1155 ();
 sg13g2_fill_2 FILLER_8_1163 ();
 sg13g2_fill_1 FILLER_8_1165 ();
 sg13g2_fill_8 FILLER_9_0 ();
 sg13g2_fill_8 FILLER_9_8 ();
 sg13g2_fill_8 FILLER_9_16 ();
 sg13g2_fill_8 FILLER_9_24 ();
 sg13g2_fill_8 FILLER_9_32 ();
 sg13g2_fill_8 FILLER_9_40 ();
 sg13g2_fill_8 FILLER_9_48 ();
 sg13g2_fill_8 FILLER_9_56 ();
 sg13g2_fill_8 FILLER_9_64 ();
 sg13g2_fill_8 FILLER_9_72 ();
 sg13g2_fill_8 FILLER_9_80 ();
 sg13g2_fill_8 FILLER_9_88 ();
 sg13g2_fill_8 FILLER_9_96 ();
 sg13g2_fill_8 FILLER_9_104 ();
 sg13g2_fill_8 FILLER_9_112 ();
 sg13g2_fill_8 FILLER_9_120 ();
 sg13g2_fill_8 FILLER_9_128 ();
 sg13g2_fill_8 FILLER_9_136 ();
 sg13g2_fill_4 FILLER_9_144 ();
 sg13g2_fill_1 FILLER_9_148 ();
 sg13g2_fill_2 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_156 ();
 sg13g2_fill_8 FILLER_9_160 ();
 sg13g2_fill_4 FILLER_9_168 ();
 sg13g2_fill_1 FILLER_9_198 ();
 sg13g2_fill_8 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_233 ();
 sg13g2_fill_4 FILLER_9_239 ();
 sg13g2_fill_2 FILLER_9_243 ();
 sg13g2_fill_1 FILLER_9_245 ();
 sg13g2_fill_4 FILLER_9_272 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_8 FILLER_9_286 ();
 sg13g2_fill_8 FILLER_9_294 ();
 sg13g2_fill_8 FILLER_9_352 ();
 sg13g2_fill_8 FILLER_9_360 ();
 sg13g2_fill_8 FILLER_9_368 ();
 sg13g2_fill_8 FILLER_9_384 ();
 sg13g2_fill_4 FILLER_9_392 ();
 sg13g2_fill_1 FILLER_9_396 ();
 sg13g2_fill_1 FILLER_9_410 ();
 sg13g2_fill_1 FILLER_9_496 ();
 sg13g2_fill_1 FILLER_9_508 ();
 sg13g2_fill_8 FILLER_9_539 ();
 sg13g2_fill_8 FILLER_9_547 ();
 sg13g2_fill_8 FILLER_9_555 ();
 sg13g2_fill_8 FILLER_9_563 ();
 sg13g2_fill_8 FILLER_9_571 ();
 sg13g2_fill_8 FILLER_9_579 ();
 sg13g2_fill_8 FILLER_9_587 ();
 sg13g2_fill_8 FILLER_9_595 ();
 sg13g2_fill_8 FILLER_9_603 ();
 sg13g2_fill_8 FILLER_9_611 ();
 sg13g2_fill_8 FILLER_9_619 ();
 sg13g2_fill_8 FILLER_9_627 ();
 sg13g2_fill_8 FILLER_9_635 ();
 sg13g2_fill_8 FILLER_9_643 ();
 sg13g2_fill_8 FILLER_9_651 ();
 sg13g2_fill_8 FILLER_9_659 ();
 sg13g2_fill_8 FILLER_9_667 ();
 sg13g2_fill_8 FILLER_9_675 ();
 sg13g2_fill_8 FILLER_9_683 ();
 sg13g2_fill_8 FILLER_9_691 ();
 sg13g2_fill_8 FILLER_9_699 ();
 sg13g2_fill_8 FILLER_9_707 ();
 sg13g2_fill_8 FILLER_9_715 ();
 sg13g2_fill_8 FILLER_9_723 ();
 sg13g2_fill_8 FILLER_9_731 ();
 sg13g2_fill_8 FILLER_9_739 ();
 sg13g2_fill_8 FILLER_9_747 ();
 sg13g2_fill_8 FILLER_9_755 ();
 sg13g2_fill_8 FILLER_9_763 ();
 sg13g2_fill_8 FILLER_9_771 ();
 sg13g2_fill_8 FILLER_9_779 ();
 sg13g2_fill_8 FILLER_9_787 ();
 sg13g2_fill_8 FILLER_9_795 ();
 sg13g2_fill_8 FILLER_9_803 ();
 sg13g2_fill_8 FILLER_9_811 ();
 sg13g2_fill_8 FILLER_9_819 ();
 sg13g2_fill_8 FILLER_9_827 ();
 sg13g2_fill_8 FILLER_9_835 ();
 sg13g2_fill_8 FILLER_9_843 ();
 sg13g2_fill_8 FILLER_9_851 ();
 sg13g2_fill_8 FILLER_9_859 ();
 sg13g2_fill_8 FILLER_9_867 ();
 sg13g2_fill_8 FILLER_9_875 ();
 sg13g2_fill_8 FILLER_9_883 ();
 sg13g2_fill_8 FILLER_9_891 ();
 sg13g2_fill_8 FILLER_9_899 ();
 sg13g2_fill_8 FILLER_9_907 ();
 sg13g2_fill_8 FILLER_9_915 ();
 sg13g2_fill_8 FILLER_9_923 ();
 sg13g2_fill_8 FILLER_9_931 ();
 sg13g2_fill_8 FILLER_9_939 ();
 sg13g2_fill_8 FILLER_9_947 ();
 sg13g2_fill_8 FILLER_9_955 ();
 sg13g2_fill_8 FILLER_9_963 ();
 sg13g2_fill_8 FILLER_9_971 ();
 sg13g2_fill_8 FILLER_9_979 ();
 sg13g2_fill_8 FILLER_9_987 ();
 sg13g2_fill_8 FILLER_9_995 ();
 sg13g2_fill_8 FILLER_9_1003 ();
 sg13g2_fill_8 FILLER_9_1011 ();
 sg13g2_fill_8 FILLER_9_1019 ();
 sg13g2_fill_8 FILLER_9_1027 ();
 sg13g2_fill_8 FILLER_9_1035 ();
 sg13g2_fill_8 FILLER_9_1043 ();
 sg13g2_fill_8 FILLER_9_1051 ();
 sg13g2_fill_8 FILLER_9_1059 ();
 sg13g2_fill_8 FILLER_9_1067 ();
 sg13g2_fill_8 FILLER_9_1075 ();
 sg13g2_fill_8 FILLER_9_1083 ();
 sg13g2_fill_8 FILLER_9_1091 ();
 sg13g2_fill_8 FILLER_9_1099 ();
 sg13g2_fill_8 FILLER_9_1107 ();
 sg13g2_fill_8 FILLER_9_1115 ();
 sg13g2_fill_8 FILLER_9_1123 ();
 sg13g2_fill_8 FILLER_9_1131 ();
 sg13g2_fill_8 FILLER_9_1139 ();
 sg13g2_fill_8 FILLER_9_1147 ();
 sg13g2_fill_8 FILLER_9_1155 ();
 sg13g2_fill_2 FILLER_9_1163 ();
 sg13g2_fill_1 FILLER_9_1165 ();
 sg13g2_fill_8 FILLER_10_0 ();
 sg13g2_fill_8 FILLER_10_8 ();
 sg13g2_fill_8 FILLER_10_16 ();
 sg13g2_fill_8 FILLER_10_24 ();
 sg13g2_fill_8 FILLER_10_32 ();
 sg13g2_fill_8 FILLER_10_40 ();
 sg13g2_fill_8 FILLER_10_48 ();
 sg13g2_fill_8 FILLER_10_56 ();
 sg13g2_fill_8 FILLER_10_64 ();
 sg13g2_fill_8 FILLER_10_72 ();
 sg13g2_fill_8 FILLER_10_80 ();
 sg13g2_fill_4 FILLER_10_88 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_fill_4 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_8 FILLER_10_209 ();
 sg13g2_fill_1 FILLER_10_236 ();
 sg13g2_fill_8 FILLER_10_266 ();
 sg13g2_fill_8 FILLER_10_274 ();
 sg13g2_fill_4 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_8 FILLER_10_348 ();
 sg13g2_fill_8 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_fill_4 FILLER_10_392 ();
 sg13g2_fill_8 FILLER_10_466 ();
 sg13g2_fill_4 FILLER_10_474 ();
 sg13g2_fill_1 FILLER_10_478 ();
 sg13g2_fill_8 FILLER_10_510 ();
 sg13g2_fill_8 FILLER_10_529 ();
 sg13g2_fill_8 FILLER_10_537 ();
 sg13g2_fill_8 FILLER_10_545 ();
 sg13g2_fill_8 FILLER_10_553 ();
 sg13g2_fill_8 FILLER_10_561 ();
 sg13g2_fill_8 FILLER_10_569 ();
 sg13g2_fill_8 FILLER_10_577 ();
 sg13g2_fill_8 FILLER_10_585 ();
 sg13g2_fill_8 FILLER_10_593 ();
 sg13g2_fill_8 FILLER_10_601 ();
 sg13g2_fill_8 FILLER_10_609 ();
 sg13g2_fill_8 FILLER_10_617 ();
 sg13g2_fill_8 FILLER_10_625 ();
 sg13g2_fill_8 FILLER_10_633 ();
 sg13g2_fill_8 FILLER_10_641 ();
 sg13g2_fill_8 FILLER_10_649 ();
 sg13g2_fill_8 FILLER_10_657 ();
 sg13g2_fill_8 FILLER_10_665 ();
 sg13g2_fill_8 FILLER_10_673 ();
 sg13g2_fill_8 FILLER_10_681 ();
 sg13g2_fill_8 FILLER_10_689 ();
 sg13g2_fill_8 FILLER_10_697 ();
 sg13g2_fill_8 FILLER_10_705 ();
 sg13g2_fill_8 FILLER_10_713 ();
 sg13g2_fill_8 FILLER_10_721 ();
 sg13g2_fill_8 FILLER_10_729 ();
 sg13g2_fill_8 FILLER_10_737 ();
 sg13g2_fill_8 FILLER_10_745 ();
 sg13g2_fill_8 FILLER_10_753 ();
 sg13g2_fill_8 FILLER_10_761 ();
 sg13g2_fill_8 FILLER_10_769 ();
 sg13g2_fill_8 FILLER_10_777 ();
 sg13g2_fill_8 FILLER_10_785 ();
 sg13g2_fill_8 FILLER_10_793 ();
 sg13g2_fill_8 FILLER_10_801 ();
 sg13g2_fill_8 FILLER_10_809 ();
 sg13g2_fill_8 FILLER_10_817 ();
 sg13g2_fill_8 FILLER_10_825 ();
 sg13g2_fill_8 FILLER_10_833 ();
 sg13g2_fill_8 FILLER_10_841 ();
 sg13g2_fill_8 FILLER_10_849 ();
 sg13g2_fill_8 FILLER_10_857 ();
 sg13g2_fill_8 FILLER_10_865 ();
 sg13g2_fill_8 FILLER_10_873 ();
 sg13g2_fill_8 FILLER_10_881 ();
 sg13g2_fill_8 FILLER_10_889 ();
 sg13g2_fill_8 FILLER_10_897 ();
 sg13g2_fill_8 FILLER_10_905 ();
 sg13g2_fill_8 FILLER_10_913 ();
 sg13g2_fill_8 FILLER_10_921 ();
 sg13g2_fill_8 FILLER_10_929 ();
 sg13g2_fill_8 FILLER_10_937 ();
 sg13g2_fill_8 FILLER_10_945 ();
 sg13g2_fill_8 FILLER_10_953 ();
 sg13g2_fill_8 FILLER_10_961 ();
 sg13g2_fill_8 FILLER_10_969 ();
 sg13g2_fill_8 FILLER_10_977 ();
 sg13g2_fill_8 FILLER_10_985 ();
 sg13g2_fill_8 FILLER_10_993 ();
 sg13g2_fill_8 FILLER_10_1001 ();
 sg13g2_fill_8 FILLER_10_1009 ();
 sg13g2_fill_8 FILLER_10_1017 ();
 sg13g2_fill_8 FILLER_10_1025 ();
 sg13g2_fill_8 FILLER_10_1033 ();
 sg13g2_fill_8 FILLER_10_1041 ();
 sg13g2_fill_8 FILLER_10_1049 ();
 sg13g2_fill_8 FILLER_10_1057 ();
 sg13g2_fill_8 FILLER_10_1065 ();
 sg13g2_fill_8 FILLER_10_1073 ();
 sg13g2_fill_8 FILLER_10_1081 ();
 sg13g2_fill_8 FILLER_10_1089 ();
 sg13g2_fill_8 FILLER_10_1097 ();
 sg13g2_fill_8 FILLER_10_1105 ();
 sg13g2_fill_8 FILLER_10_1113 ();
 sg13g2_fill_8 FILLER_10_1121 ();
 sg13g2_fill_8 FILLER_10_1129 ();
 sg13g2_fill_8 FILLER_10_1137 ();
 sg13g2_fill_8 FILLER_10_1145 ();
 sg13g2_fill_8 FILLER_10_1153 ();
 sg13g2_fill_4 FILLER_10_1161 ();
 sg13g2_fill_1 FILLER_10_1165 ();
 sg13g2_fill_8 FILLER_11_0 ();
 sg13g2_fill_8 FILLER_11_8 ();
 sg13g2_fill_8 FILLER_11_16 ();
 sg13g2_fill_8 FILLER_11_24 ();
 sg13g2_fill_8 FILLER_11_32 ();
 sg13g2_fill_8 FILLER_11_40 ();
 sg13g2_fill_8 FILLER_11_48 ();
 sg13g2_fill_1 FILLER_11_82 ();
 sg13g2_fill_8 FILLER_11_125 ();
 sg13g2_fill_8 FILLER_11_133 ();
 sg13g2_fill_2 FILLER_11_141 ();
 sg13g2_fill_4 FILLER_11_188 ();
 sg13g2_fill_2 FILLER_11_192 ();
 sg13g2_fill_8 FILLER_11_199 ();
 sg13g2_fill_4 FILLER_11_258 ();
 sg13g2_fill_8 FILLER_11_283 ();
 sg13g2_fill_8 FILLER_11_291 ();
 sg13g2_fill_2 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_301 ();
 sg13g2_fill_8 FILLER_11_316 ();
 sg13g2_fill_4 FILLER_11_324 ();
 sg13g2_fill_2 FILLER_11_328 ();
 sg13g2_fill_1 FILLER_11_330 ();
 sg13g2_fill_4 FILLER_11_399 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_434 ();
 sg13g2_fill_8 FILLER_11_462 ();
 sg13g2_fill_8 FILLER_11_470 ();
 sg13g2_fill_8 FILLER_11_478 ();
 sg13g2_fill_8 FILLER_11_501 ();
 sg13g2_fill_8 FILLER_11_509 ();
 sg13g2_fill_2 FILLER_11_517 ();
 sg13g2_fill_1 FILLER_11_519 ();
 sg13g2_fill_1 FILLER_11_530 ();
 sg13g2_fill_1 FILLER_11_536 ();
 sg13g2_fill_8 FILLER_11_563 ();
 sg13g2_fill_8 FILLER_11_571 ();
 sg13g2_fill_8 FILLER_11_579 ();
 sg13g2_fill_8 FILLER_11_587 ();
 sg13g2_fill_8 FILLER_11_595 ();
 sg13g2_fill_8 FILLER_11_603 ();
 sg13g2_fill_8 FILLER_11_611 ();
 sg13g2_fill_8 FILLER_11_619 ();
 sg13g2_fill_8 FILLER_11_627 ();
 sg13g2_fill_8 FILLER_11_635 ();
 sg13g2_fill_8 FILLER_11_643 ();
 sg13g2_fill_8 FILLER_11_651 ();
 sg13g2_fill_8 FILLER_11_659 ();
 sg13g2_fill_8 FILLER_11_667 ();
 sg13g2_fill_8 FILLER_11_675 ();
 sg13g2_fill_8 FILLER_11_683 ();
 sg13g2_fill_8 FILLER_11_691 ();
 sg13g2_fill_8 FILLER_11_699 ();
 sg13g2_fill_8 FILLER_11_707 ();
 sg13g2_fill_8 FILLER_11_715 ();
 sg13g2_fill_8 FILLER_11_723 ();
 sg13g2_fill_8 FILLER_11_731 ();
 sg13g2_fill_8 FILLER_11_739 ();
 sg13g2_fill_8 FILLER_11_747 ();
 sg13g2_fill_8 FILLER_11_755 ();
 sg13g2_fill_8 FILLER_11_763 ();
 sg13g2_fill_8 FILLER_11_771 ();
 sg13g2_fill_8 FILLER_11_779 ();
 sg13g2_fill_8 FILLER_11_787 ();
 sg13g2_fill_8 FILLER_11_795 ();
 sg13g2_fill_8 FILLER_11_803 ();
 sg13g2_fill_8 FILLER_11_811 ();
 sg13g2_fill_8 FILLER_11_819 ();
 sg13g2_fill_8 FILLER_11_827 ();
 sg13g2_fill_8 FILLER_11_835 ();
 sg13g2_fill_8 FILLER_11_843 ();
 sg13g2_fill_8 FILLER_11_851 ();
 sg13g2_fill_8 FILLER_11_859 ();
 sg13g2_fill_8 FILLER_11_867 ();
 sg13g2_fill_8 FILLER_11_875 ();
 sg13g2_fill_8 FILLER_11_883 ();
 sg13g2_fill_8 FILLER_11_891 ();
 sg13g2_fill_8 FILLER_11_899 ();
 sg13g2_fill_8 FILLER_11_907 ();
 sg13g2_fill_8 FILLER_11_915 ();
 sg13g2_fill_8 FILLER_11_923 ();
 sg13g2_fill_8 FILLER_11_931 ();
 sg13g2_fill_8 FILLER_11_939 ();
 sg13g2_fill_8 FILLER_11_947 ();
 sg13g2_fill_8 FILLER_11_955 ();
 sg13g2_fill_8 FILLER_11_963 ();
 sg13g2_fill_8 FILLER_11_971 ();
 sg13g2_fill_8 FILLER_11_979 ();
 sg13g2_fill_8 FILLER_11_987 ();
 sg13g2_fill_8 FILLER_11_995 ();
 sg13g2_fill_8 FILLER_11_1003 ();
 sg13g2_fill_8 FILLER_11_1011 ();
 sg13g2_fill_8 FILLER_11_1019 ();
 sg13g2_fill_8 FILLER_11_1027 ();
 sg13g2_fill_8 FILLER_11_1035 ();
 sg13g2_fill_8 FILLER_11_1043 ();
 sg13g2_fill_8 FILLER_11_1051 ();
 sg13g2_fill_8 FILLER_11_1059 ();
 sg13g2_fill_8 FILLER_11_1067 ();
 sg13g2_fill_8 FILLER_11_1075 ();
 sg13g2_fill_8 FILLER_11_1083 ();
 sg13g2_fill_8 FILLER_11_1091 ();
 sg13g2_fill_8 FILLER_11_1099 ();
 sg13g2_fill_8 FILLER_11_1107 ();
 sg13g2_fill_8 FILLER_11_1115 ();
 sg13g2_fill_8 FILLER_11_1123 ();
 sg13g2_fill_8 FILLER_11_1131 ();
 sg13g2_fill_8 FILLER_11_1139 ();
 sg13g2_fill_8 FILLER_11_1147 ();
 sg13g2_fill_8 FILLER_11_1155 ();
 sg13g2_fill_2 FILLER_11_1163 ();
 sg13g2_fill_1 FILLER_11_1165 ();
 sg13g2_fill_8 FILLER_12_0 ();
 sg13g2_fill_8 FILLER_12_8 ();
 sg13g2_fill_8 FILLER_12_16 ();
 sg13g2_fill_8 FILLER_12_24 ();
 sg13g2_fill_4 FILLER_12_32 ();
 sg13g2_fill_2 FILLER_12_36 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_96 ();
 sg13g2_fill_2 FILLER_12_103 ();
 sg13g2_fill_8 FILLER_12_108 ();
 sg13g2_fill_8 FILLER_12_116 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_8 FILLER_12_245 ();
 sg13g2_fill_8 FILLER_12_253 ();
 sg13g2_fill_4 FILLER_12_261 ();
 sg13g2_fill_8 FILLER_12_286 ();
 sg13g2_fill_8 FILLER_12_294 ();
 sg13g2_fill_8 FILLER_12_310 ();
 sg13g2_fill_8 FILLER_12_318 ();
 sg13g2_fill_8 FILLER_12_326 ();
 sg13g2_fill_8 FILLER_12_334 ();
 sg13g2_fill_1 FILLER_12_342 ();
 sg13g2_fill_2 FILLER_12_402 ();
 sg13g2_fill_2 FILLER_12_414 ();
 sg13g2_fill_8 FILLER_12_419 ();
 sg13g2_fill_2 FILLER_12_469 ();
 sg13g2_fill_8 FILLER_12_505 ();
 sg13g2_fill_4 FILLER_12_513 ();
 sg13g2_fill_2 FILLER_12_527 ();
 sg13g2_fill_1 FILLER_12_529 ();
 sg13g2_fill_8 FILLER_12_561 ();
 sg13g2_fill_8 FILLER_12_569 ();
 sg13g2_fill_8 FILLER_12_577 ();
 sg13g2_fill_8 FILLER_12_585 ();
 sg13g2_fill_8 FILLER_12_593 ();
 sg13g2_fill_8 FILLER_12_601 ();
 sg13g2_fill_8 FILLER_12_609 ();
 sg13g2_fill_8 FILLER_12_617 ();
 sg13g2_fill_8 FILLER_12_625 ();
 sg13g2_fill_8 FILLER_12_633 ();
 sg13g2_fill_8 FILLER_12_641 ();
 sg13g2_fill_8 FILLER_12_649 ();
 sg13g2_fill_8 FILLER_12_657 ();
 sg13g2_fill_8 FILLER_12_665 ();
 sg13g2_fill_8 FILLER_12_673 ();
 sg13g2_fill_8 FILLER_12_681 ();
 sg13g2_fill_8 FILLER_12_689 ();
 sg13g2_fill_8 FILLER_12_697 ();
 sg13g2_fill_8 FILLER_12_705 ();
 sg13g2_fill_8 FILLER_12_713 ();
 sg13g2_fill_8 FILLER_12_721 ();
 sg13g2_fill_8 FILLER_12_729 ();
 sg13g2_fill_8 FILLER_12_737 ();
 sg13g2_fill_8 FILLER_12_745 ();
 sg13g2_fill_8 FILLER_12_753 ();
 sg13g2_fill_8 FILLER_12_761 ();
 sg13g2_fill_8 FILLER_12_769 ();
 sg13g2_fill_8 FILLER_12_777 ();
 sg13g2_fill_8 FILLER_12_785 ();
 sg13g2_fill_8 FILLER_12_793 ();
 sg13g2_fill_8 FILLER_12_801 ();
 sg13g2_fill_8 FILLER_12_809 ();
 sg13g2_fill_8 FILLER_12_817 ();
 sg13g2_fill_8 FILLER_12_825 ();
 sg13g2_fill_8 FILLER_12_833 ();
 sg13g2_fill_8 FILLER_12_841 ();
 sg13g2_fill_8 FILLER_12_849 ();
 sg13g2_fill_8 FILLER_12_857 ();
 sg13g2_fill_8 FILLER_12_865 ();
 sg13g2_fill_8 FILLER_12_873 ();
 sg13g2_fill_8 FILLER_12_881 ();
 sg13g2_fill_8 FILLER_12_889 ();
 sg13g2_fill_8 FILLER_12_897 ();
 sg13g2_fill_8 FILLER_12_905 ();
 sg13g2_fill_8 FILLER_12_913 ();
 sg13g2_fill_8 FILLER_12_921 ();
 sg13g2_fill_8 FILLER_12_929 ();
 sg13g2_fill_8 FILLER_12_937 ();
 sg13g2_fill_8 FILLER_12_945 ();
 sg13g2_fill_8 FILLER_12_953 ();
 sg13g2_fill_8 FILLER_12_961 ();
 sg13g2_fill_8 FILLER_12_969 ();
 sg13g2_fill_8 FILLER_12_977 ();
 sg13g2_fill_8 FILLER_12_985 ();
 sg13g2_fill_8 FILLER_12_993 ();
 sg13g2_fill_8 FILLER_12_1001 ();
 sg13g2_fill_8 FILLER_12_1009 ();
 sg13g2_fill_8 FILLER_12_1017 ();
 sg13g2_fill_8 FILLER_12_1025 ();
 sg13g2_fill_8 FILLER_12_1033 ();
 sg13g2_fill_8 FILLER_12_1041 ();
 sg13g2_fill_8 FILLER_12_1049 ();
 sg13g2_fill_8 FILLER_12_1057 ();
 sg13g2_fill_8 FILLER_12_1065 ();
 sg13g2_fill_8 FILLER_12_1073 ();
 sg13g2_fill_8 FILLER_12_1081 ();
 sg13g2_fill_8 FILLER_12_1089 ();
 sg13g2_fill_8 FILLER_12_1097 ();
 sg13g2_fill_8 FILLER_12_1105 ();
 sg13g2_fill_8 FILLER_12_1113 ();
 sg13g2_fill_8 FILLER_12_1121 ();
 sg13g2_fill_8 FILLER_12_1129 ();
 sg13g2_fill_8 FILLER_12_1137 ();
 sg13g2_fill_8 FILLER_12_1145 ();
 sg13g2_fill_8 FILLER_12_1153 ();
 sg13g2_fill_4 FILLER_12_1161 ();
 sg13g2_fill_1 FILLER_12_1165 ();
 sg13g2_fill_8 FILLER_13_0 ();
 sg13g2_fill_8 FILLER_13_8 ();
 sg13g2_fill_8 FILLER_13_16 ();
 sg13g2_fill_2 FILLER_13_24 ();
 sg13g2_fill_1 FILLER_13_26 ();
 sg13g2_fill_4 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_97 ();
 sg13g2_fill_8 FILLER_13_119 ();
 sg13g2_fill_8 FILLER_13_127 ();
 sg13g2_fill_8 FILLER_13_135 ();
 sg13g2_fill_8 FILLER_13_143 ();
 sg13g2_fill_8 FILLER_13_151 ();
 sg13g2_fill_8 FILLER_13_159 ();
 sg13g2_fill_8 FILLER_13_167 ();
 sg13g2_fill_8 FILLER_13_175 ();
 sg13g2_fill_8 FILLER_13_183 ();
 sg13g2_fill_4 FILLER_13_191 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_4 FILLER_13_237 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_8 FILLER_13_346 ();
 sg13g2_fill_4 FILLER_13_354 ();
 sg13g2_fill_2 FILLER_13_358 ();
 sg13g2_fill_1 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_399 ();
 sg13g2_fill_4 FILLER_13_432 ();
 sg13g2_fill_2 FILLER_13_436 ();
 sg13g2_fill_4 FILLER_13_459 ();
 sg13g2_fill_8 FILLER_13_515 ();
 sg13g2_fill_8 FILLER_13_523 ();
 sg13g2_fill_2 FILLER_13_537 ();
 sg13g2_fill_8 FILLER_13_570 ();
 sg13g2_fill_8 FILLER_13_578 ();
 sg13g2_fill_8 FILLER_13_586 ();
 sg13g2_fill_8 FILLER_13_594 ();
 sg13g2_fill_8 FILLER_13_602 ();
 sg13g2_fill_8 FILLER_13_610 ();
 sg13g2_fill_8 FILLER_13_618 ();
 sg13g2_fill_8 FILLER_13_626 ();
 sg13g2_fill_8 FILLER_13_634 ();
 sg13g2_fill_8 FILLER_13_642 ();
 sg13g2_fill_8 FILLER_13_650 ();
 sg13g2_fill_8 FILLER_13_658 ();
 sg13g2_fill_8 FILLER_13_666 ();
 sg13g2_fill_8 FILLER_13_674 ();
 sg13g2_fill_8 FILLER_13_682 ();
 sg13g2_fill_8 FILLER_13_690 ();
 sg13g2_fill_8 FILLER_13_698 ();
 sg13g2_fill_8 FILLER_13_706 ();
 sg13g2_fill_8 FILLER_13_714 ();
 sg13g2_fill_8 FILLER_13_722 ();
 sg13g2_fill_8 FILLER_13_730 ();
 sg13g2_fill_8 FILLER_13_738 ();
 sg13g2_fill_8 FILLER_13_746 ();
 sg13g2_fill_8 FILLER_13_754 ();
 sg13g2_fill_8 FILLER_13_762 ();
 sg13g2_fill_8 FILLER_13_770 ();
 sg13g2_fill_8 FILLER_13_778 ();
 sg13g2_fill_8 FILLER_13_786 ();
 sg13g2_fill_8 FILLER_13_794 ();
 sg13g2_fill_8 FILLER_13_802 ();
 sg13g2_fill_8 FILLER_13_810 ();
 sg13g2_fill_8 FILLER_13_818 ();
 sg13g2_fill_8 FILLER_13_826 ();
 sg13g2_fill_8 FILLER_13_834 ();
 sg13g2_fill_8 FILLER_13_842 ();
 sg13g2_fill_8 FILLER_13_850 ();
 sg13g2_fill_8 FILLER_13_858 ();
 sg13g2_fill_8 FILLER_13_866 ();
 sg13g2_fill_8 FILLER_13_874 ();
 sg13g2_fill_8 FILLER_13_882 ();
 sg13g2_fill_8 FILLER_13_890 ();
 sg13g2_fill_8 FILLER_13_898 ();
 sg13g2_fill_8 FILLER_13_906 ();
 sg13g2_fill_8 FILLER_13_914 ();
 sg13g2_fill_8 FILLER_13_922 ();
 sg13g2_fill_8 FILLER_13_930 ();
 sg13g2_fill_8 FILLER_13_938 ();
 sg13g2_fill_8 FILLER_13_946 ();
 sg13g2_fill_8 FILLER_13_954 ();
 sg13g2_fill_8 FILLER_13_962 ();
 sg13g2_fill_8 FILLER_13_970 ();
 sg13g2_fill_8 FILLER_13_978 ();
 sg13g2_fill_8 FILLER_13_986 ();
 sg13g2_fill_8 FILLER_13_994 ();
 sg13g2_fill_8 FILLER_13_1002 ();
 sg13g2_fill_8 FILLER_13_1010 ();
 sg13g2_fill_8 FILLER_13_1018 ();
 sg13g2_fill_8 FILLER_13_1026 ();
 sg13g2_fill_8 FILLER_13_1034 ();
 sg13g2_fill_8 FILLER_13_1042 ();
 sg13g2_fill_8 FILLER_13_1050 ();
 sg13g2_fill_8 FILLER_13_1058 ();
 sg13g2_fill_8 FILLER_13_1066 ();
 sg13g2_fill_8 FILLER_13_1074 ();
 sg13g2_fill_8 FILLER_13_1082 ();
 sg13g2_fill_8 FILLER_13_1090 ();
 sg13g2_fill_8 FILLER_13_1098 ();
 sg13g2_fill_8 FILLER_13_1106 ();
 sg13g2_fill_8 FILLER_13_1114 ();
 sg13g2_fill_8 FILLER_13_1122 ();
 sg13g2_fill_8 FILLER_13_1130 ();
 sg13g2_fill_8 FILLER_13_1138 ();
 sg13g2_fill_8 FILLER_13_1146 ();
 sg13g2_fill_8 FILLER_13_1154 ();
 sg13g2_fill_4 FILLER_13_1162 ();
 sg13g2_fill_8 FILLER_14_0 ();
 sg13g2_fill_8 FILLER_14_8 ();
 sg13g2_fill_8 FILLER_14_16 ();
 sg13g2_fill_8 FILLER_14_24 ();
 sg13g2_fill_8 FILLER_14_32 ();
 sg13g2_fill_8 FILLER_14_40 ();
 sg13g2_fill_8 FILLER_14_48 ();
 sg13g2_fill_2 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_58 ();
 sg13g2_fill_4 FILLER_14_62 ();
 sg13g2_fill_1 FILLER_14_104 ();
 sg13g2_fill_8 FILLER_14_126 ();
 sg13g2_fill_4 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_fill_8 FILLER_14_188 ();
 sg13g2_fill_8 FILLER_14_196 ();
 sg13g2_fill_8 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_fill_8 FILLER_14_222 ();
 sg13g2_fill_4 FILLER_14_230 ();
 sg13g2_fill_2 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_242 ();
 sg13g2_fill_8 FILLER_14_249 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_fill_2 FILLER_14_300 ();
 sg13g2_fill_1 FILLER_14_302 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_fill_8 FILLER_14_380 ();
 sg13g2_fill_8 FILLER_14_388 ();
 sg13g2_fill_4 FILLER_14_396 ();
 sg13g2_fill_2 FILLER_14_400 ();
 sg13g2_fill_1 FILLER_14_402 ();
 sg13g2_fill_8 FILLER_14_408 ();
 sg13g2_fill_8 FILLER_14_416 ();
 sg13g2_fill_2 FILLER_14_453 ();
 sg13g2_fill_1 FILLER_14_455 ();
 sg13g2_fill_1 FILLER_14_466 ();
 sg13g2_fill_8 FILLER_14_481 ();
 sg13g2_fill_1 FILLER_14_489 ();
 sg13g2_fill_8 FILLER_14_532 ();
 sg13g2_fill_8 FILLER_14_540 ();
 sg13g2_fill_8 FILLER_14_584 ();
 sg13g2_fill_8 FILLER_14_592 ();
 sg13g2_fill_8 FILLER_14_600 ();
 sg13g2_fill_8 FILLER_14_608 ();
 sg13g2_fill_8 FILLER_14_616 ();
 sg13g2_fill_8 FILLER_14_624 ();
 sg13g2_fill_8 FILLER_14_632 ();
 sg13g2_fill_8 FILLER_14_640 ();
 sg13g2_fill_8 FILLER_14_648 ();
 sg13g2_fill_8 FILLER_14_656 ();
 sg13g2_fill_8 FILLER_14_664 ();
 sg13g2_fill_8 FILLER_14_672 ();
 sg13g2_fill_8 FILLER_14_680 ();
 sg13g2_fill_8 FILLER_14_688 ();
 sg13g2_fill_8 FILLER_14_696 ();
 sg13g2_fill_8 FILLER_14_704 ();
 sg13g2_fill_8 FILLER_14_712 ();
 sg13g2_fill_8 FILLER_14_720 ();
 sg13g2_fill_8 FILLER_14_728 ();
 sg13g2_fill_8 FILLER_14_736 ();
 sg13g2_fill_8 FILLER_14_744 ();
 sg13g2_fill_8 FILLER_14_752 ();
 sg13g2_fill_8 FILLER_14_760 ();
 sg13g2_fill_8 FILLER_14_768 ();
 sg13g2_fill_8 FILLER_14_776 ();
 sg13g2_fill_8 FILLER_14_784 ();
 sg13g2_fill_8 FILLER_14_792 ();
 sg13g2_fill_8 FILLER_14_800 ();
 sg13g2_fill_8 FILLER_14_808 ();
 sg13g2_fill_8 FILLER_14_816 ();
 sg13g2_fill_8 FILLER_14_824 ();
 sg13g2_fill_8 FILLER_14_832 ();
 sg13g2_fill_8 FILLER_14_840 ();
 sg13g2_fill_8 FILLER_14_848 ();
 sg13g2_fill_8 FILLER_14_856 ();
 sg13g2_fill_8 FILLER_14_864 ();
 sg13g2_fill_8 FILLER_14_872 ();
 sg13g2_fill_8 FILLER_14_880 ();
 sg13g2_fill_8 FILLER_14_888 ();
 sg13g2_fill_8 FILLER_14_896 ();
 sg13g2_fill_8 FILLER_14_904 ();
 sg13g2_fill_8 FILLER_14_912 ();
 sg13g2_fill_8 FILLER_14_920 ();
 sg13g2_fill_8 FILLER_14_928 ();
 sg13g2_fill_8 FILLER_14_936 ();
 sg13g2_fill_8 FILLER_14_944 ();
 sg13g2_fill_8 FILLER_14_952 ();
 sg13g2_fill_8 FILLER_14_960 ();
 sg13g2_fill_8 FILLER_14_968 ();
 sg13g2_fill_8 FILLER_14_976 ();
 sg13g2_fill_8 FILLER_14_984 ();
 sg13g2_fill_8 FILLER_14_992 ();
 sg13g2_fill_8 FILLER_14_1000 ();
 sg13g2_fill_8 FILLER_14_1008 ();
 sg13g2_fill_8 FILLER_14_1016 ();
 sg13g2_fill_8 FILLER_14_1024 ();
 sg13g2_fill_8 FILLER_14_1032 ();
 sg13g2_fill_8 FILLER_14_1040 ();
 sg13g2_fill_8 FILLER_14_1048 ();
 sg13g2_fill_8 FILLER_14_1056 ();
 sg13g2_fill_8 FILLER_14_1064 ();
 sg13g2_fill_8 FILLER_14_1072 ();
 sg13g2_fill_8 FILLER_14_1080 ();
 sg13g2_fill_8 FILLER_14_1088 ();
 sg13g2_fill_8 FILLER_14_1096 ();
 sg13g2_fill_8 FILLER_14_1104 ();
 sg13g2_fill_8 FILLER_14_1112 ();
 sg13g2_fill_8 FILLER_14_1120 ();
 sg13g2_fill_8 FILLER_14_1128 ();
 sg13g2_fill_8 FILLER_14_1136 ();
 sg13g2_fill_8 FILLER_14_1144 ();
 sg13g2_fill_8 FILLER_14_1152 ();
 sg13g2_fill_4 FILLER_14_1160 ();
 sg13g2_fill_2 FILLER_14_1164 ();
 sg13g2_fill_8 FILLER_15_0 ();
 sg13g2_fill_8 FILLER_15_8 ();
 sg13g2_fill_8 FILLER_15_16 ();
 sg13g2_fill_8 FILLER_15_24 ();
 sg13g2_fill_8 FILLER_15_32 ();
 sg13g2_fill_8 FILLER_15_40 ();
 sg13g2_fill_8 FILLER_15_74 ();
 sg13g2_fill_4 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_fill_4 FILLER_15_135 ();
 sg13g2_fill_2 FILLER_15_139 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_fill_8 FILLER_15_263 ();
 sg13g2_fill_8 FILLER_15_271 ();
 sg13g2_fill_4 FILLER_15_279 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_fill_8 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_4 FILLER_15_357 ();
 sg13g2_fill_1 FILLER_15_361 ();
 sg13g2_fill_8 FILLER_15_392 ();
 sg13g2_fill_8 FILLER_15_400 ();
 sg13g2_fill_8 FILLER_15_408 ();
 sg13g2_fill_8 FILLER_15_416 ();
 sg13g2_fill_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_15_438 ();
 sg13g2_fill_2 FILLER_15_445 ();
 sg13g2_fill_1 FILLER_15_447 ();
 sg13g2_fill_8 FILLER_15_481 ();
 sg13g2_fill_8 FILLER_15_489 ();
 sg13g2_fill_8 FILLER_15_497 ();
 sg13g2_fill_4 FILLER_15_505 ();
 sg13g2_fill_2 FILLER_15_509 ();
 sg13g2_fill_1 FILLER_15_511 ();
 sg13g2_fill_8 FILLER_15_544 ();
 sg13g2_fill_8 FILLER_15_552 ();
 sg13g2_fill_8 FILLER_15_586 ();
 sg13g2_fill_8 FILLER_15_594 ();
 sg13g2_fill_8 FILLER_15_602 ();
 sg13g2_fill_8 FILLER_15_610 ();
 sg13g2_fill_8 FILLER_15_618 ();
 sg13g2_fill_8 FILLER_15_626 ();
 sg13g2_fill_8 FILLER_15_634 ();
 sg13g2_fill_8 FILLER_15_642 ();
 sg13g2_fill_8 FILLER_15_650 ();
 sg13g2_fill_8 FILLER_15_658 ();
 sg13g2_fill_8 FILLER_15_666 ();
 sg13g2_fill_8 FILLER_15_674 ();
 sg13g2_fill_8 FILLER_15_682 ();
 sg13g2_fill_8 FILLER_15_690 ();
 sg13g2_fill_8 FILLER_15_698 ();
 sg13g2_fill_8 FILLER_15_706 ();
 sg13g2_fill_8 FILLER_15_714 ();
 sg13g2_fill_8 FILLER_15_722 ();
 sg13g2_fill_8 FILLER_15_730 ();
 sg13g2_fill_8 FILLER_15_738 ();
 sg13g2_fill_8 FILLER_15_746 ();
 sg13g2_fill_8 FILLER_15_754 ();
 sg13g2_fill_8 FILLER_15_762 ();
 sg13g2_fill_8 FILLER_15_770 ();
 sg13g2_fill_8 FILLER_15_778 ();
 sg13g2_fill_8 FILLER_15_786 ();
 sg13g2_fill_8 FILLER_15_794 ();
 sg13g2_fill_8 FILLER_15_802 ();
 sg13g2_fill_8 FILLER_15_810 ();
 sg13g2_fill_8 FILLER_15_818 ();
 sg13g2_fill_8 FILLER_15_826 ();
 sg13g2_fill_8 FILLER_15_834 ();
 sg13g2_fill_8 FILLER_15_842 ();
 sg13g2_fill_8 FILLER_15_850 ();
 sg13g2_fill_8 FILLER_15_858 ();
 sg13g2_fill_8 FILLER_15_866 ();
 sg13g2_fill_8 FILLER_15_874 ();
 sg13g2_fill_8 FILLER_15_882 ();
 sg13g2_fill_8 FILLER_15_890 ();
 sg13g2_fill_8 FILLER_15_898 ();
 sg13g2_fill_8 FILLER_15_906 ();
 sg13g2_fill_8 FILLER_15_914 ();
 sg13g2_fill_8 FILLER_15_922 ();
 sg13g2_fill_8 FILLER_15_930 ();
 sg13g2_fill_8 FILLER_15_938 ();
 sg13g2_fill_8 FILLER_15_946 ();
 sg13g2_fill_8 FILLER_15_954 ();
 sg13g2_fill_8 FILLER_15_962 ();
 sg13g2_fill_8 FILLER_15_970 ();
 sg13g2_fill_8 FILLER_15_978 ();
 sg13g2_fill_8 FILLER_15_986 ();
 sg13g2_fill_8 FILLER_15_994 ();
 sg13g2_fill_8 FILLER_15_1002 ();
 sg13g2_fill_8 FILLER_15_1010 ();
 sg13g2_fill_8 FILLER_15_1018 ();
 sg13g2_fill_8 FILLER_15_1026 ();
 sg13g2_fill_8 FILLER_15_1034 ();
 sg13g2_fill_8 FILLER_15_1042 ();
 sg13g2_fill_8 FILLER_15_1050 ();
 sg13g2_fill_8 FILLER_15_1058 ();
 sg13g2_fill_8 FILLER_15_1066 ();
 sg13g2_fill_8 FILLER_15_1074 ();
 sg13g2_fill_8 FILLER_15_1082 ();
 sg13g2_fill_8 FILLER_15_1090 ();
 sg13g2_fill_8 FILLER_15_1098 ();
 sg13g2_fill_8 FILLER_15_1106 ();
 sg13g2_fill_8 FILLER_15_1114 ();
 sg13g2_fill_8 FILLER_15_1122 ();
 sg13g2_fill_8 FILLER_15_1130 ();
 sg13g2_fill_8 FILLER_15_1138 ();
 sg13g2_fill_8 FILLER_15_1146 ();
 sg13g2_fill_8 FILLER_15_1154 ();
 sg13g2_fill_4 FILLER_15_1162 ();
 sg13g2_fill_8 FILLER_16_0 ();
 sg13g2_fill_8 FILLER_16_8 ();
 sg13g2_fill_8 FILLER_16_16 ();
 sg13g2_fill_8 FILLER_16_24 ();
 sg13g2_fill_4 FILLER_16_32 ();
 sg13g2_fill_2 FILLER_16_36 ();
 sg13g2_fill_1 FILLER_16_38 ();
 sg13g2_fill_4 FILLER_16_105 ();
 sg13g2_fill_2 FILLER_16_109 ();
 sg13g2_fill_1 FILLER_16_111 ();
 sg13g2_fill_4 FILLER_16_134 ();
 sg13g2_fill_2 FILLER_16_138 ();
 sg13g2_fill_8 FILLER_16_163 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_229 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_246 ();
 sg13g2_fill_8 FILLER_16_273 ();
 sg13g2_fill_8 FILLER_16_281 ();
 sg13g2_fill_8 FILLER_16_289 ();
 sg13g2_fill_4 FILLER_16_297 ();
 sg13g2_fill_8 FILLER_16_310 ();
 sg13g2_fill_8 FILLER_16_318 ();
 sg13g2_fill_4 FILLER_16_326 ();
 sg13g2_fill_2 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_4 FILLER_16_339 ();
 sg13g2_fill_2 FILLER_16_343 ();
 sg13g2_fill_8 FILLER_16_348 ();
 sg13g2_fill_8 FILLER_16_356 ();
 sg13g2_fill_4 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_368 ();
 sg13g2_fill_8 FILLER_16_375 ();
 sg13g2_fill_8 FILLER_16_383 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_4 FILLER_16_418 ();
 sg13g2_fill_2 FILLER_16_422 ();
 sg13g2_fill_8 FILLER_16_427 ();
 sg13g2_fill_8 FILLER_16_435 ();
 sg13g2_fill_8 FILLER_16_443 ();
 sg13g2_fill_2 FILLER_16_451 ();
 sg13g2_fill_4 FILLER_16_458 ();
 sg13g2_fill_2 FILLER_16_462 ();
 sg13g2_fill_4 FILLER_16_490 ();
 sg13g2_fill_2 FILLER_16_494 ();
 sg13g2_fill_1 FILLER_16_496 ();
 sg13g2_fill_8 FILLER_16_518 ();
 sg13g2_fill_4 FILLER_16_526 ();
 sg13g2_fill_2 FILLER_16_551 ();
 sg13g2_fill_1 FILLER_16_568 ();
 sg13g2_fill_8 FILLER_16_600 ();
 sg13g2_fill_8 FILLER_16_608 ();
 sg13g2_fill_8 FILLER_16_616 ();
 sg13g2_fill_8 FILLER_16_624 ();
 sg13g2_fill_8 FILLER_16_632 ();
 sg13g2_fill_8 FILLER_16_640 ();
 sg13g2_fill_8 FILLER_16_648 ();
 sg13g2_fill_8 FILLER_16_656 ();
 sg13g2_fill_8 FILLER_16_664 ();
 sg13g2_fill_8 FILLER_16_672 ();
 sg13g2_fill_8 FILLER_16_680 ();
 sg13g2_fill_8 FILLER_16_688 ();
 sg13g2_fill_8 FILLER_16_696 ();
 sg13g2_fill_8 FILLER_16_704 ();
 sg13g2_fill_8 FILLER_16_712 ();
 sg13g2_fill_8 FILLER_16_720 ();
 sg13g2_fill_8 FILLER_16_728 ();
 sg13g2_fill_8 FILLER_16_736 ();
 sg13g2_fill_8 FILLER_16_744 ();
 sg13g2_fill_8 FILLER_16_752 ();
 sg13g2_fill_8 FILLER_16_760 ();
 sg13g2_fill_8 FILLER_16_768 ();
 sg13g2_fill_8 FILLER_16_776 ();
 sg13g2_fill_8 FILLER_16_784 ();
 sg13g2_fill_8 FILLER_16_792 ();
 sg13g2_fill_8 FILLER_16_800 ();
 sg13g2_fill_8 FILLER_16_808 ();
 sg13g2_fill_8 FILLER_16_816 ();
 sg13g2_fill_8 FILLER_16_824 ();
 sg13g2_fill_8 FILLER_16_832 ();
 sg13g2_fill_8 FILLER_16_840 ();
 sg13g2_fill_8 FILLER_16_848 ();
 sg13g2_fill_8 FILLER_16_856 ();
 sg13g2_fill_8 FILLER_16_864 ();
 sg13g2_fill_8 FILLER_16_872 ();
 sg13g2_fill_8 FILLER_16_880 ();
 sg13g2_fill_8 FILLER_16_888 ();
 sg13g2_fill_8 FILLER_16_896 ();
 sg13g2_fill_8 FILLER_16_904 ();
 sg13g2_fill_8 FILLER_16_912 ();
 sg13g2_fill_8 FILLER_16_920 ();
 sg13g2_fill_8 FILLER_16_928 ();
 sg13g2_fill_8 FILLER_16_936 ();
 sg13g2_fill_8 FILLER_16_944 ();
 sg13g2_fill_8 FILLER_16_952 ();
 sg13g2_fill_8 FILLER_16_960 ();
 sg13g2_fill_8 FILLER_16_968 ();
 sg13g2_fill_8 FILLER_16_976 ();
 sg13g2_fill_8 FILLER_16_984 ();
 sg13g2_fill_8 FILLER_16_992 ();
 sg13g2_fill_8 FILLER_16_1000 ();
 sg13g2_fill_8 FILLER_16_1008 ();
 sg13g2_fill_8 FILLER_16_1016 ();
 sg13g2_fill_8 FILLER_16_1024 ();
 sg13g2_fill_8 FILLER_16_1032 ();
 sg13g2_fill_8 FILLER_16_1040 ();
 sg13g2_fill_8 FILLER_16_1048 ();
 sg13g2_fill_8 FILLER_16_1056 ();
 sg13g2_fill_8 FILLER_16_1064 ();
 sg13g2_fill_8 FILLER_16_1072 ();
 sg13g2_fill_8 FILLER_16_1080 ();
 sg13g2_fill_8 FILLER_16_1088 ();
 sg13g2_fill_8 FILLER_16_1096 ();
 sg13g2_fill_8 FILLER_16_1104 ();
 sg13g2_fill_8 FILLER_16_1112 ();
 sg13g2_fill_8 FILLER_16_1120 ();
 sg13g2_fill_8 FILLER_16_1128 ();
 sg13g2_fill_8 FILLER_16_1136 ();
 sg13g2_fill_8 FILLER_16_1144 ();
 sg13g2_fill_8 FILLER_16_1152 ();
 sg13g2_fill_4 FILLER_16_1160 ();
 sg13g2_fill_2 FILLER_16_1164 ();
 sg13g2_fill_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_8 ();
 sg13g2_fill_2 FILLER_17_35 ();
 sg13g2_fill_1 FILLER_17_37 ();
 sg13g2_fill_8 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_77 ();
 sg13g2_fill_2 FILLER_17_88 ();
 sg13g2_fill_8 FILLER_17_96 ();
 sg13g2_fill_8 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_8 FILLER_17_118 ();
 sg13g2_fill_8 FILLER_17_126 ();
 sg13g2_fill_4 FILLER_17_134 ();
 sg13g2_fill_4 FILLER_17_143 ();
 sg13g2_fill_2 FILLER_17_147 ();
 sg13g2_fill_1 FILLER_17_149 ();
 sg13g2_fill_4 FILLER_17_155 ();
 sg13g2_fill_2 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_fill_8 FILLER_17_174 ();
 sg13g2_fill_1 FILLER_17_182 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_237 ();
 sg13g2_fill_8 FILLER_17_244 ();
 sg13g2_fill_2 FILLER_17_252 ();
 sg13g2_fill_1 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_1 FILLER_17_289 ();
 sg13g2_fill_4 FILLER_17_320 ();
 sg13g2_fill_2 FILLER_17_345 ();
 sg13g2_fill_1 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_1 FILLER_17_378 ();
 sg13g2_fill_2 FILLER_17_394 ();
 sg13g2_fill_4 FILLER_17_456 ();
 sg13g2_fill_4 FILLER_17_501 ();
 sg13g2_fill_2 FILLER_17_505 ();
 sg13g2_fill_8 FILLER_17_528 ();
 sg13g2_fill_2 FILLER_17_536 ();
 sg13g2_fill_2 FILLER_17_569 ();
 sg13g2_fill_2 FILLER_17_576 ();
 sg13g2_fill_8 FILLER_17_583 ();
 sg13g2_fill_8 FILLER_17_591 ();
 sg13g2_fill_8 FILLER_17_599 ();
 sg13g2_fill_8 FILLER_17_607 ();
 sg13g2_fill_8 FILLER_17_615 ();
 sg13g2_fill_8 FILLER_17_623 ();
 sg13g2_fill_8 FILLER_17_631 ();
 sg13g2_fill_8 FILLER_17_639 ();
 sg13g2_fill_8 FILLER_17_647 ();
 sg13g2_fill_8 FILLER_17_655 ();
 sg13g2_fill_8 FILLER_17_663 ();
 sg13g2_fill_8 FILLER_17_671 ();
 sg13g2_fill_8 FILLER_17_679 ();
 sg13g2_fill_8 FILLER_17_687 ();
 sg13g2_fill_8 FILLER_17_695 ();
 sg13g2_fill_8 FILLER_17_703 ();
 sg13g2_fill_8 FILLER_17_711 ();
 sg13g2_fill_8 FILLER_17_719 ();
 sg13g2_fill_8 FILLER_17_727 ();
 sg13g2_fill_8 FILLER_17_735 ();
 sg13g2_fill_8 FILLER_17_743 ();
 sg13g2_fill_8 FILLER_17_751 ();
 sg13g2_fill_8 FILLER_17_759 ();
 sg13g2_fill_8 FILLER_17_767 ();
 sg13g2_fill_8 FILLER_17_775 ();
 sg13g2_fill_8 FILLER_17_783 ();
 sg13g2_fill_8 FILLER_17_791 ();
 sg13g2_fill_8 FILLER_17_799 ();
 sg13g2_fill_8 FILLER_17_807 ();
 sg13g2_fill_8 FILLER_17_815 ();
 sg13g2_fill_8 FILLER_17_823 ();
 sg13g2_fill_8 FILLER_17_831 ();
 sg13g2_fill_8 FILLER_17_839 ();
 sg13g2_fill_8 FILLER_17_847 ();
 sg13g2_fill_8 FILLER_17_855 ();
 sg13g2_fill_8 FILLER_17_863 ();
 sg13g2_fill_8 FILLER_17_871 ();
 sg13g2_fill_8 FILLER_17_879 ();
 sg13g2_fill_8 FILLER_17_887 ();
 sg13g2_fill_8 FILLER_17_895 ();
 sg13g2_fill_8 FILLER_17_903 ();
 sg13g2_fill_8 FILLER_17_911 ();
 sg13g2_fill_8 FILLER_17_919 ();
 sg13g2_fill_8 FILLER_17_927 ();
 sg13g2_fill_8 FILLER_17_935 ();
 sg13g2_fill_8 FILLER_17_943 ();
 sg13g2_fill_8 FILLER_17_951 ();
 sg13g2_fill_8 FILLER_17_959 ();
 sg13g2_fill_8 FILLER_17_967 ();
 sg13g2_fill_8 FILLER_17_975 ();
 sg13g2_fill_8 FILLER_17_983 ();
 sg13g2_fill_8 FILLER_17_991 ();
 sg13g2_fill_8 FILLER_17_999 ();
 sg13g2_fill_8 FILLER_17_1007 ();
 sg13g2_fill_8 FILLER_17_1015 ();
 sg13g2_fill_8 FILLER_17_1023 ();
 sg13g2_fill_8 FILLER_17_1031 ();
 sg13g2_fill_8 FILLER_17_1039 ();
 sg13g2_fill_8 FILLER_17_1047 ();
 sg13g2_fill_8 FILLER_17_1055 ();
 sg13g2_fill_8 FILLER_17_1063 ();
 sg13g2_fill_8 FILLER_17_1071 ();
 sg13g2_fill_8 FILLER_17_1079 ();
 sg13g2_fill_8 FILLER_17_1087 ();
 sg13g2_fill_8 FILLER_17_1095 ();
 sg13g2_fill_8 FILLER_17_1103 ();
 sg13g2_fill_8 FILLER_17_1111 ();
 sg13g2_fill_8 FILLER_17_1119 ();
 sg13g2_fill_8 FILLER_17_1127 ();
 sg13g2_fill_8 FILLER_17_1135 ();
 sg13g2_fill_8 FILLER_17_1143 ();
 sg13g2_fill_8 FILLER_17_1151 ();
 sg13g2_fill_4 FILLER_17_1159 ();
 sg13g2_fill_2 FILLER_17_1163 ();
 sg13g2_fill_1 FILLER_17_1165 ();
 sg13g2_fill_8 FILLER_18_0 ();
 sg13g2_fill_8 FILLER_18_8 ();
 sg13g2_fill_8 FILLER_18_16 ();
 sg13g2_fill_8 FILLER_18_24 ();
 sg13g2_fill_8 FILLER_18_32 ();
 sg13g2_fill_8 FILLER_18_40 ();
 sg13g2_fill_8 FILLER_18_48 ();
 sg13g2_fill_8 FILLER_18_56 ();
 sg13g2_fill_8 FILLER_18_64 ();
 sg13g2_fill_2 FILLER_18_72 ();
 sg13g2_fill_8 FILLER_18_99 ();
 sg13g2_fill_8 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_4 FILLER_18_121 ();
 sg13g2_fill_8 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_4 FILLER_18_220 ();
 sg13g2_fill_8 FILLER_18_228 ();
 sg13g2_fill_8 FILLER_18_236 ();
 sg13g2_fill_4 FILLER_18_244 ();
 sg13g2_fill_4 FILLER_18_251 ();
 sg13g2_fill_8 FILLER_18_260 ();
 sg13g2_fill_8 FILLER_18_268 ();
 sg13g2_fill_8 FILLER_18_276 ();
 sg13g2_fill_8 FILLER_18_284 ();
 sg13g2_fill_4 FILLER_18_292 ();
 sg13g2_fill_8 FILLER_18_351 ();
 sg13g2_fill_4 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_fill_4 FILLER_18_419 ();
 sg13g2_fill_4 FILLER_18_433 ();
 sg13g2_fill_4 FILLER_18_440 ();
 sg13g2_fill_4 FILLER_18_470 ();
 sg13g2_fill_1 FILLER_18_477 ();
 sg13g2_fill_2 FILLER_18_483 ();
 sg13g2_fill_8 FILLER_18_530 ();
 sg13g2_fill_4 FILLER_18_542 ();
 sg13g2_fill_8 FILLER_18_552 ();
 sg13g2_fill_8 FILLER_18_560 ();
 sg13g2_fill_8 FILLER_18_602 ();
 sg13g2_fill_8 FILLER_18_610 ();
 sg13g2_fill_8 FILLER_18_618 ();
 sg13g2_fill_8 FILLER_18_626 ();
 sg13g2_fill_8 FILLER_18_634 ();
 sg13g2_fill_8 FILLER_18_642 ();
 sg13g2_fill_8 FILLER_18_650 ();
 sg13g2_fill_8 FILLER_18_658 ();
 sg13g2_fill_8 FILLER_18_666 ();
 sg13g2_fill_8 FILLER_18_674 ();
 sg13g2_fill_8 FILLER_18_682 ();
 sg13g2_fill_8 FILLER_18_690 ();
 sg13g2_fill_8 FILLER_18_698 ();
 sg13g2_fill_8 FILLER_18_706 ();
 sg13g2_fill_8 FILLER_18_714 ();
 sg13g2_fill_8 FILLER_18_722 ();
 sg13g2_fill_8 FILLER_18_730 ();
 sg13g2_fill_8 FILLER_18_738 ();
 sg13g2_fill_8 FILLER_18_746 ();
 sg13g2_fill_8 FILLER_18_754 ();
 sg13g2_fill_8 FILLER_18_762 ();
 sg13g2_fill_8 FILLER_18_770 ();
 sg13g2_fill_8 FILLER_18_778 ();
 sg13g2_fill_8 FILLER_18_786 ();
 sg13g2_fill_8 FILLER_18_794 ();
 sg13g2_fill_8 FILLER_18_802 ();
 sg13g2_fill_8 FILLER_18_810 ();
 sg13g2_fill_8 FILLER_18_818 ();
 sg13g2_fill_8 FILLER_18_826 ();
 sg13g2_fill_8 FILLER_18_834 ();
 sg13g2_fill_8 FILLER_18_842 ();
 sg13g2_fill_8 FILLER_18_850 ();
 sg13g2_fill_8 FILLER_18_858 ();
 sg13g2_fill_8 FILLER_18_866 ();
 sg13g2_fill_8 FILLER_18_874 ();
 sg13g2_fill_8 FILLER_18_882 ();
 sg13g2_fill_8 FILLER_18_890 ();
 sg13g2_fill_8 FILLER_18_898 ();
 sg13g2_fill_8 FILLER_18_906 ();
 sg13g2_fill_8 FILLER_18_914 ();
 sg13g2_fill_8 FILLER_18_922 ();
 sg13g2_fill_8 FILLER_18_930 ();
 sg13g2_fill_8 FILLER_18_938 ();
 sg13g2_fill_8 FILLER_18_946 ();
 sg13g2_fill_8 FILLER_18_954 ();
 sg13g2_fill_8 FILLER_18_962 ();
 sg13g2_fill_8 FILLER_18_970 ();
 sg13g2_fill_8 FILLER_18_978 ();
 sg13g2_fill_8 FILLER_18_986 ();
 sg13g2_fill_8 FILLER_18_994 ();
 sg13g2_fill_8 FILLER_18_1002 ();
 sg13g2_fill_8 FILLER_18_1010 ();
 sg13g2_fill_8 FILLER_18_1018 ();
 sg13g2_fill_8 FILLER_18_1026 ();
 sg13g2_fill_8 FILLER_18_1034 ();
 sg13g2_fill_8 FILLER_18_1042 ();
 sg13g2_fill_8 FILLER_18_1050 ();
 sg13g2_fill_8 FILLER_18_1058 ();
 sg13g2_fill_8 FILLER_18_1066 ();
 sg13g2_fill_8 FILLER_18_1074 ();
 sg13g2_fill_8 FILLER_18_1082 ();
 sg13g2_fill_8 FILLER_18_1090 ();
 sg13g2_fill_8 FILLER_18_1098 ();
 sg13g2_fill_8 FILLER_18_1106 ();
 sg13g2_fill_8 FILLER_18_1114 ();
 sg13g2_fill_8 FILLER_18_1122 ();
 sg13g2_fill_8 FILLER_18_1130 ();
 sg13g2_fill_8 FILLER_18_1138 ();
 sg13g2_fill_8 FILLER_18_1146 ();
 sg13g2_fill_8 FILLER_18_1154 ();
 sg13g2_fill_4 FILLER_18_1162 ();
 sg13g2_fill_8 FILLER_19_0 ();
 sg13g2_fill_8 FILLER_19_8 ();
 sg13g2_fill_8 FILLER_19_16 ();
 sg13g2_fill_4 FILLER_19_24 ();
 sg13g2_fill_4 FILLER_19_65 ();
 sg13g2_fill_2 FILLER_19_69 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_fill_4 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_104 ();
 sg13g2_fill_1 FILLER_19_110 ();
 sg13g2_fill_8 FILLER_19_141 ();
 sg13g2_fill_4 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_fill_2 FILLER_19_186 ();
 sg13g2_fill_2 FILLER_19_217 ();
 sg13g2_fill_4 FILLER_19_227 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_fill_1 FILLER_19_233 ();
 sg13g2_fill_2 FILLER_19_239 ();
 sg13g2_fill_8 FILLER_19_247 ();
 sg13g2_fill_4 FILLER_19_255 ();
 sg13g2_fill_8 FILLER_19_285 ();
 sg13g2_fill_8 FILLER_19_293 ();
 sg13g2_fill_4 FILLER_19_301 ();
 sg13g2_fill_2 FILLER_19_305 ();
 sg13g2_fill_4 FILLER_19_313 ();
 sg13g2_fill_2 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_319 ();
 sg13g2_fill_8 FILLER_19_333 ();
 sg13g2_fill_4 FILLER_19_341 ();
 sg13g2_fill_2 FILLER_19_345 ();
 sg13g2_fill_1 FILLER_19_347 ();
 sg13g2_fill_8 FILLER_19_353 ();
 sg13g2_fill_8 FILLER_19_461 ();
 sg13g2_fill_8 FILLER_19_469 ();
 sg13g2_fill_8 FILLER_19_477 ();
 sg13g2_fill_8 FILLER_19_485 ();
 sg13g2_fill_4 FILLER_19_493 ();
 sg13g2_fill_8 FILLER_19_505 ();
 sg13g2_fill_2 FILLER_19_513 ();
 sg13g2_fill_8 FILLER_19_526 ();
 sg13g2_fill_8 FILLER_19_534 ();
 sg13g2_fill_8 FILLER_19_542 ();
 sg13g2_fill_8 FILLER_19_550 ();
 sg13g2_fill_8 FILLER_19_558 ();
 sg13g2_fill_4 FILLER_19_566 ();
 sg13g2_fill_8 FILLER_19_595 ();
 sg13g2_fill_8 FILLER_19_603 ();
 sg13g2_fill_8 FILLER_19_611 ();
 sg13g2_fill_8 FILLER_19_619 ();
 sg13g2_fill_8 FILLER_19_627 ();
 sg13g2_fill_8 FILLER_19_635 ();
 sg13g2_fill_8 FILLER_19_643 ();
 sg13g2_fill_8 FILLER_19_651 ();
 sg13g2_fill_8 FILLER_19_659 ();
 sg13g2_fill_8 FILLER_19_667 ();
 sg13g2_fill_8 FILLER_19_675 ();
 sg13g2_fill_8 FILLER_19_683 ();
 sg13g2_fill_8 FILLER_19_691 ();
 sg13g2_fill_8 FILLER_19_699 ();
 sg13g2_fill_8 FILLER_19_707 ();
 sg13g2_fill_8 FILLER_19_715 ();
 sg13g2_fill_8 FILLER_19_723 ();
 sg13g2_fill_8 FILLER_19_731 ();
 sg13g2_fill_8 FILLER_19_739 ();
 sg13g2_fill_8 FILLER_19_747 ();
 sg13g2_fill_8 FILLER_19_755 ();
 sg13g2_fill_8 FILLER_19_763 ();
 sg13g2_fill_8 FILLER_19_771 ();
 sg13g2_fill_8 FILLER_19_779 ();
 sg13g2_fill_8 FILLER_19_787 ();
 sg13g2_fill_8 FILLER_19_795 ();
 sg13g2_fill_8 FILLER_19_803 ();
 sg13g2_fill_8 FILLER_19_811 ();
 sg13g2_fill_8 FILLER_19_819 ();
 sg13g2_fill_8 FILLER_19_827 ();
 sg13g2_fill_8 FILLER_19_835 ();
 sg13g2_fill_8 FILLER_19_843 ();
 sg13g2_fill_8 FILLER_19_851 ();
 sg13g2_fill_8 FILLER_19_859 ();
 sg13g2_fill_8 FILLER_19_867 ();
 sg13g2_fill_8 FILLER_19_875 ();
 sg13g2_fill_8 FILLER_19_883 ();
 sg13g2_fill_8 FILLER_19_891 ();
 sg13g2_fill_8 FILLER_19_899 ();
 sg13g2_fill_8 FILLER_19_907 ();
 sg13g2_fill_8 FILLER_19_915 ();
 sg13g2_fill_8 FILLER_19_923 ();
 sg13g2_fill_8 FILLER_19_931 ();
 sg13g2_fill_8 FILLER_19_939 ();
 sg13g2_fill_8 FILLER_19_947 ();
 sg13g2_fill_8 FILLER_19_955 ();
 sg13g2_fill_8 FILLER_19_963 ();
 sg13g2_fill_8 FILLER_19_971 ();
 sg13g2_fill_8 FILLER_19_979 ();
 sg13g2_fill_8 FILLER_19_987 ();
 sg13g2_fill_8 FILLER_19_995 ();
 sg13g2_fill_8 FILLER_19_1003 ();
 sg13g2_fill_8 FILLER_19_1011 ();
 sg13g2_fill_8 FILLER_19_1019 ();
 sg13g2_fill_8 FILLER_19_1027 ();
 sg13g2_fill_8 FILLER_19_1035 ();
 sg13g2_fill_8 FILLER_19_1043 ();
 sg13g2_fill_8 FILLER_19_1051 ();
 sg13g2_fill_8 FILLER_19_1059 ();
 sg13g2_fill_8 FILLER_19_1067 ();
 sg13g2_fill_8 FILLER_19_1075 ();
 sg13g2_fill_8 FILLER_19_1083 ();
 sg13g2_fill_8 FILLER_19_1091 ();
 sg13g2_fill_8 FILLER_19_1099 ();
 sg13g2_fill_8 FILLER_19_1107 ();
 sg13g2_fill_8 FILLER_19_1115 ();
 sg13g2_fill_8 FILLER_19_1123 ();
 sg13g2_fill_8 FILLER_19_1131 ();
 sg13g2_fill_8 FILLER_19_1139 ();
 sg13g2_fill_8 FILLER_19_1147 ();
 sg13g2_fill_8 FILLER_19_1155 ();
 sg13g2_fill_2 FILLER_19_1163 ();
 sg13g2_fill_1 FILLER_19_1165 ();
 sg13g2_fill_8 FILLER_20_0 ();
 sg13g2_fill_8 FILLER_20_8 ();
 sg13g2_fill_8 FILLER_20_16 ();
 sg13g2_fill_4 FILLER_20_24 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_8 FILLER_20_184 ();
 sg13g2_fill_4 FILLER_20_192 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_198 ();
 sg13g2_fill_4 FILLER_20_203 ();
 sg13g2_fill_1 FILLER_20_207 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_fill_4 FILLER_20_241 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_8 FILLER_20_289 ();
 sg13g2_fill_8 FILLER_20_297 ();
 sg13g2_fill_8 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_313 ();
 sg13g2_fill_4 FILLER_20_326 ();
 sg13g2_fill_2 FILLER_20_335 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_fill_8 FILLER_20_372 ();
 sg13g2_fill_8 FILLER_20_380 ();
 sg13g2_fill_8 FILLER_20_388 ();
 sg13g2_fill_2 FILLER_20_396 ();
 sg13g2_fill_1 FILLER_20_398 ();
 sg13g2_fill_4 FILLER_20_403 ();
 sg13g2_fill_1 FILLER_20_407 ();
 sg13g2_fill_8 FILLER_20_414 ();
 sg13g2_fill_1 FILLER_20_422 ();
 sg13g2_fill_2 FILLER_20_443 ();
 sg13g2_fill_8 FILLER_20_470 ();
 sg13g2_fill_4 FILLER_20_478 ();
 sg13g2_fill_1 FILLER_20_482 ();
 sg13g2_fill_2 FILLER_20_488 ();
 sg13g2_fill_8 FILLER_20_494 ();
 sg13g2_fill_8 FILLER_20_502 ();
 sg13g2_fill_8 FILLER_20_510 ();
 sg13g2_fill_4 FILLER_20_518 ();
 sg13g2_fill_1 FILLER_20_522 ();
 sg13g2_fill_1 FILLER_20_536 ();
 sg13g2_fill_8 FILLER_20_563 ();
 sg13g2_fill_8 FILLER_20_571 ();
 sg13g2_fill_8 FILLER_20_579 ();
 sg13g2_fill_8 FILLER_20_587 ();
 sg13g2_fill_8 FILLER_20_595 ();
 sg13g2_fill_8 FILLER_20_603 ();
 sg13g2_fill_8 FILLER_20_611 ();
 sg13g2_fill_8 FILLER_20_619 ();
 sg13g2_fill_8 FILLER_20_627 ();
 sg13g2_fill_8 FILLER_20_635 ();
 sg13g2_fill_8 FILLER_20_643 ();
 sg13g2_fill_8 FILLER_20_651 ();
 sg13g2_fill_8 FILLER_20_659 ();
 sg13g2_fill_8 FILLER_20_667 ();
 sg13g2_fill_8 FILLER_20_675 ();
 sg13g2_fill_8 FILLER_20_683 ();
 sg13g2_fill_8 FILLER_20_691 ();
 sg13g2_fill_8 FILLER_20_699 ();
 sg13g2_fill_8 FILLER_20_707 ();
 sg13g2_fill_8 FILLER_20_715 ();
 sg13g2_fill_8 FILLER_20_723 ();
 sg13g2_fill_8 FILLER_20_731 ();
 sg13g2_fill_8 FILLER_20_739 ();
 sg13g2_fill_8 FILLER_20_747 ();
 sg13g2_fill_8 FILLER_20_755 ();
 sg13g2_fill_8 FILLER_20_763 ();
 sg13g2_fill_8 FILLER_20_771 ();
 sg13g2_fill_8 FILLER_20_779 ();
 sg13g2_fill_8 FILLER_20_787 ();
 sg13g2_fill_8 FILLER_20_795 ();
 sg13g2_fill_8 FILLER_20_803 ();
 sg13g2_fill_8 FILLER_20_811 ();
 sg13g2_fill_8 FILLER_20_819 ();
 sg13g2_fill_8 FILLER_20_827 ();
 sg13g2_fill_8 FILLER_20_835 ();
 sg13g2_fill_8 FILLER_20_843 ();
 sg13g2_fill_8 FILLER_20_851 ();
 sg13g2_fill_8 FILLER_20_859 ();
 sg13g2_fill_8 FILLER_20_867 ();
 sg13g2_fill_8 FILLER_20_875 ();
 sg13g2_fill_8 FILLER_20_883 ();
 sg13g2_fill_8 FILLER_20_891 ();
 sg13g2_fill_8 FILLER_20_899 ();
 sg13g2_fill_8 FILLER_20_907 ();
 sg13g2_fill_8 FILLER_20_915 ();
 sg13g2_fill_8 FILLER_20_923 ();
 sg13g2_fill_8 FILLER_20_931 ();
 sg13g2_fill_8 FILLER_20_939 ();
 sg13g2_fill_8 FILLER_20_947 ();
 sg13g2_fill_8 FILLER_20_955 ();
 sg13g2_fill_8 FILLER_20_963 ();
 sg13g2_fill_8 FILLER_20_971 ();
 sg13g2_fill_8 FILLER_20_979 ();
 sg13g2_fill_8 FILLER_20_987 ();
 sg13g2_fill_8 FILLER_20_995 ();
 sg13g2_fill_8 FILLER_20_1003 ();
 sg13g2_fill_8 FILLER_20_1011 ();
 sg13g2_fill_8 FILLER_20_1019 ();
 sg13g2_fill_8 FILLER_20_1027 ();
 sg13g2_fill_8 FILLER_20_1035 ();
 sg13g2_fill_8 FILLER_20_1043 ();
 sg13g2_fill_8 FILLER_20_1051 ();
 sg13g2_fill_8 FILLER_20_1059 ();
 sg13g2_fill_8 FILLER_20_1067 ();
 sg13g2_fill_8 FILLER_20_1075 ();
 sg13g2_fill_8 FILLER_20_1083 ();
 sg13g2_fill_8 FILLER_20_1091 ();
 sg13g2_fill_8 FILLER_20_1099 ();
 sg13g2_fill_8 FILLER_20_1107 ();
 sg13g2_fill_8 FILLER_20_1115 ();
 sg13g2_fill_8 FILLER_20_1123 ();
 sg13g2_fill_8 FILLER_20_1131 ();
 sg13g2_fill_8 FILLER_20_1139 ();
 sg13g2_fill_8 FILLER_20_1147 ();
 sg13g2_fill_8 FILLER_20_1155 ();
 sg13g2_fill_2 FILLER_20_1163 ();
 sg13g2_fill_1 FILLER_20_1165 ();
 sg13g2_fill_8 FILLER_21_0 ();
 sg13g2_fill_8 FILLER_21_8 ();
 sg13g2_fill_8 FILLER_21_16 ();
 sg13g2_fill_8 FILLER_21_24 ();
 sg13g2_fill_1 FILLER_21_36 ();
 sg13g2_fill_2 FILLER_21_45 ();
 sg13g2_fill_8 FILLER_21_60 ();
 sg13g2_fill_4 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_fill_4 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_113 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_fill_4 FILLER_21_130 ();
 sg13g2_fill_4 FILLER_21_140 ();
 sg13g2_fill_8 FILLER_21_172 ();
 sg13g2_fill_4 FILLER_21_180 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_4 FILLER_21_228 ();
 sg13g2_fill_1 FILLER_21_232 ();
 sg13g2_fill_8 FILLER_21_236 ();
 sg13g2_fill_2 FILLER_21_244 ();
 sg13g2_fill_8 FILLER_21_267 ();
 sg13g2_fill_8 FILLER_21_275 ();
 sg13g2_fill_4 FILLER_21_283 ();
 sg13g2_fill_2 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_314 ();
 sg13g2_fill_4 FILLER_21_346 ();
 sg13g2_fill_2 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_352 ();
 sg13g2_fill_8 FILLER_21_361 ();
 sg13g2_fill_8 FILLER_21_369 ();
 sg13g2_fill_4 FILLER_21_377 ();
 sg13g2_fill_2 FILLER_21_381 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_21_461 ();
 sg13g2_fill_1 FILLER_21_473 ();
 sg13g2_fill_1 FILLER_21_514 ();
 sg13g2_fill_2 FILLER_21_541 ();
 sg13g2_fill_1 FILLER_21_543 ();
 sg13g2_fill_8 FILLER_21_596 ();
 sg13g2_fill_8 FILLER_21_604 ();
 sg13g2_fill_8 FILLER_21_612 ();
 sg13g2_fill_8 FILLER_21_620 ();
 sg13g2_fill_8 FILLER_21_628 ();
 sg13g2_fill_8 FILLER_21_636 ();
 sg13g2_fill_8 FILLER_21_644 ();
 sg13g2_fill_8 FILLER_21_652 ();
 sg13g2_fill_8 FILLER_21_660 ();
 sg13g2_fill_8 FILLER_21_668 ();
 sg13g2_fill_8 FILLER_21_676 ();
 sg13g2_fill_8 FILLER_21_684 ();
 sg13g2_fill_8 FILLER_21_692 ();
 sg13g2_fill_8 FILLER_21_700 ();
 sg13g2_fill_8 FILLER_21_708 ();
 sg13g2_fill_8 FILLER_21_716 ();
 sg13g2_fill_8 FILLER_21_724 ();
 sg13g2_fill_8 FILLER_21_732 ();
 sg13g2_fill_8 FILLER_21_740 ();
 sg13g2_fill_8 FILLER_21_748 ();
 sg13g2_fill_8 FILLER_21_756 ();
 sg13g2_fill_8 FILLER_21_764 ();
 sg13g2_fill_8 FILLER_21_772 ();
 sg13g2_fill_8 FILLER_21_780 ();
 sg13g2_fill_8 FILLER_21_788 ();
 sg13g2_fill_8 FILLER_21_796 ();
 sg13g2_fill_8 FILLER_21_804 ();
 sg13g2_fill_8 FILLER_21_812 ();
 sg13g2_fill_8 FILLER_21_820 ();
 sg13g2_fill_8 FILLER_21_828 ();
 sg13g2_fill_8 FILLER_21_836 ();
 sg13g2_fill_8 FILLER_21_844 ();
 sg13g2_fill_8 FILLER_21_852 ();
 sg13g2_fill_8 FILLER_21_860 ();
 sg13g2_fill_8 FILLER_21_868 ();
 sg13g2_fill_8 FILLER_21_876 ();
 sg13g2_fill_8 FILLER_21_884 ();
 sg13g2_fill_8 FILLER_21_892 ();
 sg13g2_fill_8 FILLER_21_900 ();
 sg13g2_fill_8 FILLER_21_908 ();
 sg13g2_fill_8 FILLER_21_916 ();
 sg13g2_fill_8 FILLER_21_924 ();
 sg13g2_fill_8 FILLER_21_932 ();
 sg13g2_fill_8 FILLER_21_940 ();
 sg13g2_fill_8 FILLER_21_948 ();
 sg13g2_fill_8 FILLER_21_956 ();
 sg13g2_fill_8 FILLER_21_964 ();
 sg13g2_fill_8 FILLER_21_972 ();
 sg13g2_fill_8 FILLER_21_980 ();
 sg13g2_fill_8 FILLER_21_988 ();
 sg13g2_fill_8 FILLER_21_996 ();
 sg13g2_fill_8 FILLER_21_1004 ();
 sg13g2_fill_8 FILLER_21_1012 ();
 sg13g2_fill_8 FILLER_21_1020 ();
 sg13g2_fill_8 FILLER_21_1028 ();
 sg13g2_fill_8 FILLER_21_1036 ();
 sg13g2_fill_8 FILLER_21_1044 ();
 sg13g2_fill_8 FILLER_21_1052 ();
 sg13g2_fill_8 FILLER_21_1060 ();
 sg13g2_fill_8 FILLER_21_1068 ();
 sg13g2_fill_8 FILLER_21_1076 ();
 sg13g2_fill_8 FILLER_21_1084 ();
 sg13g2_fill_8 FILLER_21_1092 ();
 sg13g2_fill_8 FILLER_21_1100 ();
 sg13g2_fill_8 FILLER_21_1108 ();
 sg13g2_fill_8 FILLER_21_1116 ();
 sg13g2_fill_8 FILLER_21_1124 ();
 sg13g2_fill_8 FILLER_21_1132 ();
 sg13g2_fill_8 FILLER_21_1140 ();
 sg13g2_fill_8 FILLER_21_1148 ();
 sg13g2_fill_8 FILLER_21_1156 ();
 sg13g2_fill_2 FILLER_21_1164 ();
 sg13g2_fill_8 FILLER_22_0 ();
 sg13g2_fill_8 FILLER_22_8 ();
 sg13g2_fill_8 FILLER_22_16 ();
 sg13g2_fill_8 FILLER_22_64 ();
 sg13g2_fill_8 FILLER_22_72 ();
 sg13g2_fill_8 FILLER_22_80 ();
 sg13g2_fill_8 FILLER_22_88 ();
 sg13g2_fill_8 FILLER_22_96 ();
 sg13g2_fill_4 FILLER_22_104 ();
 sg13g2_fill_2 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_110 ();
 sg13g2_fill_8 FILLER_22_116 ();
 sg13g2_fill_4 FILLER_22_124 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_130 ();
 sg13g2_fill_8 FILLER_22_136 ();
 sg13g2_fill_8 FILLER_22_144 ();
 sg13g2_fill_8 FILLER_22_152 ();
 sg13g2_fill_4 FILLER_22_160 ();
 sg13g2_fill_2 FILLER_22_164 ();
 sg13g2_fill_4 FILLER_22_174 ();
 sg13g2_fill_2 FILLER_22_178 ();
 sg13g2_fill_1 FILLER_22_180 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_4 FILLER_22_218 ();
 sg13g2_fill_8 FILLER_22_280 ();
 sg13g2_fill_4 FILLER_22_288 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_8 FILLER_22_346 ();
 sg13g2_fill_8 FILLER_22_354 ();
 sg13g2_fill_4 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_366 ();
 sg13g2_fill_4 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_379 ();
 sg13g2_fill_4 FILLER_22_386 ();
 sg13g2_fill_8 FILLER_22_396 ();
 sg13g2_fill_1 FILLER_22_409 ();
 sg13g2_fill_2 FILLER_22_413 ();
 sg13g2_fill_1 FILLER_22_415 ();
 sg13g2_fill_1 FILLER_22_452 ();
 sg13g2_fill_2 FILLER_22_484 ();
 sg13g2_fill_4 FILLER_22_512 ();
 sg13g2_fill_1 FILLER_22_568 ();
 sg13g2_fill_8 FILLER_22_600 ();
 sg13g2_fill_8 FILLER_22_608 ();
 sg13g2_fill_8 FILLER_22_616 ();
 sg13g2_fill_8 FILLER_22_624 ();
 sg13g2_fill_8 FILLER_22_632 ();
 sg13g2_fill_8 FILLER_22_640 ();
 sg13g2_fill_8 FILLER_22_648 ();
 sg13g2_fill_8 FILLER_22_656 ();
 sg13g2_fill_8 FILLER_22_664 ();
 sg13g2_fill_8 FILLER_22_672 ();
 sg13g2_fill_8 FILLER_22_680 ();
 sg13g2_fill_8 FILLER_22_688 ();
 sg13g2_fill_8 FILLER_22_696 ();
 sg13g2_fill_8 FILLER_22_704 ();
 sg13g2_fill_8 FILLER_22_712 ();
 sg13g2_fill_8 FILLER_22_720 ();
 sg13g2_fill_8 FILLER_22_728 ();
 sg13g2_fill_8 FILLER_22_736 ();
 sg13g2_fill_8 FILLER_22_744 ();
 sg13g2_fill_8 FILLER_22_752 ();
 sg13g2_fill_8 FILLER_22_760 ();
 sg13g2_fill_8 FILLER_22_768 ();
 sg13g2_fill_8 FILLER_22_776 ();
 sg13g2_fill_8 FILLER_22_784 ();
 sg13g2_fill_8 FILLER_22_792 ();
 sg13g2_fill_8 FILLER_22_800 ();
 sg13g2_fill_8 FILLER_22_808 ();
 sg13g2_fill_8 FILLER_22_816 ();
 sg13g2_fill_8 FILLER_22_824 ();
 sg13g2_fill_8 FILLER_22_832 ();
 sg13g2_fill_8 FILLER_22_840 ();
 sg13g2_fill_8 FILLER_22_848 ();
 sg13g2_fill_8 FILLER_22_856 ();
 sg13g2_fill_8 FILLER_22_864 ();
 sg13g2_fill_8 FILLER_22_872 ();
 sg13g2_fill_8 FILLER_22_880 ();
 sg13g2_fill_8 FILLER_22_888 ();
 sg13g2_fill_8 FILLER_22_896 ();
 sg13g2_fill_8 FILLER_22_904 ();
 sg13g2_fill_8 FILLER_22_912 ();
 sg13g2_fill_8 FILLER_22_920 ();
 sg13g2_fill_8 FILLER_22_928 ();
 sg13g2_fill_8 FILLER_22_936 ();
 sg13g2_fill_8 FILLER_22_944 ();
 sg13g2_fill_8 FILLER_22_952 ();
 sg13g2_fill_8 FILLER_22_960 ();
 sg13g2_fill_8 FILLER_22_968 ();
 sg13g2_fill_8 FILLER_22_976 ();
 sg13g2_fill_8 FILLER_22_984 ();
 sg13g2_fill_8 FILLER_22_992 ();
 sg13g2_fill_8 FILLER_22_1000 ();
 sg13g2_fill_8 FILLER_22_1008 ();
 sg13g2_fill_8 FILLER_22_1016 ();
 sg13g2_fill_8 FILLER_22_1024 ();
 sg13g2_fill_8 FILLER_22_1032 ();
 sg13g2_fill_8 FILLER_22_1040 ();
 sg13g2_fill_8 FILLER_22_1048 ();
 sg13g2_fill_8 FILLER_22_1056 ();
 sg13g2_fill_8 FILLER_22_1064 ();
 sg13g2_fill_8 FILLER_22_1072 ();
 sg13g2_fill_8 FILLER_22_1080 ();
 sg13g2_fill_8 FILLER_22_1088 ();
 sg13g2_fill_8 FILLER_22_1096 ();
 sg13g2_fill_8 FILLER_22_1104 ();
 sg13g2_fill_8 FILLER_22_1112 ();
 sg13g2_fill_8 FILLER_22_1120 ();
 sg13g2_fill_8 FILLER_22_1128 ();
 sg13g2_fill_8 FILLER_22_1136 ();
 sg13g2_fill_8 FILLER_22_1144 ();
 sg13g2_fill_8 FILLER_22_1152 ();
 sg13g2_fill_4 FILLER_22_1160 ();
 sg13g2_fill_2 FILLER_22_1164 ();
 sg13g2_fill_8 FILLER_23_0 ();
 sg13g2_fill_8 FILLER_23_8 ();
 sg13g2_fill_4 FILLER_23_16 ();
 sg13g2_fill_1 FILLER_23_20 ();
 sg13g2_fill_2 FILLER_23_29 ();
 sg13g2_fill_2 FILLER_23_41 ();
 sg13g2_fill_1 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_70 ();
 sg13g2_fill_8 FILLER_23_92 ();
 sg13g2_fill_8 FILLER_23_100 ();
 sg13g2_fill_1 FILLER_23_108 ();
 sg13g2_fill_4 FILLER_23_114 ();
 sg13g2_fill_2 FILLER_23_118 ();
 sg13g2_fill_8 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_144 ();
 sg13g2_fill_2 FILLER_23_166 ();
 sg13g2_fill_8 FILLER_23_182 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_8 FILLER_23_210 ();
 sg13g2_fill_4 FILLER_23_218 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_1 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_325 ();
 sg13g2_fill_2 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_359 ();
 sg13g2_fill_1 FILLER_23_368 ();
 sg13g2_fill_1 FILLER_23_421 ();
 sg13g2_fill_8 FILLER_23_453 ();
 sg13g2_fill_4 FILLER_23_461 ();
 sg13g2_fill_2 FILLER_23_465 ();
 sg13g2_fill_1 FILLER_23_467 ();
 sg13g2_fill_8 FILLER_23_472 ();
 sg13g2_fill_4 FILLER_23_480 ();
 sg13g2_fill_2 FILLER_23_484 ();
 sg13g2_fill_4 FILLER_23_510 ();
 sg13g2_fill_2 FILLER_23_514 ();
 sg13g2_fill_1 FILLER_23_516 ();
 sg13g2_fill_2 FILLER_23_553 ();
 sg13g2_fill_8 FILLER_23_585 ();
 sg13g2_fill_8 FILLER_23_593 ();
 sg13g2_fill_8 FILLER_23_601 ();
 sg13g2_fill_8 FILLER_23_609 ();
 sg13g2_fill_8 FILLER_23_617 ();
 sg13g2_fill_8 FILLER_23_625 ();
 sg13g2_fill_8 FILLER_23_633 ();
 sg13g2_fill_8 FILLER_23_641 ();
 sg13g2_fill_8 FILLER_23_649 ();
 sg13g2_fill_8 FILLER_23_657 ();
 sg13g2_fill_8 FILLER_23_665 ();
 sg13g2_fill_8 FILLER_23_673 ();
 sg13g2_fill_8 FILLER_23_681 ();
 sg13g2_fill_8 FILLER_23_689 ();
 sg13g2_fill_8 FILLER_23_697 ();
 sg13g2_fill_8 FILLER_23_705 ();
 sg13g2_fill_8 FILLER_23_713 ();
 sg13g2_fill_8 FILLER_23_721 ();
 sg13g2_fill_8 FILLER_23_729 ();
 sg13g2_fill_8 FILLER_23_737 ();
 sg13g2_fill_8 FILLER_23_745 ();
 sg13g2_fill_8 FILLER_23_753 ();
 sg13g2_fill_8 FILLER_23_761 ();
 sg13g2_fill_8 FILLER_23_769 ();
 sg13g2_fill_8 FILLER_23_777 ();
 sg13g2_fill_8 FILLER_23_785 ();
 sg13g2_fill_8 FILLER_23_793 ();
 sg13g2_fill_8 FILLER_23_801 ();
 sg13g2_fill_8 FILLER_23_809 ();
 sg13g2_fill_8 FILLER_23_817 ();
 sg13g2_fill_8 FILLER_23_825 ();
 sg13g2_fill_8 FILLER_23_833 ();
 sg13g2_fill_8 FILLER_23_841 ();
 sg13g2_fill_8 FILLER_23_849 ();
 sg13g2_fill_8 FILLER_23_857 ();
 sg13g2_fill_8 FILLER_23_865 ();
 sg13g2_fill_8 FILLER_23_873 ();
 sg13g2_fill_8 FILLER_23_881 ();
 sg13g2_fill_8 FILLER_23_889 ();
 sg13g2_fill_8 FILLER_23_897 ();
 sg13g2_fill_8 FILLER_23_905 ();
 sg13g2_fill_8 FILLER_23_913 ();
 sg13g2_fill_8 FILLER_23_921 ();
 sg13g2_fill_8 FILLER_23_929 ();
 sg13g2_fill_8 FILLER_23_937 ();
 sg13g2_fill_8 FILLER_23_945 ();
 sg13g2_fill_8 FILLER_23_953 ();
 sg13g2_fill_8 FILLER_23_961 ();
 sg13g2_fill_8 FILLER_23_969 ();
 sg13g2_fill_8 FILLER_23_977 ();
 sg13g2_fill_8 FILLER_23_985 ();
 sg13g2_fill_8 FILLER_23_993 ();
 sg13g2_fill_8 FILLER_23_1001 ();
 sg13g2_fill_8 FILLER_23_1009 ();
 sg13g2_fill_8 FILLER_23_1017 ();
 sg13g2_fill_8 FILLER_23_1025 ();
 sg13g2_fill_8 FILLER_23_1033 ();
 sg13g2_fill_8 FILLER_23_1041 ();
 sg13g2_fill_8 FILLER_23_1049 ();
 sg13g2_fill_8 FILLER_23_1057 ();
 sg13g2_fill_8 FILLER_23_1065 ();
 sg13g2_fill_8 FILLER_23_1073 ();
 sg13g2_fill_8 FILLER_23_1081 ();
 sg13g2_fill_8 FILLER_23_1089 ();
 sg13g2_fill_8 FILLER_23_1097 ();
 sg13g2_fill_8 FILLER_23_1105 ();
 sg13g2_fill_8 FILLER_23_1113 ();
 sg13g2_fill_8 FILLER_23_1121 ();
 sg13g2_fill_8 FILLER_23_1129 ();
 sg13g2_fill_8 FILLER_23_1137 ();
 sg13g2_fill_8 FILLER_23_1145 ();
 sg13g2_fill_8 FILLER_23_1153 ();
 sg13g2_fill_4 FILLER_23_1161 ();
 sg13g2_fill_1 FILLER_23_1165 ();
 sg13g2_fill_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_34 ();
 sg13g2_fill_8 FILLER_24_61 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_8 FILLER_24_144 ();
 sg13g2_fill_4 FILLER_24_152 ();
 sg13g2_fill_2 FILLER_24_156 ();
 sg13g2_fill_1 FILLER_24_158 ();
 sg13g2_fill_8 FILLER_24_190 ();
 sg13g2_fill_8 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_211 ();
 sg13g2_fill_8 FILLER_24_218 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_8 FILLER_24_231 ();
 sg13g2_fill_8 FILLER_24_239 ();
 sg13g2_fill_2 FILLER_24_247 ();
 sg13g2_fill_2 FILLER_24_254 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_8 FILLER_24_265 ();
 sg13g2_fill_8 FILLER_24_273 ();
 sg13g2_fill_8 FILLER_24_281 ();
 sg13g2_fill_4 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_fill_2 FILLER_24_312 ();
 sg13g2_fill_1 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_336 ();
 sg13g2_fill_4 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_354 ();
 sg13g2_fill_8 FILLER_24_381 ();
 sg13g2_fill_4 FILLER_24_389 ();
 sg13g2_fill_8 FILLER_24_447 ();
 sg13g2_fill_8 FILLER_24_460 ();
 sg13g2_fill_8 FILLER_24_468 ();
 sg13g2_fill_8 FILLER_24_476 ();
 sg13g2_fill_8 FILLER_24_484 ();
 sg13g2_fill_8 FILLER_24_492 ();
 sg13g2_fill_8 FILLER_24_500 ();
 sg13g2_fill_8 FILLER_24_508 ();
 sg13g2_fill_8 FILLER_24_516 ();
 sg13g2_fill_4 FILLER_24_524 ();
 sg13g2_fill_1 FILLER_24_528 ();
 sg13g2_fill_4 FILLER_24_559 ();
 sg13g2_fill_2 FILLER_24_563 ();
 sg13g2_fill_8 FILLER_24_578 ();
 sg13g2_fill_8 FILLER_24_586 ();
 sg13g2_fill_8 FILLER_24_594 ();
 sg13g2_fill_8 FILLER_24_602 ();
 sg13g2_fill_8 FILLER_24_610 ();
 sg13g2_fill_8 FILLER_24_618 ();
 sg13g2_fill_8 FILLER_24_626 ();
 sg13g2_fill_8 FILLER_24_634 ();
 sg13g2_fill_8 FILLER_24_642 ();
 sg13g2_fill_8 FILLER_24_650 ();
 sg13g2_fill_8 FILLER_24_658 ();
 sg13g2_fill_8 FILLER_24_666 ();
 sg13g2_fill_8 FILLER_24_674 ();
 sg13g2_fill_8 FILLER_24_682 ();
 sg13g2_fill_8 FILLER_24_690 ();
 sg13g2_fill_8 FILLER_24_698 ();
 sg13g2_fill_8 FILLER_24_706 ();
 sg13g2_fill_8 FILLER_24_714 ();
 sg13g2_fill_8 FILLER_24_722 ();
 sg13g2_fill_8 FILLER_24_730 ();
 sg13g2_fill_8 FILLER_24_738 ();
 sg13g2_fill_8 FILLER_24_746 ();
 sg13g2_fill_8 FILLER_24_754 ();
 sg13g2_fill_8 FILLER_24_762 ();
 sg13g2_fill_8 FILLER_24_770 ();
 sg13g2_fill_8 FILLER_24_778 ();
 sg13g2_fill_8 FILLER_24_786 ();
 sg13g2_fill_8 FILLER_24_794 ();
 sg13g2_fill_8 FILLER_24_802 ();
 sg13g2_fill_8 FILLER_24_810 ();
 sg13g2_fill_8 FILLER_24_818 ();
 sg13g2_fill_8 FILLER_24_826 ();
 sg13g2_fill_8 FILLER_24_834 ();
 sg13g2_fill_8 FILLER_24_842 ();
 sg13g2_fill_8 FILLER_24_850 ();
 sg13g2_fill_8 FILLER_24_858 ();
 sg13g2_fill_8 FILLER_24_866 ();
 sg13g2_fill_8 FILLER_24_874 ();
 sg13g2_fill_8 FILLER_24_882 ();
 sg13g2_fill_8 FILLER_24_890 ();
 sg13g2_fill_8 FILLER_24_898 ();
 sg13g2_fill_8 FILLER_24_906 ();
 sg13g2_fill_8 FILLER_24_914 ();
 sg13g2_fill_8 FILLER_24_922 ();
 sg13g2_fill_8 FILLER_24_930 ();
 sg13g2_fill_8 FILLER_24_938 ();
 sg13g2_fill_8 FILLER_24_946 ();
 sg13g2_fill_8 FILLER_24_954 ();
 sg13g2_fill_8 FILLER_24_962 ();
 sg13g2_fill_8 FILLER_24_970 ();
 sg13g2_fill_8 FILLER_24_978 ();
 sg13g2_fill_8 FILLER_24_986 ();
 sg13g2_fill_8 FILLER_24_994 ();
 sg13g2_fill_8 FILLER_24_1002 ();
 sg13g2_fill_8 FILLER_24_1010 ();
 sg13g2_fill_8 FILLER_24_1018 ();
 sg13g2_fill_8 FILLER_24_1026 ();
 sg13g2_fill_8 FILLER_24_1034 ();
 sg13g2_fill_8 FILLER_24_1042 ();
 sg13g2_fill_8 FILLER_24_1050 ();
 sg13g2_fill_8 FILLER_24_1058 ();
 sg13g2_fill_8 FILLER_24_1066 ();
 sg13g2_fill_8 FILLER_24_1074 ();
 sg13g2_fill_8 FILLER_24_1082 ();
 sg13g2_fill_8 FILLER_24_1090 ();
 sg13g2_fill_8 FILLER_24_1098 ();
 sg13g2_fill_8 FILLER_24_1106 ();
 sg13g2_fill_8 FILLER_24_1114 ();
 sg13g2_fill_8 FILLER_24_1122 ();
 sg13g2_fill_8 FILLER_24_1130 ();
 sg13g2_fill_8 FILLER_24_1138 ();
 sg13g2_fill_8 FILLER_24_1146 ();
 sg13g2_fill_8 FILLER_24_1154 ();
 sg13g2_fill_4 FILLER_24_1162 ();
 sg13g2_fill_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_fill_8 FILLER_25_32 ();
 sg13g2_fill_4 FILLER_25_40 ();
 sg13g2_fill_2 FILLER_25_44 ();
 sg13g2_fill_8 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_104 ();
 sg13g2_fill_8 FILLER_25_188 ();
 sg13g2_fill_4 FILLER_25_196 ();
 sg13g2_fill_4 FILLER_25_226 ();
 sg13g2_fill_8 FILLER_25_268 ();
 sg13g2_fill_8 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_fill_8 FILLER_25_288 ();
 sg13g2_fill_8 FILLER_25_296 ();
 sg13g2_fill_4 FILLER_25_304 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_fill_8 FILLER_25_315 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_8 FILLER_25_347 ();
 sg13g2_fill_8 FILLER_25_355 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_fill_4 FILLER_25_456 ();
 sg13g2_fill_2 FILLER_25_477 ();
 sg13g2_fill_8 FILLER_25_510 ();
 sg13g2_fill_1 FILLER_25_533 ();
 sg13g2_fill_2 FILLER_25_560 ();
 sg13g2_fill_8 FILLER_25_588 ();
 sg13g2_fill_8 FILLER_25_596 ();
 sg13g2_fill_8 FILLER_25_604 ();
 sg13g2_fill_8 FILLER_25_612 ();
 sg13g2_fill_8 FILLER_25_620 ();
 sg13g2_fill_8 FILLER_25_628 ();
 sg13g2_fill_8 FILLER_25_636 ();
 sg13g2_fill_8 FILLER_25_644 ();
 sg13g2_fill_8 FILLER_25_652 ();
 sg13g2_fill_8 FILLER_25_660 ();
 sg13g2_fill_8 FILLER_25_668 ();
 sg13g2_fill_8 FILLER_25_676 ();
 sg13g2_fill_8 FILLER_25_684 ();
 sg13g2_fill_8 FILLER_25_692 ();
 sg13g2_fill_8 FILLER_25_700 ();
 sg13g2_fill_8 FILLER_25_708 ();
 sg13g2_fill_8 FILLER_25_716 ();
 sg13g2_fill_8 FILLER_25_724 ();
 sg13g2_fill_8 FILLER_25_732 ();
 sg13g2_fill_8 FILLER_25_740 ();
 sg13g2_fill_8 FILLER_25_748 ();
 sg13g2_fill_8 FILLER_25_756 ();
 sg13g2_fill_8 FILLER_25_764 ();
 sg13g2_fill_8 FILLER_25_772 ();
 sg13g2_fill_8 FILLER_25_780 ();
 sg13g2_fill_8 FILLER_25_788 ();
 sg13g2_fill_8 FILLER_25_796 ();
 sg13g2_fill_8 FILLER_25_804 ();
 sg13g2_fill_8 FILLER_25_812 ();
 sg13g2_fill_8 FILLER_25_820 ();
 sg13g2_fill_8 FILLER_25_828 ();
 sg13g2_fill_8 FILLER_25_836 ();
 sg13g2_fill_8 FILLER_25_844 ();
 sg13g2_fill_8 FILLER_25_852 ();
 sg13g2_fill_8 FILLER_25_860 ();
 sg13g2_fill_8 FILLER_25_868 ();
 sg13g2_fill_8 FILLER_25_876 ();
 sg13g2_fill_8 FILLER_25_884 ();
 sg13g2_fill_8 FILLER_25_892 ();
 sg13g2_fill_8 FILLER_25_900 ();
 sg13g2_fill_8 FILLER_25_908 ();
 sg13g2_fill_8 FILLER_25_916 ();
 sg13g2_fill_8 FILLER_25_924 ();
 sg13g2_fill_8 FILLER_25_932 ();
 sg13g2_fill_8 FILLER_25_940 ();
 sg13g2_fill_8 FILLER_25_948 ();
 sg13g2_fill_8 FILLER_25_956 ();
 sg13g2_fill_8 FILLER_25_964 ();
 sg13g2_fill_8 FILLER_25_972 ();
 sg13g2_fill_8 FILLER_25_980 ();
 sg13g2_fill_8 FILLER_25_988 ();
 sg13g2_fill_8 FILLER_25_996 ();
 sg13g2_fill_8 FILLER_25_1004 ();
 sg13g2_fill_8 FILLER_25_1012 ();
 sg13g2_fill_8 FILLER_25_1020 ();
 sg13g2_fill_8 FILLER_25_1028 ();
 sg13g2_fill_8 FILLER_25_1036 ();
 sg13g2_fill_8 FILLER_25_1044 ();
 sg13g2_fill_8 FILLER_25_1052 ();
 sg13g2_fill_8 FILLER_25_1060 ();
 sg13g2_fill_8 FILLER_25_1068 ();
 sg13g2_fill_8 FILLER_25_1076 ();
 sg13g2_fill_8 FILLER_25_1084 ();
 sg13g2_fill_8 FILLER_25_1092 ();
 sg13g2_fill_8 FILLER_25_1100 ();
 sg13g2_fill_8 FILLER_25_1108 ();
 sg13g2_fill_8 FILLER_25_1116 ();
 sg13g2_fill_8 FILLER_25_1124 ();
 sg13g2_fill_8 FILLER_25_1132 ();
 sg13g2_fill_8 FILLER_25_1140 ();
 sg13g2_fill_8 FILLER_25_1148 ();
 sg13g2_fill_8 FILLER_25_1156 ();
 sg13g2_fill_2 FILLER_25_1164 ();
 sg13g2_fill_8 FILLER_26_0 ();
 sg13g2_fill_8 FILLER_26_8 ();
 sg13g2_fill_2 FILLER_26_16 ();
 sg13g2_fill_8 FILLER_26_36 ();
 sg13g2_fill_4 FILLER_26_44 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_4 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_4 FILLER_26_200 ();
 sg13g2_fill_1 FILLER_26_204 ();
 sg13g2_fill_2 FILLER_26_209 ();
 sg13g2_fill_1 FILLER_26_247 ();
 sg13g2_fill_8 FILLER_26_256 ();
 sg13g2_fill_8 FILLER_26_298 ();
 sg13g2_fill_8 FILLER_26_306 ();
 sg13g2_fill_4 FILLER_26_314 ();
 sg13g2_fill_2 FILLER_26_318 ();
 sg13g2_fill_8 FILLER_26_354 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_371 ();
 sg13g2_fill_8 FILLER_26_403 ();
 sg13g2_fill_8 FILLER_26_411 ();
 sg13g2_fill_4 FILLER_26_419 ();
 sg13g2_fill_1 FILLER_26_423 ();
 sg13g2_fill_2 FILLER_26_461 ();
 sg13g2_fill_2 FILLER_26_510 ();
 sg13g2_fill_2 FILLER_26_563 ();
 sg13g2_fill_8 FILLER_26_604 ();
 sg13g2_fill_8 FILLER_26_612 ();
 sg13g2_fill_8 FILLER_26_620 ();
 sg13g2_fill_8 FILLER_26_628 ();
 sg13g2_fill_8 FILLER_26_636 ();
 sg13g2_fill_8 FILLER_26_644 ();
 sg13g2_fill_8 FILLER_26_652 ();
 sg13g2_fill_8 FILLER_26_660 ();
 sg13g2_fill_8 FILLER_26_668 ();
 sg13g2_fill_8 FILLER_26_676 ();
 sg13g2_fill_8 FILLER_26_684 ();
 sg13g2_fill_8 FILLER_26_692 ();
 sg13g2_fill_8 FILLER_26_700 ();
 sg13g2_fill_8 FILLER_26_708 ();
 sg13g2_fill_8 FILLER_26_716 ();
 sg13g2_fill_8 FILLER_26_724 ();
 sg13g2_fill_8 FILLER_26_732 ();
 sg13g2_fill_8 FILLER_26_740 ();
 sg13g2_fill_8 FILLER_26_748 ();
 sg13g2_fill_8 FILLER_26_756 ();
 sg13g2_fill_8 FILLER_26_764 ();
 sg13g2_fill_8 FILLER_26_772 ();
 sg13g2_fill_8 FILLER_26_780 ();
 sg13g2_fill_8 FILLER_26_788 ();
 sg13g2_fill_8 FILLER_26_796 ();
 sg13g2_fill_8 FILLER_26_804 ();
 sg13g2_fill_8 FILLER_26_812 ();
 sg13g2_fill_8 FILLER_26_820 ();
 sg13g2_fill_8 FILLER_26_828 ();
 sg13g2_fill_8 FILLER_26_836 ();
 sg13g2_fill_8 FILLER_26_844 ();
 sg13g2_fill_8 FILLER_26_852 ();
 sg13g2_fill_8 FILLER_26_860 ();
 sg13g2_fill_8 FILLER_26_868 ();
 sg13g2_fill_8 FILLER_26_876 ();
 sg13g2_fill_8 FILLER_26_884 ();
 sg13g2_fill_8 FILLER_26_892 ();
 sg13g2_fill_8 FILLER_26_900 ();
 sg13g2_fill_8 FILLER_26_908 ();
 sg13g2_fill_8 FILLER_26_916 ();
 sg13g2_fill_8 FILLER_26_924 ();
 sg13g2_fill_8 FILLER_26_932 ();
 sg13g2_fill_8 FILLER_26_940 ();
 sg13g2_fill_8 FILLER_26_948 ();
 sg13g2_fill_8 FILLER_26_956 ();
 sg13g2_fill_8 FILLER_26_964 ();
 sg13g2_fill_8 FILLER_26_972 ();
 sg13g2_fill_8 FILLER_26_980 ();
 sg13g2_fill_8 FILLER_26_988 ();
 sg13g2_fill_8 FILLER_26_996 ();
 sg13g2_fill_8 FILLER_26_1004 ();
 sg13g2_fill_8 FILLER_26_1012 ();
 sg13g2_fill_8 FILLER_26_1020 ();
 sg13g2_fill_8 FILLER_26_1028 ();
 sg13g2_fill_8 FILLER_26_1036 ();
 sg13g2_fill_8 FILLER_26_1044 ();
 sg13g2_fill_8 FILLER_26_1052 ();
 sg13g2_fill_8 FILLER_26_1060 ();
 sg13g2_fill_8 FILLER_26_1068 ();
 sg13g2_fill_8 FILLER_26_1076 ();
 sg13g2_fill_8 FILLER_26_1084 ();
 sg13g2_fill_8 FILLER_26_1092 ();
 sg13g2_fill_8 FILLER_26_1100 ();
 sg13g2_fill_8 FILLER_26_1108 ();
 sg13g2_fill_8 FILLER_26_1116 ();
 sg13g2_fill_8 FILLER_26_1124 ();
 sg13g2_fill_8 FILLER_26_1132 ();
 sg13g2_fill_8 FILLER_26_1140 ();
 sg13g2_fill_8 FILLER_26_1148 ();
 sg13g2_fill_8 FILLER_26_1156 ();
 sg13g2_fill_2 FILLER_26_1164 ();
 sg13g2_fill_8 FILLER_27_0 ();
 sg13g2_fill_8 FILLER_27_8 ();
 sg13g2_fill_4 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_32 ();
 sg13g2_fill_4 FILLER_27_41 ();
 sg13g2_fill_8 FILLER_27_53 ();
 sg13g2_fill_2 FILLER_27_82 ();
 sg13g2_fill_1 FILLER_27_84 ();
 sg13g2_fill_4 FILLER_27_91 ();
 sg13g2_fill_4 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_124 ();
 sg13g2_fill_2 FILLER_27_131 ();
 sg13g2_fill_8 FILLER_27_136 ();
 sg13g2_fill_8 FILLER_27_144 ();
 sg13g2_fill_8 FILLER_27_152 ();
 sg13g2_fill_4 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_8 FILLER_27_172 ();
 sg13g2_fill_4 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_4 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_8 FILLER_27_226 ();
 sg13g2_fill_8 FILLER_27_234 ();
 sg13g2_fill_8 FILLER_27_242 ();
 sg13g2_fill_8 FILLER_27_250 ();
 sg13g2_fill_4 FILLER_27_258 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_fill_1 FILLER_27_269 ();
 sg13g2_fill_4 FILLER_27_273 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_fill_4 FILLER_27_288 ();
 sg13g2_fill_4 FILLER_27_318 ();
 sg13g2_fill_1 FILLER_27_322 ();
 sg13g2_fill_4 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_1 FILLER_27_386 ();
 sg13g2_fill_8 FILLER_27_421 ();
 sg13g2_fill_4 FILLER_27_429 ();
 sg13g2_fill_2 FILLER_27_433 ();
 sg13g2_fill_8 FILLER_27_440 ();
 sg13g2_fill_4 FILLER_27_448 ();
 sg13g2_fill_2 FILLER_27_452 ();
 sg13g2_fill_2 FILLER_27_485 ();
 sg13g2_fill_4 FILLER_27_493 ();
 sg13g2_fill_2 FILLER_27_497 ();
 sg13g2_fill_1 FILLER_27_527 ();
 sg13g2_fill_8 FILLER_27_534 ();
 sg13g2_fill_8 FILLER_27_542 ();
 sg13g2_fill_4 FILLER_27_550 ();
 sg13g2_fill_2 FILLER_27_554 ();
 sg13g2_fill_1 FILLER_27_556 ();
 sg13g2_fill_8 FILLER_27_567 ();
 sg13g2_fill_2 FILLER_27_575 ();
 sg13g2_fill_1 FILLER_27_608 ();
 sg13g2_fill_8 FILLER_27_639 ();
 sg13g2_fill_8 FILLER_27_655 ();
 sg13g2_fill_8 FILLER_27_663 ();
 sg13g2_fill_8 FILLER_27_671 ();
 sg13g2_fill_4 FILLER_27_679 ();
 sg13g2_fill_2 FILLER_27_683 ();
 sg13g2_fill_1 FILLER_27_685 ();
 sg13g2_fill_8 FILLER_27_694 ();
 sg13g2_fill_8 FILLER_27_702 ();
 sg13g2_fill_8 FILLER_27_710 ();
 sg13g2_fill_8 FILLER_27_718 ();
 sg13g2_fill_8 FILLER_27_726 ();
 sg13g2_fill_8 FILLER_27_734 ();
 sg13g2_fill_8 FILLER_27_742 ();
 sg13g2_fill_8 FILLER_27_750 ();
 sg13g2_fill_8 FILLER_27_758 ();
 sg13g2_fill_8 FILLER_27_766 ();
 sg13g2_fill_8 FILLER_27_774 ();
 sg13g2_fill_8 FILLER_27_782 ();
 sg13g2_fill_8 FILLER_27_790 ();
 sg13g2_fill_8 FILLER_27_798 ();
 sg13g2_fill_8 FILLER_27_806 ();
 sg13g2_fill_8 FILLER_27_814 ();
 sg13g2_fill_8 FILLER_27_822 ();
 sg13g2_fill_8 FILLER_27_830 ();
 sg13g2_fill_8 FILLER_27_838 ();
 sg13g2_fill_8 FILLER_27_846 ();
 sg13g2_fill_8 FILLER_27_854 ();
 sg13g2_fill_8 FILLER_27_862 ();
 sg13g2_fill_8 FILLER_27_870 ();
 sg13g2_fill_8 FILLER_27_878 ();
 sg13g2_fill_8 FILLER_27_886 ();
 sg13g2_fill_8 FILLER_27_894 ();
 sg13g2_fill_8 FILLER_27_902 ();
 sg13g2_fill_8 FILLER_27_910 ();
 sg13g2_fill_8 FILLER_27_918 ();
 sg13g2_fill_8 FILLER_27_926 ();
 sg13g2_fill_8 FILLER_27_934 ();
 sg13g2_fill_8 FILLER_27_942 ();
 sg13g2_fill_8 FILLER_27_950 ();
 sg13g2_fill_8 FILLER_27_958 ();
 sg13g2_fill_8 FILLER_27_966 ();
 sg13g2_fill_8 FILLER_27_974 ();
 sg13g2_fill_8 FILLER_27_982 ();
 sg13g2_fill_8 FILLER_27_990 ();
 sg13g2_fill_8 FILLER_27_998 ();
 sg13g2_fill_8 FILLER_27_1006 ();
 sg13g2_fill_8 FILLER_27_1014 ();
 sg13g2_fill_8 FILLER_27_1022 ();
 sg13g2_fill_8 FILLER_27_1030 ();
 sg13g2_fill_8 FILLER_27_1038 ();
 sg13g2_fill_8 FILLER_27_1046 ();
 sg13g2_fill_8 FILLER_27_1054 ();
 sg13g2_fill_8 FILLER_27_1062 ();
 sg13g2_fill_8 FILLER_27_1070 ();
 sg13g2_fill_8 FILLER_27_1078 ();
 sg13g2_fill_8 FILLER_27_1086 ();
 sg13g2_fill_8 FILLER_27_1094 ();
 sg13g2_fill_8 FILLER_27_1102 ();
 sg13g2_fill_8 FILLER_27_1110 ();
 sg13g2_fill_8 FILLER_27_1118 ();
 sg13g2_fill_8 FILLER_27_1126 ();
 sg13g2_fill_8 FILLER_27_1134 ();
 sg13g2_fill_8 FILLER_27_1142 ();
 sg13g2_fill_8 FILLER_27_1150 ();
 sg13g2_fill_8 FILLER_27_1158 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_8 FILLER_28_34 ();
 sg13g2_fill_8 FILLER_28_42 ();
 sg13g2_fill_8 FILLER_28_50 ();
 sg13g2_fill_8 FILLER_28_58 ();
 sg13g2_fill_8 FILLER_28_66 ();
 sg13g2_fill_2 FILLER_28_74 ();
 sg13g2_fill_8 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_93 ();
 sg13g2_fill_8 FILLER_28_120 ();
 sg13g2_fill_4 FILLER_28_128 ();
 sg13g2_fill_2 FILLER_28_132 ();
 sg13g2_fill_8 FILLER_28_142 ();
 sg13g2_fill_8 FILLER_28_150 ();
 sg13g2_fill_2 FILLER_28_158 ();
 sg13g2_fill_1 FILLER_28_160 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_8 FILLER_28_203 ();
 sg13g2_fill_4 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_8 FILLER_28_349 ();
 sg13g2_fill_8 FILLER_28_357 ();
 sg13g2_fill_4 FILLER_28_365 ();
 sg13g2_fill_1 FILLER_28_369 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_fill_4 FILLER_28_387 ();
 sg13g2_fill_2 FILLER_28_399 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_441 ();
 sg13g2_fill_2 FILLER_28_467 ();
 sg13g2_fill_8 FILLER_28_472 ();
 sg13g2_fill_2 FILLER_28_480 ();
 sg13g2_fill_1 FILLER_28_482 ();
 sg13g2_fill_8 FILLER_28_515 ();
 sg13g2_fill_4 FILLER_28_523 ();
 sg13g2_fill_2 FILLER_28_559 ();
 sg13g2_fill_8 FILLER_28_566 ();
 sg13g2_fill_8 FILLER_28_574 ();
 sg13g2_fill_8 FILLER_28_582 ();
 sg13g2_fill_8 FILLER_28_590 ();
 sg13g2_fill_4 FILLER_28_598 ();
 sg13g2_fill_2 FILLER_28_602 ();
 sg13g2_fill_1 FILLER_28_604 ();
 sg13g2_fill_1 FILLER_28_635 ();
 sg13g2_fill_8 FILLER_28_662 ();
 sg13g2_fill_2 FILLER_28_670 ();
 sg13g2_fill_1 FILLER_28_672 ();
 sg13g2_fill_8 FILLER_28_699 ();
 sg13g2_fill_8 FILLER_28_717 ();
 sg13g2_fill_8 FILLER_28_725 ();
 sg13g2_fill_8 FILLER_28_733 ();
 sg13g2_fill_8 FILLER_28_741 ();
 sg13g2_fill_8 FILLER_28_749 ();
 sg13g2_fill_4 FILLER_28_757 ();
 sg13g2_fill_1 FILLER_28_761 ();
 sg13g2_fill_8 FILLER_28_766 ();
 sg13g2_fill_8 FILLER_28_774 ();
 sg13g2_fill_8 FILLER_28_782 ();
 sg13g2_fill_8 FILLER_28_790 ();
 sg13g2_fill_8 FILLER_28_798 ();
 sg13g2_fill_8 FILLER_28_806 ();
 sg13g2_fill_8 FILLER_28_814 ();
 sg13g2_fill_8 FILLER_28_822 ();
 sg13g2_fill_8 FILLER_28_830 ();
 sg13g2_fill_8 FILLER_28_838 ();
 sg13g2_fill_8 FILLER_28_846 ();
 sg13g2_fill_8 FILLER_28_854 ();
 sg13g2_fill_8 FILLER_28_862 ();
 sg13g2_fill_8 FILLER_28_870 ();
 sg13g2_fill_8 FILLER_28_878 ();
 sg13g2_fill_8 FILLER_28_886 ();
 sg13g2_fill_8 FILLER_28_894 ();
 sg13g2_fill_8 FILLER_28_902 ();
 sg13g2_fill_8 FILLER_28_910 ();
 sg13g2_fill_8 FILLER_28_918 ();
 sg13g2_fill_8 FILLER_28_926 ();
 sg13g2_fill_8 FILLER_28_934 ();
 sg13g2_fill_8 FILLER_28_942 ();
 sg13g2_fill_8 FILLER_28_950 ();
 sg13g2_fill_8 FILLER_28_958 ();
 sg13g2_fill_8 FILLER_28_966 ();
 sg13g2_fill_8 FILLER_28_974 ();
 sg13g2_fill_8 FILLER_28_982 ();
 sg13g2_fill_8 FILLER_28_990 ();
 sg13g2_fill_8 FILLER_28_998 ();
 sg13g2_fill_8 FILLER_28_1006 ();
 sg13g2_fill_8 FILLER_28_1014 ();
 sg13g2_fill_8 FILLER_28_1022 ();
 sg13g2_fill_8 FILLER_28_1030 ();
 sg13g2_fill_8 FILLER_28_1038 ();
 sg13g2_fill_8 FILLER_28_1046 ();
 sg13g2_fill_8 FILLER_28_1054 ();
 sg13g2_fill_8 FILLER_28_1062 ();
 sg13g2_fill_8 FILLER_28_1070 ();
 sg13g2_fill_8 FILLER_28_1078 ();
 sg13g2_fill_8 FILLER_28_1086 ();
 sg13g2_fill_8 FILLER_28_1094 ();
 sg13g2_fill_8 FILLER_28_1102 ();
 sg13g2_fill_8 FILLER_28_1110 ();
 sg13g2_fill_8 FILLER_28_1118 ();
 sg13g2_fill_8 FILLER_28_1126 ();
 sg13g2_fill_8 FILLER_28_1134 ();
 sg13g2_fill_8 FILLER_28_1142 ();
 sg13g2_fill_8 FILLER_28_1150 ();
 sg13g2_fill_8 FILLER_28_1158 ();
 sg13g2_fill_8 FILLER_29_0 ();
 sg13g2_fill_8 FILLER_29_8 ();
 sg13g2_fill_8 FILLER_29_16 ();
 sg13g2_fill_2 FILLER_29_24 ();
 sg13g2_fill_8 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_74 ();
 sg13g2_fill_1 FILLER_29_80 ();
 sg13g2_fill_8 FILLER_29_90 ();
 sg13g2_fill_4 FILLER_29_98 ();
 sg13g2_fill_4 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_4 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_159 ();
 sg13g2_fill_1 FILLER_29_161 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_4 FILLER_29_172 ();
 sg13g2_fill_1 FILLER_29_176 ();
 sg13g2_fill_8 FILLER_29_180 ();
 sg13g2_fill_4 FILLER_29_188 ();
 sg13g2_fill_1 FILLER_29_192 ();
 sg13g2_fill_8 FILLER_29_235 ();
 sg13g2_fill_8 FILLER_29_248 ();
 sg13g2_fill_2 FILLER_29_256 ();
 sg13g2_fill_4 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_269 ();
 sg13g2_fill_8 FILLER_29_296 ();
 sg13g2_fill_2 FILLER_29_304 ();
 sg13g2_fill_8 FILLER_29_331 ();
 sg13g2_fill_8 FILLER_29_339 ();
 sg13g2_fill_4 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_351 ();
 sg13g2_fill_1 FILLER_29_353 ();
 sg13g2_fill_8 FILLER_29_367 ();
 sg13g2_fill_8 FILLER_29_375 ();
 sg13g2_fill_8 FILLER_29_383 ();
 sg13g2_fill_8 FILLER_29_391 ();
 sg13g2_fill_8 FILLER_29_399 ();
 sg13g2_fill_8 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_29_415 ();
 sg13g2_fill_4 FILLER_29_419 ();
 sg13g2_fill_1 FILLER_29_423 ();
 sg13g2_fill_8 FILLER_29_429 ();
 sg13g2_fill_8 FILLER_29_437 ();
 sg13g2_fill_2 FILLER_29_445 ();
 sg13g2_fill_1 FILLER_29_447 ();
 sg13g2_fill_1 FILLER_29_466 ();
 sg13g2_fill_8 FILLER_29_472 ();
 sg13g2_fill_8 FILLER_29_480 ();
 sg13g2_fill_8 FILLER_29_488 ();
 sg13g2_fill_8 FILLER_29_496 ();
 sg13g2_fill_8 FILLER_29_504 ();
 sg13g2_fill_4 FILLER_29_512 ();
 sg13g2_fill_2 FILLER_29_516 ();
 sg13g2_fill_1 FILLER_29_552 ();
 sg13g2_fill_8 FILLER_29_572 ();
 sg13g2_fill_8 FILLER_29_580 ();
 sg13g2_fill_8 FILLER_29_588 ();
 sg13g2_fill_2 FILLER_29_596 ();
 sg13g2_fill_8 FILLER_29_624 ();
 sg13g2_fill_4 FILLER_29_632 ();
 sg13g2_fill_1 FILLER_29_636 ();
 sg13g2_fill_8 FILLER_29_663 ();
 sg13g2_fill_4 FILLER_29_671 ();
 sg13g2_fill_2 FILLER_29_675 ();
 sg13g2_fill_1 FILLER_29_677 ();
 sg13g2_fill_4 FILLER_29_704 ();
 sg13g2_fill_2 FILLER_29_708 ();
 sg13g2_fill_1 FILLER_29_710 ();
 sg13g2_fill_8 FILLER_29_737 ();
 sg13g2_fill_4 FILLER_29_745 ();
 sg13g2_fill_8 FILLER_29_785 ();
 sg13g2_fill_4 FILLER_29_793 ();
 sg13g2_fill_2 FILLER_29_797 ();
 sg13g2_fill_8 FILLER_29_807 ();
 sg13g2_fill_8 FILLER_29_815 ();
 sg13g2_fill_8 FILLER_29_823 ();
 sg13g2_fill_8 FILLER_29_831 ();
 sg13g2_fill_8 FILLER_29_839 ();
 sg13g2_fill_8 FILLER_29_847 ();
 sg13g2_fill_8 FILLER_29_855 ();
 sg13g2_fill_8 FILLER_29_863 ();
 sg13g2_fill_8 FILLER_29_871 ();
 sg13g2_fill_8 FILLER_29_879 ();
 sg13g2_fill_8 FILLER_29_887 ();
 sg13g2_fill_8 FILLER_29_895 ();
 sg13g2_fill_8 FILLER_29_903 ();
 sg13g2_fill_8 FILLER_29_911 ();
 sg13g2_fill_8 FILLER_29_919 ();
 sg13g2_fill_8 FILLER_29_927 ();
 sg13g2_fill_8 FILLER_29_935 ();
 sg13g2_fill_8 FILLER_29_943 ();
 sg13g2_fill_8 FILLER_29_951 ();
 sg13g2_fill_8 FILLER_29_959 ();
 sg13g2_fill_8 FILLER_29_967 ();
 sg13g2_fill_8 FILLER_29_975 ();
 sg13g2_fill_8 FILLER_29_983 ();
 sg13g2_fill_8 FILLER_29_991 ();
 sg13g2_fill_8 FILLER_29_999 ();
 sg13g2_fill_8 FILLER_29_1007 ();
 sg13g2_fill_8 FILLER_29_1015 ();
 sg13g2_fill_8 FILLER_29_1023 ();
 sg13g2_fill_8 FILLER_29_1031 ();
 sg13g2_fill_8 FILLER_29_1039 ();
 sg13g2_fill_8 FILLER_29_1047 ();
 sg13g2_fill_8 FILLER_29_1055 ();
 sg13g2_fill_8 FILLER_29_1063 ();
 sg13g2_fill_8 FILLER_29_1071 ();
 sg13g2_fill_8 FILLER_29_1079 ();
 sg13g2_fill_8 FILLER_29_1087 ();
 sg13g2_fill_8 FILLER_29_1095 ();
 sg13g2_fill_8 FILLER_29_1103 ();
 sg13g2_fill_8 FILLER_29_1111 ();
 sg13g2_fill_8 FILLER_29_1119 ();
 sg13g2_fill_8 FILLER_29_1127 ();
 sg13g2_fill_8 FILLER_29_1135 ();
 sg13g2_fill_8 FILLER_29_1143 ();
 sg13g2_fill_8 FILLER_29_1151 ();
 sg13g2_fill_4 FILLER_29_1159 ();
 sg13g2_fill_2 FILLER_29_1163 ();
 sg13g2_fill_1 FILLER_29_1165 ();
 sg13g2_fill_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_fill_4 FILLER_30_36 ();
 sg13g2_fill_2 FILLER_30_40 ();
 sg13g2_fill_1 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_48 ();
 sg13g2_fill_2 FILLER_30_76 ();
 sg13g2_fill_8 FILLER_30_87 ();
 sg13g2_fill_8 FILLER_30_95 ();
 sg13g2_fill_8 FILLER_30_103 ();
 sg13g2_fill_4 FILLER_30_111 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_160 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_8 FILLER_30_214 ();
 sg13g2_fill_8 FILLER_30_222 ();
 sg13g2_fill_8 FILLER_30_230 ();
 sg13g2_fill_2 FILLER_30_238 ();
 sg13g2_fill_8 FILLER_30_253 ();
 sg13g2_fill_8 FILLER_30_261 ();
 sg13g2_fill_8 FILLER_30_269 ();
 sg13g2_fill_8 FILLER_30_277 ();
 sg13g2_fill_4 FILLER_30_285 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_fill_8 FILLER_30_294 ();
 sg13g2_fill_8 FILLER_30_302 ();
 sg13g2_fill_8 FILLER_30_310 ();
 sg13g2_fill_1 FILLER_30_318 ();
 sg13g2_fill_4 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_349 ();
 sg13g2_fill_8 FILLER_30_363 ();
 sg13g2_fill_4 FILLER_30_371 ();
 sg13g2_fill_2 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_377 ();
 sg13g2_fill_8 FILLER_30_386 ();
 sg13g2_fill_4 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_fill_4 FILLER_30_404 ();
 sg13g2_fill_2 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_425 ();
 sg13g2_fill_4 FILLER_30_483 ();
 sg13g2_fill_2 FILLER_30_487 ();
 sg13g2_fill_8 FILLER_30_493 ();
 sg13g2_fill_4 FILLER_30_501 ();
 sg13g2_fill_1 FILLER_30_514 ();
 sg13g2_fill_2 FILLER_30_546 ();
 sg13g2_fill_1 FILLER_30_548 ();
 sg13g2_fill_2 FILLER_30_553 ();
 sg13g2_fill_1 FILLER_30_555 ();
 sg13g2_fill_2 FILLER_30_561 ();
 sg13g2_fill_1 FILLER_30_568 ();
 sg13g2_fill_8 FILLER_30_575 ();
 sg13g2_fill_8 FILLER_30_591 ();
 sg13g2_fill_4 FILLER_30_599 ();
 sg13g2_fill_2 FILLER_30_603 ();
 sg13g2_fill_1 FILLER_30_605 ();
 sg13g2_fill_8 FILLER_30_614 ();
 sg13g2_fill_8 FILLER_30_622 ();
 sg13g2_fill_8 FILLER_30_630 ();
 sg13g2_fill_8 FILLER_30_638 ();
 sg13g2_fill_2 FILLER_30_646 ();
 sg13g2_fill_8 FILLER_30_703 ();
 sg13g2_fill_1 FILLER_30_711 ();
 sg13g2_fill_8 FILLER_30_738 ();
 sg13g2_fill_2 FILLER_30_746 ();
 sg13g2_fill_1 FILLER_30_753 ();
 sg13g2_fill_8 FILLER_30_785 ();
 sg13g2_fill_8 FILLER_30_793 ();
 sg13g2_fill_2 FILLER_30_801 ();
 sg13g2_fill_1 FILLER_30_803 ();
 sg13g2_fill_2 FILLER_30_824 ();
 sg13g2_fill_8 FILLER_30_831 ();
 sg13g2_fill_2 FILLER_30_839 ();
 sg13g2_fill_1 FILLER_30_841 ();
 sg13g2_fill_2 FILLER_30_847 ();
 sg13g2_fill_8 FILLER_30_901 ();
 sg13g2_fill_8 FILLER_30_909 ();
 sg13g2_fill_8 FILLER_30_917 ();
 sg13g2_fill_8 FILLER_30_925 ();
 sg13g2_fill_8 FILLER_30_933 ();
 sg13g2_fill_8 FILLER_30_941 ();
 sg13g2_fill_8 FILLER_30_949 ();
 sg13g2_fill_8 FILLER_30_957 ();
 sg13g2_fill_8 FILLER_30_965 ();
 sg13g2_fill_8 FILLER_30_973 ();
 sg13g2_fill_8 FILLER_30_981 ();
 sg13g2_fill_8 FILLER_30_989 ();
 sg13g2_fill_8 FILLER_30_997 ();
 sg13g2_fill_8 FILLER_30_1005 ();
 sg13g2_fill_8 FILLER_30_1013 ();
 sg13g2_fill_8 FILLER_30_1021 ();
 sg13g2_fill_8 FILLER_30_1029 ();
 sg13g2_fill_8 FILLER_30_1037 ();
 sg13g2_fill_8 FILLER_30_1045 ();
 sg13g2_fill_8 FILLER_30_1053 ();
 sg13g2_fill_8 FILLER_30_1061 ();
 sg13g2_fill_8 FILLER_30_1069 ();
 sg13g2_fill_8 FILLER_30_1077 ();
 sg13g2_fill_8 FILLER_30_1085 ();
 sg13g2_fill_8 FILLER_30_1093 ();
 sg13g2_fill_8 FILLER_30_1101 ();
 sg13g2_fill_8 FILLER_30_1109 ();
 sg13g2_fill_8 FILLER_30_1117 ();
 sg13g2_fill_8 FILLER_30_1125 ();
 sg13g2_fill_8 FILLER_30_1133 ();
 sg13g2_fill_8 FILLER_30_1141 ();
 sg13g2_fill_8 FILLER_30_1149 ();
 sg13g2_fill_8 FILLER_30_1157 ();
 sg13g2_fill_1 FILLER_30_1165 ();
 sg13g2_fill_8 FILLER_31_0 ();
 sg13g2_fill_8 FILLER_31_8 ();
 sg13g2_fill_2 FILLER_31_16 ();
 sg13g2_fill_1 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_29 ();
 sg13g2_fill_8 FILLER_31_62 ();
 sg13g2_fill_4 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_76 ();
 sg13g2_fill_4 FILLER_31_98 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_4 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_132 ();
 sg13g2_fill_4 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_fill_4 FILLER_31_195 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_8 FILLER_31_210 ();
 sg13g2_fill_8 FILLER_31_218 ();
 sg13g2_fill_4 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_241 ();
 sg13g2_fill_8 FILLER_31_269 ();
 sg13g2_fill_8 FILLER_31_277 ();
 sg13g2_fill_8 FILLER_31_285 ();
 sg13g2_fill_8 FILLER_31_293 ();
 sg13g2_fill_2 FILLER_31_301 ();
 sg13g2_fill_2 FILLER_31_311 ();
 sg13g2_fill_4 FILLER_31_318 ();
 sg13g2_fill_8 FILLER_31_326 ();
 sg13g2_fill_8 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_342 ();
 sg13g2_fill_4 FILLER_31_357 ();
 sg13g2_fill_2 FILLER_31_361 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_fill_4 FILLER_31_390 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_4 FILLER_31_403 ();
 sg13g2_fill_1 FILLER_31_433 ();
 sg13g2_fill_2 FILLER_31_561 ();
 sg13g2_fill_4 FILLER_31_569 ();
 sg13g2_fill_2 FILLER_31_573 ();
 sg13g2_fill_1 FILLER_31_575 ();
 sg13g2_fill_2 FILLER_31_593 ();
 sg13g2_fill_8 FILLER_31_624 ();
 sg13g2_fill_4 FILLER_31_632 ();
 sg13g2_fill_2 FILLER_31_636 ();
 sg13g2_fill_2 FILLER_31_650 ();
 sg13g2_fill_1 FILLER_31_652 ();
 sg13g2_fill_8 FILLER_31_658 ();
 sg13g2_fill_8 FILLER_31_666 ();
 sg13g2_fill_8 FILLER_31_681 ();
 sg13g2_fill_4 FILLER_31_689 ();
 sg13g2_fill_2 FILLER_31_693 ();
 sg13g2_fill_4 FILLER_31_698 ();
 sg13g2_fill_1 FILLER_31_702 ();
 sg13g2_fill_1 FILLER_31_733 ();
 sg13g2_fill_8 FILLER_31_745 ();
 sg13g2_fill_2 FILLER_31_753 ();
 sg13g2_fill_1 FILLER_31_768 ();
 sg13g2_fill_8 FILLER_31_795 ();
 sg13g2_fill_1 FILLER_31_803 ();
 sg13g2_fill_2 FILLER_31_819 ();
 sg13g2_fill_1 FILLER_31_821 ();
 sg13g2_fill_8 FILLER_31_890 ();
 sg13g2_fill_4 FILLER_31_898 ();
 sg13g2_fill_8 FILLER_31_911 ();
 sg13g2_fill_4 FILLER_31_919 ();
 sg13g2_fill_1 FILLER_31_923 ();
 sg13g2_fill_8 FILLER_31_934 ();
 sg13g2_fill_8 FILLER_31_942 ();
 sg13g2_fill_8 FILLER_31_950 ();
 sg13g2_fill_8 FILLER_31_958 ();
 sg13g2_fill_8 FILLER_31_966 ();
 sg13g2_fill_8 FILLER_31_974 ();
 sg13g2_fill_8 FILLER_31_982 ();
 sg13g2_fill_8 FILLER_31_990 ();
 sg13g2_fill_8 FILLER_31_998 ();
 sg13g2_fill_8 FILLER_31_1006 ();
 sg13g2_fill_8 FILLER_31_1014 ();
 sg13g2_fill_8 FILLER_31_1022 ();
 sg13g2_fill_8 FILLER_31_1030 ();
 sg13g2_fill_8 FILLER_31_1038 ();
 sg13g2_fill_8 FILLER_31_1046 ();
 sg13g2_fill_8 FILLER_31_1054 ();
 sg13g2_fill_8 FILLER_31_1062 ();
 sg13g2_fill_8 FILLER_31_1070 ();
 sg13g2_fill_8 FILLER_31_1078 ();
 sg13g2_fill_8 FILLER_31_1086 ();
 sg13g2_fill_8 FILLER_31_1094 ();
 sg13g2_fill_8 FILLER_31_1102 ();
 sg13g2_fill_8 FILLER_31_1110 ();
 sg13g2_fill_8 FILLER_31_1118 ();
 sg13g2_fill_8 FILLER_31_1126 ();
 sg13g2_fill_8 FILLER_31_1134 ();
 sg13g2_fill_8 FILLER_31_1142 ();
 sg13g2_fill_8 FILLER_31_1150 ();
 sg13g2_fill_8 FILLER_31_1158 ();
 sg13g2_fill_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_6 ();
 sg13g2_fill_8 FILLER_32_36 ();
 sg13g2_fill_8 FILLER_32_44 ();
 sg13g2_fill_4 FILLER_32_52 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_fill_8 FILLER_32_153 ();
 sg13g2_fill_1 FILLER_32_161 ();
 sg13g2_fill_8 FILLER_32_167 ();
 sg13g2_fill_4 FILLER_32_175 ();
 sg13g2_fill_8 FILLER_32_190 ();
 sg13g2_fill_8 FILLER_32_198 ();
 sg13g2_fill_8 FILLER_32_206 ();
 sg13g2_fill_8 FILLER_32_214 ();
 sg13g2_fill_8 FILLER_32_233 ();
 sg13g2_fill_8 FILLER_32_241 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_8 FILLER_32_304 ();
 sg13g2_fill_8 FILLER_32_312 ();
 sg13g2_fill_8 FILLER_32_320 ();
 sg13g2_fill_8 FILLER_32_328 ();
 sg13g2_fill_8 FILLER_32_336 ();
 sg13g2_fill_2 FILLER_32_344 ();
 sg13g2_fill_8 FILLER_32_414 ();
 sg13g2_fill_8 FILLER_32_422 ();
 sg13g2_fill_2 FILLER_32_430 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_4 FILLER_32_438 ();
 sg13g2_fill_2 FILLER_32_442 ();
 sg13g2_fill_1 FILLER_32_444 ();
 sg13g2_fill_4 FILLER_32_471 ();
 sg13g2_fill_2 FILLER_32_496 ();
 sg13g2_fill_1 FILLER_32_498 ();
 sg13g2_fill_2 FILLER_32_509 ();
 sg13g2_fill_1 FILLER_32_511 ();
 sg13g2_fill_4 FILLER_32_515 ();
 sg13g2_fill_2 FILLER_32_519 ();
 sg13g2_fill_2 FILLER_32_552 ();
 sg13g2_fill_1 FILLER_32_554 ();
 sg13g2_fill_4 FILLER_32_566 ();
 sg13g2_fill_1 FILLER_32_570 ();
 sg13g2_fill_8 FILLER_32_575 ();
 sg13g2_fill_4 FILLER_32_583 ();
 sg13g2_fill_4 FILLER_32_592 ();
 sg13g2_fill_2 FILLER_32_596 ();
 sg13g2_fill_1 FILLER_32_598 ();
 sg13g2_fill_4 FILLER_32_624 ();
 sg13g2_fill_2 FILLER_32_628 ();
 sg13g2_fill_1 FILLER_32_630 ();
 sg13g2_fill_1 FILLER_32_636 ();
 sg13g2_fill_2 FILLER_32_642 ();
 sg13g2_fill_2 FILLER_32_664 ();
 sg13g2_fill_8 FILLER_32_681 ();
 sg13g2_fill_8 FILLER_32_689 ();
 sg13g2_fill_4 FILLER_32_697 ();
 sg13g2_fill_2 FILLER_32_701 ();
 sg13g2_fill_4 FILLER_32_742 ();
 sg13g2_fill_2 FILLER_32_746 ();
 sg13g2_fill_8 FILLER_32_753 ();
 sg13g2_fill_8 FILLER_32_761 ();
 sg13g2_fill_2 FILLER_32_769 ();
 sg13g2_fill_1 FILLER_32_771 ();
 sg13g2_fill_4 FILLER_32_782 ();
 sg13g2_fill_1 FILLER_32_786 ();
 sg13g2_fill_8 FILLER_32_791 ();
 sg13g2_fill_4 FILLER_32_799 ();
 sg13g2_fill_8 FILLER_32_828 ();
 sg13g2_fill_8 FILLER_32_836 ();
 sg13g2_fill_4 FILLER_32_844 ();
 sg13g2_fill_2 FILLER_32_848 ();
 sg13g2_fill_2 FILLER_32_855 ();
 sg13g2_fill_2 FILLER_32_863 ();
 sg13g2_fill_1 FILLER_32_865 ();
 sg13g2_fill_8 FILLER_32_879 ();
 sg13g2_fill_4 FILLER_32_887 ();
 sg13g2_fill_8 FILLER_32_947 ();
 sg13g2_fill_8 FILLER_32_955 ();
 sg13g2_fill_8 FILLER_32_963 ();
 sg13g2_fill_8 FILLER_32_971 ();
 sg13g2_fill_8 FILLER_32_979 ();
 sg13g2_fill_8 FILLER_32_987 ();
 sg13g2_fill_8 FILLER_32_995 ();
 sg13g2_fill_8 FILLER_32_1003 ();
 sg13g2_fill_8 FILLER_32_1011 ();
 sg13g2_fill_8 FILLER_32_1019 ();
 sg13g2_fill_8 FILLER_32_1027 ();
 sg13g2_fill_8 FILLER_32_1035 ();
 sg13g2_fill_8 FILLER_32_1043 ();
 sg13g2_fill_8 FILLER_32_1051 ();
 sg13g2_fill_8 FILLER_32_1059 ();
 sg13g2_fill_8 FILLER_32_1067 ();
 sg13g2_fill_8 FILLER_32_1075 ();
 sg13g2_fill_8 FILLER_32_1083 ();
 sg13g2_fill_8 FILLER_32_1091 ();
 sg13g2_fill_8 FILLER_32_1099 ();
 sg13g2_fill_8 FILLER_32_1107 ();
 sg13g2_fill_8 FILLER_32_1115 ();
 sg13g2_fill_8 FILLER_32_1123 ();
 sg13g2_fill_8 FILLER_32_1131 ();
 sg13g2_fill_8 FILLER_32_1139 ();
 sg13g2_fill_8 FILLER_32_1147 ();
 sg13g2_fill_8 FILLER_32_1155 ();
 sg13g2_fill_2 FILLER_32_1163 ();
 sg13g2_fill_1 FILLER_32_1165 ();
 sg13g2_fill_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_fill_1 FILLER_33_6 ();
 sg13g2_fill_4 FILLER_33_38 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_fill_8 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_99 ();
 sg13g2_fill_1 FILLER_33_101 ();
 sg13g2_fill_2 FILLER_33_118 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_8 FILLER_33_176 ();
 sg13g2_fill_8 FILLER_33_184 ();
 sg13g2_fill_8 FILLER_33_192 ();
 sg13g2_fill_8 FILLER_33_200 ();
 sg13g2_fill_8 FILLER_33_208 ();
 sg13g2_fill_2 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_fill_4 FILLER_33_279 ();
 sg13g2_fill_4 FILLER_33_287 ();
 sg13g2_fill_8 FILLER_33_297 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_4 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_341 ();
 sg13g2_fill_1 FILLER_33_343 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_8 FILLER_33_403 ();
 sg13g2_fill_8 FILLER_33_411 ();
 sg13g2_fill_8 FILLER_33_419 ();
 sg13g2_fill_8 FILLER_33_427 ();
 sg13g2_fill_8 FILLER_33_435 ();
 sg13g2_fill_8 FILLER_33_443 ();
 sg13g2_fill_8 FILLER_33_451 ();
 sg13g2_fill_8 FILLER_33_459 ();
 sg13g2_fill_1 FILLER_33_467 ();
 sg13g2_fill_2 FILLER_33_491 ();
 sg13g2_fill_1 FILLER_33_493 ();
 sg13g2_fill_1 FILLER_33_499 ();
 sg13g2_fill_4 FILLER_33_505 ();
 sg13g2_fill_1 FILLER_33_509 ();
 sg13g2_fill_8 FILLER_33_516 ();
 sg13g2_fill_4 FILLER_33_524 ();
 sg13g2_fill_8 FILLER_33_533 ();
 sg13g2_fill_4 FILLER_33_541 ();
 sg13g2_fill_2 FILLER_33_545 ();
 sg13g2_fill_4 FILLER_33_555 ();
 sg13g2_fill_2 FILLER_33_559 ();
 sg13g2_fill_1 FILLER_33_561 ();
 sg13g2_fill_8 FILLER_33_566 ();
 sg13g2_fill_8 FILLER_33_574 ();
 sg13g2_fill_1 FILLER_33_582 ();
 sg13g2_fill_4 FILLER_33_588 ();
 sg13g2_fill_2 FILLER_33_592 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_2 FILLER_33_612 ();
 sg13g2_fill_4 FILLER_33_626 ();
 sg13g2_fill_2 FILLER_33_630 ();
 sg13g2_fill_4 FILLER_33_638 ();
 sg13g2_fill_1 FILLER_33_642 ();
 sg13g2_fill_8 FILLER_33_663 ();
 sg13g2_fill_8 FILLER_33_671 ();
 sg13g2_fill_8 FILLER_33_679 ();
 sg13g2_fill_2 FILLER_33_687 ();
 sg13g2_fill_1 FILLER_33_689 ();
 sg13g2_fill_8 FILLER_33_695 ();
 sg13g2_fill_4 FILLER_33_703 ();
 sg13g2_fill_2 FILLER_33_707 ();
 sg13g2_fill_1 FILLER_33_709 ();
 sg13g2_fill_1 FILLER_33_724 ();
 sg13g2_fill_8 FILLER_33_730 ();
 sg13g2_fill_8 FILLER_33_738 ();
 sg13g2_fill_8 FILLER_33_746 ();
 sg13g2_fill_8 FILLER_33_754 ();
 sg13g2_fill_4 FILLER_33_762 ();
 sg13g2_fill_2 FILLER_33_766 ();
 sg13g2_fill_4 FILLER_33_798 ();
 sg13g2_fill_1 FILLER_33_802 ();
 sg13g2_fill_8 FILLER_33_826 ();
 sg13g2_fill_4 FILLER_33_834 ();
 sg13g2_fill_8 FILLER_33_846 ();
 sg13g2_fill_4 FILLER_33_854 ();
 sg13g2_fill_4 FILLER_33_868 ();
 sg13g2_fill_2 FILLER_33_872 ();
 sg13g2_fill_2 FILLER_33_903 ();
 sg13g2_fill_2 FILLER_33_935 ();
 sg13g2_fill_8 FILLER_33_945 ();
 sg13g2_fill_8 FILLER_33_953 ();
 sg13g2_fill_8 FILLER_33_961 ();
 sg13g2_fill_8 FILLER_33_969 ();
 sg13g2_fill_8 FILLER_33_977 ();
 sg13g2_fill_8 FILLER_33_985 ();
 sg13g2_fill_8 FILLER_33_993 ();
 sg13g2_fill_8 FILLER_33_1001 ();
 sg13g2_fill_8 FILLER_33_1009 ();
 sg13g2_fill_8 FILLER_33_1017 ();
 sg13g2_fill_8 FILLER_33_1025 ();
 sg13g2_fill_8 FILLER_33_1033 ();
 sg13g2_fill_8 FILLER_33_1041 ();
 sg13g2_fill_8 FILLER_33_1049 ();
 sg13g2_fill_8 FILLER_33_1057 ();
 sg13g2_fill_8 FILLER_33_1065 ();
 sg13g2_fill_8 FILLER_33_1073 ();
 sg13g2_fill_8 FILLER_33_1081 ();
 sg13g2_fill_8 FILLER_33_1089 ();
 sg13g2_fill_8 FILLER_33_1097 ();
 sg13g2_fill_8 FILLER_33_1105 ();
 sg13g2_fill_8 FILLER_33_1113 ();
 sg13g2_fill_8 FILLER_33_1121 ();
 sg13g2_fill_8 FILLER_33_1129 ();
 sg13g2_fill_8 FILLER_33_1137 ();
 sg13g2_fill_8 FILLER_33_1145 ();
 sg13g2_fill_8 FILLER_33_1153 ();
 sg13g2_fill_4 FILLER_33_1161 ();
 sg13g2_fill_1 FILLER_33_1165 ();
 sg13g2_fill_8 FILLER_34_0 ();
 sg13g2_fill_4 FILLER_34_8 ();
 sg13g2_fill_1 FILLER_34_12 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_fill_8 FILLER_34_59 ();
 sg13g2_fill_4 FILLER_34_67 ();
 sg13g2_fill_8 FILLER_34_86 ();
 sg13g2_fill_8 FILLER_34_94 ();
 sg13g2_fill_4 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_fill_4 FILLER_34_166 ();
 sg13g2_fill_4 FILLER_34_200 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_8 FILLER_34_240 ();
 sg13g2_fill_8 FILLER_34_248 ();
 sg13g2_fill_4 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_348 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_372 ();
 sg13g2_fill_4 FILLER_34_407 ();
 sg13g2_fill_2 FILLER_34_411 ();
 sg13g2_fill_1 FILLER_34_413 ();
 sg13g2_fill_4 FILLER_34_453 ();
 sg13g2_fill_2 FILLER_34_457 ();
 sg13g2_fill_8 FILLER_34_465 ();
 sg13g2_fill_8 FILLER_34_473 ();
 sg13g2_fill_8 FILLER_34_501 ();
 sg13g2_fill_8 FILLER_34_509 ();
 sg13g2_fill_4 FILLER_34_517 ();
 sg13g2_fill_4 FILLER_34_533 ();
 sg13g2_fill_2 FILLER_34_537 ();
 sg13g2_fill_4 FILLER_34_544 ();
 sg13g2_fill_1 FILLER_34_560 ();
 sg13g2_fill_4 FILLER_34_573 ();
 sg13g2_fill_4 FILLER_34_582 ();
 sg13g2_fill_2 FILLER_34_586 ();
 sg13g2_fill_4 FILLER_34_594 ();
 sg13g2_fill_2 FILLER_34_598 ();
 sg13g2_fill_1 FILLER_34_600 ();
 sg13g2_fill_2 FILLER_34_606 ();
 sg13g2_fill_1 FILLER_34_608 ();
 sg13g2_fill_2 FILLER_34_617 ();
 sg13g2_fill_1 FILLER_34_619 ();
 sg13g2_fill_1 FILLER_34_634 ();
 sg13g2_fill_8 FILLER_34_640 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_fill_1 FILLER_34_663 ();
 sg13g2_fill_2 FILLER_34_694 ();
 sg13g2_fill_1 FILLER_34_696 ();
 sg13g2_fill_8 FILLER_34_728 ();
 sg13g2_fill_2 FILLER_34_768 ();
 sg13g2_fill_2 FILLER_34_800 ();
 sg13g2_fill_2 FILLER_34_807 ();
 sg13g2_fill_8 FILLER_34_828 ();
 sg13g2_fill_8 FILLER_34_836 ();
 sg13g2_fill_2 FILLER_34_854 ();
 sg13g2_fill_4 FILLER_34_865 ();
 sg13g2_fill_2 FILLER_34_869 ();
 sg13g2_fill_8 FILLER_34_892 ();
 sg13g2_fill_2 FILLER_34_900 ();
 sg13g2_fill_8 FILLER_34_945 ();
 sg13g2_fill_8 FILLER_34_953 ();
 sg13g2_fill_8 FILLER_34_961 ();
 sg13g2_fill_8 FILLER_34_969 ();
 sg13g2_fill_8 FILLER_34_977 ();
 sg13g2_fill_8 FILLER_34_985 ();
 sg13g2_fill_8 FILLER_34_993 ();
 sg13g2_fill_8 FILLER_34_1001 ();
 sg13g2_fill_8 FILLER_34_1009 ();
 sg13g2_fill_8 FILLER_34_1017 ();
 sg13g2_fill_8 FILLER_34_1025 ();
 sg13g2_fill_8 FILLER_34_1033 ();
 sg13g2_fill_8 FILLER_34_1041 ();
 sg13g2_fill_8 FILLER_34_1049 ();
 sg13g2_fill_8 FILLER_34_1057 ();
 sg13g2_fill_8 FILLER_34_1065 ();
 sg13g2_fill_8 FILLER_34_1073 ();
 sg13g2_fill_8 FILLER_34_1081 ();
 sg13g2_fill_8 FILLER_34_1089 ();
 sg13g2_fill_8 FILLER_34_1097 ();
 sg13g2_fill_8 FILLER_34_1105 ();
 sg13g2_fill_8 FILLER_34_1113 ();
 sg13g2_fill_8 FILLER_34_1121 ();
 sg13g2_fill_8 FILLER_34_1129 ();
 sg13g2_fill_8 FILLER_34_1137 ();
 sg13g2_fill_8 FILLER_34_1145 ();
 sg13g2_fill_8 FILLER_34_1153 ();
 sg13g2_fill_4 FILLER_34_1161 ();
 sg13g2_fill_1 FILLER_34_1165 ();
 sg13g2_fill_8 FILLER_35_0 ();
 sg13g2_fill_4 FILLER_35_8 ();
 sg13g2_fill_8 FILLER_35_16 ();
 sg13g2_fill_8 FILLER_35_24 ();
 sg13g2_fill_8 FILLER_35_32 ();
 sg13g2_fill_8 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_73 ();
 sg13g2_fill_8 FILLER_35_79 ();
 sg13g2_fill_8 FILLER_35_87 ();
 sg13g2_fill_4 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_2 FILLER_35_131 ();
 sg13g2_fill_1 FILLER_35_133 ();
 sg13g2_fill_8 FILLER_35_155 ();
 sg13g2_fill_8 FILLER_35_163 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_4 FILLER_35_245 ();
 sg13g2_fill_1 FILLER_35_249 ();
 sg13g2_fill_2 FILLER_35_277 ();
 sg13g2_fill_1 FILLER_35_279 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_fill_4 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_320 ();
 sg13g2_fill_4 FILLER_35_325 ();
 sg13g2_fill_2 FILLER_35_335 ();
 sg13g2_fill_1 FILLER_35_337 ();
 sg13g2_fill_2 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_401 ();
 sg13g2_fill_4 FILLER_35_440 ();
 sg13g2_fill_2 FILLER_35_444 ();
 sg13g2_fill_1 FILLER_35_472 ();
 sg13g2_fill_4 FILLER_35_479 ();
 sg13g2_fill_2 FILLER_35_489 ();
 sg13g2_fill_2 FILLER_35_499 ();
 sg13g2_fill_2 FILLER_35_509 ();
 sg13g2_fill_8 FILLER_35_517 ();
 sg13g2_fill_8 FILLER_35_525 ();
 sg13g2_fill_8 FILLER_35_533 ();
 sg13g2_fill_8 FILLER_35_541 ();
 sg13g2_fill_4 FILLER_35_549 ();
 sg13g2_fill_1 FILLER_35_553 ();
 sg13g2_fill_8 FILLER_35_593 ();
 sg13g2_fill_8 FILLER_35_601 ();
 sg13g2_fill_4 FILLER_35_609 ();
 sg13g2_fill_2 FILLER_35_613 ();
 sg13g2_fill_1 FILLER_35_615 ();
 sg13g2_fill_4 FILLER_35_630 ();
 sg13g2_fill_2 FILLER_35_634 ();
 sg13g2_fill_4 FILLER_35_650 ();
 sg13g2_fill_2 FILLER_35_654 ();
 sg13g2_fill_1 FILLER_35_656 ();
 sg13g2_fill_2 FILLER_35_724 ();
 sg13g2_fill_2 FILLER_35_770 ();
 sg13g2_fill_4 FILLER_35_798 ();
 sg13g2_fill_4 FILLER_35_827 ();
 sg13g2_fill_2 FILLER_35_831 ();
 sg13g2_fill_1 FILLER_35_842 ();
 sg13g2_fill_1 FILLER_35_848 ();
 sg13g2_fill_1 FILLER_35_870 ();
 sg13g2_fill_2 FILLER_35_876 ();
 sg13g2_fill_8 FILLER_35_892 ();
 sg13g2_fill_8 FILLER_35_900 ();
 sg13g2_fill_4 FILLER_35_908 ();
 sg13g2_fill_1 FILLER_35_912 ();
 sg13g2_fill_2 FILLER_35_918 ();
 sg13g2_fill_8 FILLER_35_936 ();
 sg13g2_fill_8 FILLER_35_944 ();
 sg13g2_fill_8 FILLER_35_952 ();
 sg13g2_fill_8 FILLER_35_960 ();
 sg13g2_fill_8 FILLER_35_968 ();
 sg13g2_fill_8 FILLER_35_976 ();
 sg13g2_fill_8 FILLER_35_984 ();
 sg13g2_fill_8 FILLER_35_992 ();
 sg13g2_fill_8 FILLER_35_1000 ();
 sg13g2_fill_8 FILLER_35_1008 ();
 sg13g2_fill_8 FILLER_35_1016 ();
 sg13g2_fill_8 FILLER_35_1024 ();
 sg13g2_fill_8 FILLER_35_1032 ();
 sg13g2_fill_8 FILLER_35_1040 ();
 sg13g2_fill_8 FILLER_35_1048 ();
 sg13g2_fill_8 FILLER_35_1056 ();
 sg13g2_fill_8 FILLER_35_1064 ();
 sg13g2_fill_8 FILLER_35_1072 ();
 sg13g2_fill_8 FILLER_35_1080 ();
 sg13g2_fill_8 FILLER_35_1088 ();
 sg13g2_fill_8 FILLER_35_1096 ();
 sg13g2_fill_8 FILLER_35_1104 ();
 sg13g2_fill_8 FILLER_35_1112 ();
 sg13g2_fill_8 FILLER_35_1120 ();
 sg13g2_fill_8 FILLER_35_1128 ();
 sg13g2_fill_8 FILLER_35_1136 ();
 sg13g2_fill_8 FILLER_35_1144 ();
 sg13g2_fill_8 FILLER_35_1152 ();
 sg13g2_fill_4 FILLER_35_1160 ();
 sg13g2_fill_2 FILLER_35_1164 ();
 sg13g2_fill_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_2 FILLER_36_19 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_fill_2 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_78 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_fill_8 FILLER_36_122 ();
 sg13g2_fill_4 FILLER_36_130 ();
 sg13g2_fill_8 FILLER_36_155 ();
 sg13g2_fill_8 FILLER_36_163 ();
 sg13g2_fill_8 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_4 FILLER_36_189 ();
 sg13g2_fill_8 FILLER_36_202 ();
 sg13g2_fill_2 FILLER_36_210 ();
 sg13g2_fill_8 FILLER_36_221 ();
 sg13g2_fill_8 FILLER_36_229 ();
 sg13g2_fill_4 FILLER_36_237 ();
 sg13g2_fill_2 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_243 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_fill_1 FILLER_36_309 ();
 sg13g2_fill_4 FILLER_36_333 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_4 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_2 FILLER_36_384 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_4 FILLER_36_401 ();
 sg13g2_fill_4 FILLER_36_410 ();
 sg13g2_fill_1 FILLER_36_419 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_fill_2 FILLER_36_435 ();
 sg13g2_fill_1 FILLER_36_437 ();
 sg13g2_fill_4 FILLER_36_442 ();
 sg13g2_fill_1 FILLER_36_446 ();
 sg13g2_fill_8 FILLER_36_452 ();
 sg13g2_fill_8 FILLER_36_460 ();
 sg13g2_fill_8 FILLER_36_468 ();
 sg13g2_fill_4 FILLER_36_476 ();
 sg13g2_fill_2 FILLER_36_480 ();
 sg13g2_fill_4 FILLER_36_495 ();
 sg13g2_fill_8 FILLER_36_509 ();
 sg13g2_fill_8 FILLER_36_530 ();
 sg13g2_fill_4 FILLER_36_538 ();
 sg13g2_fill_2 FILLER_36_542 ();
 sg13g2_fill_1 FILLER_36_560 ();
 sg13g2_fill_8 FILLER_36_566 ();
 sg13g2_fill_8 FILLER_36_574 ();
 sg13g2_fill_1 FILLER_36_582 ();
 sg13g2_fill_4 FILLER_36_588 ();
 sg13g2_fill_2 FILLER_36_592 ();
 sg13g2_fill_8 FILLER_36_599 ();
 sg13g2_fill_8 FILLER_36_607 ();
 sg13g2_fill_8 FILLER_36_615 ();
 sg13g2_fill_8 FILLER_36_623 ();
 sg13g2_fill_2 FILLER_36_631 ();
 sg13g2_fill_8 FILLER_36_638 ();
 sg13g2_fill_1 FILLER_36_646 ();
 sg13g2_fill_2 FILLER_36_652 ();
 sg13g2_fill_8 FILLER_36_659 ();
 sg13g2_fill_1 FILLER_36_667 ();
 sg13g2_fill_2 FILLER_36_713 ();
 sg13g2_fill_2 FILLER_36_725 ();
 sg13g2_fill_2 FILLER_36_732 ();
 sg13g2_fill_4 FILLER_36_739 ();
 sg13g2_fill_2 FILLER_36_743 ();
 sg13g2_fill_8 FILLER_36_756 ();
 sg13g2_fill_8 FILLER_36_795 ();
 sg13g2_fill_8 FILLER_36_803 ();
 sg13g2_fill_2 FILLER_36_811 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_fill_1 FILLER_36_819 ();
 sg13g2_fill_8 FILLER_36_824 ();
 sg13g2_fill_1 FILLER_36_832 ();
 sg13g2_fill_1 FILLER_36_838 ();
 sg13g2_fill_8 FILLER_36_864 ();
 sg13g2_fill_4 FILLER_36_872 ();
 sg13g2_fill_2 FILLER_36_876 ();
 sg13g2_fill_1 FILLER_36_884 ();
 sg13g2_fill_8 FILLER_36_891 ();
 sg13g2_fill_4 FILLER_36_899 ();
 sg13g2_fill_1 FILLER_36_907 ();
 sg13g2_fill_8 FILLER_36_935 ();
 sg13g2_fill_8 FILLER_36_943 ();
 sg13g2_fill_8 FILLER_36_951 ();
 sg13g2_fill_8 FILLER_36_959 ();
 sg13g2_fill_8 FILLER_36_967 ();
 sg13g2_fill_8 FILLER_36_975 ();
 sg13g2_fill_8 FILLER_36_983 ();
 sg13g2_fill_8 FILLER_36_991 ();
 sg13g2_fill_8 FILLER_36_999 ();
 sg13g2_fill_8 FILLER_36_1007 ();
 sg13g2_fill_8 FILLER_36_1015 ();
 sg13g2_fill_8 FILLER_36_1023 ();
 sg13g2_fill_8 FILLER_36_1031 ();
 sg13g2_fill_8 FILLER_36_1039 ();
 sg13g2_fill_8 FILLER_36_1047 ();
 sg13g2_fill_8 FILLER_36_1055 ();
 sg13g2_fill_8 FILLER_36_1063 ();
 sg13g2_fill_8 FILLER_36_1071 ();
 sg13g2_fill_8 FILLER_36_1079 ();
 sg13g2_fill_8 FILLER_36_1087 ();
 sg13g2_fill_8 FILLER_36_1095 ();
 sg13g2_fill_8 FILLER_36_1103 ();
 sg13g2_fill_8 FILLER_36_1111 ();
 sg13g2_fill_8 FILLER_36_1119 ();
 sg13g2_fill_8 FILLER_36_1127 ();
 sg13g2_fill_8 FILLER_36_1135 ();
 sg13g2_fill_8 FILLER_36_1143 ();
 sg13g2_fill_8 FILLER_36_1151 ();
 sg13g2_fill_4 FILLER_36_1159 ();
 sg13g2_fill_2 FILLER_36_1163 ();
 sg13g2_fill_1 FILLER_36_1165 ();
 sg13g2_fill_8 FILLER_37_0 ();
 sg13g2_fill_4 FILLER_37_8 ();
 sg13g2_fill_2 FILLER_37_12 ();
 sg13g2_fill_4 FILLER_37_102 ();
 sg13g2_fill_2 FILLER_37_106 ();
 sg13g2_fill_8 FILLER_37_119 ();
 sg13g2_fill_8 FILLER_37_127 ();
 sg13g2_fill_8 FILLER_37_156 ();
 sg13g2_fill_8 FILLER_37_164 ();
 sg13g2_fill_4 FILLER_37_172 ();
 sg13g2_fill_2 FILLER_37_176 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_198 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_2 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_fill_8 FILLER_37_286 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_fill_8 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_326 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_8 FILLER_37_342 ();
 sg13g2_fill_8 FILLER_37_350 ();
 sg13g2_fill_1 FILLER_37_358 ();
 sg13g2_fill_2 FILLER_37_373 ();
 sg13g2_fill_1 FILLER_37_375 ();
 sg13g2_fill_8 FILLER_37_407 ();
 sg13g2_fill_1 FILLER_37_415 ();
 sg13g2_fill_1 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_435 ();
 sg13g2_fill_8 FILLER_37_463 ();
 sg13g2_fill_8 FILLER_37_471 ();
 sg13g2_fill_2 FILLER_37_479 ();
 sg13g2_fill_1 FILLER_37_481 ();
 sg13g2_fill_8 FILLER_37_495 ();
 sg13g2_fill_1 FILLER_37_503 ();
 sg13g2_fill_2 FILLER_37_512 ();
 sg13g2_fill_4 FILLER_37_543 ();
 sg13g2_fill_1 FILLER_37_547 ();
 sg13g2_fill_4 FILLER_37_558 ();
 sg13g2_fill_1 FILLER_37_562 ();
 sg13g2_fill_8 FILLER_37_567 ();
 sg13g2_fill_1 FILLER_37_575 ();
 sg13g2_fill_4 FILLER_37_586 ();
 sg13g2_fill_4 FILLER_37_622 ();
 sg13g2_fill_2 FILLER_37_626 ();
 sg13g2_fill_1 FILLER_37_628 ();
 sg13g2_fill_8 FILLER_37_663 ();
 sg13g2_fill_4 FILLER_37_671 ();
 sg13g2_fill_2 FILLER_37_675 ();
 sg13g2_fill_1 FILLER_37_677 ();
 sg13g2_fill_8 FILLER_37_683 ();
 sg13g2_fill_1 FILLER_37_691 ();
 sg13g2_fill_8 FILLER_37_695 ();
 sg13g2_fill_8 FILLER_37_703 ();
 sg13g2_fill_8 FILLER_37_711 ();
 sg13g2_fill_8 FILLER_37_719 ();
 sg13g2_fill_2 FILLER_37_727 ();
 sg13g2_fill_8 FILLER_37_760 ();
 sg13g2_fill_1 FILLER_37_768 ();
 sg13g2_fill_8 FILLER_37_778 ();
 sg13g2_fill_8 FILLER_37_786 ();
 sg13g2_fill_8 FILLER_37_794 ();
 sg13g2_fill_8 FILLER_37_802 ();
 sg13g2_fill_8 FILLER_37_810 ();
 sg13g2_fill_8 FILLER_37_818 ();
 sg13g2_fill_2 FILLER_37_826 ();
 sg13g2_fill_8 FILLER_37_833 ();
 sg13g2_fill_4 FILLER_37_841 ();
 sg13g2_fill_1 FILLER_37_845 ();
 sg13g2_fill_2 FILLER_37_855 ();
 sg13g2_fill_1 FILLER_37_857 ();
 sg13g2_fill_8 FILLER_37_892 ();
 sg13g2_fill_2 FILLER_37_900 ();
 sg13g2_fill_1 FILLER_37_902 ();
 sg13g2_fill_1 FILLER_37_909 ();
 sg13g2_fill_1 FILLER_37_925 ();
 sg13g2_fill_4 FILLER_37_930 ();
 sg13g2_fill_8 FILLER_37_945 ();
 sg13g2_fill_8 FILLER_37_953 ();
 sg13g2_fill_8 FILLER_37_961 ();
 sg13g2_fill_8 FILLER_37_969 ();
 sg13g2_fill_8 FILLER_37_977 ();
 sg13g2_fill_8 FILLER_37_985 ();
 sg13g2_fill_8 FILLER_37_993 ();
 sg13g2_fill_8 FILLER_37_1001 ();
 sg13g2_fill_8 FILLER_37_1009 ();
 sg13g2_fill_8 FILLER_37_1017 ();
 sg13g2_fill_8 FILLER_37_1025 ();
 sg13g2_fill_8 FILLER_37_1033 ();
 sg13g2_fill_8 FILLER_37_1041 ();
 sg13g2_fill_8 FILLER_37_1049 ();
 sg13g2_fill_8 FILLER_37_1057 ();
 sg13g2_fill_8 FILLER_37_1065 ();
 sg13g2_fill_8 FILLER_37_1073 ();
 sg13g2_fill_8 FILLER_37_1081 ();
 sg13g2_fill_8 FILLER_37_1089 ();
 sg13g2_fill_8 FILLER_37_1097 ();
 sg13g2_fill_8 FILLER_37_1105 ();
 sg13g2_fill_8 FILLER_37_1113 ();
 sg13g2_fill_8 FILLER_37_1121 ();
 sg13g2_fill_8 FILLER_37_1129 ();
 sg13g2_fill_8 FILLER_37_1137 ();
 sg13g2_fill_8 FILLER_37_1145 ();
 sg13g2_fill_8 FILLER_37_1153 ();
 sg13g2_fill_4 FILLER_37_1161 ();
 sg13g2_fill_1 FILLER_37_1165 ();
 sg13g2_fill_2 FILLER_38_29 ();
 sg13g2_fill_2 FILLER_38_36 ();
 sg13g2_fill_8 FILLER_38_41 ();
 sg13g2_fill_8 FILLER_38_49 ();
 sg13g2_fill_8 FILLER_38_57 ();
 sg13g2_fill_8 FILLER_38_65 ();
 sg13g2_fill_4 FILLER_38_73 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_fill_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_100 ();
 sg13g2_fill_8 FILLER_38_105 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_144 ();
 sg13g2_fill_1 FILLER_38_148 ();
 sg13g2_fill_8 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_8 FILLER_38_225 ();
 sg13g2_fill_1 FILLER_38_233 ();
 sg13g2_fill_4 FILLER_38_239 ();
 sg13g2_fill_8 FILLER_38_256 ();
 sg13g2_fill_4 FILLER_38_264 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_270 ();
 sg13g2_fill_8 FILLER_38_280 ();
 sg13g2_fill_8 FILLER_38_288 ();
 sg13g2_fill_4 FILLER_38_296 ();
 sg13g2_fill_8 FILLER_38_305 ();
 sg13g2_fill_8 FILLER_38_313 ();
 sg13g2_fill_8 FILLER_38_321 ();
 sg13g2_fill_2 FILLER_38_329 ();
 sg13g2_fill_1 FILLER_38_331 ();
 sg13g2_fill_4 FILLER_38_340 ();
 sg13g2_fill_2 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_354 ();
 sg13g2_fill_4 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_373 ();
 sg13g2_fill_8 FILLER_38_403 ();
 sg13g2_fill_4 FILLER_38_411 ();
 sg13g2_fill_1 FILLER_38_428 ();
 sg13g2_fill_1 FILLER_38_443 ();
 sg13g2_fill_8 FILLER_38_475 ();
 sg13g2_fill_4 FILLER_38_483 ();
 sg13g2_fill_8 FILLER_38_495 ();
 sg13g2_fill_2 FILLER_38_503 ();
 sg13g2_fill_1 FILLER_38_505 ();
 sg13g2_fill_2 FILLER_38_527 ();
 sg13g2_fill_2 FILLER_38_542 ();
 sg13g2_fill_1 FILLER_38_544 ();
 sg13g2_fill_8 FILLER_38_551 ();
 sg13g2_fill_1 FILLER_38_559 ();
 sg13g2_fill_1 FILLER_38_593 ();
 sg13g2_fill_2 FILLER_38_616 ();
 sg13g2_fill_1 FILLER_38_626 ();
 sg13g2_fill_2 FILLER_38_650 ();
 sg13g2_fill_4 FILLER_38_660 ();
 sg13g2_fill_2 FILLER_38_664 ();
 sg13g2_fill_4 FILLER_38_723 ();
 sg13g2_fill_1 FILLER_38_727 ();
 sg13g2_fill_8 FILLER_38_732 ();
 sg13g2_fill_2 FILLER_38_740 ();
 sg13g2_fill_8 FILLER_38_746 ();
 sg13g2_fill_8 FILLER_38_754 ();
 sg13g2_fill_4 FILLER_38_762 ();
 sg13g2_fill_4 FILLER_38_771 ();
 sg13g2_fill_1 FILLER_38_775 ();
 sg13g2_fill_8 FILLER_38_780 ();
 sg13g2_fill_8 FILLER_38_788 ();
 sg13g2_fill_2 FILLER_38_796 ();
 sg13g2_fill_1 FILLER_38_798 ();
 sg13g2_fill_8 FILLER_38_834 ();
 sg13g2_fill_2 FILLER_38_842 ();
 sg13g2_fill_1 FILLER_38_844 ();
 sg13g2_fill_2 FILLER_38_869 ();
 sg13g2_fill_4 FILLER_38_907 ();
 sg13g2_fill_2 FILLER_38_911 ();
 sg13g2_fill_2 FILLER_38_935 ();
 sg13g2_fill_1 FILLER_38_937 ();
 sg13g2_fill_8 FILLER_38_950 ();
 sg13g2_fill_8 FILLER_38_958 ();
 sg13g2_fill_8 FILLER_38_966 ();
 sg13g2_fill_8 FILLER_38_974 ();
 sg13g2_fill_8 FILLER_38_982 ();
 sg13g2_fill_8 FILLER_38_990 ();
 sg13g2_fill_8 FILLER_38_998 ();
 sg13g2_fill_8 FILLER_38_1006 ();
 sg13g2_fill_8 FILLER_38_1014 ();
 sg13g2_fill_8 FILLER_38_1022 ();
 sg13g2_fill_8 FILLER_38_1030 ();
 sg13g2_fill_8 FILLER_38_1038 ();
 sg13g2_fill_8 FILLER_38_1046 ();
 sg13g2_fill_8 FILLER_38_1054 ();
 sg13g2_fill_8 FILLER_38_1062 ();
 sg13g2_fill_8 FILLER_38_1070 ();
 sg13g2_fill_8 FILLER_38_1078 ();
 sg13g2_fill_8 FILLER_38_1086 ();
 sg13g2_fill_8 FILLER_38_1094 ();
 sg13g2_fill_8 FILLER_38_1102 ();
 sg13g2_fill_8 FILLER_38_1110 ();
 sg13g2_fill_8 FILLER_38_1118 ();
 sg13g2_fill_8 FILLER_38_1126 ();
 sg13g2_fill_8 FILLER_38_1134 ();
 sg13g2_fill_8 FILLER_38_1142 ();
 sg13g2_fill_8 FILLER_38_1150 ();
 sg13g2_fill_8 FILLER_38_1158 ();
 sg13g2_fill_8 FILLER_39_0 ();
 sg13g2_fill_8 FILLER_39_8 ();
 sg13g2_fill_2 FILLER_39_16 ();
 sg13g2_fill_1 FILLER_39_18 ();
 sg13g2_fill_4 FILLER_39_22 ();
 sg13g2_fill_1 FILLER_39_26 ();
 sg13g2_fill_8 FILLER_39_35 ();
 sg13g2_fill_2 FILLER_39_43 ();
 sg13g2_fill_1 FILLER_39_45 ();
 sg13g2_fill_1 FILLER_39_51 ();
 sg13g2_fill_8 FILLER_39_104 ();
 sg13g2_fill_8 FILLER_39_112 ();
 sg13g2_fill_8 FILLER_39_120 ();
 sg13g2_fill_8 FILLER_39_128 ();
 sg13g2_fill_8 FILLER_39_136 ();
 sg13g2_fill_8 FILLER_39_144 ();
 sg13g2_fill_8 FILLER_39_152 ();
 sg13g2_fill_8 FILLER_39_160 ();
 sg13g2_fill_8 FILLER_39_168 ();
 sg13g2_fill_4 FILLER_39_176 ();
 sg13g2_fill_2 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_182 ();
 sg13g2_fill_4 FILLER_39_188 ();
 sg13g2_fill_2 FILLER_39_192 ();
 sg13g2_fill_1 FILLER_39_194 ();
 sg13g2_fill_4 FILLER_39_220 ();
 sg13g2_fill_1 FILLER_39_224 ();
 sg13g2_fill_8 FILLER_39_259 ();
 sg13g2_fill_2 FILLER_39_286 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_8 FILLER_39_323 ();
 sg13g2_fill_8 FILLER_39_331 ();
 sg13g2_fill_2 FILLER_39_370 ();
 sg13g2_fill_1 FILLER_39_372 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_fill_2 FILLER_39_389 ();
 sg13g2_fill_2 FILLER_39_396 ();
 sg13g2_fill_4 FILLER_39_403 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_39_414 ();
 sg13g2_fill_1 FILLER_39_416 ();
 sg13g2_fill_1 FILLER_39_422 ();
 sg13g2_fill_8 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_440 ();
 sg13g2_fill_1 FILLER_39_442 ();
 sg13g2_fill_8 FILLER_39_453 ();
 sg13g2_fill_8 FILLER_39_461 ();
 sg13g2_fill_4 FILLER_39_469 ();
 sg13g2_fill_2 FILLER_39_473 ();
 sg13g2_fill_8 FILLER_39_503 ();
 sg13g2_fill_1 FILLER_39_511 ();
 sg13g2_fill_8 FILLER_39_519 ();
 sg13g2_fill_8 FILLER_39_527 ();
 sg13g2_fill_4 FILLER_39_545 ();
 sg13g2_fill_2 FILLER_39_549 ();
 sg13g2_fill_1 FILLER_39_551 ();
 sg13g2_fill_2 FILLER_39_557 ();
 sg13g2_fill_4 FILLER_39_565 ();
 sg13g2_fill_2 FILLER_39_582 ();
 sg13g2_fill_1 FILLER_39_584 ();
 sg13g2_fill_4 FILLER_39_590 ();
 sg13g2_fill_1 FILLER_39_594 ();
 sg13g2_fill_2 FILLER_39_599 ();
 sg13g2_fill_1 FILLER_39_601 ();
 sg13g2_fill_2 FILLER_39_610 ();
 sg13g2_fill_1 FILLER_39_612 ();
 sg13g2_fill_4 FILLER_39_617 ();
 sg13g2_fill_2 FILLER_39_626 ();
 sg13g2_fill_8 FILLER_39_650 ();
 sg13g2_fill_2 FILLER_39_658 ();
 sg13g2_fill_1 FILLER_39_660 ();
 sg13g2_fill_8 FILLER_39_665 ();
 sg13g2_fill_4 FILLER_39_673 ();
 sg13g2_fill_2 FILLER_39_677 ();
 sg13g2_fill_1 FILLER_39_679 ();
 sg13g2_fill_2 FILLER_39_683 ();
 sg13g2_fill_1 FILLER_39_685 ();
 sg13g2_fill_2 FILLER_39_719 ();
 sg13g2_fill_1 FILLER_39_721 ();
 sg13g2_fill_2 FILLER_39_732 ();
 sg13g2_fill_1 FILLER_39_734 ();
 sg13g2_fill_2 FILLER_39_761 ();
 sg13g2_fill_8 FILLER_39_794 ();
 sg13g2_fill_4 FILLER_39_802 ();
 sg13g2_fill_2 FILLER_39_806 ();
 sg13g2_fill_8 FILLER_39_837 ();
 sg13g2_fill_2 FILLER_39_845 ();
 sg13g2_fill_1 FILLER_39_847 ();
 sg13g2_fill_2 FILLER_39_868 ();
 sg13g2_fill_2 FILLER_39_891 ();
 sg13g2_fill_2 FILLER_39_899 ();
 sg13g2_fill_4 FILLER_39_922 ();
 sg13g2_fill_8 FILLER_39_953 ();
 sg13g2_fill_8 FILLER_39_961 ();
 sg13g2_fill_8 FILLER_39_969 ();
 sg13g2_fill_8 FILLER_39_977 ();
 sg13g2_fill_8 FILLER_39_985 ();
 sg13g2_fill_8 FILLER_39_993 ();
 sg13g2_fill_8 FILLER_39_1001 ();
 sg13g2_fill_8 FILLER_39_1009 ();
 sg13g2_fill_8 FILLER_39_1017 ();
 sg13g2_fill_8 FILLER_39_1025 ();
 sg13g2_fill_8 FILLER_39_1033 ();
 sg13g2_fill_8 FILLER_39_1041 ();
 sg13g2_fill_8 FILLER_39_1049 ();
 sg13g2_fill_8 FILLER_39_1057 ();
 sg13g2_fill_8 FILLER_39_1065 ();
 sg13g2_fill_8 FILLER_39_1073 ();
 sg13g2_fill_8 FILLER_39_1081 ();
 sg13g2_fill_8 FILLER_39_1089 ();
 sg13g2_fill_8 FILLER_39_1097 ();
 sg13g2_fill_8 FILLER_39_1105 ();
 sg13g2_fill_8 FILLER_39_1113 ();
 sg13g2_fill_8 FILLER_39_1121 ();
 sg13g2_fill_8 FILLER_39_1129 ();
 sg13g2_fill_8 FILLER_39_1137 ();
 sg13g2_fill_8 FILLER_39_1145 ();
 sg13g2_fill_8 FILLER_39_1153 ();
 sg13g2_fill_4 FILLER_39_1161 ();
 sg13g2_fill_1 FILLER_39_1165 ();
 sg13g2_fill_8 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_8 ();
 sg13g2_fill_1 FILLER_40_61 ();
 sg13g2_fill_8 FILLER_40_108 ();
 sg13g2_fill_8 FILLER_40_116 ();
 sg13g2_fill_2 FILLER_40_124 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_fill_8 FILLER_40_140 ();
 sg13g2_fill_8 FILLER_40_148 ();
 sg13g2_fill_4 FILLER_40_156 ();
 sg13g2_fill_2 FILLER_40_160 ();
 sg13g2_fill_1 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_194 ();
 sg13g2_fill_2 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_214 ();
 sg13g2_fill_8 FILLER_40_220 ();
 sg13g2_fill_2 FILLER_40_228 ();
 sg13g2_fill_4 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_239 ();
 sg13g2_fill_8 FILLER_40_245 ();
 sg13g2_fill_4 FILLER_40_253 ();
 sg13g2_fill_2 FILLER_40_257 ();
 sg13g2_fill_1 FILLER_40_259 ();
 sg13g2_fill_2 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_fill_4 FILLER_40_303 ();
 sg13g2_fill_1 FILLER_40_307 ();
 sg13g2_fill_4 FILLER_40_313 ();
 sg13g2_fill_4 FILLER_40_325 ();
 sg13g2_fill_4 FILLER_40_363 ();
 sg13g2_fill_1 FILLER_40_367 ();
 sg13g2_fill_2 FILLER_40_373 ();
 sg13g2_fill_1 FILLER_40_375 ();
 sg13g2_fill_8 FILLER_40_420 ();
 sg13g2_fill_4 FILLER_40_428 ();
 sg13g2_fill_2 FILLER_40_432 ();
 sg13g2_fill_1 FILLER_40_434 ();
 sg13g2_fill_4 FILLER_40_444 ();
 sg13g2_fill_2 FILLER_40_474 ();
 sg13g2_fill_8 FILLER_40_510 ();
 sg13g2_fill_4 FILLER_40_518 ();
 sg13g2_fill_2 FILLER_40_522 ();
 sg13g2_fill_1 FILLER_40_524 ();
 sg13g2_fill_1 FILLER_40_548 ();
 sg13g2_fill_1 FILLER_40_560 ();
 sg13g2_fill_4 FILLER_40_570 ();
 sg13g2_fill_8 FILLER_40_589 ();
 sg13g2_fill_4 FILLER_40_597 ();
 sg13g2_fill_2 FILLER_40_601 ();
 sg13g2_fill_1 FILLER_40_603 ();
 sg13g2_fill_8 FILLER_40_610 ();
 sg13g2_fill_8 FILLER_40_618 ();
 sg13g2_fill_4 FILLER_40_631 ();
 sg13g2_fill_2 FILLER_40_635 ();
 sg13g2_fill_4 FILLER_40_646 ();
 sg13g2_fill_1 FILLER_40_650 ();
 sg13g2_fill_1 FILLER_40_656 ();
 sg13g2_fill_8 FILLER_40_662 ();
 sg13g2_fill_1 FILLER_40_686 ();
 sg13g2_fill_1 FILLER_40_717 ();
 sg13g2_fill_2 FILLER_40_728 ();
 sg13g2_fill_1 FILLER_40_735 ();
 sg13g2_fill_8 FILLER_40_792 ();
 sg13g2_fill_4 FILLER_40_800 ();
 sg13g2_fill_8 FILLER_40_833 ();
 sg13g2_fill_2 FILLER_40_841 ();
 sg13g2_fill_1 FILLER_40_843 ();
 sg13g2_fill_2 FILLER_40_861 ();
 sg13g2_fill_1 FILLER_40_863 ();
 sg13g2_fill_8 FILLER_40_887 ();
 sg13g2_fill_4 FILLER_40_895 ();
 sg13g2_fill_1 FILLER_40_899 ();
 sg13g2_fill_2 FILLER_40_905 ();
 sg13g2_fill_4 FILLER_40_917 ();
 sg13g2_fill_2 FILLER_40_921 ();
 sg13g2_fill_1 FILLER_40_923 ();
 sg13g2_fill_8 FILLER_40_944 ();
 sg13g2_fill_8 FILLER_40_952 ();
 sg13g2_fill_8 FILLER_40_960 ();
 sg13g2_fill_8 FILLER_40_968 ();
 sg13g2_fill_8 FILLER_40_976 ();
 sg13g2_fill_8 FILLER_40_984 ();
 sg13g2_fill_8 FILLER_40_992 ();
 sg13g2_fill_8 FILLER_40_1000 ();
 sg13g2_fill_8 FILLER_40_1008 ();
 sg13g2_fill_8 FILLER_40_1016 ();
 sg13g2_fill_8 FILLER_40_1024 ();
 sg13g2_fill_8 FILLER_40_1032 ();
 sg13g2_fill_8 FILLER_40_1040 ();
 sg13g2_fill_8 FILLER_40_1048 ();
 sg13g2_fill_8 FILLER_40_1056 ();
 sg13g2_fill_8 FILLER_40_1064 ();
 sg13g2_fill_8 FILLER_40_1072 ();
 sg13g2_fill_8 FILLER_40_1080 ();
 sg13g2_fill_8 FILLER_40_1088 ();
 sg13g2_fill_8 FILLER_40_1096 ();
 sg13g2_fill_8 FILLER_40_1104 ();
 sg13g2_fill_8 FILLER_40_1112 ();
 sg13g2_fill_8 FILLER_40_1120 ();
 sg13g2_fill_8 FILLER_40_1128 ();
 sg13g2_fill_8 FILLER_40_1136 ();
 sg13g2_fill_8 FILLER_40_1144 ();
 sg13g2_fill_8 FILLER_40_1152 ();
 sg13g2_fill_4 FILLER_40_1160 ();
 sg13g2_fill_2 FILLER_40_1164 ();
 sg13g2_fill_8 FILLER_41_39 ();
 sg13g2_fill_8 FILLER_41_47 ();
 sg13g2_fill_4 FILLER_41_55 ();
 sg13g2_fill_2 FILLER_41_59 ();
 sg13g2_fill_1 FILLER_41_66 ();
 sg13g2_fill_1 FILLER_41_88 ();
 sg13g2_fill_2 FILLER_41_120 ();
 sg13g2_fill_1 FILLER_41_161 ();
 sg13g2_fill_4 FILLER_41_208 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_fill_2 FILLER_41_229 ();
 sg13g2_fill_1 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_242 ();
 sg13g2_fill_8 FILLER_41_252 ();
 sg13g2_fill_8 FILLER_41_260 ();
 sg13g2_fill_2 FILLER_41_268 ();
 sg13g2_fill_8 FILLER_41_290 ();
 sg13g2_fill_8 FILLER_41_298 ();
 sg13g2_fill_1 FILLER_41_337 ();
 sg13g2_fill_8 FILLER_41_343 ();
 sg13g2_fill_8 FILLER_41_351 ();
 sg13g2_fill_8 FILLER_41_359 ();
 sg13g2_fill_8 FILLER_41_367 ();
 sg13g2_fill_8 FILLER_41_375 ();
 sg13g2_fill_1 FILLER_41_383 ();
 sg13g2_fill_2 FILLER_41_398 ();
 sg13g2_fill_8 FILLER_41_405 ();
 sg13g2_fill_8 FILLER_41_413 ();
 sg13g2_fill_4 FILLER_41_421 ();
 sg13g2_fill_1 FILLER_41_425 ();
 sg13g2_fill_4 FILLER_41_434 ();
 sg13g2_fill_4 FILLER_41_474 ();
 sg13g2_fill_1 FILLER_41_483 ();
 sg13g2_fill_8 FILLER_41_489 ();
 sg13g2_fill_1 FILLER_41_497 ();
 sg13g2_fill_4 FILLER_41_503 ();
 sg13g2_fill_1 FILLER_41_513 ();
 sg13g2_fill_4 FILLER_41_521 ();
 sg13g2_fill_1 FILLER_41_529 ();
 sg13g2_fill_1 FILLER_41_567 ();
 sg13g2_fill_4 FILLER_41_581 ();
 sg13g2_fill_2 FILLER_41_589 ();
 sg13g2_fill_8 FILLER_41_596 ();
 sg13g2_fill_1 FILLER_41_604 ();
 sg13g2_fill_8 FILLER_41_611 ();
 sg13g2_fill_2 FILLER_41_619 ();
 sg13g2_fill_4 FILLER_41_625 ();
 sg13g2_fill_1 FILLER_41_629 ();
 sg13g2_fill_2 FILLER_41_635 ();
 sg13g2_fill_2 FILLER_41_645 ();
 sg13g2_fill_1 FILLER_41_647 ();
 sg13g2_fill_8 FILLER_41_671 ();
 sg13g2_fill_2 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_684 ();
 sg13g2_fill_8 FILLER_41_693 ();
 sg13g2_fill_8 FILLER_41_701 ();
 sg13g2_fill_2 FILLER_41_709 ();
 sg13g2_fill_1 FILLER_41_711 ();
 sg13g2_fill_4 FILLER_41_715 ();
 sg13g2_fill_1 FILLER_41_719 ();
 sg13g2_fill_2 FILLER_41_751 ();
 sg13g2_fill_4 FILLER_41_788 ();
 sg13g2_fill_1 FILLER_41_792 ();
 sg13g2_fill_8 FILLER_41_797 ();
 sg13g2_fill_8 FILLER_41_810 ();
 sg13g2_fill_1 FILLER_41_818 ();
 sg13g2_fill_8 FILLER_41_823 ();
 sg13g2_fill_8 FILLER_41_831 ();
 sg13g2_fill_1 FILLER_41_839 ();
 sg13g2_fill_8 FILLER_41_859 ();
 sg13g2_fill_2 FILLER_41_867 ();
 sg13g2_fill_1 FILLER_41_869 ();
 sg13g2_fill_8 FILLER_41_873 ();
 sg13g2_fill_8 FILLER_41_885 ();
 sg13g2_fill_8 FILLER_41_893 ();
 sg13g2_fill_8 FILLER_41_901 ();
 sg13g2_fill_4 FILLER_41_909 ();
 sg13g2_fill_2 FILLER_41_913 ();
 sg13g2_fill_4 FILLER_41_919 ();
 sg13g2_fill_1 FILLER_41_923 ();
 sg13g2_fill_8 FILLER_41_945 ();
 sg13g2_fill_8 FILLER_41_953 ();
 sg13g2_fill_8 FILLER_41_961 ();
 sg13g2_fill_8 FILLER_41_969 ();
 sg13g2_fill_8 FILLER_41_977 ();
 sg13g2_fill_8 FILLER_41_985 ();
 sg13g2_fill_8 FILLER_41_993 ();
 sg13g2_fill_8 FILLER_41_1001 ();
 sg13g2_fill_8 FILLER_41_1009 ();
 sg13g2_fill_8 FILLER_41_1017 ();
 sg13g2_fill_8 FILLER_41_1025 ();
 sg13g2_fill_8 FILLER_41_1033 ();
 sg13g2_fill_8 FILLER_41_1041 ();
 sg13g2_fill_8 FILLER_41_1049 ();
 sg13g2_fill_8 FILLER_41_1057 ();
 sg13g2_fill_8 FILLER_41_1065 ();
 sg13g2_fill_8 FILLER_41_1073 ();
 sg13g2_fill_8 FILLER_41_1081 ();
 sg13g2_fill_8 FILLER_41_1089 ();
 sg13g2_fill_8 FILLER_41_1097 ();
 sg13g2_fill_8 FILLER_41_1105 ();
 sg13g2_fill_8 FILLER_41_1113 ();
 sg13g2_fill_8 FILLER_41_1121 ();
 sg13g2_fill_8 FILLER_41_1129 ();
 sg13g2_fill_8 FILLER_41_1137 ();
 sg13g2_fill_8 FILLER_41_1145 ();
 sg13g2_fill_8 FILLER_41_1153 ();
 sg13g2_fill_4 FILLER_41_1161 ();
 sg13g2_fill_1 FILLER_41_1165 ();
 sg13g2_fill_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_8 ();
 sg13g2_fill_8 FILLER_42_28 ();
 sg13g2_fill_8 FILLER_42_36 ();
 sg13g2_fill_4 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_48 ();
 sg13g2_fill_1 FILLER_42_50 ();
 sg13g2_fill_8 FILLER_42_77 ();
 sg13g2_fill_8 FILLER_42_85 ();
 sg13g2_fill_4 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_97 ();
 sg13g2_fill_4 FILLER_42_117 ();
 sg13g2_fill_8 FILLER_42_147 ();
 sg13g2_fill_8 FILLER_42_155 ();
 sg13g2_fill_8 FILLER_42_163 ();
 sg13g2_fill_4 FILLER_42_171 ();
 sg13g2_fill_2 FILLER_42_175 ();
 sg13g2_fill_1 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_198 ();
 sg13g2_fill_2 FILLER_42_210 ();
 sg13g2_fill_1 FILLER_42_212 ();
 sg13g2_fill_8 FILLER_42_218 ();
 sg13g2_fill_8 FILLER_42_226 ();
 sg13g2_fill_8 FILLER_42_234 ();
 sg13g2_fill_4 FILLER_42_255 ();
 sg13g2_fill_2 FILLER_42_259 ();
 sg13g2_fill_8 FILLER_42_266 ();
 sg13g2_fill_8 FILLER_42_274 ();
 sg13g2_fill_8 FILLER_42_282 ();
 sg13g2_fill_8 FILLER_42_290 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_1 FILLER_42_300 ();
 sg13g2_fill_2 FILLER_42_331 ();
 sg13g2_fill_1 FILLER_42_333 ();
 sg13g2_fill_2 FILLER_42_347 ();
 sg13g2_fill_2 FILLER_42_359 ();
 sg13g2_fill_2 FILLER_42_366 ();
 sg13g2_fill_1 FILLER_42_368 ();
 sg13g2_fill_8 FILLER_42_374 ();
 sg13g2_fill_4 FILLER_42_382 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_fill_8 FILLER_42_404 ();
 sg13g2_fill_4 FILLER_42_412 ();
 sg13g2_fill_2 FILLER_42_416 ();
 sg13g2_fill_1 FILLER_42_418 ();
 sg13g2_fill_2 FILLER_42_432 ();
 sg13g2_fill_1 FILLER_42_434 ();
 sg13g2_fill_2 FILLER_42_450 ();
 sg13g2_fill_8 FILLER_42_477 ();
 sg13g2_fill_2 FILLER_42_485 ();
 sg13g2_fill_1 FILLER_42_487 ();
 sg13g2_fill_2 FILLER_42_493 ();
 sg13g2_fill_1 FILLER_42_502 ();
 sg13g2_fill_2 FILLER_42_509 ();
 sg13g2_fill_2 FILLER_42_520 ();
 sg13g2_fill_1 FILLER_42_530 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_600 ();
 sg13g2_fill_1 FILLER_42_606 ();
 sg13g2_fill_1 FILLER_42_615 ();
 sg13g2_fill_4 FILLER_42_631 ();
 sg13g2_fill_2 FILLER_42_645 ();
 sg13g2_fill_8 FILLER_42_652 ();
 sg13g2_fill_8 FILLER_42_668 ();
 sg13g2_fill_8 FILLER_42_676 ();
 sg13g2_fill_8 FILLER_42_684 ();
 sg13g2_fill_8 FILLER_42_692 ();
 sg13g2_fill_8 FILLER_42_700 ();
 sg13g2_fill_4 FILLER_42_708 ();
 sg13g2_fill_8 FILLER_42_742 ();
 sg13g2_fill_1 FILLER_42_750 ();
 sg13g2_fill_8 FILLER_42_755 ();
 sg13g2_fill_8 FILLER_42_763 ();
 sg13g2_fill_1 FILLER_42_771 ();
 sg13g2_fill_8 FILLER_42_780 ();
 sg13g2_fill_8 FILLER_42_788 ();
 sg13g2_fill_1 FILLER_42_796 ();
 sg13g2_fill_8 FILLER_42_802 ();
 sg13g2_fill_8 FILLER_42_810 ();
 sg13g2_fill_8 FILLER_42_818 ();
 sg13g2_fill_8 FILLER_42_826 ();
 sg13g2_fill_4 FILLER_42_834 ();
 sg13g2_fill_1 FILLER_42_843 ();
 sg13g2_fill_8 FILLER_42_857 ();
 sg13g2_fill_8 FILLER_42_865 ();
 sg13g2_fill_4 FILLER_42_873 ();
 sg13g2_fill_1 FILLER_42_877 ();
 sg13g2_fill_4 FILLER_42_900 ();
 sg13g2_fill_2 FILLER_42_904 ();
 sg13g2_fill_1 FILLER_42_918 ();
 sg13g2_fill_2 FILLER_42_925 ();
 sg13g2_fill_1 FILLER_42_927 ();
 sg13g2_fill_8 FILLER_42_952 ();
 sg13g2_fill_8 FILLER_42_960 ();
 sg13g2_fill_8 FILLER_42_968 ();
 sg13g2_fill_8 FILLER_42_976 ();
 sg13g2_fill_8 FILLER_42_984 ();
 sg13g2_fill_8 FILLER_42_992 ();
 sg13g2_fill_8 FILLER_42_1000 ();
 sg13g2_fill_8 FILLER_42_1008 ();
 sg13g2_fill_8 FILLER_42_1016 ();
 sg13g2_fill_8 FILLER_42_1024 ();
 sg13g2_fill_8 FILLER_42_1032 ();
 sg13g2_fill_8 FILLER_42_1040 ();
 sg13g2_fill_8 FILLER_42_1048 ();
 sg13g2_fill_8 FILLER_42_1056 ();
 sg13g2_fill_8 FILLER_42_1064 ();
 sg13g2_fill_8 FILLER_42_1072 ();
 sg13g2_fill_8 FILLER_42_1080 ();
 sg13g2_fill_8 FILLER_42_1088 ();
 sg13g2_fill_8 FILLER_42_1096 ();
 sg13g2_fill_8 FILLER_42_1104 ();
 sg13g2_fill_8 FILLER_42_1112 ();
 sg13g2_fill_8 FILLER_42_1120 ();
 sg13g2_fill_8 FILLER_42_1128 ();
 sg13g2_fill_8 FILLER_42_1136 ();
 sg13g2_fill_8 FILLER_42_1144 ();
 sg13g2_fill_8 FILLER_42_1152 ();
 sg13g2_fill_4 FILLER_42_1160 ();
 sg13g2_fill_2 FILLER_42_1164 ();
 sg13g2_fill_4 FILLER_43_0 ();
 sg13g2_fill_2 FILLER_43_4 ();
 sg13g2_fill_1 FILLER_43_6 ();
 sg13g2_fill_2 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_fill_8 FILLER_43_69 ();
 sg13g2_fill_8 FILLER_43_77 ();
 sg13g2_fill_8 FILLER_43_85 ();
 sg13g2_fill_4 FILLER_43_93 ();
 sg13g2_fill_2 FILLER_43_97 ();
 sg13g2_fill_8 FILLER_43_104 ();
 sg13g2_fill_8 FILLER_43_112 ();
 sg13g2_fill_4 FILLER_43_120 ();
 sg13g2_fill_8 FILLER_43_137 ();
 sg13g2_fill_8 FILLER_43_145 ();
 sg13g2_fill_8 FILLER_43_153 ();
 sg13g2_fill_8 FILLER_43_161 ();
 sg13g2_fill_8 FILLER_43_169 ();
 sg13g2_fill_2 FILLER_43_177 ();
 sg13g2_fill_8 FILLER_43_187 ();
 sg13g2_fill_2 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_207 ();
 sg13g2_fill_8 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_4 FILLER_43_235 ();
 sg13g2_fill_2 FILLER_43_239 ();
 sg13g2_fill_1 FILLER_43_241 ();
 sg13g2_fill_4 FILLER_43_252 ();
 sg13g2_fill_1 FILLER_43_264 ();
 sg13g2_fill_8 FILLER_43_275 ();
 sg13g2_fill_2 FILLER_43_283 ();
 sg13g2_fill_1 FILLER_43_285 ();
 sg13g2_fill_2 FILLER_43_326 ();
 sg13g2_fill_1 FILLER_43_328 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_fill_4 FILLER_43_369 ();
 sg13g2_fill_1 FILLER_43_386 ();
 sg13g2_fill_8 FILLER_43_413 ();
 sg13g2_fill_1 FILLER_43_421 ();
 sg13g2_fill_2 FILLER_43_427 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_fill_1 FILLER_43_440 ();
 sg13g2_fill_2 FILLER_43_449 ();
 sg13g2_fill_1 FILLER_43_451 ();
 sg13g2_fill_8 FILLER_43_461 ();
 sg13g2_fill_4 FILLER_43_469 ();
 sg13g2_fill_1 FILLER_43_473 ();
 sg13g2_fill_2 FILLER_43_489 ();
 sg13g2_fill_1 FILLER_43_522 ();
 sg13g2_fill_1 FILLER_43_527 ();
 sg13g2_fill_1 FILLER_43_539 ();
 sg13g2_fill_1 FILLER_43_544 ();
 sg13g2_fill_2 FILLER_43_559 ();
 sg13g2_fill_1 FILLER_43_566 ();
 sg13g2_fill_1 FILLER_43_608 ();
 sg13g2_fill_2 FILLER_43_632 ();
 sg13g2_fill_1 FILLER_43_634 ();
 sg13g2_fill_1 FILLER_43_641 ();
 sg13g2_fill_1 FILLER_43_647 ();
 sg13g2_fill_4 FILLER_43_667 ();
 sg13g2_fill_1 FILLER_43_671 ();
 sg13g2_fill_4 FILLER_43_681 ();
 sg13g2_fill_1 FILLER_43_685 ();
 sg13g2_fill_2 FILLER_43_689 ();
 sg13g2_fill_4 FILLER_43_699 ();
 sg13g2_fill_1 FILLER_43_703 ();
 sg13g2_fill_8 FILLER_43_715 ();
 sg13g2_fill_4 FILLER_43_723 ();
 sg13g2_fill_2 FILLER_43_727 ();
 sg13g2_fill_1 FILLER_43_734 ();
 sg13g2_fill_8 FILLER_43_739 ();
 sg13g2_fill_8 FILLER_43_747 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_fill_1 FILLER_43_757 ();
 sg13g2_fill_2 FILLER_43_824 ();
 sg13g2_fill_8 FILLER_43_834 ();
 sg13g2_fill_4 FILLER_43_842 ();
 sg13g2_fill_4 FILLER_43_852 ();
 sg13g2_fill_2 FILLER_43_856 ();
 sg13g2_fill_4 FILLER_43_863 ();
 sg13g2_fill_1 FILLER_43_904 ();
 sg13g2_fill_2 FILLER_43_911 ();
 sg13g2_fill_1 FILLER_43_938 ();
 sg13g2_fill_8 FILLER_43_948 ();
 sg13g2_fill_8 FILLER_43_956 ();
 sg13g2_fill_8 FILLER_43_964 ();
 sg13g2_fill_8 FILLER_43_972 ();
 sg13g2_fill_8 FILLER_43_980 ();
 sg13g2_fill_8 FILLER_43_988 ();
 sg13g2_fill_8 FILLER_43_996 ();
 sg13g2_fill_8 FILLER_43_1004 ();
 sg13g2_fill_8 FILLER_43_1012 ();
 sg13g2_fill_8 FILLER_43_1020 ();
 sg13g2_fill_8 FILLER_43_1028 ();
 sg13g2_fill_8 FILLER_43_1036 ();
 sg13g2_fill_8 FILLER_43_1044 ();
 sg13g2_fill_8 FILLER_43_1052 ();
 sg13g2_fill_8 FILLER_43_1060 ();
 sg13g2_fill_8 FILLER_43_1068 ();
 sg13g2_fill_8 FILLER_43_1076 ();
 sg13g2_fill_8 FILLER_43_1084 ();
 sg13g2_fill_8 FILLER_43_1092 ();
 sg13g2_fill_8 FILLER_43_1100 ();
 sg13g2_fill_8 FILLER_43_1108 ();
 sg13g2_fill_8 FILLER_43_1116 ();
 sg13g2_fill_8 FILLER_43_1124 ();
 sg13g2_fill_8 FILLER_43_1132 ();
 sg13g2_fill_8 FILLER_43_1140 ();
 sg13g2_fill_8 FILLER_43_1148 ();
 sg13g2_fill_8 FILLER_43_1156 ();
 sg13g2_fill_2 FILLER_43_1164 ();
 sg13g2_fill_8 FILLER_44_0 ();
 sg13g2_fill_4 FILLER_44_8 ();
 sg13g2_fill_1 FILLER_44_12 ();
 sg13g2_fill_8 FILLER_44_21 ();
 sg13g2_fill_4 FILLER_44_29 ();
 sg13g2_fill_8 FILLER_44_36 ();
 sg13g2_fill_4 FILLER_44_44 ();
 sg13g2_fill_2 FILLER_44_48 ();
 sg13g2_fill_1 FILLER_44_50 ();
 sg13g2_fill_8 FILLER_44_72 ();
 sg13g2_fill_4 FILLER_44_80 ();
 sg13g2_fill_8 FILLER_44_109 ();
 sg13g2_fill_8 FILLER_44_117 ();
 sg13g2_fill_4 FILLER_44_125 ();
 sg13g2_fill_2 FILLER_44_129 ();
 sg13g2_fill_2 FILLER_44_135 ();
 sg13g2_fill_1 FILLER_44_137 ();
 sg13g2_fill_8 FILLER_44_190 ();
 sg13g2_fill_2 FILLER_44_198 ();
 sg13g2_fill_1 FILLER_44_200 ();
 sg13g2_fill_8 FILLER_44_212 ();
 sg13g2_fill_4 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_237 ();
 sg13g2_fill_4 FILLER_44_249 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_fill_2 FILLER_44_298 ();
 sg13g2_fill_1 FILLER_44_300 ();
 sg13g2_fill_1 FILLER_44_319 ();
 sg13g2_fill_8 FILLER_44_325 ();
 sg13g2_fill_8 FILLER_44_343 ();
 sg13g2_fill_2 FILLER_44_351 ();
 sg13g2_fill_8 FILLER_44_358 ();
 sg13g2_fill_4 FILLER_44_366 ();
 sg13g2_fill_8 FILLER_44_401 ();
 sg13g2_fill_8 FILLER_44_409 ();
 sg13g2_fill_8 FILLER_44_417 ();
 sg13g2_fill_1 FILLER_44_425 ();
 sg13g2_fill_4 FILLER_44_455 ();
 sg13g2_fill_2 FILLER_44_459 ();
 sg13g2_fill_1 FILLER_44_461 ();
 sg13g2_fill_4 FILLER_44_468 ();
 sg13g2_fill_2 FILLER_44_481 ();
 sg13g2_fill_4 FILLER_44_533 ();
 sg13g2_fill_4 FILLER_44_540 ();
 sg13g2_fill_2 FILLER_44_548 ();
 sg13g2_fill_1 FILLER_44_550 ();
 sg13g2_fill_4 FILLER_44_555 ();
 sg13g2_fill_2 FILLER_44_559 ();
 sg13g2_fill_8 FILLER_44_566 ();
 sg13g2_fill_2 FILLER_44_574 ();
 sg13g2_fill_1 FILLER_44_581 ();
 sg13g2_fill_8 FILLER_44_601 ();
 sg13g2_fill_4 FILLER_44_609 ();
 sg13g2_fill_2 FILLER_44_613 ();
 sg13g2_fill_1 FILLER_44_615 ();
 sg13g2_fill_8 FILLER_44_621 ();
 sg13g2_fill_2 FILLER_44_629 ();
 sg13g2_fill_1 FILLER_44_631 ();
 sg13g2_fill_2 FILLER_44_671 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_fill_4 FILLER_44_726 ();
 sg13g2_fill_4 FILLER_44_756 ();
 sg13g2_fill_1 FILLER_44_760 ();
 sg13g2_fill_8 FILLER_44_799 ();
 sg13g2_fill_4 FILLER_44_807 ();
 sg13g2_fill_1 FILLER_44_811 ();
 sg13g2_fill_4 FILLER_44_833 ();
 sg13g2_fill_2 FILLER_44_847 ();
 sg13g2_fill_1 FILLER_44_849 ();
 sg13g2_fill_4 FILLER_44_871 ();
 sg13g2_fill_1 FILLER_44_880 ();
 sg13g2_fill_1 FILLER_44_896 ();
 sg13g2_fill_2 FILLER_44_906 ();
 sg13g2_fill_8 FILLER_44_912 ();
 sg13g2_fill_1 FILLER_44_920 ();
 sg13g2_fill_8 FILLER_44_950 ();
 sg13g2_fill_8 FILLER_44_958 ();
 sg13g2_fill_8 FILLER_44_966 ();
 sg13g2_fill_8 FILLER_44_974 ();
 sg13g2_fill_8 FILLER_44_982 ();
 sg13g2_fill_8 FILLER_44_990 ();
 sg13g2_fill_8 FILLER_44_998 ();
 sg13g2_fill_8 FILLER_44_1006 ();
 sg13g2_fill_8 FILLER_44_1014 ();
 sg13g2_fill_8 FILLER_44_1022 ();
 sg13g2_fill_8 FILLER_44_1030 ();
 sg13g2_fill_8 FILLER_44_1038 ();
 sg13g2_fill_8 FILLER_44_1046 ();
 sg13g2_fill_8 FILLER_44_1054 ();
 sg13g2_fill_8 FILLER_44_1062 ();
 sg13g2_fill_8 FILLER_44_1070 ();
 sg13g2_fill_8 FILLER_44_1078 ();
 sg13g2_fill_8 FILLER_44_1086 ();
 sg13g2_fill_8 FILLER_44_1094 ();
 sg13g2_fill_8 FILLER_44_1102 ();
 sg13g2_fill_8 FILLER_44_1110 ();
 sg13g2_fill_8 FILLER_44_1118 ();
 sg13g2_fill_8 FILLER_44_1126 ();
 sg13g2_fill_8 FILLER_44_1134 ();
 sg13g2_fill_8 FILLER_44_1142 ();
 sg13g2_fill_8 FILLER_44_1150 ();
 sg13g2_fill_8 FILLER_44_1158 ();
 sg13g2_fill_1 FILLER_45_51 ();
 sg13g2_fill_8 FILLER_45_78 ();
 sg13g2_fill_8 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_120 ();
 sg13g2_fill_4 FILLER_45_173 ();
 sg13g2_fill_2 FILLER_45_177 ();
 sg13g2_fill_1 FILLER_45_179 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_fill_2 FILLER_45_195 ();
 sg13g2_fill_1 FILLER_45_197 ();
 sg13g2_fill_1 FILLER_45_221 ();
 sg13g2_fill_4 FILLER_45_258 ();
 sg13g2_fill_4 FILLER_45_271 ();
 sg13g2_fill_1 FILLER_45_275 ();
 sg13g2_fill_1 FILLER_45_301 ();
 sg13g2_fill_4 FILLER_45_307 ();
 sg13g2_fill_1 FILLER_45_311 ();
 sg13g2_fill_8 FILLER_45_321 ();
 sg13g2_fill_2 FILLER_45_329 ();
 sg13g2_fill_1 FILLER_45_331 ();
 sg13g2_fill_4 FILLER_45_340 ();
 sg13g2_fill_8 FILLER_45_352 ();
 sg13g2_fill_4 FILLER_45_360 ();
 sg13g2_fill_2 FILLER_45_364 ();
 sg13g2_fill_8 FILLER_45_381 ();
 sg13g2_fill_4 FILLER_45_389 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_fill_8 FILLER_45_403 ();
 sg13g2_fill_4 FILLER_45_411 ();
 sg13g2_fill_1 FILLER_45_415 ();
 sg13g2_fill_1 FILLER_45_441 ();
 sg13g2_fill_1 FILLER_45_452 ();
 sg13g2_fill_1 FILLER_45_479 ();
 sg13g2_fill_2 FILLER_45_500 ();
 sg13g2_fill_1 FILLER_45_502 ();
 sg13g2_fill_2 FILLER_45_527 ();
 sg13g2_fill_8 FILLER_45_537 ();
 sg13g2_fill_4 FILLER_45_545 ();
 sg13g2_fill_2 FILLER_45_549 ();
 sg13g2_fill_2 FILLER_45_555 ();
 sg13g2_fill_1 FILLER_45_557 ();
 sg13g2_fill_8 FILLER_45_571 ();
 sg13g2_fill_4 FILLER_45_579 ();
 sg13g2_fill_2 FILLER_45_583 ();
 sg13g2_fill_8 FILLER_45_595 ();
 sg13g2_fill_4 FILLER_45_603 ();
 sg13g2_fill_2 FILLER_45_607 ();
 sg13g2_fill_1 FILLER_45_609 ();
 sg13g2_fill_4 FILLER_45_616 ();
 sg13g2_fill_2 FILLER_45_620 ();
 sg13g2_fill_1 FILLER_45_622 ();
 sg13g2_fill_4 FILLER_45_639 ();
 sg13g2_fill_2 FILLER_45_643 ();
 sg13g2_fill_4 FILLER_45_669 ();
 sg13g2_fill_8 FILLER_45_677 ();
 sg13g2_fill_2 FILLER_45_685 ();
 sg13g2_fill_2 FILLER_45_693 ();
 sg13g2_fill_1 FILLER_45_695 ();
 sg13g2_fill_2 FILLER_45_722 ();
 sg13g2_fill_2 FILLER_45_766 ();
 sg13g2_fill_1 FILLER_45_768 ();
 sg13g2_fill_4 FILLER_45_773 ();
 sg13g2_fill_1 FILLER_45_777 ();
 sg13g2_fill_1 FILLER_45_791 ();
 sg13g2_fill_8 FILLER_45_827 ();
 sg13g2_fill_2 FILLER_45_835 ();
 sg13g2_fill_1 FILLER_45_837 ();
 sg13g2_fill_2 FILLER_45_843 ();
 sg13g2_fill_4 FILLER_45_855 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_8 FILLER_45_866 ();
 sg13g2_fill_2 FILLER_45_874 ();
 sg13g2_fill_2 FILLER_45_887 ();
 sg13g2_fill_1 FILLER_45_889 ();
 sg13g2_fill_2 FILLER_45_895 ();
 sg13g2_fill_8 FILLER_45_902 ();
 sg13g2_fill_4 FILLER_45_910 ();
 sg13g2_fill_2 FILLER_45_914 ();
 sg13g2_fill_1 FILLER_45_916 ();
 sg13g2_fill_8 FILLER_45_946 ();
 sg13g2_fill_8 FILLER_45_954 ();
 sg13g2_fill_8 FILLER_45_962 ();
 sg13g2_fill_8 FILLER_45_970 ();
 sg13g2_fill_8 FILLER_45_978 ();
 sg13g2_fill_8 FILLER_45_986 ();
 sg13g2_fill_8 FILLER_45_994 ();
 sg13g2_fill_8 FILLER_45_1002 ();
 sg13g2_fill_8 FILLER_45_1010 ();
 sg13g2_fill_8 FILLER_45_1018 ();
 sg13g2_fill_8 FILLER_45_1026 ();
 sg13g2_fill_8 FILLER_45_1034 ();
 sg13g2_fill_8 FILLER_45_1042 ();
 sg13g2_fill_8 FILLER_45_1050 ();
 sg13g2_fill_8 FILLER_45_1058 ();
 sg13g2_fill_8 FILLER_45_1066 ();
 sg13g2_fill_8 FILLER_45_1074 ();
 sg13g2_fill_8 FILLER_45_1082 ();
 sg13g2_fill_8 FILLER_45_1090 ();
 sg13g2_fill_8 FILLER_45_1098 ();
 sg13g2_fill_8 FILLER_45_1106 ();
 sg13g2_fill_8 FILLER_45_1114 ();
 sg13g2_fill_8 FILLER_45_1122 ();
 sg13g2_fill_8 FILLER_45_1130 ();
 sg13g2_fill_8 FILLER_45_1138 ();
 sg13g2_fill_8 FILLER_45_1146 ();
 sg13g2_fill_8 FILLER_45_1154 ();
 sg13g2_fill_4 FILLER_45_1162 ();
 sg13g2_fill_8 FILLER_46_0 ();
 sg13g2_fill_8 FILLER_46_8 ();
 sg13g2_fill_2 FILLER_46_16 ();
 sg13g2_fill_8 FILLER_46_44 ();
 sg13g2_fill_4 FILLER_46_52 ();
 sg13g2_fill_2 FILLER_46_98 ();
 sg13g2_fill_8 FILLER_46_108 ();
 sg13g2_fill_8 FILLER_46_116 ();
 sg13g2_fill_4 FILLER_46_124 ();
 sg13g2_fill_1 FILLER_46_128 ();
 sg13g2_fill_2 FILLER_46_134 ();
 sg13g2_fill_2 FILLER_46_202 ();
 sg13g2_fill_8 FILLER_46_209 ();
 sg13g2_fill_4 FILLER_46_217 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_fill_2 FILLER_46_226 ();
 sg13g2_fill_2 FILLER_46_233 ();
 sg13g2_fill_8 FILLER_46_249 ();
 sg13g2_fill_8 FILLER_46_257 ();
 sg13g2_fill_8 FILLER_46_265 ();
 sg13g2_fill_4 FILLER_46_273 ();
 sg13g2_fill_2 FILLER_46_285 ();
 sg13g2_fill_8 FILLER_46_323 ();
 sg13g2_fill_4 FILLER_46_331 ();
 sg13g2_fill_2 FILLER_46_335 ();
 sg13g2_fill_8 FILLER_46_365 ();
 sg13g2_fill_2 FILLER_46_378 ();
 sg13g2_fill_4 FILLER_46_389 ();
 sg13g2_fill_2 FILLER_46_393 ();
 sg13g2_fill_2 FILLER_46_421 ();
 sg13g2_fill_1 FILLER_46_423 ();
 sg13g2_fill_4 FILLER_46_490 ();
 sg13g2_fill_8 FILLER_46_534 ();
 sg13g2_fill_8 FILLER_46_542 ();
 sg13g2_fill_2 FILLER_46_550 ();
 sg13g2_fill_1 FILLER_46_552 ();
 sg13g2_fill_8 FILLER_46_568 ();
 sg13g2_fill_2 FILLER_46_576 ();
 sg13g2_fill_8 FILLER_46_592 ();
 sg13g2_fill_1 FILLER_46_614 ();
 sg13g2_fill_8 FILLER_46_620 ();
 sg13g2_fill_4 FILLER_46_628 ();
 sg13g2_fill_2 FILLER_46_632 ();
 sg13g2_fill_2 FILLER_46_639 ();
 sg13g2_fill_1 FILLER_46_641 ();
 sg13g2_fill_4 FILLER_46_648 ();
 sg13g2_fill_1 FILLER_46_652 ();
 sg13g2_fill_2 FILLER_46_656 ();
 sg13g2_fill_1 FILLER_46_658 ();
 sg13g2_fill_8 FILLER_46_663 ();
 sg13g2_fill_8 FILLER_46_671 ();
 sg13g2_fill_8 FILLER_46_679 ();
 sg13g2_fill_8 FILLER_46_687 ();
 sg13g2_fill_1 FILLER_46_695 ();
 sg13g2_fill_4 FILLER_46_701 ();
 sg13g2_fill_2 FILLER_46_705 ();
 sg13g2_fill_1 FILLER_46_707 ();
 sg13g2_fill_8 FILLER_46_712 ();
 sg13g2_fill_2 FILLER_46_720 ();
 sg13g2_fill_1 FILLER_46_732 ();
 sg13g2_fill_8 FILLER_46_758 ();
 sg13g2_fill_8 FILLER_46_770 ();
 sg13g2_fill_2 FILLER_46_778 ();
 sg13g2_fill_8 FILLER_46_810 ();
 sg13g2_fill_8 FILLER_46_818 ();
 sg13g2_fill_4 FILLER_46_826 ();
 sg13g2_fill_2 FILLER_46_830 ();
 sg13g2_fill_1 FILLER_46_840 ();
 sg13g2_fill_4 FILLER_46_856 ();
 sg13g2_fill_8 FILLER_46_865 ();
 sg13g2_fill_8 FILLER_46_873 ();
 sg13g2_fill_1 FILLER_46_881 ();
 sg13g2_fill_2 FILLER_46_891 ();
 sg13g2_fill_1 FILLER_46_893 ();
 sg13g2_fill_2 FILLER_46_913 ();
 sg13g2_fill_1 FILLER_46_929 ();
 sg13g2_fill_8 FILLER_46_950 ();
 sg13g2_fill_8 FILLER_46_958 ();
 sg13g2_fill_8 FILLER_46_966 ();
 sg13g2_fill_8 FILLER_46_974 ();
 sg13g2_fill_8 FILLER_46_982 ();
 sg13g2_fill_8 FILLER_46_990 ();
 sg13g2_fill_8 FILLER_46_998 ();
 sg13g2_fill_8 FILLER_46_1006 ();
 sg13g2_fill_8 FILLER_46_1014 ();
 sg13g2_fill_8 FILLER_46_1022 ();
 sg13g2_fill_8 FILLER_46_1030 ();
 sg13g2_fill_8 FILLER_46_1038 ();
 sg13g2_fill_8 FILLER_46_1046 ();
 sg13g2_fill_8 FILLER_46_1054 ();
 sg13g2_fill_8 FILLER_46_1062 ();
 sg13g2_fill_8 FILLER_46_1070 ();
 sg13g2_fill_8 FILLER_46_1078 ();
 sg13g2_fill_8 FILLER_46_1086 ();
 sg13g2_fill_8 FILLER_46_1094 ();
 sg13g2_fill_8 FILLER_46_1102 ();
 sg13g2_fill_8 FILLER_46_1110 ();
 sg13g2_fill_8 FILLER_46_1118 ();
 sg13g2_fill_8 FILLER_46_1126 ();
 sg13g2_fill_8 FILLER_46_1134 ();
 sg13g2_fill_8 FILLER_46_1142 ();
 sg13g2_fill_8 FILLER_46_1150 ();
 sg13g2_fill_8 FILLER_46_1158 ();
 sg13g2_fill_8 FILLER_47_0 ();
 sg13g2_fill_8 FILLER_47_8 ();
 sg13g2_fill_8 FILLER_47_16 ();
 sg13g2_fill_2 FILLER_47_24 ();
 sg13g2_fill_8 FILLER_47_36 ();
 sg13g2_fill_8 FILLER_47_44 ();
 sg13g2_fill_8 FILLER_47_52 ();
 sg13g2_fill_8 FILLER_47_60 ();
 sg13g2_fill_8 FILLER_47_68 ();
 sg13g2_fill_2 FILLER_47_76 ();
 sg13g2_fill_4 FILLER_47_99 ();
 sg13g2_fill_1 FILLER_47_103 ();
 sg13g2_fill_4 FILLER_47_114 ();
 sg13g2_fill_8 FILLER_47_144 ();
 sg13g2_fill_8 FILLER_47_152 ();
 sg13g2_fill_4 FILLER_47_160 ();
 sg13g2_fill_4 FILLER_47_190 ();
 sg13g2_fill_2 FILLER_47_194 ();
 sg13g2_fill_2 FILLER_47_211 ();
 sg13g2_fill_2 FILLER_47_223 ();
 sg13g2_fill_1 FILLER_47_225 ();
 sg13g2_fill_8 FILLER_47_236 ();
 sg13g2_fill_8 FILLER_47_244 ();
 sg13g2_fill_2 FILLER_47_252 ();
 sg13g2_fill_1 FILLER_47_254 ();
 sg13g2_fill_8 FILLER_47_286 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_fill_8 FILLER_47_300 ();
 sg13g2_fill_4 FILLER_47_308 ();
 sg13g2_fill_4 FILLER_47_325 ();
 sg13g2_fill_1 FILLER_47_329 ();
 sg13g2_fill_1 FILLER_47_340 ();
 sg13g2_fill_4 FILLER_47_367 ();
 sg13g2_fill_8 FILLER_47_411 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_fill_1 FILLER_47_421 ();
 sg13g2_fill_2 FILLER_47_427 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_fill_2 FILLER_47_435 ();
 sg13g2_fill_4 FILLER_47_442 ();
 sg13g2_fill_2 FILLER_47_446 ();
 sg13g2_fill_8 FILLER_47_457 ();
 sg13g2_fill_8 FILLER_47_465 ();
 sg13g2_fill_8 FILLER_47_473 ();
 sg13g2_fill_8 FILLER_47_481 ();
 sg13g2_fill_4 FILLER_47_533 ();
 sg13g2_fill_2 FILLER_47_537 ();
 sg13g2_fill_2 FILLER_47_547 ();
 sg13g2_fill_1 FILLER_47_549 ();
 sg13g2_fill_4 FILLER_47_572 ();
 sg13g2_fill_2 FILLER_47_576 ();
 sg13g2_fill_2 FILLER_47_583 ();
 sg13g2_fill_8 FILLER_47_595 ();
 sg13g2_fill_4 FILLER_47_603 ();
 sg13g2_fill_2 FILLER_47_607 ();
 sg13g2_fill_4 FILLER_47_629 ();
 sg13g2_fill_2 FILLER_47_633 ();
 sg13g2_fill_1 FILLER_47_635 ();
 sg13g2_fill_8 FILLER_47_652 ();
 sg13g2_fill_8 FILLER_47_660 ();
 sg13g2_fill_8 FILLER_47_668 ();
 sg13g2_fill_2 FILLER_47_676 ();
 sg13g2_fill_8 FILLER_47_681 ();
 sg13g2_fill_2 FILLER_47_689 ();
 sg13g2_fill_8 FILLER_47_700 ();
 sg13g2_fill_4 FILLER_47_708 ();
 sg13g2_fill_1 FILLER_47_712 ();
 sg13g2_fill_8 FILLER_47_723 ();
 sg13g2_fill_2 FILLER_47_731 ();
 sg13g2_fill_1 FILLER_47_733 ();
 sg13g2_fill_8 FILLER_47_741 ();
 sg13g2_fill_1 FILLER_47_754 ();
 sg13g2_fill_8 FILLER_47_784 ();
 sg13g2_fill_8 FILLER_47_792 ();
 sg13g2_fill_8 FILLER_47_800 ();
 sg13g2_fill_8 FILLER_47_808 ();
 sg13g2_fill_8 FILLER_47_816 ();
 sg13g2_fill_8 FILLER_47_824 ();
 sg13g2_fill_8 FILLER_47_832 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_fill_1 FILLER_47_872 ();
 sg13g2_fill_2 FILLER_47_878 ();
 sg13g2_fill_2 FILLER_47_920 ();
 sg13g2_fill_2 FILLER_47_927 ();
 sg13g2_fill_8 FILLER_47_952 ();
 sg13g2_fill_8 FILLER_47_960 ();
 sg13g2_fill_8 FILLER_47_968 ();
 sg13g2_fill_8 FILLER_47_976 ();
 sg13g2_fill_8 FILLER_47_984 ();
 sg13g2_fill_8 FILLER_47_992 ();
 sg13g2_fill_8 FILLER_47_1000 ();
 sg13g2_fill_8 FILLER_47_1008 ();
 sg13g2_fill_8 FILLER_47_1016 ();
 sg13g2_fill_8 FILLER_47_1024 ();
 sg13g2_fill_8 FILLER_47_1032 ();
 sg13g2_fill_8 FILLER_47_1040 ();
 sg13g2_fill_8 FILLER_47_1048 ();
 sg13g2_fill_8 FILLER_47_1056 ();
 sg13g2_fill_8 FILLER_47_1064 ();
 sg13g2_fill_8 FILLER_47_1072 ();
 sg13g2_fill_8 FILLER_47_1080 ();
 sg13g2_fill_8 FILLER_47_1088 ();
 sg13g2_fill_8 FILLER_47_1096 ();
 sg13g2_fill_8 FILLER_47_1104 ();
 sg13g2_fill_8 FILLER_47_1112 ();
 sg13g2_fill_8 FILLER_47_1120 ();
 sg13g2_fill_8 FILLER_47_1128 ();
 sg13g2_fill_8 FILLER_47_1136 ();
 sg13g2_fill_8 FILLER_47_1144 ();
 sg13g2_fill_8 FILLER_47_1152 ();
 sg13g2_fill_4 FILLER_47_1160 ();
 sg13g2_fill_2 FILLER_47_1164 ();
 sg13g2_fill_1 FILLER_48_29 ();
 sg13g2_fill_4 FILLER_48_36 ();
 sg13g2_fill_2 FILLER_48_40 ();
 sg13g2_fill_1 FILLER_48_42 ();
 sg13g2_fill_4 FILLER_48_90 ();
 sg13g2_fill_1 FILLER_48_94 ();
 sg13g2_fill_1 FILLER_48_100 ();
 sg13g2_fill_8 FILLER_48_109 ();
 sg13g2_fill_8 FILLER_48_117 ();
 sg13g2_fill_4 FILLER_48_125 ();
 sg13g2_fill_1 FILLER_48_129 ();
 sg13g2_fill_8 FILLER_48_159 ();
 sg13g2_fill_8 FILLER_48_167 ();
 sg13g2_fill_8 FILLER_48_175 ();
 sg13g2_fill_8 FILLER_48_183 ();
 sg13g2_fill_8 FILLER_48_191 ();
 sg13g2_fill_2 FILLER_48_199 ();
 sg13g2_fill_2 FILLER_48_247 ();
 sg13g2_fill_1 FILLER_48_249 ();
 sg13g2_fill_2 FILLER_48_263 ();
 sg13g2_fill_4 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_4 FILLER_48_284 ();
 sg13g2_fill_4 FILLER_48_298 ();
 sg13g2_fill_1 FILLER_48_302 ();
 sg13g2_fill_8 FILLER_48_313 ();
 sg13g2_fill_4 FILLER_48_321 ();
 sg13g2_fill_2 FILLER_48_325 ();
 sg13g2_fill_2 FILLER_48_338 ();
 sg13g2_fill_8 FILLER_48_344 ();
 sg13g2_fill_8 FILLER_48_352 ();
 sg13g2_fill_8 FILLER_48_360 ();
 sg13g2_fill_2 FILLER_48_368 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_4 FILLER_48_386 ();
 sg13g2_fill_2 FILLER_48_390 ();
 sg13g2_fill_1 FILLER_48_397 ();
 sg13g2_fill_8 FILLER_48_413 ();
 sg13g2_fill_8 FILLER_48_421 ();
 sg13g2_fill_8 FILLER_48_429 ();
 sg13g2_fill_4 FILLER_48_437 ();
 sg13g2_fill_1 FILLER_48_441 ();
 sg13g2_fill_2 FILLER_48_450 ();
 sg13g2_fill_1 FILLER_48_452 ();
 sg13g2_fill_8 FILLER_48_458 ();
 sg13g2_fill_8 FILLER_48_466 ();
 sg13g2_fill_4 FILLER_48_474 ();
 sg13g2_fill_2 FILLER_48_478 ();
 sg13g2_fill_1 FILLER_48_480 ();
 sg13g2_fill_8 FILLER_48_485 ();
 sg13g2_fill_2 FILLER_48_493 ();
 sg13g2_fill_2 FILLER_48_509 ();
 sg13g2_fill_1 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_550 ();
 sg13g2_fill_1 FILLER_48_556 ();
 sg13g2_fill_4 FILLER_48_561 ();
 sg13g2_fill_1 FILLER_48_565 ();
 sg13g2_fill_2 FILLER_48_596 ();
 sg13g2_fill_1 FILLER_48_598 ();
 sg13g2_fill_4 FILLER_48_610 ();
 sg13g2_fill_2 FILLER_48_619 ();
 sg13g2_fill_1 FILLER_48_626 ();
 sg13g2_fill_1 FILLER_48_632 ();
 sg13g2_fill_2 FILLER_48_654 ();
 sg13g2_fill_1 FILLER_48_656 ();
 sg13g2_fill_2 FILLER_48_663 ();
 sg13g2_fill_8 FILLER_48_755 ();
 sg13g2_fill_8 FILLER_48_763 ();
 sg13g2_fill_8 FILLER_48_771 ();
 sg13g2_fill_2 FILLER_48_779 ();
 sg13g2_fill_1 FILLER_48_781 ();
 sg13g2_fill_4 FILLER_48_812 ();
 sg13g2_fill_8 FILLER_48_829 ();
 sg13g2_fill_8 FILLER_48_837 ();
 sg13g2_fill_1 FILLER_48_845 ();
 sg13g2_fill_2 FILLER_48_850 ();
 sg13g2_fill_1 FILLER_48_852 ();
 sg13g2_fill_1 FILLER_48_863 ();
 sg13g2_fill_2 FILLER_48_869 ();
 sg13g2_fill_1 FILLER_48_871 ();
 sg13g2_fill_4 FILLER_48_877 ();
 sg13g2_fill_4 FILLER_48_895 ();
 sg13g2_fill_2 FILLER_48_924 ();
 sg13g2_fill_8 FILLER_48_947 ();
 sg13g2_fill_8 FILLER_48_955 ();
 sg13g2_fill_8 FILLER_48_963 ();
 sg13g2_fill_8 FILLER_48_971 ();
 sg13g2_fill_8 FILLER_48_979 ();
 sg13g2_fill_8 FILLER_48_987 ();
 sg13g2_fill_8 FILLER_48_995 ();
 sg13g2_fill_8 FILLER_48_1003 ();
 sg13g2_fill_8 FILLER_48_1011 ();
 sg13g2_fill_8 FILLER_48_1019 ();
 sg13g2_fill_8 FILLER_48_1027 ();
 sg13g2_fill_8 FILLER_48_1035 ();
 sg13g2_fill_8 FILLER_48_1043 ();
 sg13g2_fill_8 FILLER_48_1051 ();
 sg13g2_fill_8 FILLER_48_1059 ();
 sg13g2_fill_8 FILLER_48_1067 ();
 sg13g2_fill_8 FILLER_48_1075 ();
 sg13g2_fill_8 FILLER_48_1083 ();
 sg13g2_fill_8 FILLER_48_1091 ();
 sg13g2_fill_8 FILLER_48_1099 ();
 sg13g2_fill_8 FILLER_48_1107 ();
 sg13g2_fill_8 FILLER_48_1115 ();
 sg13g2_fill_8 FILLER_48_1123 ();
 sg13g2_fill_8 FILLER_48_1131 ();
 sg13g2_fill_8 FILLER_48_1139 ();
 sg13g2_fill_8 FILLER_48_1147 ();
 sg13g2_fill_8 FILLER_48_1155 ();
 sg13g2_fill_2 FILLER_48_1163 ();
 sg13g2_fill_1 FILLER_48_1165 ();
 sg13g2_fill_4 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_4 ();
 sg13g2_fill_4 FILLER_49_40 ();
 sg13g2_fill_8 FILLER_49_76 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_fill_8 FILLER_49_117 ();
 sg13g2_fill_8 FILLER_49_125 ();
 sg13g2_fill_4 FILLER_49_133 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_fill_8 FILLER_49_159 ();
 sg13g2_fill_4 FILLER_49_167 ();
 sg13g2_fill_2 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_198 ();
 sg13g2_fill_1 FILLER_49_200 ();
 sg13g2_fill_4 FILLER_49_266 ();
 sg13g2_fill_2 FILLER_49_270 ();
 sg13g2_fill_1 FILLER_49_272 ();
 sg13g2_fill_2 FILLER_49_295 ();
 sg13g2_fill_2 FILLER_49_313 ();
 sg13g2_fill_1 FILLER_49_315 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_8 FILLER_49_343 ();
 sg13g2_fill_8 FILLER_49_351 ();
 sg13g2_fill_1 FILLER_49_359 ();
 sg13g2_fill_4 FILLER_49_375 ();
 sg13g2_fill_4 FILLER_49_384 ();
 sg13g2_fill_1 FILLER_49_388 ();
 sg13g2_fill_2 FILLER_49_432 ();
 sg13g2_fill_1 FILLER_49_434 ();
 sg13g2_fill_8 FILLER_49_480 ();
 sg13g2_fill_4 FILLER_49_488 ();
 sg13g2_fill_1 FILLER_49_492 ();
 sg13g2_fill_2 FILLER_49_512 ();
 sg13g2_fill_8 FILLER_49_530 ();
 sg13g2_fill_4 FILLER_49_538 ();
 sg13g2_fill_2 FILLER_49_542 ();
 sg13g2_fill_8 FILLER_49_548 ();
 sg13g2_fill_4 FILLER_49_556 ();
 sg13g2_fill_8 FILLER_49_569 ();
 sg13g2_fill_2 FILLER_49_577 ();
 sg13g2_fill_1 FILLER_49_579 ();
 sg13g2_fill_2 FILLER_49_593 ();
 sg13g2_fill_1 FILLER_49_595 ();
 sg13g2_fill_2 FILLER_49_600 ();
 sg13g2_fill_1 FILLER_49_602 ();
 sg13g2_fill_4 FILLER_49_609 ();
 sg13g2_fill_2 FILLER_49_646 ();
 sg13g2_fill_1 FILLER_49_648 ();
 sg13g2_fill_8 FILLER_49_661 ();
 sg13g2_fill_8 FILLER_49_669 ();
 sg13g2_fill_4 FILLER_49_677 ();
 sg13g2_fill_8 FILLER_49_685 ();
 sg13g2_fill_8 FILLER_49_693 ();
 sg13g2_fill_8 FILLER_49_701 ();
 sg13g2_fill_4 FILLER_49_709 ();
 sg13g2_fill_2 FILLER_49_713 ();
 sg13g2_fill_1 FILLER_49_715 ();
 sg13g2_fill_2 FILLER_49_726 ();
 sg13g2_fill_8 FILLER_49_799 ();
 sg13g2_fill_1 FILLER_49_807 ();
 sg13g2_fill_8 FILLER_49_832 ();
 sg13g2_fill_4 FILLER_49_845 ();
 sg13g2_fill_1 FILLER_49_849 ();
 sg13g2_fill_4 FILLER_49_857 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_8 FILLER_49_882 ();
 sg13g2_fill_4 FILLER_49_890 ();
 sg13g2_fill_8 FILLER_49_908 ();
 sg13g2_fill_4 FILLER_49_916 ();
 sg13g2_fill_1 FILLER_49_920 ();
 sg13g2_fill_8 FILLER_49_925 ();
 sg13g2_fill_1 FILLER_49_933 ();
 sg13g2_fill_8 FILLER_49_942 ();
 sg13g2_fill_8 FILLER_49_950 ();
 sg13g2_fill_8 FILLER_49_958 ();
 sg13g2_fill_8 FILLER_49_966 ();
 sg13g2_fill_8 FILLER_49_974 ();
 sg13g2_fill_8 FILLER_49_982 ();
 sg13g2_fill_8 FILLER_49_990 ();
 sg13g2_fill_8 FILLER_49_998 ();
 sg13g2_fill_8 FILLER_49_1006 ();
 sg13g2_fill_8 FILLER_49_1014 ();
 sg13g2_fill_8 FILLER_49_1022 ();
 sg13g2_fill_8 FILLER_49_1030 ();
 sg13g2_fill_8 FILLER_49_1038 ();
 sg13g2_fill_8 FILLER_49_1046 ();
 sg13g2_fill_8 FILLER_49_1054 ();
 sg13g2_fill_8 FILLER_49_1062 ();
 sg13g2_fill_8 FILLER_49_1070 ();
 sg13g2_fill_8 FILLER_49_1078 ();
 sg13g2_fill_8 FILLER_49_1086 ();
 sg13g2_fill_8 FILLER_49_1094 ();
 sg13g2_fill_8 FILLER_49_1102 ();
 sg13g2_fill_8 FILLER_49_1110 ();
 sg13g2_fill_8 FILLER_49_1118 ();
 sg13g2_fill_8 FILLER_49_1126 ();
 sg13g2_fill_8 FILLER_49_1134 ();
 sg13g2_fill_8 FILLER_49_1142 ();
 sg13g2_fill_8 FILLER_49_1150 ();
 sg13g2_fill_8 FILLER_49_1158 ();
 sg13g2_fill_8 FILLER_50_0 ();
 sg13g2_fill_4 FILLER_50_8 ();
 sg13g2_fill_2 FILLER_50_12 ();
 sg13g2_fill_8 FILLER_50_29 ();
 sg13g2_fill_8 FILLER_50_37 ();
 sg13g2_fill_1 FILLER_50_45 ();
 sg13g2_fill_8 FILLER_50_66 ();
 sg13g2_fill_2 FILLER_50_74 ();
 sg13g2_fill_1 FILLER_50_76 ();
 sg13g2_fill_8 FILLER_50_136 ();
 sg13g2_fill_8 FILLER_50_165 ();
 sg13g2_fill_8 FILLER_50_173 ();
 sg13g2_fill_8 FILLER_50_181 ();
 sg13g2_fill_2 FILLER_50_189 ();
 sg13g2_fill_1 FILLER_50_191 ();
 sg13g2_fill_8 FILLER_50_197 ();
 sg13g2_fill_4 FILLER_50_205 ();
 sg13g2_fill_1 FILLER_50_209 ();
 sg13g2_fill_2 FILLER_50_215 ();
 sg13g2_fill_4 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_232 ();
 sg13g2_fill_1 FILLER_50_234 ();
 sg13g2_fill_4 FILLER_50_244 ();
 sg13g2_fill_2 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_250 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_fill_4 FILLER_50_266 ();
 sg13g2_fill_1 FILLER_50_270 ();
 sg13g2_fill_2 FILLER_50_289 ();
 sg13g2_fill_1 FILLER_50_291 ();
 sg13g2_fill_4 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_326 ();
 sg13g2_fill_4 FILLER_50_332 ();
 sg13g2_fill_2 FILLER_50_336 ();
 sg13g2_fill_1 FILLER_50_338 ();
 sg13g2_fill_2 FILLER_50_344 ();
 sg13g2_fill_4 FILLER_50_351 ();
 sg13g2_fill_1 FILLER_50_355 ();
 sg13g2_fill_2 FILLER_50_369 ();
 sg13g2_fill_1 FILLER_50_371 ();
 sg13g2_fill_1 FILLER_50_377 ();
 sg13g2_fill_8 FILLER_50_388 ();
 sg13g2_fill_4 FILLER_50_402 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_4 FILLER_50_452 ();
 sg13g2_fill_2 FILLER_50_456 ();
 sg13g2_fill_1 FILLER_50_458 ();
 sg13g2_fill_8 FILLER_50_465 ();
 sg13g2_fill_4 FILLER_50_473 ();
 sg13g2_fill_1 FILLER_50_477 ();
 sg13g2_fill_2 FILLER_50_504 ();
 sg13g2_fill_1 FILLER_50_506 ();
 sg13g2_fill_8 FILLER_50_522 ();
 sg13g2_fill_4 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_534 ();
 sg13g2_fill_8 FILLER_50_560 ();
 sg13g2_fill_4 FILLER_50_568 ();
 sg13g2_fill_4 FILLER_50_577 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_fill_2 FILLER_50_588 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_8 FILLER_50_603 ();
 sg13g2_fill_2 FILLER_50_611 ();
 sg13g2_fill_4 FILLER_50_633 ();
 sg13g2_fill_2 FILLER_50_647 ();
 sg13g2_fill_8 FILLER_50_654 ();
 sg13g2_fill_8 FILLER_50_662 ();
 sg13g2_fill_8 FILLER_50_670 ();
 sg13g2_fill_2 FILLER_50_678 ();
 sg13g2_fill_1 FILLER_50_680 ();
 sg13g2_fill_4 FILLER_50_690 ();
 sg13g2_fill_1 FILLER_50_694 ();
 sg13g2_fill_4 FILLER_50_713 ();
 sg13g2_fill_2 FILLER_50_717 ();
 sg13g2_fill_2 FILLER_50_749 ();
 sg13g2_fill_4 FILLER_50_756 ();
 sg13g2_fill_1 FILLER_50_760 ();
 sg13g2_fill_8 FILLER_50_800 ();
 sg13g2_fill_2 FILLER_50_808 ();
 sg13g2_fill_1 FILLER_50_810 ();
 sg13g2_fill_1 FILLER_50_816 ();
 sg13g2_fill_4 FILLER_50_833 ();
 sg13g2_fill_1 FILLER_50_837 ();
 sg13g2_fill_8 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_864 ();
 sg13g2_fill_1 FILLER_50_866 ();
 sg13g2_fill_4 FILLER_50_902 ();
 sg13g2_fill_2 FILLER_50_906 ();
 sg13g2_fill_1 FILLER_50_908 ();
 sg13g2_fill_8 FILLER_50_914 ();
 sg13g2_fill_4 FILLER_50_922 ();
 sg13g2_fill_2 FILLER_50_926 ();
 sg13g2_fill_1 FILLER_50_928 ();
 sg13g2_fill_8 FILLER_50_934 ();
 sg13g2_fill_8 FILLER_50_942 ();
 sg13g2_fill_8 FILLER_50_950 ();
 sg13g2_fill_8 FILLER_50_958 ();
 sg13g2_fill_8 FILLER_50_966 ();
 sg13g2_fill_8 FILLER_50_974 ();
 sg13g2_fill_8 FILLER_50_982 ();
 sg13g2_fill_8 FILLER_50_990 ();
 sg13g2_fill_8 FILLER_50_998 ();
 sg13g2_fill_8 FILLER_50_1006 ();
 sg13g2_fill_8 FILLER_50_1014 ();
 sg13g2_fill_8 FILLER_50_1022 ();
 sg13g2_fill_8 FILLER_50_1030 ();
 sg13g2_fill_8 FILLER_50_1038 ();
 sg13g2_fill_8 FILLER_50_1046 ();
 sg13g2_fill_8 FILLER_50_1054 ();
 sg13g2_fill_8 FILLER_50_1062 ();
 sg13g2_fill_8 FILLER_50_1070 ();
 sg13g2_fill_8 FILLER_50_1078 ();
 sg13g2_fill_8 FILLER_50_1086 ();
 sg13g2_fill_8 FILLER_50_1094 ();
 sg13g2_fill_8 FILLER_50_1102 ();
 sg13g2_fill_8 FILLER_50_1110 ();
 sg13g2_fill_8 FILLER_50_1118 ();
 sg13g2_fill_8 FILLER_50_1126 ();
 sg13g2_fill_8 FILLER_50_1134 ();
 sg13g2_fill_8 FILLER_50_1142 ();
 sg13g2_fill_8 FILLER_50_1150 ();
 sg13g2_fill_8 FILLER_50_1158 ();
 sg13g2_fill_8 FILLER_51_0 ();
 sg13g2_fill_4 FILLER_51_8 ();
 sg13g2_fill_2 FILLER_51_12 ();
 sg13g2_fill_4 FILLER_51_19 ();
 sg13g2_fill_2 FILLER_51_23 ();
 sg13g2_fill_8 FILLER_51_29 ();
 sg13g2_fill_8 FILLER_51_37 ();
 sg13g2_fill_2 FILLER_51_45 ();
 sg13g2_fill_1 FILLER_51_47 ();
 sg13g2_fill_2 FILLER_51_52 ();
 sg13g2_fill_8 FILLER_51_60 ();
 sg13g2_fill_8 FILLER_51_71 ();
 sg13g2_fill_8 FILLER_51_79 ();
 sg13g2_fill_1 FILLER_51_143 ();
 sg13g2_fill_4 FILLER_51_188 ();
 sg13g2_fill_2 FILLER_51_202 ();
 sg13g2_fill_2 FILLER_51_209 ();
 sg13g2_fill_8 FILLER_51_223 ();
 sg13g2_fill_4 FILLER_51_231 ();
 sg13g2_fill_2 FILLER_51_235 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_fill_2 FILLER_51_243 ();
 sg13g2_fill_1 FILLER_51_245 ();
 sg13g2_fill_1 FILLER_51_340 ();
 sg13g2_fill_2 FILLER_51_375 ();
 sg13g2_fill_4 FILLER_51_387 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_fill_1 FILLER_51_409 ();
 sg13g2_fill_2 FILLER_51_423 ();
 sg13g2_fill_8 FILLER_51_451 ();
 sg13g2_fill_8 FILLER_51_459 ();
 sg13g2_fill_8 FILLER_51_467 ();
 sg13g2_fill_1 FILLER_51_475 ();
 sg13g2_fill_2 FILLER_51_484 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_fill_8 FILLER_51_527 ();
 sg13g2_fill_2 FILLER_51_561 ();
 sg13g2_fill_1 FILLER_51_579 ();
 sg13g2_fill_8 FILLER_51_590 ();
 sg13g2_fill_8 FILLER_51_598 ();
 sg13g2_fill_1 FILLER_51_606 ();
 sg13g2_fill_8 FILLER_51_625 ();
 sg13g2_fill_8 FILLER_51_633 ();
 sg13g2_fill_8 FILLER_51_645 ();
 sg13g2_fill_8 FILLER_51_653 ();
 sg13g2_fill_4 FILLER_51_661 ();
 sg13g2_fill_2 FILLER_51_665 ();
 sg13g2_fill_1 FILLER_51_667 ();
 sg13g2_fill_4 FILLER_51_674 ();
 sg13g2_fill_4 FILLER_51_691 ();
 sg13g2_fill_1 FILLER_51_695 ();
 sg13g2_fill_8 FILLER_51_722 ();
 sg13g2_fill_8 FILLER_51_741 ();
 sg13g2_fill_4 FILLER_51_749 ();
 sg13g2_fill_8 FILLER_51_807 ();
 sg13g2_fill_4 FILLER_51_815 ();
 sg13g2_fill_2 FILLER_51_819 ();
 sg13g2_fill_1 FILLER_51_821 ();
 sg13g2_fill_8 FILLER_51_827 ();
 sg13g2_fill_8 FILLER_51_835 ();
 sg13g2_fill_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_861 ();
 sg13g2_fill_1 FILLER_51_863 ();
 sg13g2_fill_8 FILLER_51_872 ();
 sg13g2_fill_4 FILLER_51_880 ();
 sg13g2_fill_2 FILLER_51_884 ();
 sg13g2_fill_1 FILLER_51_886 ();
 sg13g2_fill_8 FILLER_51_892 ();
 sg13g2_fill_2 FILLER_51_900 ();
 sg13g2_fill_4 FILLER_51_917 ();
 sg13g2_fill_2 FILLER_51_921 ();
 sg13g2_fill_8 FILLER_51_928 ();
 sg13g2_fill_8 FILLER_51_936 ();
 sg13g2_fill_8 FILLER_51_944 ();
 sg13g2_fill_8 FILLER_51_952 ();
 sg13g2_fill_8 FILLER_51_960 ();
 sg13g2_fill_8 FILLER_51_968 ();
 sg13g2_fill_8 FILLER_51_976 ();
 sg13g2_fill_8 FILLER_51_984 ();
 sg13g2_fill_8 FILLER_51_992 ();
 sg13g2_fill_8 FILLER_51_1000 ();
 sg13g2_fill_8 FILLER_51_1008 ();
 sg13g2_fill_8 FILLER_51_1016 ();
 sg13g2_fill_8 FILLER_51_1024 ();
 sg13g2_fill_8 FILLER_51_1032 ();
 sg13g2_fill_8 FILLER_51_1040 ();
 sg13g2_fill_8 FILLER_51_1048 ();
 sg13g2_fill_8 FILLER_51_1056 ();
 sg13g2_fill_8 FILLER_51_1064 ();
 sg13g2_fill_8 FILLER_51_1072 ();
 sg13g2_fill_8 FILLER_51_1080 ();
 sg13g2_fill_8 FILLER_51_1088 ();
 sg13g2_fill_8 FILLER_51_1096 ();
 sg13g2_fill_8 FILLER_51_1104 ();
 sg13g2_fill_8 FILLER_51_1112 ();
 sg13g2_fill_8 FILLER_51_1120 ();
 sg13g2_fill_8 FILLER_51_1128 ();
 sg13g2_fill_8 FILLER_51_1136 ();
 sg13g2_fill_8 FILLER_51_1144 ();
 sg13g2_fill_8 FILLER_51_1152 ();
 sg13g2_fill_4 FILLER_51_1160 ();
 sg13g2_fill_2 FILLER_51_1164 ();
 sg13g2_fill_8 FILLER_52_0 ();
 sg13g2_fill_4 FILLER_52_8 ();
 sg13g2_fill_1 FILLER_52_12 ();
 sg13g2_fill_2 FILLER_52_22 ();
 sg13g2_fill_4 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_36 ();
 sg13g2_fill_2 FILLER_52_68 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_fill_1 FILLER_52_93 ();
 sg13g2_fill_2 FILLER_52_104 ();
 sg13g2_fill_1 FILLER_52_106 ();
 sg13g2_fill_4 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_116 ();
 sg13g2_fill_8 FILLER_52_132 ();
 sg13g2_fill_8 FILLER_52_140 ();
 sg13g2_fill_8 FILLER_52_148 ();
 sg13g2_fill_8 FILLER_52_156 ();
 sg13g2_fill_8 FILLER_52_164 ();
 sg13g2_fill_8 FILLER_52_172 ();
 sg13g2_fill_8 FILLER_52_180 ();
 sg13g2_fill_2 FILLER_52_188 ();
 sg13g2_fill_8 FILLER_52_216 ();
 sg13g2_fill_4 FILLER_52_224 ();
 sg13g2_fill_2 FILLER_52_228 ();
 sg13g2_fill_2 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_247 ();
 sg13g2_fill_8 FILLER_52_253 ();
 sg13g2_fill_8 FILLER_52_261 ();
 sg13g2_fill_8 FILLER_52_269 ();
 sg13g2_fill_8 FILLER_52_277 ();
 sg13g2_fill_2 FILLER_52_285 ();
 sg13g2_fill_8 FILLER_52_293 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_fill_1 FILLER_52_303 ();
 sg13g2_fill_4 FILLER_52_315 ();
 sg13g2_fill_1 FILLER_52_319 ();
 sg13g2_fill_8 FILLER_52_325 ();
 sg13g2_fill_4 FILLER_52_350 ();
 sg13g2_fill_2 FILLER_52_354 ();
 sg13g2_fill_8 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_422 ();
 sg13g2_fill_2 FILLER_52_427 ();
 sg13g2_fill_1 FILLER_52_442 ();
 sg13g2_fill_4 FILLER_52_486 ();
 sg13g2_fill_2 FILLER_52_490 ();
 sg13g2_fill_1 FILLER_52_492 ();
 sg13g2_fill_8 FILLER_52_534 ();
 sg13g2_fill_8 FILLER_52_599 ();
 sg13g2_fill_8 FILLER_52_607 ();
 sg13g2_fill_8 FILLER_52_615 ();
 sg13g2_fill_8 FILLER_52_623 ();
 sg13g2_fill_8 FILLER_52_631 ();
 sg13g2_fill_4 FILLER_52_639 ();
 sg13g2_fill_2 FILLER_52_643 ();
 sg13g2_fill_1 FILLER_52_645 ();
 sg13g2_fill_2 FILLER_52_672 ();
 sg13g2_fill_2 FILLER_52_700 ();
 sg13g2_fill_1 FILLER_52_727 ();
 sg13g2_fill_8 FILLER_52_769 ();
 sg13g2_fill_4 FILLER_52_777 ();
 sg13g2_fill_2 FILLER_52_781 ();
 sg13g2_fill_8 FILLER_52_821 ();
 sg13g2_fill_4 FILLER_52_829 ();
 sg13g2_fill_2 FILLER_52_833 ();
 sg13g2_fill_4 FILLER_52_839 ();
 sg13g2_fill_2 FILLER_52_843 ();
 sg13g2_fill_8 FILLER_52_873 ();
 sg13g2_fill_4 FILLER_52_881 ();
 sg13g2_fill_1 FILLER_52_885 ();
 sg13g2_fill_8 FILLER_52_911 ();
 sg13g2_fill_8 FILLER_52_919 ();
 sg13g2_fill_2 FILLER_52_927 ();
 sg13g2_fill_8 FILLER_52_948 ();
 sg13g2_fill_8 FILLER_52_956 ();
 sg13g2_fill_8 FILLER_52_964 ();
 sg13g2_fill_8 FILLER_52_972 ();
 sg13g2_fill_8 FILLER_52_980 ();
 sg13g2_fill_8 FILLER_52_988 ();
 sg13g2_fill_8 FILLER_52_996 ();
 sg13g2_fill_8 FILLER_52_1004 ();
 sg13g2_fill_8 FILLER_52_1012 ();
 sg13g2_fill_8 FILLER_52_1020 ();
 sg13g2_fill_8 FILLER_52_1028 ();
 sg13g2_fill_8 FILLER_52_1036 ();
 sg13g2_fill_8 FILLER_52_1044 ();
 sg13g2_fill_8 FILLER_52_1052 ();
 sg13g2_fill_8 FILLER_52_1060 ();
 sg13g2_fill_8 FILLER_52_1068 ();
 sg13g2_fill_8 FILLER_52_1076 ();
 sg13g2_fill_8 FILLER_52_1084 ();
 sg13g2_fill_8 FILLER_52_1092 ();
 sg13g2_fill_8 FILLER_52_1100 ();
 sg13g2_fill_8 FILLER_52_1108 ();
 sg13g2_fill_8 FILLER_52_1116 ();
 sg13g2_fill_8 FILLER_52_1124 ();
 sg13g2_fill_8 FILLER_52_1132 ();
 sg13g2_fill_8 FILLER_52_1140 ();
 sg13g2_fill_8 FILLER_52_1148 ();
 sg13g2_fill_8 FILLER_52_1156 ();
 sg13g2_fill_2 FILLER_52_1164 ();
 sg13g2_fill_8 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_8 ();
 sg13g2_fill_2 FILLER_53_41 ();
 sg13g2_fill_1 FILLER_53_43 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_fill_8 FILLER_53_92 ();
 sg13g2_fill_1 FILLER_53_105 ();
 sg13g2_fill_8 FILLER_53_109 ();
 sg13g2_fill_4 FILLER_53_117 ();
 sg13g2_fill_2 FILLER_53_121 ();
 sg13g2_fill_8 FILLER_53_140 ();
 sg13g2_fill_8 FILLER_53_148 ();
 sg13g2_fill_8 FILLER_53_156 ();
 sg13g2_fill_4 FILLER_53_164 ();
 sg13g2_fill_2 FILLER_53_168 ();
 sg13g2_fill_1 FILLER_53_170 ();
 sg13g2_fill_2 FILLER_53_202 ();
 sg13g2_fill_2 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_211 ();
 sg13g2_fill_4 FILLER_53_250 ();
 sg13g2_fill_8 FILLER_53_258 ();
 sg13g2_fill_2 FILLER_53_266 ();
 sg13g2_fill_1 FILLER_53_268 ();
 sg13g2_fill_8 FILLER_53_294 ();
 sg13g2_fill_8 FILLER_53_302 ();
 sg13g2_fill_8 FILLER_53_310 ();
 sg13g2_fill_8 FILLER_53_318 ();
 sg13g2_fill_8 FILLER_53_326 ();
 sg13g2_fill_8 FILLER_53_334 ();
 sg13g2_fill_8 FILLER_53_342 ();
 sg13g2_fill_8 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_358 ();
 sg13g2_fill_8 FILLER_53_364 ();
 sg13g2_fill_8 FILLER_53_372 ();
 sg13g2_fill_4 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_384 ();
 sg13g2_fill_8 FILLER_53_390 ();
 sg13g2_fill_8 FILLER_53_398 ();
 sg13g2_fill_8 FILLER_53_406 ();
 sg13g2_fill_4 FILLER_53_414 ();
 sg13g2_fill_2 FILLER_53_426 ();
 sg13g2_fill_2 FILLER_53_437 ();
 sg13g2_fill_1 FILLER_53_439 ();
 sg13g2_fill_4 FILLER_53_466 ();
 sg13g2_fill_2 FILLER_53_470 ();
 sg13g2_fill_8 FILLER_53_480 ();
 sg13g2_fill_8 FILLER_53_488 ();
 sg13g2_fill_2 FILLER_53_496 ();
 sg13g2_fill_1 FILLER_53_498 ();
 sg13g2_fill_2 FILLER_53_513 ();
 sg13g2_fill_1 FILLER_53_515 ();
 sg13g2_fill_4 FILLER_53_529 ();
 sg13g2_fill_2 FILLER_53_533 ();
 sg13g2_fill_4 FILLER_53_564 ();
 sg13g2_fill_2 FILLER_53_568 ();
 sg13g2_fill_1 FILLER_53_570 ();
 sg13g2_fill_4 FILLER_53_727 ();
 sg13g2_fill_8 FILLER_53_745 ();
 sg13g2_fill_4 FILLER_53_753 ();
 sg13g2_fill_2 FILLER_53_783 ();
 sg13g2_fill_1 FILLER_53_785 ();
 sg13g2_fill_2 FILLER_53_827 ();
 sg13g2_fill_1 FILLER_53_829 ();
 sg13g2_fill_8 FILLER_53_834 ();
 sg13g2_fill_4 FILLER_53_842 ();
 sg13g2_fill_1 FILLER_53_846 ();
 sg13g2_fill_8 FILLER_53_852 ();
 sg13g2_fill_8 FILLER_53_860 ();
 sg13g2_fill_8 FILLER_53_868 ();
 sg13g2_fill_4 FILLER_53_876 ();
 sg13g2_fill_2 FILLER_53_880 ();
 sg13g2_fill_4 FILLER_53_886 ();
 sg13g2_fill_2 FILLER_53_890 ();
 sg13g2_fill_1 FILLER_53_892 ();
 sg13g2_fill_2 FILLER_53_904 ();
 sg13g2_fill_8 FILLER_53_914 ();
 sg13g2_fill_8 FILLER_53_922 ();
 sg13g2_fill_8 FILLER_53_930 ();
 sg13g2_fill_8 FILLER_53_938 ();
 sg13g2_fill_8 FILLER_53_946 ();
 sg13g2_fill_8 FILLER_53_954 ();
 sg13g2_fill_8 FILLER_53_962 ();
 sg13g2_fill_8 FILLER_53_970 ();
 sg13g2_fill_8 FILLER_53_978 ();
 sg13g2_fill_8 FILLER_53_986 ();
 sg13g2_fill_8 FILLER_53_994 ();
 sg13g2_fill_8 FILLER_53_1002 ();
 sg13g2_fill_8 FILLER_53_1010 ();
 sg13g2_fill_8 FILLER_53_1018 ();
 sg13g2_fill_8 FILLER_53_1026 ();
 sg13g2_fill_8 FILLER_53_1034 ();
 sg13g2_fill_8 FILLER_53_1042 ();
 sg13g2_fill_8 FILLER_53_1050 ();
 sg13g2_fill_8 FILLER_53_1058 ();
 sg13g2_fill_8 FILLER_53_1066 ();
 sg13g2_fill_8 FILLER_53_1074 ();
 sg13g2_fill_8 FILLER_53_1082 ();
 sg13g2_fill_8 FILLER_53_1090 ();
 sg13g2_fill_8 FILLER_53_1098 ();
 sg13g2_fill_8 FILLER_53_1106 ();
 sg13g2_fill_8 FILLER_53_1114 ();
 sg13g2_fill_8 FILLER_53_1122 ();
 sg13g2_fill_8 FILLER_53_1130 ();
 sg13g2_fill_8 FILLER_53_1138 ();
 sg13g2_fill_8 FILLER_53_1146 ();
 sg13g2_fill_8 FILLER_53_1154 ();
 sg13g2_fill_4 FILLER_53_1162 ();
 sg13g2_fill_2 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_2 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_2 FILLER_54_89 ();
 sg13g2_fill_1 FILLER_54_91 ();
 sg13g2_fill_8 FILLER_54_170 ();
 sg13g2_fill_8 FILLER_54_178 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_fill_2 FILLER_54_202 ();
 sg13g2_fill_2 FILLER_54_218 ();
 sg13g2_fill_1 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_239 ();
 sg13g2_fill_2 FILLER_54_246 ();
 sg13g2_fill_8 FILLER_54_267 ();
 sg13g2_fill_8 FILLER_54_275 ();
 sg13g2_fill_2 FILLER_54_283 ();
 sg13g2_fill_1 FILLER_54_289 ();
 sg13g2_fill_8 FILLER_54_326 ();
 sg13g2_fill_4 FILLER_54_334 ();
 sg13g2_fill_4 FILLER_54_351 ();
 sg13g2_fill_1 FILLER_54_393 ();
 sg13g2_fill_1 FILLER_54_399 ();
 sg13g2_fill_2 FILLER_54_405 ();
 sg13g2_fill_1 FILLER_54_416 ();
 sg13g2_fill_8 FILLER_54_432 ();
 sg13g2_fill_4 FILLER_54_440 ();
 sg13g2_fill_2 FILLER_54_444 ();
 sg13g2_fill_1 FILLER_54_471 ();
 sg13g2_fill_2 FILLER_54_480 ();
 sg13g2_fill_8 FILLER_54_490 ();
 sg13g2_fill_8 FILLER_54_498 ();
 sg13g2_fill_8 FILLER_54_506 ();
 sg13g2_fill_8 FILLER_54_514 ();
 sg13g2_fill_8 FILLER_54_522 ();
 sg13g2_fill_8 FILLER_54_530 ();
 sg13g2_fill_4 FILLER_54_538 ();
 sg13g2_fill_8 FILLER_54_564 ();
 sg13g2_fill_8 FILLER_54_572 ();
 sg13g2_fill_8 FILLER_54_580 ();
 sg13g2_fill_1 FILLER_54_602 ();
 sg13g2_fill_2 FILLER_54_614 ();
 sg13g2_fill_1 FILLER_54_616 ();
 sg13g2_fill_4 FILLER_54_626 ();
 sg13g2_fill_2 FILLER_54_630 ();
 sg13g2_fill_1 FILLER_54_632 ();
 sg13g2_fill_2 FILLER_54_644 ();
 sg13g2_fill_1 FILLER_54_646 ();
 sg13g2_fill_4 FILLER_54_679 ();
 sg13g2_fill_2 FILLER_54_683 ();
 sg13g2_fill_4 FILLER_54_693 ();
 sg13g2_fill_1 FILLER_54_697 ();
 sg13g2_fill_2 FILLER_54_727 ();
 sg13g2_fill_4 FILLER_54_768 ();
 sg13g2_fill_8 FILLER_54_776 ();
 sg13g2_fill_8 FILLER_54_784 ();
 sg13g2_fill_8 FILLER_54_792 ();
 sg13g2_fill_8 FILLER_54_800 ();
 sg13g2_fill_4 FILLER_54_808 ();
 sg13g2_fill_8 FILLER_54_816 ();
 sg13g2_fill_8 FILLER_54_824 ();
 sg13g2_fill_4 FILLER_54_832 ();
 sg13g2_fill_8 FILLER_54_862 ();
 sg13g2_fill_8 FILLER_54_870 ();
 sg13g2_fill_8 FILLER_54_878 ();
 sg13g2_fill_8 FILLER_54_886 ();
 sg13g2_fill_8 FILLER_54_894 ();
 sg13g2_fill_8 FILLER_54_902 ();
 sg13g2_fill_8 FILLER_54_910 ();
 sg13g2_fill_8 FILLER_54_918 ();
 sg13g2_fill_8 FILLER_54_926 ();
 sg13g2_fill_8 FILLER_54_934 ();
 sg13g2_fill_8 FILLER_54_942 ();
 sg13g2_fill_8 FILLER_54_950 ();
 sg13g2_fill_8 FILLER_54_958 ();
 sg13g2_fill_8 FILLER_54_966 ();
 sg13g2_fill_8 FILLER_54_974 ();
 sg13g2_fill_8 FILLER_54_982 ();
 sg13g2_fill_8 FILLER_54_990 ();
 sg13g2_fill_8 FILLER_54_998 ();
 sg13g2_fill_8 FILLER_54_1006 ();
 sg13g2_fill_8 FILLER_54_1014 ();
 sg13g2_fill_8 FILLER_54_1022 ();
 sg13g2_fill_8 FILLER_54_1030 ();
 sg13g2_fill_8 FILLER_54_1038 ();
 sg13g2_fill_8 FILLER_54_1046 ();
 sg13g2_fill_8 FILLER_54_1054 ();
 sg13g2_fill_8 FILLER_54_1062 ();
 sg13g2_fill_8 FILLER_54_1070 ();
 sg13g2_fill_8 FILLER_54_1078 ();
 sg13g2_fill_8 FILLER_54_1086 ();
 sg13g2_fill_8 FILLER_54_1094 ();
 sg13g2_fill_8 FILLER_54_1102 ();
 sg13g2_fill_8 FILLER_54_1110 ();
 sg13g2_fill_8 FILLER_54_1118 ();
 sg13g2_fill_8 FILLER_54_1126 ();
 sg13g2_fill_8 FILLER_54_1134 ();
 sg13g2_fill_8 FILLER_54_1142 ();
 sg13g2_fill_8 FILLER_54_1150 ();
 sg13g2_fill_8 FILLER_54_1158 ();
 sg13g2_fill_8 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_8 ();
 sg13g2_fill_8 FILLER_55_42 ();
 sg13g2_fill_4 FILLER_55_50 ();
 sg13g2_fill_1 FILLER_55_54 ();
 sg13g2_fill_8 FILLER_55_106 ();
 sg13g2_fill_1 FILLER_55_114 ();
 sg13g2_fill_2 FILLER_55_159 ();
 sg13g2_fill_2 FILLER_55_195 ();
 sg13g2_fill_1 FILLER_55_197 ();
 sg13g2_fill_4 FILLER_55_215 ();
 sg13g2_fill_2 FILLER_55_219 ();
 sg13g2_fill_1 FILLER_55_236 ();
 sg13g2_fill_1 FILLER_55_252 ();
 sg13g2_fill_2 FILLER_55_261 ();
 sg13g2_fill_4 FILLER_55_273 ();
 sg13g2_fill_2 FILLER_55_277 ();
 sg13g2_fill_2 FILLER_55_311 ();
 sg13g2_fill_4 FILLER_55_323 ();
 sg13g2_fill_2 FILLER_55_327 ();
 sg13g2_fill_8 FILLER_55_355 ();
 sg13g2_fill_4 FILLER_55_363 ();
 sg13g2_fill_1 FILLER_55_367 ();
 sg13g2_fill_2 FILLER_55_403 ();
 sg13g2_fill_1 FILLER_55_405 ();
 sg13g2_fill_2 FILLER_55_414 ();
 sg13g2_fill_1 FILLER_55_416 ();
 sg13g2_fill_1 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_440 ();
 sg13g2_fill_2 FILLER_55_459 ();
 sg13g2_fill_1 FILLER_55_461 ();
 sg13g2_fill_2 FILLER_55_478 ();
 sg13g2_fill_8 FILLER_55_501 ();
 sg13g2_fill_4 FILLER_55_509 ();
 sg13g2_fill_2 FILLER_55_513 ();
 sg13g2_fill_8 FILLER_55_530 ();
 sg13g2_fill_1 FILLER_55_538 ();
 sg13g2_fill_4 FILLER_55_571 ();
 sg13g2_fill_2 FILLER_55_575 ();
 sg13g2_fill_1 FILLER_55_577 ();
 sg13g2_fill_2 FILLER_55_634 ();
 sg13g2_fill_1 FILLER_55_636 ();
 sg13g2_fill_8 FILLER_55_668 ();
 sg13g2_fill_8 FILLER_55_676 ();
 sg13g2_fill_8 FILLER_55_684 ();
 sg13g2_fill_8 FILLER_55_692 ();
 sg13g2_fill_2 FILLER_55_700 ();
 sg13g2_fill_8 FILLER_55_761 ();
 sg13g2_fill_8 FILLER_55_769 ();
 sg13g2_fill_2 FILLER_55_777 ();
 sg13g2_fill_4 FILLER_55_783 ();
 sg13g2_fill_2 FILLER_55_787 ();
 sg13g2_fill_8 FILLER_55_793 ();
 sg13g2_fill_8 FILLER_55_801 ();
 sg13g2_fill_8 FILLER_55_809 ();
 sg13g2_fill_8 FILLER_55_821 ();
 sg13g2_fill_8 FILLER_55_833 ();
 sg13g2_fill_4 FILLER_55_841 ();
 sg13g2_fill_1 FILLER_55_845 ();
 sg13g2_fill_2 FILLER_55_851 ();
 sg13g2_fill_1 FILLER_55_853 ();
 sg13g2_fill_1 FILLER_55_858 ();
 sg13g2_fill_8 FILLER_55_875 ();
 sg13g2_fill_8 FILLER_55_883 ();
 sg13g2_fill_8 FILLER_55_891 ();
 sg13g2_fill_8 FILLER_55_899 ();
 sg13g2_fill_8 FILLER_55_907 ();
 sg13g2_fill_8 FILLER_55_915 ();
 sg13g2_fill_8 FILLER_55_923 ();
 sg13g2_fill_8 FILLER_55_931 ();
 sg13g2_fill_8 FILLER_55_939 ();
 sg13g2_fill_8 FILLER_55_947 ();
 sg13g2_fill_8 FILLER_55_955 ();
 sg13g2_fill_8 FILLER_55_963 ();
 sg13g2_fill_8 FILLER_55_971 ();
 sg13g2_fill_8 FILLER_55_979 ();
 sg13g2_fill_8 FILLER_55_987 ();
 sg13g2_fill_8 FILLER_55_995 ();
 sg13g2_fill_8 FILLER_55_1003 ();
 sg13g2_fill_8 FILLER_55_1011 ();
 sg13g2_fill_8 FILLER_55_1019 ();
 sg13g2_fill_8 FILLER_55_1027 ();
 sg13g2_fill_8 FILLER_55_1035 ();
 sg13g2_fill_8 FILLER_55_1043 ();
 sg13g2_fill_8 FILLER_55_1051 ();
 sg13g2_fill_8 FILLER_55_1059 ();
 sg13g2_fill_8 FILLER_55_1067 ();
 sg13g2_fill_8 FILLER_55_1075 ();
 sg13g2_fill_8 FILLER_55_1083 ();
 sg13g2_fill_8 FILLER_55_1091 ();
 sg13g2_fill_8 FILLER_55_1099 ();
 sg13g2_fill_8 FILLER_55_1107 ();
 sg13g2_fill_8 FILLER_55_1115 ();
 sg13g2_fill_8 FILLER_55_1123 ();
 sg13g2_fill_8 FILLER_55_1131 ();
 sg13g2_fill_8 FILLER_55_1139 ();
 sg13g2_fill_8 FILLER_55_1147 ();
 sg13g2_fill_8 FILLER_55_1155 ();
 sg13g2_fill_2 FILLER_55_1163 ();
 sg13g2_fill_1 FILLER_55_1165 ();
 sg13g2_fill_8 FILLER_56_0 ();
 sg13g2_fill_8 FILLER_56_8 ();
 sg13g2_fill_4 FILLER_56_16 ();
 sg13g2_fill_2 FILLER_56_20 ();
 sg13g2_fill_1 FILLER_56_22 ();
 sg13g2_fill_4 FILLER_56_32 ();
 sg13g2_fill_2 FILLER_56_36 ();
 sg13g2_fill_1 FILLER_56_38 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_8 FILLER_56_72 ();
 sg13g2_fill_8 FILLER_56_80 ();
 sg13g2_fill_8 FILLER_56_88 ();
 sg13g2_fill_8 FILLER_56_96 ();
 sg13g2_fill_8 FILLER_56_104 ();
 sg13g2_fill_2 FILLER_56_112 ();
 sg13g2_fill_1 FILLER_56_114 ();
 sg13g2_fill_1 FILLER_56_141 ();
 sg13g2_fill_8 FILLER_56_147 ();
 sg13g2_fill_8 FILLER_56_155 ();
 sg13g2_fill_2 FILLER_56_163 ();
 sg13g2_fill_1 FILLER_56_165 ();
 sg13g2_fill_2 FILLER_56_207 ();
 sg13g2_fill_1 FILLER_56_209 ();
 sg13g2_fill_4 FILLER_56_243 ();
 sg13g2_fill_2 FILLER_56_281 ();
 sg13g2_fill_1 FILLER_56_283 ();
 sg13g2_fill_8 FILLER_56_316 ();
 sg13g2_fill_8 FILLER_56_324 ();
 sg13g2_fill_4 FILLER_56_332 ();
 sg13g2_fill_2 FILLER_56_336 ();
 sg13g2_fill_2 FILLER_56_357 ();
 sg13g2_fill_1 FILLER_56_359 ();
 sg13g2_fill_4 FILLER_56_377 ();
 sg13g2_fill_2 FILLER_56_381 ();
 sg13g2_fill_8 FILLER_56_388 ();
 sg13g2_fill_1 FILLER_56_402 ();
 sg13g2_fill_4 FILLER_56_440 ();
 sg13g2_fill_2 FILLER_56_444 ();
 sg13g2_fill_4 FILLER_56_451 ();
 sg13g2_fill_8 FILLER_56_461 ();
 sg13g2_fill_8 FILLER_56_469 ();
 sg13g2_fill_4 FILLER_56_477 ();
 sg13g2_fill_2 FILLER_56_481 ();
 sg13g2_fill_8 FILLER_56_492 ();
 sg13g2_fill_4 FILLER_56_500 ();
 sg13g2_fill_2 FILLER_56_504 ();
 sg13g2_fill_1 FILLER_56_532 ();
 sg13g2_fill_1 FILLER_56_590 ();
 sg13g2_fill_2 FILLER_56_639 ();
 sg13g2_fill_8 FILLER_56_700 ();
 sg13g2_fill_8 FILLER_56_708 ();
 sg13g2_fill_1 FILLER_56_716 ();
 sg13g2_fill_8 FILLER_56_742 ();
 sg13g2_fill_4 FILLER_56_750 ();
 sg13g2_fill_2 FILLER_56_754 ();
 sg13g2_fill_2 FILLER_56_801 ();
 sg13g2_fill_8 FILLER_56_837 ();
 sg13g2_fill_1 FILLER_56_845 ();
 sg13g2_fill_8 FILLER_56_856 ();
 sg13g2_fill_4 FILLER_56_864 ();
 sg13g2_fill_1 FILLER_56_868 ();
 sg13g2_fill_8 FILLER_56_906 ();
 sg13g2_fill_8 FILLER_56_914 ();
 sg13g2_fill_8 FILLER_56_922 ();
 sg13g2_fill_8 FILLER_56_930 ();
 sg13g2_fill_8 FILLER_56_938 ();
 sg13g2_fill_8 FILLER_56_946 ();
 sg13g2_fill_8 FILLER_56_954 ();
 sg13g2_fill_8 FILLER_56_962 ();
 sg13g2_fill_8 FILLER_56_970 ();
 sg13g2_fill_8 FILLER_56_978 ();
 sg13g2_fill_8 FILLER_56_986 ();
 sg13g2_fill_8 FILLER_56_994 ();
 sg13g2_fill_8 FILLER_56_1002 ();
 sg13g2_fill_8 FILLER_56_1010 ();
 sg13g2_fill_8 FILLER_56_1018 ();
 sg13g2_fill_8 FILLER_56_1026 ();
 sg13g2_fill_8 FILLER_56_1034 ();
 sg13g2_fill_8 FILLER_56_1042 ();
 sg13g2_fill_8 FILLER_56_1050 ();
 sg13g2_fill_8 FILLER_56_1058 ();
 sg13g2_fill_8 FILLER_56_1066 ();
 sg13g2_fill_8 FILLER_56_1074 ();
 sg13g2_fill_8 FILLER_56_1082 ();
 sg13g2_fill_8 FILLER_56_1090 ();
 sg13g2_fill_8 FILLER_56_1098 ();
 sg13g2_fill_8 FILLER_56_1106 ();
 sg13g2_fill_8 FILLER_56_1114 ();
 sg13g2_fill_8 FILLER_56_1122 ();
 sg13g2_fill_8 FILLER_56_1130 ();
 sg13g2_fill_8 FILLER_56_1138 ();
 sg13g2_fill_8 FILLER_56_1146 ();
 sg13g2_fill_8 FILLER_56_1154 ();
 sg13g2_fill_4 FILLER_56_1162 ();
 sg13g2_fill_8 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_8 ();
 sg13g2_fill_2 FILLER_57_17 ();
 sg13g2_fill_1 FILLER_57_19 ();
 sg13g2_fill_8 FILLER_57_28 ();
 sg13g2_fill_8 FILLER_57_36 ();
 sg13g2_fill_1 FILLER_57_44 ();
 sg13g2_fill_8 FILLER_57_83 ();
 sg13g2_fill_4 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_fill_8 FILLER_57_105 ();
 sg13g2_fill_2 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_124 ();
 sg13g2_fill_1 FILLER_57_126 ();
 sg13g2_fill_4 FILLER_57_133 ();
 sg13g2_fill_2 FILLER_57_137 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_fill_8 FILLER_57_145 ();
 sg13g2_fill_8 FILLER_57_153 ();
 sg13g2_fill_8 FILLER_57_161 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_fill_2 FILLER_57_212 ();
 sg13g2_fill_1 FILLER_57_214 ();
 sg13g2_fill_8 FILLER_57_234 ();
 sg13g2_fill_4 FILLER_57_242 ();
 sg13g2_fill_2 FILLER_57_246 ();
 sg13g2_fill_4 FILLER_57_279 ();
 sg13g2_fill_2 FILLER_57_291 ();
 sg13g2_fill_1 FILLER_57_293 ();
 sg13g2_fill_2 FILLER_57_299 ();
 sg13g2_fill_1 FILLER_57_301 ();
 sg13g2_fill_1 FILLER_57_311 ();
 sg13g2_fill_4 FILLER_57_338 ();
 sg13g2_fill_2 FILLER_57_342 ();
 sg13g2_fill_8 FILLER_57_380 ();
 sg13g2_fill_8 FILLER_57_388 ();
 sg13g2_fill_8 FILLER_57_396 ();
 sg13g2_fill_4 FILLER_57_421 ();
 sg13g2_fill_8 FILLER_57_461 ();
 sg13g2_fill_4 FILLER_57_475 ();
 sg13g2_fill_1 FILLER_57_479 ();
 sg13g2_fill_4 FILLER_57_485 ();
 sg13g2_fill_1 FILLER_57_489 ();
 sg13g2_fill_4 FILLER_57_499 ();
 sg13g2_fill_2 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_510 ();
 sg13g2_fill_2 FILLER_57_522 ();
 sg13g2_fill_1 FILLER_57_524 ();
 sg13g2_fill_4 FILLER_57_569 ();
 sg13g2_fill_1 FILLER_57_573 ();
 sg13g2_fill_2 FILLER_57_635 ();
 sg13g2_fill_1 FILLER_57_637 ();
 sg13g2_fill_8 FILLER_57_697 ();
 sg13g2_fill_1 FILLER_57_705 ();
 sg13g2_fill_8 FILLER_57_761 ();
 sg13g2_fill_4 FILLER_57_769 ();
 sg13g2_fill_2 FILLER_57_804 ();
 sg13g2_fill_4 FILLER_57_837 ();
 sg13g2_fill_4 FILLER_57_863 ();
 sg13g2_fill_1 FILLER_57_867 ();
 sg13g2_fill_4 FILLER_57_894 ();
 sg13g2_fill_1 FILLER_57_898 ();
 sg13g2_fill_8 FILLER_57_936 ();
 sg13g2_fill_8 FILLER_57_944 ();
 sg13g2_fill_8 FILLER_57_952 ();
 sg13g2_fill_8 FILLER_57_960 ();
 sg13g2_fill_8 FILLER_57_968 ();
 sg13g2_fill_8 FILLER_57_976 ();
 sg13g2_fill_8 FILLER_57_984 ();
 sg13g2_fill_8 FILLER_57_992 ();
 sg13g2_fill_8 FILLER_57_1000 ();
 sg13g2_fill_8 FILLER_57_1008 ();
 sg13g2_fill_8 FILLER_57_1016 ();
 sg13g2_fill_8 FILLER_57_1024 ();
 sg13g2_fill_8 FILLER_57_1032 ();
 sg13g2_fill_8 FILLER_57_1040 ();
 sg13g2_fill_8 FILLER_57_1048 ();
 sg13g2_fill_8 FILLER_57_1056 ();
 sg13g2_fill_8 FILLER_57_1064 ();
 sg13g2_fill_8 FILLER_57_1072 ();
 sg13g2_fill_8 FILLER_57_1080 ();
 sg13g2_fill_8 FILLER_57_1088 ();
 sg13g2_fill_8 FILLER_57_1096 ();
 sg13g2_fill_8 FILLER_57_1104 ();
 sg13g2_fill_8 FILLER_57_1112 ();
 sg13g2_fill_8 FILLER_57_1120 ();
 sg13g2_fill_8 FILLER_57_1128 ();
 sg13g2_fill_8 FILLER_57_1136 ();
 sg13g2_fill_8 FILLER_57_1144 ();
 sg13g2_fill_8 FILLER_57_1152 ();
 sg13g2_fill_4 FILLER_57_1160 ();
 sg13g2_fill_2 FILLER_57_1164 ();
 sg13g2_fill_8 FILLER_58_0 ();
 sg13g2_fill_8 FILLER_58_39 ();
 sg13g2_fill_8 FILLER_58_47 ();
 sg13g2_fill_4 FILLER_58_61 ();
 sg13g2_fill_4 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_82 ();
 sg13g2_fill_2 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_145 ();
 sg13g2_fill_8 FILLER_58_172 ();
 sg13g2_fill_4 FILLER_58_180 ();
 sg13g2_fill_2 FILLER_58_184 ();
 sg13g2_fill_1 FILLER_58_186 ();
 sg13g2_fill_4 FILLER_58_213 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_fill_4 FILLER_58_248 ();
 sg13g2_fill_2 FILLER_58_252 ();
 sg13g2_fill_1 FILLER_58_254 ();
 sg13g2_fill_4 FILLER_58_281 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_292 ();
 sg13g2_fill_8 FILLER_58_324 ();
 sg13g2_fill_8 FILLER_58_332 ();
 sg13g2_fill_2 FILLER_58_340 ();
 sg13g2_fill_1 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_359 ();
 sg13g2_fill_2 FILLER_58_366 ();
 sg13g2_fill_8 FILLER_58_376 ();
 sg13g2_fill_2 FILLER_58_384 ();
 sg13g2_fill_1 FILLER_58_391 ();
 sg13g2_fill_4 FILLER_58_398 ();
 sg13g2_fill_2 FILLER_58_402 ();
 sg13g2_fill_1 FILLER_58_404 ();
 sg13g2_fill_8 FILLER_58_419 ();
 sg13g2_fill_8 FILLER_58_427 ();
 sg13g2_fill_8 FILLER_58_435 ();
 sg13g2_fill_8 FILLER_58_443 ();
 sg13g2_fill_2 FILLER_58_451 ();
 sg13g2_fill_1 FILLER_58_453 ();
 sg13g2_fill_8 FILLER_58_484 ();
 sg13g2_fill_2 FILLER_58_504 ();
 sg13g2_fill_2 FILLER_58_566 ();
 sg13g2_fill_1 FILLER_58_568 ();
 sg13g2_fill_4 FILLER_58_573 ();
 sg13g2_fill_2 FILLER_58_583 ();
 sg13g2_fill_1 FILLER_58_585 ();
 sg13g2_fill_4 FILLER_58_637 ();
 sg13g2_fill_2 FILLER_58_651 ();
 sg13g2_fill_1 FILLER_58_653 ();
 sg13g2_fill_4 FILLER_58_690 ();
 sg13g2_fill_1 FILLER_58_694 ();
 sg13g2_fill_2 FILLER_58_725 ();
 sg13g2_fill_8 FILLER_58_757 ();
 sg13g2_fill_8 FILLER_58_765 ();
 sg13g2_fill_4 FILLER_58_773 ();
 sg13g2_fill_2 FILLER_58_777 ();
 sg13g2_fill_2 FILLER_58_805 ();
 sg13g2_fill_1 FILLER_58_807 ();
 sg13g2_fill_2 FILLER_58_818 ();
 sg13g2_fill_1 FILLER_58_820 ();
 sg13g2_fill_4 FILLER_58_847 ();
 sg13g2_fill_4 FILLER_58_862 ();
 sg13g2_fill_1 FILLER_58_876 ();
 sg13g2_fill_2 FILLER_58_897 ();
 sg13g2_fill_8 FILLER_58_925 ();
 sg13g2_fill_8 FILLER_58_933 ();
 sg13g2_fill_8 FILLER_58_941 ();
 sg13g2_fill_8 FILLER_58_949 ();
 sg13g2_fill_8 FILLER_58_957 ();
 sg13g2_fill_8 FILLER_58_965 ();
 sg13g2_fill_8 FILLER_58_973 ();
 sg13g2_fill_8 FILLER_58_981 ();
 sg13g2_fill_8 FILLER_58_989 ();
 sg13g2_fill_8 FILLER_58_997 ();
 sg13g2_fill_8 FILLER_58_1005 ();
 sg13g2_fill_8 FILLER_58_1013 ();
 sg13g2_fill_8 FILLER_58_1021 ();
 sg13g2_fill_8 FILLER_58_1029 ();
 sg13g2_fill_8 FILLER_58_1037 ();
 sg13g2_fill_8 FILLER_58_1045 ();
 sg13g2_fill_8 FILLER_58_1053 ();
 sg13g2_fill_8 FILLER_58_1061 ();
 sg13g2_fill_8 FILLER_58_1069 ();
 sg13g2_fill_8 FILLER_58_1077 ();
 sg13g2_fill_8 FILLER_58_1085 ();
 sg13g2_fill_8 FILLER_58_1093 ();
 sg13g2_fill_8 FILLER_58_1101 ();
 sg13g2_fill_8 FILLER_58_1109 ();
 sg13g2_fill_8 FILLER_58_1117 ();
 sg13g2_fill_8 FILLER_58_1125 ();
 sg13g2_fill_8 FILLER_58_1133 ();
 sg13g2_fill_8 FILLER_58_1141 ();
 sg13g2_fill_8 FILLER_58_1149 ();
 sg13g2_fill_8 FILLER_58_1157 ();
 sg13g2_fill_1 FILLER_58_1165 ();
 sg13g2_fill_8 FILLER_59_0 ();
 sg13g2_fill_8 FILLER_59_8 ();
 sg13g2_fill_4 FILLER_59_16 ();
 sg13g2_fill_2 FILLER_59_20 ();
 sg13g2_fill_8 FILLER_59_72 ();
 sg13g2_fill_1 FILLER_59_80 ();
 sg13g2_fill_2 FILLER_59_91 ();
 sg13g2_fill_1 FILLER_59_93 ();
 sg13g2_fill_8 FILLER_59_120 ();
 sg13g2_fill_4 FILLER_59_128 ();
 sg13g2_fill_2 FILLER_59_132 ();
 sg13g2_fill_1 FILLER_59_134 ();
 sg13g2_fill_4 FILLER_59_159 ();
 sg13g2_fill_8 FILLER_59_213 ();
 sg13g2_fill_1 FILLER_59_221 ();
 sg13g2_fill_8 FILLER_59_252 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_4 FILLER_59_312 ();
 sg13g2_fill_8 FILLER_59_326 ();
 sg13g2_fill_8 FILLER_59_334 ();
 sg13g2_fill_8 FILLER_59_342 ();
 sg13g2_fill_4 FILLER_59_350 ();
 sg13g2_fill_8 FILLER_59_358 ();
 sg13g2_fill_8 FILLER_59_366 ();
 sg13g2_fill_8 FILLER_59_374 ();
 sg13g2_fill_4 FILLER_59_382 ();
 sg13g2_fill_8 FILLER_59_409 ();
 sg13g2_fill_4 FILLER_59_417 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_fill_4 FILLER_59_431 ();
 sg13g2_fill_2 FILLER_59_435 ();
 sg13g2_fill_1 FILLER_59_442 ();
 sg13g2_fill_4 FILLER_59_456 ();
 sg13g2_fill_1 FILLER_59_460 ();
 sg13g2_fill_2 FILLER_59_467 ();
 sg13g2_fill_4 FILLER_59_473 ();
 sg13g2_fill_2 FILLER_59_477 ();
 sg13g2_fill_4 FILLER_59_482 ();
 sg13g2_fill_2 FILLER_59_486 ();
 sg13g2_fill_8 FILLER_59_513 ();
 sg13g2_fill_2 FILLER_59_521 ();
 sg13g2_fill_8 FILLER_59_528 ();
 sg13g2_fill_2 FILLER_59_606 ();
 sg13g2_fill_8 FILLER_59_684 ();
 sg13g2_fill_8 FILLER_59_692 ();
 sg13g2_fill_8 FILLER_59_700 ();
 sg13g2_fill_4 FILLER_59_708 ();
 sg13g2_fill_1 FILLER_59_717 ();
 sg13g2_fill_2 FILLER_59_737 ();
 sg13g2_fill_1 FILLER_59_739 ();
 sg13g2_fill_8 FILLER_59_745 ();
 sg13g2_fill_8 FILLER_59_753 ();
 sg13g2_fill_8 FILLER_59_761 ();
 sg13g2_fill_4 FILLER_59_769 ();
 sg13g2_fill_2 FILLER_59_773 ();
 sg13g2_fill_1 FILLER_59_775 ();
 sg13g2_fill_8 FILLER_59_784 ();
 sg13g2_fill_8 FILLER_59_792 ();
 sg13g2_fill_8 FILLER_59_800 ();
 sg13g2_fill_8 FILLER_59_838 ();
 sg13g2_fill_1 FILLER_59_846 ();
 sg13g2_fill_8 FILLER_59_852 ();
 sg13g2_fill_4 FILLER_59_860 ();
 sg13g2_fill_2 FILLER_59_864 ();
 sg13g2_fill_4 FILLER_59_876 ();
 sg13g2_fill_1 FILLER_59_880 ();
 sg13g2_fill_8 FILLER_59_916 ();
 sg13g2_fill_8 FILLER_59_924 ();
 sg13g2_fill_4 FILLER_59_932 ();
 sg13g2_fill_2 FILLER_59_936 ();
 sg13g2_fill_1 FILLER_59_938 ();
 sg13g2_fill_8 FILLER_59_965 ();
 sg13g2_fill_8 FILLER_59_973 ();
 sg13g2_fill_8 FILLER_59_981 ();
 sg13g2_fill_8 FILLER_59_989 ();
 sg13g2_fill_8 FILLER_59_997 ();
 sg13g2_fill_8 FILLER_59_1005 ();
 sg13g2_fill_8 FILLER_59_1013 ();
 sg13g2_fill_8 FILLER_59_1021 ();
 sg13g2_fill_8 FILLER_59_1029 ();
 sg13g2_fill_8 FILLER_59_1037 ();
 sg13g2_fill_8 FILLER_59_1045 ();
 sg13g2_fill_8 FILLER_59_1053 ();
 sg13g2_fill_8 FILLER_59_1061 ();
 sg13g2_fill_8 FILLER_59_1069 ();
 sg13g2_fill_8 FILLER_59_1077 ();
 sg13g2_fill_8 FILLER_59_1085 ();
 sg13g2_fill_8 FILLER_59_1093 ();
 sg13g2_fill_8 FILLER_59_1101 ();
 sg13g2_fill_8 FILLER_59_1109 ();
 sg13g2_fill_8 FILLER_59_1117 ();
 sg13g2_fill_8 FILLER_59_1125 ();
 sg13g2_fill_8 FILLER_59_1133 ();
 sg13g2_fill_8 FILLER_59_1141 ();
 sg13g2_fill_8 FILLER_59_1149 ();
 sg13g2_fill_8 FILLER_59_1157 ();
 sg13g2_fill_1 FILLER_59_1165 ();
 sg13g2_fill_2 FILLER_60_38 ();
 sg13g2_fill_4 FILLER_60_66 ();
 sg13g2_fill_1 FILLER_60_70 ();
 sg13g2_fill_8 FILLER_60_79 ();
 sg13g2_fill_2 FILLER_60_87 ();
 sg13g2_fill_1 FILLER_60_102 ();
 sg13g2_fill_8 FILLER_60_108 ();
 sg13g2_fill_8 FILLER_60_116 ();
 sg13g2_fill_8 FILLER_60_124 ();
 sg13g2_fill_8 FILLER_60_153 ();
 sg13g2_fill_4 FILLER_60_161 ();
 sg13g2_fill_4 FILLER_60_186 ();
 sg13g2_fill_1 FILLER_60_190 ();
 sg13g2_fill_8 FILLER_60_204 ();
 sg13g2_fill_8 FILLER_60_212 ();
 sg13g2_fill_2 FILLER_60_220 ();
 sg13g2_fill_8 FILLER_60_227 ();
 sg13g2_fill_8 FILLER_60_235 ();
 sg13g2_fill_8 FILLER_60_243 ();
 sg13g2_fill_8 FILLER_60_251 ();
 sg13g2_fill_8 FILLER_60_259 ();
 sg13g2_fill_8 FILLER_60_267 ();
 sg13g2_fill_8 FILLER_60_275 ();
 sg13g2_fill_8 FILLER_60_283 ();
 sg13g2_fill_4 FILLER_60_291 ();
 sg13g2_fill_2 FILLER_60_295 ();
 sg13g2_fill_1 FILLER_60_297 ();
 sg13g2_fill_2 FILLER_60_316 ();
 sg13g2_fill_1 FILLER_60_318 ();
 sg13g2_fill_8 FILLER_60_366 ();
 sg13g2_fill_4 FILLER_60_374 ();
 sg13g2_fill_2 FILLER_60_378 ();
 sg13g2_fill_1 FILLER_60_380 ();
 sg13g2_fill_8 FILLER_60_386 ();
 sg13g2_fill_1 FILLER_60_394 ();
 sg13g2_fill_8 FILLER_60_419 ();
 sg13g2_fill_2 FILLER_60_427 ();
 sg13g2_fill_8 FILLER_60_449 ();
 sg13g2_fill_1 FILLER_60_457 ();
 sg13g2_fill_8 FILLER_60_489 ();
 sg13g2_fill_4 FILLER_60_497 ();
 sg13g2_fill_2 FILLER_60_501 ();
 sg13g2_fill_1 FILLER_60_503 ();
 sg13g2_fill_8 FILLER_60_520 ();
 sg13g2_fill_8 FILLER_60_528 ();
 sg13g2_fill_2 FILLER_60_536 ();
 sg13g2_fill_1 FILLER_60_538 ();
 sg13g2_fill_4 FILLER_60_545 ();
 sg13g2_fill_1 FILLER_60_549 ();
 sg13g2_fill_8 FILLER_60_563 ();
 sg13g2_fill_4 FILLER_60_609 ();
 sg13g2_fill_2 FILLER_60_613 ();
 sg13g2_fill_2 FILLER_60_626 ();
 sg13g2_fill_1 FILLER_60_628 ();
 sg13g2_fill_8 FILLER_60_655 ();
 sg13g2_fill_8 FILLER_60_663 ();
 sg13g2_fill_8 FILLER_60_671 ();
 sg13g2_fill_8 FILLER_60_679 ();
 sg13g2_fill_4 FILLER_60_687 ();
 sg13g2_fill_2 FILLER_60_691 ();
 sg13g2_fill_4 FILLER_60_698 ();
 sg13g2_fill_4 FILLER_60_706 ();
 sg13g2_fill_2 FILLER_60_710 ();
 sg13g2_fill_2 FILLER_60_721 ();
 sg13g2_fill_8 FILLER_60_778 ();
 sg13g2_fill_8 FILLER_60_786 ();
 sg13g2_fill_4 FILLER_60_794 ();
 sg13g2_fill_1 FILLER_60_798 ();
 sg13g2_fill_8 FILLER_60_833 ();
 sg13g2_fill_8 FILLER_60_841 ();
 sg13g2_fill_8 FILLER_60_849 ();
 sg13g2_fill_8 FILLER_60_857 ();
 sg13g2_fill_8 FILLER_60_891 ();
 sg13g2_fill_1 FILLER_60_899 ();
 sg13g2_fill_2 FILLER_60_926 ();
 sg13g2_fill_1 FILLER_60_928 ();
 sg13g2_fill_8 FILLER_60_976 ();
 sg13g2_fill_8 FILLER_60_984 ();
 sg13g2_fill_8 FILLER_60_992 ();
 sg13g2_fill_8 FILLER_60_1000 ();
 sg13g2_fill_8 FILLER_60_1008 ();
 sg13g2_fill_8 FILLER_60_1016 ();
 sg13g2_fill_8 FILLER_60_1024 ();
 sg13g2_fill_8 FILLER_60_1032 ();
 sg13g2_fill_8 FILLER_60_1040 ();
 sg13g2_fill_8 FILLER_60_1048 ();
 sg13g2_fill_8 FILLER_60_1056 ();
 sg13g2_fill_8 FILLER_60_1064 ();
 sg13g2_fill_8 FILLER_60_1072 ();
 sg13g2_fill_8 FILLER_60_1080 ();
 sg13g2_fill_8 FILLER_60_1088 ();
 sg13g2_fill_8 FILLER_60_1096 ();
 sg13g2_fill_8 FILLER_60_1104 ();
 sg13g2_fill_8 FILLER_60_1112 ();
 sg13g2_fill_8 FILLER_60_1120 ();
 sg13g2_fill_8 FILLER_60_1128 ();
 sg13g2_fill_8 FILLER_60_1136 ();
 sg13g2_fill_8 FILLER_60_1144 ();
 sg13g2_fill_8 FILLER_60_1152 ();
 sg13g2_fill_4 FILLER_60_1160 ();
 sg13g2_fill_2 FILLER_60_1164 ();
 sg13g2_fill_4 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_4 ();
 sg13g2_fill_4 FILLER_61_35 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_fill_4 FILLER_61_53 ();
 sg13g2_fill_8 FILLER_61_86 ();
 sg13g2_fill_8 FILLER_61_94 ();
 sg13g2_fill_8 FILLER_61_102 ();
 sg13g2_fill_4 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_114 ();
 sg13g2_fill_1 FILLER_61_116 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_4 FILLER_61_144 ();
 sg13g2_fill_1 FILLER_61_148 ();
 sg13g2_fill_8 FILLER_61_159 ();
 sg13g2_fill_4 FILLER_61_167 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_4 FILLER_61_198 ();
 sg13g2_fill_8 FILLER_61_223 ();
 sg13g2_fill_8 FILLER_61_231 ();
 sg13g2_fill_8 FILLER_61_239 ();
 sg13g2_fill_4 FILLER_61_247 ();
 sg13g2_fill_2 FILLER_61_251 ();
 sg13g2_fill_8 FILLER_61_258 ();
 sg13g2_fill_8 FILLER_61_266 ();
 sg13g2_fill_8 FILLER_61_274 ();
 sg13g2_fill_4 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_286 ();
 sg13g2_fill_4 FILLER_61_313 ();
 sg13g2_fill_8 FILLER_61_343 ();
 sg13g2_fill_1 FILLER_61_351 ();
 sg13g2_fill_2 FILLER_61_358 ();
 sg13g2_fill_1 FILLER_61_360 ();
 sg13g2_fill_8 FILLER_61_382 ();
 sg13g2_fill_8 FILLER_61_390 ();
 sg13g2_fill_2 FILLER_61_398 ();
 sg13g2_fill_1 FILLER_61_400 ();
 sg13g2_fill_8 FILLER_61_409 ();
 sg13g2_fill_8 FILLER_61_417 ();
 sg13g2_fill_4 FILLER_61_425 ();
 sg13g2_fill_2 FILLER_61_429 ();
 sg13g2_fill_4 FILLER_61_438 ();
 sg13g2_fill_1 FILLER_61_442 ();
 sg13g2_fill_4 FILLER_61_451 ();
 sg13g2_fill_2 FILLER_61_455 ();
 sg13g2_fill_1 FILLER_61_457 ();
 sg13g2_fill_1 FILLER_61_492 ();
 sg13g2_fill_8 FILLER_61_496 ();
 sg13g2_fill_2 FILLER_61_504 ();
 sg13g2_fill_4 FILLER_61_574 ();
 sg13g2_fill_8 FILLER_61_613 ();
 sg13g2_fill_2 FILLER_61_621 ();
 sg13g2_fill_1 FILLER_61_623 ();
 sg13g2_fill_2 FILLER_61_629 ();
 sg13g2_fill_2 FILLER_61_646 ();
 sg13g2_fill_1 FILLER_61_648 ();
 sg13g2_fill_4 FILLER_61_655 ();
 sg13g2_fill_1 FILLER_61_659 ();
 sg13g2_fill_4 FILLER_61_686 ();
 sg13g2_fill_2 FILLER_61_694 ();
 sg13g2_fill_2 FILLER_61_713 ();
 sg13g2_fill_1 FILLER_61_736 ();
 sg13g2_fill_8 FILLER_61_767 ();
 sg13g2_fill_2 FILLER_61_775 ();
 sg13g2_fill_1 FILLER_61_777 ();
 sg13g2_fill_8 FILLER_61_808 ();
 sg13g2_fill_8 FILLER_61_816 ();
 sg13g2_fill_2 FILLER_61_832 ();
 sg13g2_fill_4 FILLER_61_859 ();
 sg13g2_fill_2 FILLER_61_863 ();
 sg13g2_fill_8 FILLER_61_891 ();
 sg13g2_fill_1 FILLER_61_899 ();
 sg13g2_fill_8 FILLER_61_947 ();
 sg13g2_fill_8 FILLER_61_955 ();
 sg13g2_fill_8 FILLER_61_963 ();
 sg13g2_fill_8 FILLER_61_971 ();
 sg13g2_fill_8 FILLER_61_979 ();
 sg13g2_fill_8 FILLER_61_987 ();
 sg13g2_fill_8 FILLER_61_995 ();
 sg13g2_fill_8 FILLER_61_1003 ();
 sg13g2_fill_8 FILLER_61_1011 ();
 sg13g2_fill_8 FILLER_61_1019 ();
 sg13g2_fill_8 FILLER_61_1027 ();
 sg13g2_fill_8 FILLER_61_1035 ();
 sg13g2_fill_8 FILLER_61_1043 ();
 sg13g2_fill_8 FILLER_61_1051 ();
 sg13g2_fill_8 FILLER_61_1059 ();
 sg13g2_fill_8 FILLER_61_1067 ();
 sg13g2_fill_8 FILLER_61_1075 ();
 sg13g2_fill_8 FILLER_61_1083 ();
 sg13g2_fill_8 FILLER_61_1091 ();
 sg13g2_fill_8 FILLER_61_1099 ();
 sg13g2_fill_8 FILLER_61_1107 ();
 sg13g2_fill_8 FILLER_61_1115 ();
 sg13g2_fill_8 FILLER_61_1123 ();
 sg13g2_fill_8 FILLER_61_1131 ();
 sg13g2_fill_8 FILLER_61_1139 ();
 sg13g2_fill_8 FILLER_61_1147 ();
 sg13g2_fill_8 FILLER_61_1155 ();
 sg13g2_fill_2 FILLER_61_1163 ();
 sg13g2_fill_1 FILLER_61_1165 ();
 sg13g2_fill_8 FILLER_62_0 ();
 sg13g2_fill_4 FILLER_62_8 ();
 sg13g2_fill_2 FILLER_62_12 ();
 sg13g2_fill_1 FILLER_62_14 ();
 sg13g2_fill_4 FILLER_62_25 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_fill_8 FILLER_62_78 ();
 sg13g2_fill_8 FILLER_62_86 ();
 sg13g2_fill_4 FILLER_62_94 ();
 sg13g2_fill_2 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_100 ();
 sg13g2_fill_4 FILLER_62_126 ();
 sg13g2_fill_8 FILLER_62_144 ();
 sg13g2_fill_8 FILLER_62_152 ();
 sg13g2_fill_4 FILLER_62_160 ();
 sg13g2_fill_2 FILLER_62_164 ();
 sg13g2_fill_8 FILLER_62_179 ();
 sg13g2_fill_8 FILLER_62_187 ();
 sg13g2_fill_8 FILLER_62_195 ();
 sg13g2_fill_8 FILLER_62_203 ();
 sg13g2_fill_8 FILLER_62_211 ();
 sg13g2_fill_8 FILLER_62_219 ();
 sg13g2_fill_8 FILLER_62_227 ();
 sg13g2_fill_8 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_243 ();
 sg13g2_fill_8 FILLER_62_267 ();
 sg13g2_fill_8 FILLER_62_275 ();
 sg13g2_fill_2 FILLER_62_283 ();
 sg13g2_fill_1 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_312 ();
 sg13g2_fill_2 FILLER_62_319 ();
 sg13g2_fill_1 FILLER_62_321 ();
 sg13g2_fill_4 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_62_412 ();
 sg13g2_fill_1 FILLER_62_414 ();
 sg13g2_fill_8 FILLER_62_502 ();
 sg13g2_fill_8 FILLER_62_510 ();
 sg13g2_fill_8 FILLER_62_518 ();
 sg13g2_fill_8 FILLER_62_526 ();
 sg13g2_fill_4 FILLER_62_534 ();
 sg13g2_fill_1 FILLER_62_538 ();
 sg13g2_fill_4 FILLER_62_545 ();
 sg13g2_fill_2 FILLER_62_549 ();
 sg13g2_fill_8 FILLER_62_557 ();
 sg13g2_fill_2 FILLER_62_565 ();
 sg13g2_fill_1 FILLER_62_567 ();
 sg13g2_fill_4 FILLER_62_572 ();
 sg13g2_fill_2 FILLER_62_576 ();
 sg13g2_fill_1 FILLER_62_578 ();
 sg13g2_fill_1 FILLER_62_584 ();
 sg13g2_fill_4 FILLER_62_591 ();
 sg13g2_fill_8 FILLER_62_630 ();
 sg13g2_fill_4 FILLER_62_638 ();
 sg13g2_fill_2 FILLER_62_642 ();
 sg13g2_fill_1 FILLER_62_644 ();
 sg13g2_fill_4 FILLER_62_651 ();
 sg13g2_fill_1 FILLER_62_655 ();
 sg13g2_fill_8 FILLER_62_682 ();
 sg13g2_fill_8 FILLER_62_690 ();
 sg13g2_fill_8 FILLER_62_698 ();
 sg13g2_fill_4 FILLER_62_706 ();
 sg13g2_fill_1 FILLER_62_710 ();
 sg13g2_fill_1 FILLER_62_717 ();
 sg13g2_fill_8 FILLER_62_741 ();
 sg13g2_fill_1 FILLER_62_749 ();
 sg13g2_fill_4 FILLER_62_755 ();
 sg13g2_fill_2 FILLER_62_796 ();
 sg13g2_fill_4 FILLER_62_879 ();
 sg13g2_fill_2 FILLER_62_883 ();
 sg13g2_fill_1 FILLER_62_885 ();
 sg13g2_fill_8 FILLER_62_907 ();
 sg13g2_fill_8 FILLER_62_915 ();
 sg13g2_fill_8 FILLER_62_923 ();
 sg13g2_fill_8 FILLER_62_931 ();
 sg13g2_fill_4 FILLER_62_939 ();
 sg13g2_fill_8 FILLER_62_969 ();
 sg13g2_fill_8 FILLER_62_977 ();
 sg13g2_fill_8 FILLER_62_985 ();
 sg13g2_fill_8 FILLER_62_993 ();
 sg13g2_fill_8 FILLER_62_1001 ();
 sg13g2_fill_8 FILLER_62_1009 ();
 sg13g2_fill_8 FILLER_62_1017 ();
 sg13g2_fill_8 FILLER_62_1025 ();
 sg13g2_fill_8 FILLER_62_1033 ();
 sg13g2_fill_8 FILLER_62_1041 ();
 sg13g2_fill_8 FILLER_62_1049 ();
 sg13g2_fill_8 FILLER_62_1057 ();
 sg13g2_fill_8 FILLER_62_1065 ();
 sg13g2_fill_8 FILLER_62_1073 ();
 sg13g2_fill_8 FILLER_62_1081 ();
 sg13g2_fill_8 FILLER_62_1089 ();
 sg13g2_fill_8 FILLER_62_1097 ();
 sg13g2_fill_8 FILLER_62_1105 ();
 sg13g2_fill_8 FILLER_62_1113 ();
 sg13g2_fill_8 FILLER_62_1121 ();
 sg13g2_fill_8 FILLER_62_1129 ();
 sg13g2_fill_8 FILLER_62_1137 ();
 sg13g2_fill_8 FILLER_62_1145 ();
 sg13g2_fill_8 FILLER_62_1153 ();
 sg13g2_fill_4 FILLER_62_1161 ();
 sg13g2_fill_1 FILLER_62_1165 ();
 sg13g2_fill_8 FILLER_63_25 ();
 sg13g2_fill_4 FILLER_63_33 ();
 sg13g2_fill_8 FILLER_63_50 ();
 sg13g2_fill_8 FILLER_63_58 ();
 sg13g2_fill_4 FILLER_63_66 ();
 sg13g2_fill_2 FILLER_63_70 ();
 sg13g2_fill_8 FILLER_63_101 ();
 sg13g2_fill_4 FILLER_63_109 ();
 sg13g2_fill_1 FILLER_63_113 ();
 sg13g2_fill_8 FILLER_63_152 ();
 sg13g2_fill_1 FILLER_63_160 ();
 sg13g2_fill_8 FILLER_63_186 ();
 sg13g2_fill_4 FILLER_63_194 ();
 sg13g2_fill_2 FILLER_63_198 ();
 sg13g2_fill_4 FILLER_63_229 ();
 sg13g2_fill_2 FILLER_63_233 ();
 sg13g2_fill_8 FILLER_63_269 ();
 sg13g2_fill_4 FILLER_63_277 ();
 sg13g2_fill_2 FILLER_63_281 ();
 sg13g2_fill_1 FILLER_63_283 ();
 sg13g2_fill_2 FILLER_63_318 ();
 sg13g2_fill_1 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_352 ();
 sg13g2_fill_8 FILLER_63_387 ();
 sg13g2_fill_8 FILLER_63_395 ();
 sg13g2_fill_4 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_63_407 ();
 sg13g2_fill_8 FILLER_63_418 ();
 sg13g2_fill_4 FILLER_63_432 ();
 sg13g2_fill_4 FILLER_63_509 ();
 sg13g2_fill_2 FILLER_63_523 ();
 sg13g2_fill_1 FILLER_63_525 ();
 sg13g2_fill_8 FILLER_63_533 ();
 sg13g2_fill_4 FILLER_63_567 ();
 sg13g2_fill_2 FILLER_63_571 ();
 sg13g2_fill_1 FILLER_63_573 ();
 sg13g2_fill_8 FILLER_63_590 ();
 sg13g2_fill_2 FILLER_63_598 ();
 sg13g2_fill_1 FILLER_63_600 ();
 sg13g2_fill_8 FILLER_63_607 ();
 sg13g2_fill_8 FILLER_63_615 ();
 sg13g2_fill_8 FILLER_63_623 ();
 sg13g2_fill_4 FILLER_63_631 ();
 sg13g2_fill_8 FILLER_63_649 ();
 sg13g2_fill_8 FILLER_63_657 ();
 sg13g2_fill_4 FILLER_63_665 ();
 sg13g2_fill_8 FILLER_63_687 ();
 sg13g2_fill_8 FILLER_63_700 ();
 sg13g2_fill_4 FILLER_63_708 ();
 sg13g2_fill_1 FILLER_63_712 ();
 sg13g2_fill_8 FILLER_63_739 ();
 sg13g2_fill_1 FILLER_63_747 ();
 sg13g2_fill_4 FILLER_63_753 ();
 sg13g2_fill_2 FILLER_63_757 ();
 sg13g2_fill_1 FILLER_63_759 ();
 sg13g2_fill_8 FILLER_63_767 ();
 sg13g2_fill_2 FILLER_63_775 ();
 sg13g2_fill_2 FILLER_63_782 ();
 sg13g2_fill_4 FILLER_63_788 ();
 sg13g2_fill_8 FILLER_63_805 ();
 sg13g2_fill_8 FILLER_63_813 ();
 sg13g2_fill_8 FILLER_63_821 ();
 sg13g2_fill_8 FILLER_63_829 ();
 sg13g2_fill_2 FILLER_63_837 ();
 sg13g2_fill_1 FILLER_63_839 ();
 sg13g2_fill_4 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_862 ();
 sg13g2_fill_1 FILLER_63_864 ();
 sg13g2_fill_8 FILLER_63_875 ();
 sg13g2_fill_8 FILLER_63_883 ();
 sg13g2_fill_8 FILLER_63_891 ();
 sg13g2_fill_8 FILLER_63_899 ();
 sg13g2_fill_8 FILLER_63_907 ();
 sg13g2_fill_8 FILLER_63_915 ();
 sg13g2_fill_8 FILLER_63_923 ();
 sg13g2_fill_2 FILLER_63_931 ();
 sg13g2_fill_8 FILLER_63_980 ();
 sg13g2_fill_8 FILLER_63_988 ();
 sg13g2_fill_8 FILLER_63_996 ();
 sg13g2_fill_8 FILLER_63_1004 ();
 sg13g2_fill_8 FILLER_63_1012 ();
 sg13g2_fill_8 FILLER_63_1020 ();
 sg13g2_fill_8 FILLER_63_1028 ();
 sg13g2_fill_8 FILLER_63_1036 ();
 sg13g2_fill_8 FILLER_63_1044 ();
 sg13g2_fill_8 FILLER_63_1052 ();
 sg13g2_fill_8 FILLER_63_1060 ();
 sg13g2_fill_8 FILLER_63_1068 ();
 sg13g2_fill_8 FILLER_63_1076 ();
 sg13g2_fill_8 FILLER_63_1084 ();
 sg13g2_fill_8 FILLER_63_1092 ();
 sg13g2_fill_8 FILLER_63_1100 ();
 sg13g2_fill_8 FILLER_63_1108 ();
 sg13g2_fill_8 FILLER_63_1116 ();
 sg13g2_fill_8 FILLER_63_1124 ();
 sg13g2_fill_8 FILLER_63_1132 ();
 sg13g2_fill_8 FILLER_63_1140 ();
 sg13g2_fill_8 FILLER_63_1148 ();
 sg13g2_fill_8 FILLER_63_1156 ();
 sg13g2_fill_2 FILLER_63_1164 ();
 sg13g2_fill_8 FILLER_64_0 ();
 sg13g2_fill_4 FILLER_64_8 ();
 sg13g2_fill_2 FILLER_64_12 ();
 sg13g2_fill_1 FILLER_64_14 ();
 sg13g2_fill_8 FILLER_64_20 ();
 sg13g2_fill_8 FILLER_64_28 ();
 sg13g2_fill_1 FILLER_64_36 ();
 sg13g2_fill_8 FILLER_64_63 ();
 sg13g2_fill_4 FILLER_64_71 ();
 sg13g2_fill_1 FILLER_64_96 ();
 sg13g2_fill_2 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_188 ();
 sg13g2_fill_1 FILLER_64_211 ();
 sg13g2_fill_1 FILLER_64_284 ();
 sg13g2_fill_8 FILLER_64_303 ();
 sg13g2_fill_8 FILLER_64_315 ();
 sg13g2_fill_2 FILLER_64_337 ();
 sg13g2_fill_4 FILLER_64_343 ();
 sg13g2_fill_8 FILLER_64_352 ();
 sg13g2_fill_8 FILLER_64_360 ();
 sg13g2_fill_8 FILLER_64_378 ();
 sg13g2_fill_8 FILLER_64_390 ();
 sg13g2_fill_4 FILLER_64_398 ();
 sg13g2_fill_1 FILLER_64_434 ();
 sg13g2_fill_2 FILLER_64_441 ();
 sg13g2_fill_1 FILLER_64_443 ();
 sg13g2_fill_4 FILLER_64_455 ();
 sg13g2_fill_2 FILLER_64_459 ();
 sg13g2_fill_1 FILLER_64_465 ();
 sg13g2_fill_8 FILLER_64_484 ();
 sg13g2_fill_8 FILLER_64_492 ();
 sg13g2_fill_8 FILLER_64_500 ();
 sg13g2_fill_2 FILLER_64_508 ();
 sg13g2_fill_1 FILLER_64_510 ();
 sg13g2_fill_4 FILLER_64_537 ();
 sg13g2_fill_2 FILLER_64_541 ();
 sg13g2_fill_4 FILLER_64_553 ();
 sg13g2_fill_4 FILLER_64_600 ();
 sg13g2_fill_1 FILLER_64_604 ();
 sg13g2_fill_2 FILLER_64_635 ();
 sg13g2_fill_4 FILLER_64_663 ();
 sg13g2_fill_8 FILLER_64_672 ();
 sg13g2_fill_2 FILLER_64_680 ();
 sg13g2_fill_1 FILLER_64_682 ();
 sg13g2_fill_1 FILLER_64_700 ();
 sg13g2_fill_8 FILLER_64_732 ();
 sg13g2_fill_8 FILLER_64_740 ();
 sg13g2_fill_2 FILLER_64_748 ();
 sg13g2_fill_1 FILLER_64_750 ();
 sg13g2_fill_8 FILLER_64_756 ();
 sg13g2_fill_8 FILLER_64_790 ();
 sg13g2_fill_4 FILLER_64_798 ();
 sg13g2_fill_2 FILLER_64_802 ();
 sg13g2_fill_1 FILLER_64_804 ();
 sg13g2_fill_8 FILLER_64_817 ();
 sg13g2_fill_8 FILLER_64_825 ();
 sg13g2_fill_8 FILLER_64_833 ();
 sg13g2_fill_8 FILLER_64_841 ();
 sg13g2_fill_1 FILLER_64_849 ();
 sg13g2_fill_2 FILLER_64_856 ();
 sg13g2_fill_1 FILLER_64_858 ();
 sg13g2_fill_8 FILLER_64_875 ();
 sg13g2_fill_4 FILLER_64_883 ();
 sg13g2_fill_1 FILLER_64_887 ();
 sg13g2_fill_4 FILLER_64_896 ();
 sg13g2_fill_1 FILLER_64_900 ();
 sg13g2_fill_8 FILLER_64_911 ();
 sg13g2_fill_8 FILLER_64_919 ();
 sg13g2_fill_8 FILLER_64_927 ();
 sg13g2_fill_8 FILLER_64_945 ();
 sg13g2_fill_1 FILLER_64_953 ();
 sg13g2_fill_8 FILLER_64_979 ();
 sg13g2_fill_8 FILLER_64_987 ();
 sg13g2_fill_8 FILLER_64_995 ();
 sg13g2_fill_8 FILLER_64_1003 ();
 sg13g2_fill_8 FILLER_64_1011 ();
 sg13g2_fill_8 FILLER_64_1019 ();
 sg13g2_fill_8 FILLER_64_1027 ();
 sg13g2_fill_8 FILLER_64_1035 ();
 sg13g2_fill_8 FILLER_64_1043 ();
 sg13g2_fill_8 FILLER_64_1051 ();
 sg13g2_fill_8 FILLER_64_1059 ();
 sg13g2_fill_8 FILLER_64_1067 ();
 sg13g2_fill_8 FILLER_64_1075 ();
 sg13g2_fill_8 FILLER_64_1083 ();
 sg13g2_fill_8 FILLER_64_1091 ();
 sg13g2_fill_8 FILLER_64_1099 ();
 sg13g2_fill_8 FILLER_64_1107 ();
 sg13g2_fill_8 FILLER_64_1115 ();
 sg13g2_fill_8 FILLER_64_1123 ();
 sg13g2_fill_8 FILLER_64_1131 ();
 sg13g2_fill_8 FILLER_64_1139 ();
 sg13g2_fill_8 FILLER_64_1147 ();
 sg13g2_fill_8 FILLER_64_1155 ();
 sg13g2_fill_2 FILLER_64_1163 ();
 sg13g2_fill_1 FILLER_64_1165 ();
 sg13g2_fill_8 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_8 ();
 sg13g2_fill_4 FILLER_65_35 ();
 sg13g2_fill_1 FILLER_65_39 ();
 sg13g2_fill_4 FILLER_65_45 ();
 sg13g2_fill_8 FILLER_65_98 ();
 sg13g2_fill_4 FILLER_65_130 ();
 sg13g2_fill_8 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_145 ();
 sg13g2_fill_1 FILLER_65_147 ();
 sg13g2_fill_8 FILLER_65_220 ();
 sg13g2_fill_8 FILLER_65_228 ();
 sg13g2_fill_4 FILLER_65_236 ();
 sg13g2_fill_2 FILLER_65_240 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_8 FILLER_65_251 ();
 sg13g2_fill_2 FILLER_65_259 ();
 sg13g2_fill_8 FILLER_65_282 ();
 sg13g2_fill_8 FILLER_65_290 ();
 sg13g2_fill_4 FILLER_65_298 ();
 sg13g2_fill_2 FILLER_65_302 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_337 ();
 sg13g2_fill_8 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_362 ();
 sg13g2_fill_8 FILLER_65_368 ();
 sg13g2_fill_4 FILLER_65_376 ();
 sg13g2_fill_2 FILLER_65_380 ();
 sg13g2_fill_1 FILLER_65_399 ();
 sg13g2_fill_2 FILLER_65_424 ();
 sg13g2_fill_1 FILLER_65_426 ();
 sg13g2_fill_4 FILLER_65_435 ();
 sg13g2_fill_2 FILLER_65_439 ();
 sg13g2_fill_4 FILLER_65_445 ();
 sg13g2_fill_2 FILLER_65_449 ();
 sg13g2_fill_8 FILLER_65_456 ();
 sg13g2_fill_1 FILLER_65_464 ();
 sg13g2_fill_8 FILLER_65_469 ();
 sg13g2_fill_8 FILLER_65_477 ();
 sg13g2_fill_8 FILLER_65_485 ();
 sg13g2_fill_1 FILLER_65_498 ();
 sg13g2_fill_8 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_551 ();
 sg13g2_fill_4 FILLER_65_560 ();
 sg13g2_fill_2 FILLER_65_564 ();
 sg13g2_fill_4 FILLER_65_602 ();
 sg13g2_fill_2 FILLER_65_606 ();
 sg13g2_fill_1 FILLER_65_608 ();
 sg13g2_fill_4 FILLER_65_615 ();
 sg13g2_fill_4 FILLER_65_683 ();
 sg13g2_fill_8 FILLER_65_723 ();
 sg13g2_fill_8 FILLER_65_731 ();
 sg13g2_fill_8 FILLER_65_739 ();
 sg13g2_fill_8 FILLER_65_747 ();
 sg13g2_fill_8 FILLER_65_755 ();
 sg13g2_fill_2 FILLER_65_763 ();
 sg13g2_fill_8 FILLER_65_783 ();
 sg13g2_fill_8 FILLER_65_791 ();
 sg13g2_fill_1 FILLER_65_799 ();
 sg13g2_fill_2 FILLER_65_814 ();
 sg13g2_fill_2 FILLER_65_821 ();
 sg13g2_fill_1 FILLER_65_823 ();
 sg13g2_fill_1 FILLER_65_829 ();
 sg13g2_fill_8 FILLER_65_835 ();
 sg13g2_fill_4 FILLER_65_843 ();
 sg13g2_fill_2 FILLER_65_847 ();
 sg13g2_fill_2 FILLER_65_867 ();
 sg13g2_fill_4 FILLER_65_895 ();
 sg13g2_fill_2 FILLER_65_899 ();
 sg13g2_fill_4 FILLER_65_927 ();
 sg13g2_fill_8 FILLER_65_967 ();
 sg13g2_fill_8 FILLER_65_975 ();
 sg13g2_fill_8 FILLER_65_983 ();
 sg13g2_fill_8 FILLER_65_991 ();
 sg13g2_fill_8 FILLER_65_999 ();
 sg13g2_fill_8 FILLER_65_1007 ();
 sg13g2_fill_8 FILLER_65_1015 ();
 sg13g2_fill_8 FILLER_65_1023 ();
 sg13g2_fill_8 FILLER_65_1031 ();
 sg13g2_fill_8 FILLER_65_1039 ();
 sg13g2_fill_8 FILLER_65_1047 ();
 sg13g2_fill_8 FILLER_65_1055 ();
 sg13g2_fill_8 FILLER_65_1063 ();
 sg13g2_fill_8 FILLER_65_1071 ();
 sg13g2_fill_8 FILLER_65_1079 ();
 sg13g2_fill_8 FILLER_65_1087 ();
 sg13g2_fill_8 FILLER_65_1095 ();
 sg13g2_fill_8 FILLER_65_1103 ();
 sg13g2_fill_8 FILLER_65_1111 ();
 sg13g2_fill_8 FILLER_65_1119 ();
 sg13g2_fill_8 FILLER_65_1127 ();
 sg13g2_fill_8 FILLER_65_1135 ();
 sg13g2_fill_8 FILLER_65_1143 ();
 sg13g2_fill_8 FILLER_65_1151 ();
 sg13g2_fill_4 FILLER_65_1159 ();
 sg13g2_fill_2 FILLER_65_1163 ();
 sg13g2_fill_1 FILLER_65_1165 ();
 sg13g2_fill_8 FILLER_66_0 ();
 sg13g2_fill_4 FILLER_66_8 ();
 sg13g2_fill_2 FILLER_66_12 ();
 sg13g2_fill_1 FILLER_66_14 ();
 sg13g2_fill_8 FILLER_66_31 ();
 sg13g2_fill_2 FILLER_66_39 ();
 sg13g2_fill_8 FILLER_66_113 ();
 sg13g2_fill_2 FILLER_66_121 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_fill_4 FILLER_66_155 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_fill_4 FILLER_66_163 ();
 sg13g2_fill_8 FILLER_66_213 ();
 sg13g2_fill_8 FILLER_66_234 ();
 sg13g2_fill_4 FILLER_66_242 ();
 sg13g2_fill_2 FILLER_66_246 ();
 sg13g2_fill_1 FILLER_66_248 ();
 sg13g2_fill_2 FILLER_66_253 ();
 sg13g2_fill_1 FILLER_66_255 ();
 sg13g2_fill_4 FILLER_66_262 ();
 sg13g2_fill_4 FILLER_66_295 ();
 sg13g2_fill_2 FILLER_66_299 ();
 sg13g2_fill_1 FILLER_66_301 ();
 sg13g2_fill_2 FILLER_66_307 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_fill_2 FILLER_66_358 ();
 sg13g2_fill_8 FILLER_66_378 ();
 sg13g2_fill_8 FILLER_66_386 ();
 sg13g2_fill_1 FILLER_66_394 ();
 sg13g2_fill_8 FILLER_66_414 ();
 sg13g2_fill_2 FILLER_66_422 ();
 sg13g2_fill_1 FILLER_66_424 ();
 sg13g2_fill_4 FILLER_66_433 ();
 sg13g2_fill_2 FILLER_66_437 ();
 sg13g2_fill_2 FILLER_66_477 ();
 sg13g2_fill_8 FILLER_66_512 ();
 sg13g2_fill_4 FILLER_66_520 ();
 sg13g2_fill_1 FILLER_66_524 ();
 sg13g2_fill_8 FILLER_66_597 ();
 sg13g2_fill_8 FILLER_66_605 ();
 sg13g2_fill_8 FILLER_66_613 ();
 sg13g2_fill_4 FILLER_66_621 ();
 sg13g2_fill_2 FILLER_66_625 ();
 sg13g2_fill_8 FILLER_66_638 ();
 sg13g2_fill_1 FILLER_66_646 ();
 sg13g2_fill_1 FILLER_66_656 ();
 sg13g2_fill_1 FILLER_66_663 ();
 sg13g2_fill_8 FILLER_66_674 ();
 sg13g2_fill_8 FILLER_66_682 ();
 sg13g2_fill_8 FILLER_66_690 ();
 sg13g2_fill_8 FILLER_66_698 ();
 sg13g2_fill_4 FILLER_66_706 ();
 sg13g2_fill_2 FILLER_66_710 ();
 sg13g2_fill_1 FILLER_66_712 ();
 sg13g2_fill_4 FILLER_66_717 ();
 sg13g2_fill_2 FILLER_66_721 ();
 sg13g2_fill_4 FILLER_66_733 ();
 sg13g2_fill_8 FILLER_66_767 ();
 sg13g2_fill_8 FILLER_66_775 ();
 sg13g2_fill_4 FILLER_66_783 ();
 sg13g2_fill_2 FILLER_66_787 ();
 sg13g2_fill_1 FILLER_66_789 ();
 sg13g2_fill_2 FILLER_66_797 ();
 sg13g2_fill_2 FILLER_66_822 ();
 sg13g2_fill_1 FILLER_66_824 ();
 sg13g2_fill_8 FILLER_66_842 ();
 sg13g2_fill_1 FILLER_66_850 ();
 sg13g2_fill_2 FILLER_66_857 ();
 sg13g2_fill_4 FILLER_66_895 ();
 sg13g2_fill_2 FILLER_66_899 ();
 sg13g2_fill_1 FILLER_66_901 ();
 sg13g2_fill_2 FILLER_66_939 ();
 sg13g2_fill_8 FILLER_66_978 ();
 sg13g2_fill_8 FILLER_66_986 ();
 sg13g2_fill_8 FILLER_66_994 ();
 sg13g2_fill_8 FILLER_66_1002 ();
 sg13g2_fill_8 FILLER_66_1010 ();
 sg13g2_fill_8 FILLER_66_1018 ();
 sg13g2_fill_8 FILLER_66_1026 ();
 sg13g2_fill_8 FILLER_66_1034 ();
 sg13g2_fill_8 FILLER_66_1042 ();
 sg13g2_fill_8 FILLER_66_1050 ();
 sg13g2_fill_8 FILLER_66_1058 ();
 sg13g2_fill_8 FILLER_66_1066 ();
 sg13g2_fill_8 FILLER_66_1074 ();
 sg13g2_fill_8 FILLER_66_1082 ();
 sg13g2_fill_8 FILLER_66_1090 ();
 sg13g2_fill_8 FILLER_66_1098 ();
 sg13g2_fill_8 FILLER_66_1106 ();
 sg13g2_fill_8 FILLER_66_1114 ();
 sg13g2_fill_8 FILLER_66_1122 ();
 sg13g2_fill_8 FILLER_66_1130 ();
 sg13g2_fill_8 FILLER_66_1138 ();
 sg13g2_fill_8 FILLER_66_1146 ();
 sg13g2_fill_8 FILLER_66_1154 ();
 sg13g2_fill_4 FILLER_66_1162 ();
 sg13g2_fill_8 FILLER_67_0 ();
 sg13g2_fill_8 FILLER_67_34 ();
 sg13g2_fill_2 FILLER_67_73 ();
 sg13g2_fill_1 FILLER_67_75 ();
 sg13g2_fill_4 FILLER_67_84 ();
 sg13g2_fill_8 FILLER_67_93 ();
 sg13g2_fill_8 FILLER_67_101 ();
 sg13g2_fill_8 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_117 ();
 sg13g2_fill_8 FILLER_67_137 ();
 sg13g2_fill_1 FILLER_67_145 ();
 sg13g2_fill_2 FILLER_67_151 ();
 sg13g2_fill_8 FILLER_67_172 ();
 sg13g2_fill_8 FILLER_67_180 ();
 sg13g2_fill_8 FILLER_67_213 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_fill_2 FILLER_67_295 ();
 sg13g2_fill_4 FILLER_67_323 ();
 sg13g2_fill_2 FILLER_67_327 ();
 sg13g2_fill_8 FILLER_67_346 ();
 sg13g2_fill_4 FILLER_67_354 ();
 sg13g2_fill_2 FILLER_67_358 ();
 sg13g2_fill_1 FILLER_67_360 ();
 sg13g2_fill_1 FILLER_67_384 ();
 sg13g2_fill_4 FILLER_67_404 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_fill_2 FILLER_67_414 ();
 sg13g2_fill_1 FILLER_67_416 ();
 sg13g2_fill_8 FILLER_67_438 ();
 sg13g2_fill_2 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_455 ();
 sg13g2_fill_2 FILLER_67_476 ();
 sg13g2_fill_2 FILLER_67_495 ();
 sg13g2_fill_8 FILLER_67_516 ();
 sg13g2_fill_8 FILLER_67_524 ();
 sg13g2_fill_4 FILLER_67_532 ();
 sg13g2_fill_8 FILLER_67_543 ();
 sg13g2_fill_8 FILLER_67_551 ();
 sg13g2_fill_8 FILLER_67_559 ();
 sg13g2_fill_4 FILLER_67_567 ();
 sg13g2_fill_2 FILLER_67_571 ();
 sg13g2_fill_4 FILLER_67_580 ();
 sg13g2_fill_1 FILLER_67_584 ();
 sg13g2_fill_4 FILLER_67_593 ();
 sg13g2_fill_2 FILLER_67_597 ();
 sg13g2_fill_4 FILLER_67_607 ();
 sg13g2_fill_2 FILLER_67_611 ();
 sg13g2_fill_4 FILLER_67_626 ();
 sg13g2_fill_1 FILLER_67_630 ();
 sg13g2_fill_1 FILLER_67_682 ();
 sg13g2_fill_8 FILLER_67_688 ();
 sg13g2_fill_8 FILLER_67_696 ();
 sg13g2_fill_2 FILLER_67_704 ();
 sg13g2_fill_1 FILLER_67_706 ();
 sg13g2_fill_8 FILLER_67_742 ();
 sg13g2_fill_2 FILLER_67_750 ();
 sg13g2_fill_4 FILLER_67_775 ();
 sg13g2_fill_2 FILLER_67_779 ();
 sg13g2_fill_1 FILLER_67_781 ();
 sg13g2_fill_2 FILLER_67_793 ();
 sg13g2_fill_2 FILLER_67_826 ();
 sg13g2_fill_8 FILLER_67_839 ();
 sg13g2_fill_8 FILLER_67_847 ();
 sg13g2_fill_1 FILLER_67_855 ();
 sg13g2_fill_4 FILLER_67_862 ();
 sg13g2_fill_8 FILLER_67_876 ();
 sg13g2_fill_4 FILLER_67_884 ();
 sg13g2_fill_1 FILLER_67_934 ();
 sg13g2_fill_8 FILLER_67_945 ();
 sg13g2_fill_8 FILLER_67_953 ();
 sg13g2_fill_1 FILLER_67_961 ();
 sg13g2_fill_4 FILLER_67_970 ();
 sg13g2_fill_1 FILLER_67_974 ();
 sg13g2_fill_8 FILLER_67_1001 ();
 sg13g2_fill_8 FILLER_67_1009 ();
 sg13g2_fill_8 FILLER_67_1017 ();
 sg13g2_fill_8 FILLER_67_1025 ();
 sg13g2_fill_8 FILLER_67_1033 ();
 sg13g2_fill_8 FILLER_67_1041 ();
 sg13g2_fill_8 FILLER_67_1049 ();
 sg13g2_fill_8 FILLER_67_1057 ();
 sg13g2_fill_8 FILLER_67_1065 ();
 sg13g2_fill_8 FILLER_67_1073 ();
 sg13g2_fill_8 FILLER_67_1081 ();
 sg13g2_fill_8 FILLER_67_1089 ();
 sg13g2_fill_8 FILLER_67_1097 ();
 sg13g2_fill_8 FILLER_67_1105 ();
 sg13g2_fill_8 FILLER_67_1113 ();
 sg13g2_fill_8 FILLER_67_1121 ();
 sg13g2_fill_8 FILLER_67_1129 ();
 sg13g2_fill_8 FILLER_67_1137 ();
 sg13g2_fill_8 FILLER_67_1145 ();
 sg13g2_fill_8 FILLER_67_1153 ();
 sg13g2_fill_4 FILLER_67_1161 ();
 sg13g2_fill_1 FILLER_67_1165 ();
 sg13g2_fill_2 FILLER_68_69 ();
 sg13g2_fill_1 FILLER_68_71 ();
 sg13g2_fill_8 FILLER_68_98 ();
 sg13g2_fill_8 FILLER_68_106 ();
 sg13g2_fill_8 FILLER_68_114 ();
 sg13g2_fill_4 FILLER_68_122 ();
 sg13g2_fill_8 FILLER_68_131 ();
 sg13g2_fill_8 FILLER_68_139 ();
 sg13g2_fill_4 FILLER_68_147 ();
 sg13g2_fill_1 FILLER_68_151 ();
 sg13g2_fill_2 FILLER_68_219 ();
 sg13g2_fill_1 FILLER_68_221 ();
 sg13g2_fill_8 FILLER_68_248 ();
 sg13g2_fill_8 FILLER_68_256 ();
 sg13g2_fill_1 FILLER_68_264 ();
 sg13g2_fill_2 FILLER_68_305 ();
 sg13g2_fill_1 FILLER_68_307 ();
 sg13g2_fill_8 FILLER_68_314 ();
 sg13g2_fill_8 FILLER_68_322 ();
 sg13g2_fill_1 FILLER_68_330 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_8 FILLER_68_351 ();
 sg13g2_fill_4 FILLER_68_359 ();
 sg13g2_fill_2 FILLER_68_363 ();
 sg13g2_fill_1 FILLER_68_365 ();
 sg13g2_fill_2 FILLER_68_387 ();
 sg13g2_fill_1 FILLER_68_389 ();
 sg13g2_fill_1 FILLER_68_395 ();
 sg13g2_fill_2 FILLER_68_400 ();
 sg13g2_fill_4 FILLER_68_415 ();
 sg13g2_fill_2 FILLER_68_419 ();
 sg13g2_fill_1 FILLER_68_421 ();
 sg13g2_fill_8 FILLER_68_465 ();
 sg13g2_fill_8 FILLER_68_473 ();
 sg13g2_fill_8 FILLER_68_486 ();
 sg13g2_fill_1 FILLER_68_494 ();
 sg13g2_fill_8 FILLER_68_500 ();
 sg13g2_fill_4 FILLER_68_508 ();
 sg13g2_fill_2 FILLER_68_512 ();
 sg13g2_fill_1 FILLER_68_514 ();
 sg13g2_fill_2 FILLER_68_527 ();
 sg13g2_fill_8 FILLER_68_561 ();
 sg13g2_fill_8 FILLER_68_569 ();
 sg13g2_fill_8 FILLER_68_577 ();
 sg13g2_fill_8 FILLER_68_585 ();
 sg13g2_fill_8 FILLER_68_593 ();
 sg13g2_fill_4 FILLER_68_601 ();
 sg13g2_fill_2 FILLER_68_613 ();
 sg13g2_fill_1 FILLER_68_615 ();
 sg13g2_fill_4 FILLER_68_679 ();
 sg13g2_fill_2 FILLER_68_683 ();
 sg13g2_fill_8 FILLER_68_698 ();
 sg13g2_fill_2 FILLER_68_706 ();
 sg13g2_fill_1 FILLER_68_708 ();
 sg13g2_fill_2 FILLER_68_736 ();
 sg13g2_fill_1 FILLER_68_738 ();
 sg13g2_fill_4 FILLER_68_784 ();
 sg13g2_fill_1 FILLER_68_788 ();
 sg13g2_fill_1 FILLER_68_794 ();
 sg13g2_fill_8 FILLER_68_813 ();
 sg13g2_fill_8 FILLER_68_872 ();
 sg13g2_fill_8 FILLER_68_880 ();
 sg13g2_fill_8 FILLER_68_888 ();
 sg13g2_fill_4 FILLER_68_896 ();
 sg13g2_fill_2 FILLER_68_900 ();
 sg13g2_fill_8 FILLER_68_943 ();
 sg13g2_fill_8 FILLER_68_951 ();
 sg13g2_fill_8 FILLER_68_959 ();
 sg13g2_fill_8 FILLER_68_967 ();
 sg13g2_fill_8 FILLER_68_1001 ();
 sg13g2_fill_8 FILLER_68_1009 ();
 sg13g2_fill_8 FILLER_68_1017 ();
 sg13g2_fill_8 FILLER_68_1025 ();
 sg13g2_fill_8 FILLER_68_1033 ();
 sg13g2_fill_8 FILLER_68_1041 ();
 sg13g2_fill_8 FILLER_68_1049 ();
 sg13g2_fill_8 FILLER_68_1057 ();
 sg13g2_fill_8 FILLER_68_1065 ();
 sg13g2_fill_8 FILLER_68_1073 ();
 sg13g2_fill_8 FILLER_68_1081 ();
 sg13g2_fill_8 FILLER_68_1089 ();
 sg13g2_fill_8 FILLER_68_1097 ();
 sg13g2_fill_8 FILLER_68_1105 ();
 sg13g2_fill_8 FILLER_68_1113 ();
 sg13g2_fill_8 FILLER_68_1121 ();
 sg13g2_fill_8 FILLER_68_1129 ();
 sg13g2_fill_8 FILLER_68_1137 ();
 sg13g2_fill_8 FILLER_68_1145 ();
 sg13g2_fill_8 FILLER_68_1153 ();
 sg13g2_fill_4 FILLER_68_1161 ();
 sg13g2_fill_1 FILLER_68_1165 ();
 sg13g2_fill_8 FILLER_69_0 ();
 sg13g2_fill_8 FILLER_69_8 ();
 sg13g2_fill_8 FILLER_69_16 ();
 sg13g2_fill_8 FILLER_69_24 ();
 sg13g2_fill_8 FILLER_69_32 ();
 sg13g2_fill_8 FILLER_69_40 ();
 sg13g2_fill_4 FILLER_69_48 ();
 sg13g2_fill_8 FILLER_69_56 ();
 sg13g2_fill_8 FILLER_69_64 ();
 sg13g2_fill_8 FILLER_69_72 ();
 sg13g2_fill_4 FILLER_69_80 ();
 sg13g2_fill_4 FILLER_69_107 ();
 sg13g2_fill_2 FILLER_69_111 ();
 sg13g2_fill_1 FILLER_69_113 ();
 sg13g2_fill_8 FILLER_69_122 ();
 sg13g2_fill_8 FILLER_69_130 ();
 sg13g2_fill_4 FILLER_69_138 ();
 sg13g2_fill_2 FILLER_69_142 ();
 sg13g2_fill_1 FILLER_69_144 ();
 sg13g2_fill_2 FILLER_69_149 ();
 sg13g2_fill_8 FILLER_69_166 ();
 sg13g2_fill_8 FILLER_69_174 ();
 sg13g2_fill_4 FILLER_69_182 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_fill_1 FILLER_69_188 ();
 sg13g2_fill_4 FILLER_69_215 ();
 sg13g2_fill_1 FILLER_69_219 ();
 sg13g2_fill_8 FILLER_69_225 ();
 sg13g2_fill_8 FILLER_69_233 ();
 sg13g2_fill_2 FILLER_69_241 ();
 sg13g2_fill_1 FILLER_69_243 ();
 sg13g2_fill_8 FILLER_69_254 ();
 sg13g2_fill_8 FILLER_69_262 ();
 sg13g2_fill_4 FILLER_69_270 ();
 sg13g2_fill_2 FILLER_69_279 ();
 sg13g2_fill_8 FILLER_69_284 ();
 sg13g2_fill_4 FILLER_69_292 ();
 sg13g2_fill_1 FILLER_69_296 ();
 sg13g2_fill_4 FILLER_69_306 ();
 sg13g2_fill_8 FILLER_69_315 ();
 sg13g2_fill_8 FILLER_69_323 ();
 sg13g2_fill_8 FILLER_69_331 ();
 sg13g2_fill_8 FILLER_69_342 ();
 sg13g2_fill_4 FILLER_69_350 ();
 sg13g2_fill_2 FILLER_69_372 ();
 sg13g2_fill_1 FILLER_69_374 ();
 sg13g2_fill_2 FILLER_69_388 ();
 sg13g2_fill_1 FILLER_69_390 ();
 sg13g2_fill_1 FILLER_69_403 ();
 sg13g2_fill_1 FILLER_69_424 ();
 sg13g2_fill_4 FILLER_69_440 ();
 sg13g2_fill_1 FILLER_69_444 ();
 sg13g2_fill_1 FILLER_69_450 ();
 sg13g2_fill_2 FILLER_69_465 ();
 sg13g2_fill_2 FILLER_69_472 ();
 sg13g2_fill_2 FILLER_69_497 ();
 sg13g2_fill_1 FILLER_69_499 ();
 sg13g2_fill_2 FILLER_69_531 ();
 sg13g2_fill_8 FILLER_69_541 ();
 sg13g2_fill_1 FILLER_69_549 ();
 sg13g2_fill_8 FILLER_69_556 ();
 sg13g2_fill_1 FILLER_69_564 ();
 sg13g2_fill_4 FILLER_69_584 ();
 sg13g2_fill_2 FILLER_69_588 ();
 sg13g2_fill_8 FILLER_69_623 ();
 sg13g2_fill_8 FILLER_69_631 ();
 sg13g2_fill_8 FILLER_69_639 ();
 sg13g2_fill_1 FILLER_69_647 ();
 sg13g2_fill_2 FILLER_69_652 ();
 sg13g2_fill_1 FILLER_69_654 ();
 sg13g2_fill_8 FILLER_69_670 ();
 sg13g2_fill_1 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_718 ();
 sg13g2_fill_8 FILLER_69_755 ();
 sg13g2_fill_2 FILLER_69_763 ();
 sg13g2_fill_4 FILLER_69_786 ();
 sg13g2_fill_2 FILLER_69_790 ();
 sg13g2_fill_2 FILLER_69_807 ();
 sg13g2_fill_1 FILLER_69_809 ();
 sg13g2_fill_1 FILLER_69_833 ();
 sg13g2_fill_1 FILLER_69_839 ();
 sg13g2_fill_8 FILLER_69_850 ();
 sg13g2_fill_8 FILLER_69_858 ();
 sg13g2_fill_8 FILLER_69_866 ();
 sg13g2_fill_4 FILLER_69_874 ();
 sg13g2_fill_8 FILLER_69_927 ();
 sg13g2_fill_1 FILLER_69_935 ();
 sg13g2_fill_4 FILLER_69_982 ();
 sg13g2_fill_8 FILLER_69_997 ();
 sg13g2_fill_8 FILLER_69_1005 ();
 sg13g2_fill_2 FILLER_69_1013 ();
 sg13g2_fill_1 FILLER_69_1015 ();
 sg13g2_fill_8 FILLER_69_1042 ();
 sg13g2_fill_8 FILLER_69_1050 ();
 sg13g2_fill_8 FILLER_69_1058 ();
 sg13g2_fill_8 FILLER_69_1066 ();
 sg13g2_fill_8 FILLER_69_1074 ();
 sg13g2_fill_8 FILLER_69_1082 ();
 sg13g2_fill_8 FILLER_69_1090 ();
 sg13g2_fill_8 FILLER_69_1098 ();
 sg13g2_fill_8 FILLER_69_1106 ();
 sg13g2_fill_8 FILLER_69_1114 ();
 sg13g2_fill_8 FILLER_69_1122 ();
 sg13g2_fill_8 FILLER_69_1130 ();
 sg13g2_fill_8 FILLER_69_1138 ();
 sg13g2_fill_8 FILLER_69_1146 ();
 sg13g2_fill_8 FILLER_69_1154 ();
 sg13g2_fill_4 FILLER_69_1162 ();
 sg13g2_fill_4 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_4 ();
 sg13g2_fill_1 FILLER_70_6 ();
 sg13g2_fill_4 FILLER_70_23 ();
 sg13g2_fill_2 FILLER_70_27 ();
 sg13g2_fill_1 FILLER_70_34 ();
 sg13g2_fill_8 FILLER_70_38 ();
 sg13g2_fill_8 FILLER_70_46 ();
 sg13g2_fill_8 FILLER_70_54 ();
 sg13g2_fill_8 FILLER_70_62 ();
 sg13g2_fill_8 FILLER_70_70 ();
 sg13g2_fill_4 FILLER_70_78 ();
 sg13g2_fill_2 FILLER_70_82 ();
 sg13g2_fill_1 FILLER_70_84 ();
 sg13g2_fill_1 FILLER_70_91 ();
 sg13g2_fill_1 FILLER_70_141 ();
 sg13g2_fill_8 FILLER_70_174 ();
 sg13g2_fill_8 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_190 ();
 sg13g2_fill_4 FILLER_70_197 ();
 sg13g2_fill_8 FILLER_70_209 ();
 sg13g2_fill_8 FILLER_70_217 ();
 sg13g2_fill_8 FILLER_70_225 ();
 sg13g2_fill_2 FILLER_70_241 ();
 sg13g2_fill_1 FILLER_70_243 ();
 sg13g2_fill_8 FILLER_70_269 ();
 sg13g2_fill_4 FILLER_70_277 ();
 sg13g2_fill_1 FILLER_70_293 ();
 sg13g2_fill_2 FILLER_70_305 ();
 sg13g2_fill_8 FILLER_70_314 ();
 sg13g2_fill_2 FILLER_70_322 ();
 sg13g2_fill_1 FILLER_70_324 ();
 sg13g2_fill_8 FILLER_70_362 ();
 sg13g2_fill_2 FILLER_70_375 ();
 sg13g2_fill_1 FILLER_70_412 ();
 sg13g2_fill_8 FILLER_70_416 ();
 sg13g2_fill_2 FILLER_70_424 ();
 sg13g2_fill_1 FILLER_70_426 ();
 sg13g2_fill_8 FILLER_70_436 ();
 sg13g2_fill_8 FILLER_70_444 ();
 sg13g2_fill_8 FILLER_70_452 ();
 sg13g2_fill_1 FILLER_70_460 ();
 sg13g2_fill_2 FILLER_70_466 ();
 sg13g2_fill_1 FILLER_70_468 ();
 sg13g2_fill_4 FILLER_70_494 ();
 sg13g2_fill_2 FILLER_70_498 ();
 sg13g2_fill_1 FILLER_70_500 ();
 sg13g2_fill_2 FILLER_70_534 ();
 sg13g2_fill_8 FILLER_70_540 ();
 sg13g2_fill_1 FILLER_70_548 ();
 sg13g2_fill_8 FILLER_70_555 ();
 sg13g2_fill_2 FILLER_70_563 ();
 sg13g2_fill_8 FILLER_70_591 ();
 sg13g2_fill_4 FILLER_70_599 ();
 sg13g2_fill_2 FILLER_70_603 ();
 sg13g2_fill_1 FILLER_70_605 ();
 sg13g2_fill_8 FILLER_70_631 ();
 sg13g2_fill_8 FILLER_70_639 ();
 sg13g2_fill_2 FILLER_70_647 ();
 sg13g2_fill_4 FILLER_70_654 ();
 sg13g2_fill_2 FILLER_70_658 ();
 sg13g2_fill_1 FILLER_70_660 ();
 sg13g2_fill_8 FILLER_70_673 ();
 sg13g2_fill_1 FILLER_70_681 ();
 sg13g2_fill_8 FILLER_70_687 ();
 sg13g2_fill_8 FILLER_70_695 ();
 sg13g2_fill_2 FILLER_70_703 ();
 sg13g2_fill_1 FILLER_70_705 ();
 sg13g2_fill_8 FILLER_70_727 ();
 sg13g2_fill_4 FILLER_70_735 ();
 sg13g2_fill_8 FILLER_70_744 ();
 sg13g2_fill_8 FILLER_70_752 ();
 sg13g2_fill_8 FILLER_70_760 ();
 sg13g2_fill_8 FILLER_70_768 ();
 sg13g2_fill_4 FILLER_70_776 ();
 sg13g2_fill_2 FILLER_70_780 ();
 sg13g2_fill_1 FILLER_70_782 ();
 sg13g2_fill_1 FILLER_70_795 ();
 sg13g2_fill_8 FILLER_70_813 ();
 sg13g2_fill_1 FILLER_70_821 ();
 sg13g2_fill_2 FILLER_70_827 ();
 sg13g2_fill_2 FILLER_70_843 ();
 sg13g2_fill_4 FILLER_70_851 ();
 sg13g2_fill_2 FILLER_70_855 ();
 sg13g2_fill_1 FILLER_70_882 ();
 sg13g2_fill_4 FILLER_70_930 ();
 sg13g2_fill_2 FILLER_70_971 ();
 sg13g2_fill_1 FILLER_70_973 ();
 sg13g2_fill_4 FILLER_70_1000 ();
 sg13g2_fill_2 FILLER_70_1004 ();
 sg13g2_fill_8 FILLER_70_1053 ();
 sg13g2_fill_8 FILLER_70_1061 ();
 sg13g2_fill_8 FILLER_70_1069 ();
 sg13g2_fill_8 FILLER_70_1077 ();
 sg13g2_fill_8 FILLER_70_1085 ();
 sg13g2_fill_8 FILLER_70_1093 ();
 sg13g2_fill_8 FILLER_70_1101 ();
 sg13g2_fill_8 FILLER_70_1109 ();
 sg13g2_fill_8 FILLER_70_1117 ();
 sg13g2_fill_8 FILLER_70_1125 ();
 sg13g2_fill_8 FILLER_70_1133 ();
 sg13g2_fill_8 FILLER_70_1141 ();
 sg13g2_fill_8 FILLER_70_1149 ();
 sg13g2_fill_8 FILLER_70_1157 ();
 sg13g2_fill_1 FILLER_70_1165 ();
 sg13g2_fill_8 FILLER_71_0 ();
 sg13g2_fill_8 FILLER_71_8 ();
 sg13g2_fill_2 FILLER_71_16 ();
 sg13g2_fill_1 FILLER_71_18 ();
 sg13g2_fill_4 FILLER_71_45 ();
 sg13g2_fill_1 FILLER_71_49 ();
 sg13g2_fill_4 FILLER_71_55 ();
 sg13g2_fill_2 FILLER_71_59 ();
 sg13g2_fill_1 FILLER_71_61 ();
 sg13g2_fill_2 FILLER_71_93 ();
 sg13g2_fill_1 FILLER_71_95 ();
 sg13g2_fill_8 FILLER_71_100 ();
 sg13g2_fill_4 FILLER_71_108 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_4 FILLER_71_205 ();
 sg13g2_fill_8 FILLER_71_243 ();
 sg13g2_fill_2 FILLER_71_251 ();
 sg13g2_fill_8 FILLER_71_273 ();
 sg13g2_fill_4 FILLER_71_281 ();
 sg13g2_fill_2 FILLER_71_285 ();
 sg13g2_fill_1 FILLER_71_323 ();
 sg13g2_fill_8 FILLER_71_350 ();
 sg13g2_fill_4 FILLER_71_358 ();
 sg13g2_fill_4 FILLER_71_366 ();
 sg13g2_fill_1 FILLER_71_370 ();
 sg13g2_fill_2 FILLER_71_380 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_fill_4 FILLER_71_388 ();
 sg13g2_fill_2 FILLER_71_392 ();
 sg13g2_fill_1 FILLER_71_394 ();
 sg13g2_fill_2 FILLER_71_408 ();
 sg13g2_fill_2 FILLER_71_418 ();
 sg13g2_fill_2 FILLER_71_428 ();
 sg13g2_fill_2 FILLER_71_443 ();
 sg13g2_fill_4 FILLER_71_450 ();
 sg13g2_fill_2 FILLER_71_454 ();
 sg13g2_fill_1 FILLER_71_456 ();
 sg13g2_fill_1 FILLER_71_471 ();
 sg13g2_fill_1 FILLER_71_485 ();
 sg13g2_fill_1 FILLER_71_496 ();
 sg13g2_fill_2 FILLER_71_524 ();
 sg13g2_fill_8 FILLER_71_542 ();
 sg13g2_fill_4 FILLER_71_583 ();
 sg13g2_fill_2 FILLER_71_587 ();
 sg13g2_fill_8 FILLER_71_626 ();
 sg13g2_fill_8 FILLER_71_634 ();
 sg13g2_fill_1 FILLER_71_647 ();
 sg13g2_fill_4 FILLER_71_657 ();
 sg13g2_fill_2 FILLER_71_661 ();
 sg13g2_fill_1 FILLER_71_663 ();
 sg13g2_fill_1 FILLER_71_669 ();
 sg13g2_fill_4 FILLER_71_675 ();
 sg13g2_fill_2 FILLER_71_679 ();
 sg13g2_fill_1 FILLER_71_681 ();
 sg13g2_fill_4 FILLER_71_708 ();
 sg13g2_fill_2 FILLER_71_712 ();
 sg13g2_fill_1 FILLER_71_714 ();
 sg13g2_fill_8 FILLER_71_720 ();
 sg13g2_fill_8 FILLER_71_728 ();
 sg13g2_fill_8 FILLER_71_736 ();
 sg13g2_fill_2 FILLER_71_779 ();
 sg13g2_fill_1 FILLER_71_781 ();
 sg13g2_fill_2 FILLER_71_787 ();
 sg13g2_fill_1 FILLER_71_794 ();
 sg13g2_fill_2 FILLER_71_800 ();
 sg13g2_fill_1 FILLER_71_802 ();
 sg13g2_fill_4 FILLER_71_813 ();
 sg13g2_fill_2 FILLER_71_817 ();
 sg13g2_fill_1 FILLER_71_824 ();
 sg13g2_fill_1 FILLER_71_852 ();
 sg13g2_fill_8 FILLER_71_884 ();
 sg13g2_fill_4 FILLER_71_892 ();
 sg13g2_fill_2 FILLER_71_896 ();
 sg13g2_fill_8 FILLER_71_908 ();
 sg13g2_fill_8 FILLER_71_916 ();
 sg13g2_fill_4 FILLER_71_924 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_8 FILLER_71_950 ();
 sg13g2_fill_4 FILLER_71_958 ();
 sg13g2_fill_2 FILLER_71_962 ();
 sg13g2_fill_8 FILLER_71_1021 ();
 sg13g2_fill_8 FILLER_71_1029 ();
 sg13g2_fill_8 FILLER_71_1037 ();
 sg13g2_fill_8 FILLER_71_1045 ();
 sg13g2_fill_8 FILLER_71_1053 ();
 sg13g2_fill_8 FILLER_71_1061 ();
 sg13g2_fill_8 FILLER_71_1069 ();
 sg13g2_fill_8 FILLER_71_1077 ();
 sg13g2_fill_8 FILLER_71_1085 ();
 sg13g2_fill_8 FILLER_71_1093 ();
 sg13g2_fill_8 FILLER_71_1101 ();
 sg13g2_fill_8 FILLER_71_1109 ();
 sg13g2_fill_8 FILLER_71_1117 ();
 sg13g2_fill_8 FILLER_71_1125 ();
 sg13g2_fill_8 FILLER_71_1133 ();
 sg13g2_fill_8 FILLER_71_1141 ();
 sg13g2_fill_8 FILLER_71_1149 ();
 sg13g2_fill_8 FILLER_71_1157 ();
 sg13g2_fill_1 FILLER_71_1165 ();
 sg13g2_fill_4 FILLER_72_0 ();
 sg13g2_fill_4 FILLER_72_38 ();
 sg13g2_fill_2 FILLER_72_42 ();
 sg13g2_fill_1 FILLER_72_44 ();
 sg13g2_fill_2 FILLER_72_76 ();
 sg13g2_fill_1 FILLER_72_78 ();
 sg13g2_fill_4 FILLER_72_100 ();
 sg13g2_fill_1 FILLER_72_104 ();
 sg13g2_fill_8 FILLER_72_116 ();
 sg13g2_fill_4 FILLER_72_124 ();
 sg13g2_fill_2 FILLER_72_128 ();
 sg13g2_fill_1 FILLER_72_130 ();
 sg13g2_fill_2 FILLER_72_135 ();
 sg13g2_fill_1 FILLER_72_137 ();
 sg13g2_fill_8 FILLER_72_169 ();
 sg13g2_fill_8 FILLER_72_177 ();
 sg13g2_fill_2 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_196 ();
 sg13g2_fill_8 FILLER_72_230 ();
 sg13g2_fill_8 FILLER_72_238 ();
 sg13g2_fill_2 FILLER_72_246 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_fill_1 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_303 ();
 sg13g2_fill_4 FILLER_72_319 ();
 sg13g2_fill_2 FILLER_72_323 ();
 sg13g2_fill_4 FILLER_72_331 ();
 sg13g2_fill_1 FILLER_72_335 ();
 sg13g2_fill_8 FILLER_72_345 ();
 sg13g2_fill_4 FILLER_72_353 ();
 sg13g2_fill_1 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_8 FILLER_72_377 ();
 sg13g2_fill_4 FILLER_72_385 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_fill_8 FILLER_72_395 ();
 sg13g2_fill_8 FILLER_72_403 ();
 sg13g2_fill_4 FILLER_72_411 ();
 sg13g2_fill_2 FILLER_72_415 ();
 sg13g2_fill_1 FILLER_72_422 ();
 sg13g2_fill_4 FILLER_72_427 ();
 sg13g2_fill_1 FILLER_72_431 ();
 sg13g2_fill_8 FILLER_72_440 ();
 sg13g2_fill_2 FILLER_72_448 ();
 sg13g2_fill_4 FILLER_72_455 ();
 sg13g2_fill_1 FILLER_72_459 ();
 sg13g2_fill_4 FILLER_72_487 ();
 sg13g2_fill_4 FILLER_72_494 ();
 sg13g2_fill_1 FILLER_72_498 ();
 sg13g2_fill_8 FILLER_72_504 ();
 sg13g2_fill_2 FILLER_72_512 ();
 sg13g2_fill_8 FILLER_72_519 ();
 sg13g2_fill_1 FILLER_72_527 ();
 sg13g2_fill_8 FILLER_72_544 ();
 sg13g2_fill_8 FILLER_72_552 ();
 sg13g2_fill_8 FILLER_72_560 ();
 sg13g2_fill_4 FILLER_72_568 ();
 sg13g2_fill_2 FILLER_72_576 ();
 sg13g2_fill_1 FILLER_72_610 ();
 sg13g2_fill_2 FILLER_72_616 ();
 sg13g2_fill_1 FILLER_72_618 ();
 sg13g2_fill_4 FILLER_72_645 ();
 sg13g2_fill_1 FILLER_72_649 ();
 sg13g2_fill_8 FILLER_72_675 ();
 sg13g2_fill_8 FILLER_72_683 ();
 sg13g2_fill_2 FILLER_72_691 ();
 sg13g2_fill_8 FILLER_72_699 ();
 sg13g2_fill_8 FILLER_72_707 ();
 sg13g2_fill_8 FILLER_72_715 ();
 sg13g2_fill_2 FILLER_72_723 ();
 sg13g2_fill_8 FILLER_72_745 ();
 sg13g2_fill_8 FILLER_72_753 ();
 sg13g2_fill_1 FILLER_72_761 ();
 sg13g2_fill_4 FILLER_72_766 ();
 sg13g2_fill_1 FILLER_72_770 ();
 sg13g2_fill_8 FILLER_72_776 ();
 sg13g2_fill_8 FILLER_72_784 ();
 sg13g2_fill_8 FILLER_72_792 ();
 sg13g2_fill_4 FILLER_72_806 ();
 sg13g2_fill_2 FILLER_72_817 ();
 sg13g2_fill_2 FILLER_72_826 ();
 sg13g2_fill_1 FILLER_72_828 ();
 sg13g2_fill_4 FILLER_72_859 ();
 sg13g2_fill_1 FILLER_72_863 ();
 sg13g2_fill_2 FILLER_72_870 ();
 sg13g2_fill_8 FILLER_72_897 ();
 sg13g2_fill_8 FILLER_72_905 ();
 sg13g2_fill_8 FILLER_72_913 ();
 sg13g2_fill_4 FILLER_72_921 ();
 sg13g2_fill_8 FILLER_72_933 ();
 sg13g2_fill_8 FILLER_72_941 ();
 sg13g2_fill_8 FILLER_72_949 ();
 sg13g2_fill_8 FILLER_72_957 ();
 sg13g2_fill_4 FILLER_72_965 ();
 sg13g2_fill_2 FILLER_72_969 ();
 sg13g2_fill_8 FILLER_72_981 ();
 sg13g2_fill_4 FILLER_72_989 ();
 sg13g2_fill_8 FILLER_72_1044 ();
 sg13g2_fill_8 FILLER_72_1052 ();
 sg13g2_fill_8 FILLER_72_1060 ();
 sg13g2_fill_8 FILLER_72_1068 ();
 sg13g2_fill_8 FILLER_72_1076 ();
 sg13g2_fill_8 FILLER_72_1084 ();
 sg13g2_fill_8 FILLER_72_1092 ();
 sg13g2_fill_8 FILLER_72_1100 ();
 sg13g2_fill_8 FILLER_72_1108 ();
 sg13g2_fill_8 FILLER_72_1116 ();
 sg13g2_fill_8 FILLER_72_1124 ();
 sg13g2_fill_8 FILLER_72_1132 ();
 sg13g2_fill_8 FILLER_72_1140 ();
 sg13g2_fill_8 FILLER_72_1148 ();
 sg13g2_fill_8 FILLER_72_1156 ();
 sg13g2_fill_2 FILLER_72_1164 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_57 ();
 sg13g2_fill_1 FILLER_73_64 ();
 sg13g2_fill_8 FILLER_73_132 ();
 sg13g2_fill_8 FILLER_73_140 ();
 sg13g2_fill_4 FILLER_73_148 ();
 sg13g2_fill_8 FILLER_73_178 ();
 sg13g2_fill_1 FILLER_73_186 ();
 sg13g2_fill_8 FILLER_73_239 ();
 sg13g2_fill_8 FILLER_73_247 ();
 sg13g2_fill_2 FILLER_73_281 ();
 sg13g2_fill_2 FILLER_73_299 ();
 sg13g2_fill_1 FILLER_73_301 ();
 sg13g2_fill_2 FILLER_73_312 ();
 sg13g2_fill_1 FILLER_73_324 ();
 sg13g2_fill_2 FILLER_73_328 ();
 sg13g2_fill_8 FILLER_73_337 ();
 sg13g2_fill_4 FILLER_73_345 ();
 sg13g2_fill_1 FILLER_73_349 ();
 sg13g2_fill_2 FILLER_73_356 ();
 sg13g2_fill_8 FILLER_73_371 ();
 sg13g2_fill_4 FILLER_73_387 ();
 sg13g2_fill_4 FILLER_73_396 ();
 sg13g2_fill_2 FILLER_73_400 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_8 FILLER_73_453 ();
 sg13g2_fill_8 FILLER_73_465 ();
 sg13g2_fill_8 FILLER_73_473 ();
 sg13g2_fill_4 FILLER_73_481 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_fill_8 FILLER_73_526 ();
 sg13g2_fill_1 FILLER_73_534 ();
 sg13g2_fill_8 FILLER_73_553 ();
 sg13g2_fill_2 FILLER_73_561 ();
 sg13g2_fill_2 FILLER_73_572 ();
 sg13g2_fill_1 FILLER_73_574 ();
 sg13g2_fill_2 FILLER_73_610 ();
 sg13g2_fill_4 FILLER_73_623 ();
 sg13g2_fill_1 FILLER_73_627 ();
 sg13g2_fill_8 FILLER_73_670 ();
 sg13g2_fill_2 FILLER_73_678 ();
 sg13g2_fill_1 FILLER_73_680 ();
 sg13g2_fill_1 FILLER_73_684 ();
 sg13g2_fill_8 FILLER_73_715 ();
 sg13g2_fill_1 FILLER_73_723 ();
 sg13g2_fill_4 FILLER_73_735 ();
 sg13g2_fill_1 FILLER_73_739 ();
 sg13g2_fill_4 FILLER_73_778 ();
 sg13g2_fill_1 FILLER_73_782 ();
 sg13g2_fill_4 FILLER_73_797 ();
 sg13g2_fill_2 FILLER_73_801 ();
 sg13g2_fill_4 FILLER_73_819 ();
 sg13g2_fill_8 FILLER_73_867 ();
 sg13g2_fill_8 FILLER_73_875 ();
 sg13g2_fill_8 FILLER_73_887 ();
 sg13g2_fill_8 FILLER_73_895 ();
 sg13g2_fill_4 FILLER_73_903 ();
 sg13g2_fill_4 FILLER_73_917 ();
 sg13g2_fill_8 FILLER_73_957 ();
 sg13g2_fill_2 FILLER_73_965 ();
 sg13g2_fill_1 FILLER_73_975 ();
 sg13g2_fill_8 FILLER_73_984 ();
 sg13g2_fill_8 FILLER_73_992 ();
 sg13g2_fill_8 FILLER_73_1000 ();
 sg13g2_fill_8 FILLER_73_1055 ();
 sg13g2_fill_8 FILLER_73_1063 ();
 sg13g2_fill_8 FILLER_73_1071 ();
 sg13g2_fill_8 FILLER_73_1079 ();
 sg13g2_fill_8 FILLER_73_1087 ();
 sg13g2_fill_8 FILLER_73_1095 ();
 sg13g2_fill_8 FILLER_73_1103 ();
 sg13g2_fill_8 FILLER_73_1111 ();
 sg13g2_fill_8 FILLER_73_1119 ();
 sg13g2_fill_8 FILLER_73_1127 ();
 sg13g2_fill_8 FILLER_73_1135 ();
 sg13g2_fill_8 FILLER_73_1143 ();
 sg13g2_fill_8 FILLER_73_1151 ();
 sg13g2_fill_4 FILLER_73_1159 ();
 sg13g2_fill_2 FILLER_73_1163 ();
 sg13g2_fill_1 FILLER_73_1165 ();
 sg13g2_fill_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_8 ();
 sg13g2_fill_1 FILLER_74_10 ();
 sg13g2_fill_2 FILLER_74_29 ();
 sg13g2_fill_1 FILLER_74_31 ();
 sg13g2_fill_4 FILLER_74_35 ();
 sg13g2_fill_4 FILLER_74_78 ();
 sg13g2_fill_2 FILLER_74_82 ();
 sg13g2_fill_2 FILLER_74_105 ();
 sg13g2_fill_2 FILLER_74_145 ();
 sg13g2_fill_1 FILLER_74_152 ();
 sg13g2_fill_4 FILLER_74_184 ();
 sg13g2_fill_2 FILLER_74_188 ();
 sg13g2_fill_1 FILLER_74_190 ();
 sg13g2_fill_8 FILLER_74_212 ();
 sg13g2_fill_4 FILLER_74_220 ();
 sg13g2_fill_2 FILLER_74_224 ();
 sg13g2_fill_4 FILLER_74_252 ();
 sg13g2_fill_2 FILLER_74_256 ();
 sg13g2_fill_8 FILLER_74_262 ();
 sg13g2_fill_2 FILLER_74_270 ();
 sg13g2_fill_2 FILLER_74_299 ();
 sg13g2_fill_2 FILLER_74_311 ();
 sg13g2_fill_8 FILLER_74_357 ();
 sg13g2_fill_1 FILLER_74_365 ();
 sg13g2_fill_1 FILLER_74_375 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_fill_4 FILLER_74_402 ();
 sg13g2_fill_8 FILLER_74_440 ();
 sg13g2_fill_4 FILLER_74_472 ();
 sg13g2_fill_2 FILLER_74_476 ();
 sg13g2_fill_1 FILLER_74_478 ();
 sg13g2_fill_1 FILLER_74_482 ();
 sg13g2_fill_4 FILLER_74_491 ();
 sg13g2_fill_2 FILLER_74_495 ();
 sg13g2_fill_1 FILLER_74_497 ();
 sg13g2_fill_4 FILLER_74_510 ();
 sg13g2_fill_2 FILLER_74_514 ();
 sg13g2_fill_1 FILLER_74_516 ();
 sg13g2_fill_4 FILLER_74_535 ();
 sg13g2_fill_1 FILLER_74_539 ();
 sg13g2_fill_4 FILLER_74_577 ();
 sg13g2_fill_2 FILLER_74_581 ();
 sg13g2_fill_2 FILLER_74_608 ();
 sg13g2_fill_8 FILLER_74_614 ();
 sg13g2_fill_4 FILLER_74_631 ();
 sg13g2_fill_8 FILLER_74_645 ();
 sg13g2_fill_1 FILLER_74_653 ();
 sg13g2_fill_8 FILLER_74_664 ();
 sg13g2_fill_2 FILLER_74_672 ();
 sg13g2_fill_8 FILLER_74_704 ();
 sg13g2_fill_1 FILLER_74_712 ();
 sg13g2_fill_2 FILLER_74_721 ();
 sg13g2_fill_1 FILLER_74_723 ();
 sg13g2_fill_4 FILLER_74_754 ();
 sg13g2_fill_2 FILLER_74_758 ();
 sg13g2_fill_2 FILLER_74_770 ();
 sg13g2_fill_2 FILLER_74_781 ();
 sg13g2_fill_8 FILLER_74_793 ();
 sg13g2_fill_4 FILLER_74_801 ();
 sg13g2_fill_2 FILLER_74_809 ();
 sg13g2_fill_2 FILLER_74_827 ();
 sg13g2_fill_1 FILLER_74_829 ();
 sg13g2_fill_2 FILLER_74_840 ();
 sg13g2_fill_2 FILLER_74_871 ();
 sg13g2_fill_1 FILLER_74_873 ();
 sg13g2_fill_8 FILLER_74_880 ();
 sg13g2_fill_8 FILLER_74_888 ();
 sg13g2_fill_4 FILLER_74_896 ();
 sg13g2_fill_2 FILLER_74_900 ();
 sg13g2_fill_8 FILLER_74_933 ();
 sg13g2_fill_8 FILLER_74_941 ();
 sg13g2_fill_4 FILLER_74_949 ();
 sg13g2_fill_1 FILLER_74_953 ();
 sg13g2_fill_4 FILLER_74_965 ();
 sg13g2_fill_1 FILLER_74_969 ();
 sg13g2_fill_1 FILLER_74_978 ();
 sg13g2_fill_4 FILLER_74_1005 ();
 sg13g2_fill_8 FILLER_74_1029 ();
 sg13g2_fill_8 FILLER_74_1037 ();
 sg13g2_fill_8 FILLER_74_1045 ();
 sg13g2_fill_8 FILLER_74_1053 ();
 sg13g2_fill_8 FILLER_74_1061 ();
 sg13g2_fill_8 FILLER_74_1069 ();
 sg13g2_fill_8 FILLER_74_1077 ();
 sg13g2_fill_8 FILLER_74_1085 ();
 sg13g2_fill_8 FILLER_74_1093 ();
 sg13g2_fill_8 FILLER_74_1101 ();
 sg13g2_fill_8 FILLER_74_1109 ();
 sg13g2_fill_8 FILLER_74_1117 ();
 sg13g2_fill_8 FILLER_74_1125 ();
 sg13g2_fill_8 FILLER_74_1133 ();
 sg13g2_fill_8 FILLER_74_1141 ();
 sg13g2_fill_8 FILLER_74_1149 ();
 sg13g2_fill_8 FILLER_74_1157 ();
 sg13g2_fill_1 FILLER_74_1165 ();
 sg13g2_fill_8 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_8 ();
 sg13g2_fill_8 FILLER_75_22 ();
 sg13g2_fill_2 FILLER_75_30 ();
 sg13g2_fill_4 FILLER_75_62 ();
 sg13g2_fill_2 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_73 ();
 sg13g2_fill_1 FILLER_75_75 ();
 sg13g2_fill_2 FILLER_75_87 ();
 sg13g2_fill_1 FILLER_75_89 ();
 sg13g2_fill_2 FILLER_75_150 ();
 sg13g2_fill_4 FILLER_75_161 ();
 sg13g2_fill_8 FILLER_75_174 ();
 sg13g2_fill_1 FILLER_75_182 ();
 sg13g2_fill_4 FILLER_75_186 ();
 sg13g2_fill_2 FILLER_75_190 ();
 sg13g2_fill_2 FILLER_75_200 ();
 sg13g2_fill_4 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_fill_8 FILLER_75_219 ();
 sg13g2_fill_8 FILLER_75_227 ();
 sg13g2_fill_8 FILLER_75_235 ();
 sg13g2_fill_2 FILLER_75_243 ();
 sg13g2_fill_4 FILLER_75_253 ();
 sg13g2_fill_2 FILLER_75_257 ();
 sg13g2_fill_2 FILLER_75_264 ();
 sg13g2_fill_8 FILLER_75_272 ();
 sg13g2_fill_4 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_284 ();
 sg13g2_fill_1 FILLER_75_286 ();
 sg13g2_fill_8 FILLER_75_293 ();
 sg13g2_fill_4 FILLER_75_301 ();
 sg13g2_fill_1 FILLER_75_305 ();
 sg13g2_fill_8 FILLER_75_333 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_fill_4 FILLER_75_357 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_2 FILLER_75_416 ();
 sg13g2_fill_1 FILLER_75_418 ();
 sg13g2_fill_2 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_427 ();
 sg13g2_fill_2 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_447 ();
 sg13g2_fill_2 FILLER_75_465 ();
 sg13g2_fill_4 FILLER_75_485 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_fill_1 FILLER_75_526 ();
 sg13g2_fill_8 FILLER_75_583 ();
 sg13g2_fill_4 FILLER_75_591 ();
 sg13g2_fill_2 FILLER_75_595 ();
 sg13g2_fill_1 FILLER_75_597 ();
 sg13g2_fill_4 FILLER_75_603 ();
 sg13g2_fill_2 FILLER_75_607 ();
 sg13g2_fill_8 FILLER_75_614 ();
 sg13g2_fill_8 FILLER_75_622 ();
 sg13g2_fill_2 FILLER_75_630 ();
 sg13g2_fill_1 FILLER_75_632 ();
 sg13g2_fill_2 FILLER_75_675 ();
 sg13g2_fill_1 FILLER_75_677 ();
 sg13g2_fill_4 FILLER_75_689 ();
 sg13g2_fill_8 FILLER_75_749 ();
 sg13g2_fill_8 FILLER_75_757 ();
 sg13g2_fill_1 FILLER_75_765 ();
 sg13g2_fill_8 FILLER_75_779 ();
 sg13g2_fill_4 FILLER_75_787 ();
 sg13g2_fill_2 FILLER_75_791 ();
 sg13g2_fill_8 FILLER_75_805 ();
 sg13g2_fill_2 FILLER_75_813 ();
 sg13g2_fill_2 FILLER_75_847 ();
 sg13g2_fill_8 FILLER_75_857 ();
 sg13g2_fill_1 FILLER_75_865 ();
 sg13g2_fill_8 FILLER_75_872 ();
 sg13g2_fill_8 FILLER_75_880 ();
 sg13g2_fill_1 FILLER_75_888 ();
 sg13g2_fill_8 FILLER_75_895 ();
 sg13g2_fill_8 FILLER_75_903 ();
 sg13g2_fill_4 FILLER_75_911 ();
 sg13g2_fill_1 FILLER_75_915 ();
 sg13g2_fill_4 FILLER_75_924 ();
 sg13g2_fill_4 FILLER_75_964 ();
 sg13g2_fill_1 FILLER_75_968 ();
 sg13g2_fill_8 FILLER_75_1052 ();
 sg13g2_fill_8 FILLER_75_1060 ();
 sg13g2_fill_8 FILLER_75_1068 ();
 sg13g2_fill_8 FILLER_75_1076 ();
 sg13g2_fill_8 FILLER_75_1084 ();
 sg13g2_fill_8 FILLER_75_1092 ();
 sg13g2_fill_8 FILLER_75_1100 ();
 sg13g2_fill_8 FILLER_75_1108 ();
 sg13g2_fill_8 FILLER_75_1116 ();
 sg13g2_fill_8 FILLER_75_1124 ();
 sg13g2_fill_8 FILLER_75_1132 ();
 sg13g2_fill_8 FILLER_75_1140 ();
 sg13g2_fill_8 FILLER_75_1148 ();
 sg13g2_fill_8 FILLER_75_1156 ();
 sg13g2_fill_2 FILLER_75_1164 ();
 sg13g2_fill_4 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_4 ();
 sg13g2_fill_4 FILLER_76_27 ();
 sg13g2_fill_1 FILLER_76_31 ();
 sg13g2_fill_4 FILLER_76_37 ();
 sg13g2_fill_4 FILLER_76_55 ();
 sg13g2_fill_1 FILLER_76_59 ();
 sg13g2_fill_8 FILLER_76_86 ();
 sg13g2_fill_8 FILLER_76_94 ();
 sg13g2_fill_8 FILLER_76_102 ();
 sg13g2_fill_8 FILLER_76_110 ();
 sg13g2_fill_2 FILLER_76_118 ();
 sg13g2_fill_8 FILLER_76_140 ();
 sg13g2_fill_8 FILLER_76_148 ();
 sg13g2_fill_2 FILLER_76_156 ();
 sg13g2_fill_1 FILLER_76_158 ();
 sg13g2_fill_4 FILLER_76_195 ();
 sg13g2_fill_2 FILLER_76_217 ();
 sg13g2_fill_8 FILLER_76_245 ();
 sg13g2_fill_2 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_255 ();
 sg13g2_fill_4 FILLER_76_282 ();
 sg13g2_fill_8 FILLER_76_299 ();
 sg13g2_fill_1 FILLER_76_310 ();
 sg13g2_fill_2 FILLER_76_318 ();
 sg13g2_fill_8 FILLER_76_332 ();
 sg13g2_fill_8 FILLER_76_340 ();
 sg13g2_fill_8 FILLER_76_348 ();
 sg13g2_fill_8 FILLER_76_356 ();
 sg13g2_fill_8 FILLER_76_364 ();
 sg13g2_fill_8 FILLER_76_372 ();
 sg13g2_fill_4 FILLER_76_380 ();
 sg13g2_fill_2 FILLER_76_384 ();
 sg13g2_fill_1 FILLER_76_386 ();
 sg13g2_fill_4 FILLER_76_400 ();
 sg13g2_fill_1 FILLER_76_436 ();
 sg13g2_fill_2 FILLER_76_445 ();
 sg13g2_fill_1 FILLER_76_447 ();
 sg13g2_fill_8 FILLER_76_452 ();
 sg13g2_fill_2 FILLER_76_460 ();
 sg13g2_fill_1 FILLER_76_462 ();
 sg13g2_fill_1 FILLER_76_477 ();
 sg13g2_fill_1 FILLER_76_484 ();
 sg13g2_fill_2 FILLER_76_506 ();
 sg13g2_fill_1 FILLER_76_508 ();
 sg13g2_fill_4 FILLER_76_513 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_fill_2 FILLER_76_530 ();
 sg13g2_fill_4 FILLER_76_537 ();
 sg13g2_fill_2 FILLER_76_541 ();
 sg13g2_fill_1 FILLER_76_543 ();
 sg13g2_fill_8 FILLER_76_548 ();
 sg13g2_fill_4 FILLER_76_556 ();
 sg13g2_fill_8 FILLER_76_566 ();
 sg13g2_fill_8 FILLER_76_583 ();
 sg13g2_fill_1 FILLER_76_591 ();
 sg13g2_fill_1 FILLER_76_602 ();
 sg13g2_fill_1 FILLER_76_629 ();
 sg13g2_fill_8 FILLER_76_635 ();
 sg13g2_fill_8 FILLER_76_643 ();
 sg13g2_fill_4 FILLER_76_651 ();
 sg13g2_fill_2 FILLER_76_660 ();
 sg13g2_fill_4 FILLER_76_667 ();
 sg13g2_fill_2 FILLER_76_681 ();
 sg13g2_fill_1 FILLER_76_683 ();
 sg13g2_fill_8 FILLER_76_705 ();
 sg13g2_fill_2 FILLER_76_713 ();
 sg13g2_fill_4 FILLER_76_719 ();
 sg13g2_fill_2 FILLER_76_723 ();
 sg13g2_fill_8 FILLER_76_729 ();
 sg13g2_fill_8 FILLER_76_737 ();
 sg13g2_fill_8 FILLER_76_745 ();
 sg13g2_fill_4 FILLER_76_753 ();
 sg13g2_fill_8 FILLER_76_771 ();
 sg13g2_fill_8 FILLER_76_779 ();
 sg13g2_fill_8 FILLER_76_809 ();
 sg13g2_fill_8 FILLER_76_817 ();
 sg13g2_fill_1 FILLER_76_825 ();
 sg13g2_fill_1 FILLER_76_838 ();
 sg13g2_fill_8 FILLER_76_849 ();
 sg13g2_fill_8 FILLER_76_857 ();
 sg13g2_fill_1 FILLER_76_865 ();
 sg13g2_fill_8 FILLER_76_883 ();
 sg13g2_fill_8 FILLER_76_891 ();
 sg13g2_fill_8 FILLER_76_899 ();
 sg13g2_fill_2 FILLER_76_912 ();
 sg13g2_fill_1 FILLER_76_914 ();
 sg13g2_fill_8 FILLER_76_920 ();
 sg13g2_fill_2 FILLER_76_928 ();
 sg13g2_fill_8 FILLER_76_987 ();
 sg13g2_fill_2 FILLER_76_995 ();
 sg13g2_fill_4 FILLER_76_1008 ();
 sg13g2_fill_2 FILLER_76_1012 ();
 sg13g2_fill_1 FILLER_76_1014 ();
 sg13g2_fill_8 FILLER_76_1041 ();
 sg13g2_fill_8 FILLER_76_1049 ();
 sg13g2_fill_8 FILLER_76_1057 ();
 sg13g2_fill_8 FILLER_76_1065 ();
 sg13g2_fill_8 FILLER_76_1073 ();
 sg13g2_fill_8 FILLER_76_1081 ();
 sg13g2_fill_8 FILLER_76_1089 ();
 sg13g2_fill_8 FILLER_76_1097 ();
 sg13g2_fill_8 FILLER_76_1105 ();
 sg13g2_fill_8 FILLER_76_1113 ();
 sg13g2_fill_8 FILLER_76_1121 ();
 sg13g2_fill_8 FILLER_76_1129 ();
 sg13g2_fill_8 FILLER_76_1137 ();
 sg13g2_fill_8 FILLER_76_1145 ();
 sg13g2_fill_8 FILLER_76_1153 ();
 sg13g2_fill_4 FILLER_76_1161 ();
 sg13g2_fill_1 FILLER_76_1165 ();
 sg13g2_fill_4 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_32 ();
 sg13g2_fill_2 FILLER_77_64 ();
 sg13g2_fill_1 FILLER_77_66 ();
 sg13g2_fill_8 FILLER_77_71 ();
 sg13g2_fill_8 FILLER_77_100 ();
 sg13g2_fill_8 FILLER_77_108 ();
 sg13g2_fill_8 FILLER_77_116 ();
 sg13g2_fill_2 FILLER_77_124 ();
 sg13g2_fill_1 FILLER_77_126 ();
 sg13g2_fill_8 FILLER_77_137 ();
 sg13g2_fill_4 FILLER_77_145 ();
 sg13g2_fill_2 FILLER_77_149 ();
 sg13g2_fill_1 FILLER_77_151 ();
 sg13g2_fill_2 FILLER_77_162 ();
 sg13g2_fill_2 FILLER_77_174 ();
 sg13g2_fill_1 FILLER_77_176 ();
 sg13g2_fill_4 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_184 ();
 sg13g2_fill_2 FILLER_77_215 ();
 sg13g2_fill_1 FILLER_77_217 ();
 sg13g2_fill_8 FILLER_77_243 ();
 sg13g2_fill_2 FILLER_77_251 ();
 sg13g2_fill_1 FILLER_77_253 ();
 sg13g2_fill_8 FILLER_77_267 ();
 sg13g2_fill_8 FILLER_77_275 ();
 sg13g2_fill_8 FILLER_77_283 ();
 sg13g2_fill_8 FILLER_77_291 ();
 sg13g2_fill_4 FILLER_77_299 ();
 sg13g2_fill_8 FILLER_77_325 ();
 sg13g2_fill_8 FILLER_77_333 ();
 sg13g2_fill_8 FILLER_77_341 ();
 sg13g2_fill_4 FILLER_77_349 ();
 sg13g2_fill_1 FILLER_77_358 ();
 sg13g2_fill_8 FILLER_77_364 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_fill_1 FILLER_77_379 ();
 sg13g2_fill_8 FILLER_77_385 ();
 sg13g2_fill_8 FILLER_77_393 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_fill_1 FILLER_77_409 ();
 sg13g2_fill_8 FILLER_77_427 ();
 sg13g2_fill_8 FILLER_77_435 ();
 sg13g2_fill_8 FILLER_77_443 ();
 sg13g2_fill_4 FILLER_77_451 ();
 sg13g2_fill_1 FILLER_77_455 ();
 sg13g2_fill_4 FILLER_77_462 ();
 sg13g2_fill_2 FILLER_77_466 ();
 sg13g2_fill_1 FILLER_77_473 ();
 sg13g2_fill_8 FILLER_77_480 ();
 sg13g2_fill_4 FILLER_77_488 ();
 sg13g2_fill_2 FILLER_77_492 ();
 sg13g2_fill_2 FILLER_77_500 ();
 sg13g2_fill_8 FILLER_77_507 ();
 sg13g2_fill_8 FILLER_77_515 ();
 sg13g2_fill_8 FILLER_77_523 ();
 sg13g2_fill_4 FILLER_77_531 ();
 sg13g2_fill_2 FILLER_77_535 ();
 sg13g2_fill_8 FILLER_77_544 ();
 sg13g2_fill_8 FILLER_77_552 ();
 sg13g2_fill_8 FILLER_77_560 ();
 sg13g2_fill_4 FILLER_77_568 ();
 sg13g2_fill_1 FILLER_77_572 ();
 sg13g2_fill_1 FILLER_77_591 ();
 sg13g2_fill_4 FILLER_77_606 ();
 sg13g2_fill_1 FILLER_77_610 ();
 sg13g2_fill_4 FILLER_77_637 ();
 sg13g2_fill_4 FILLER_77_646 ();
 sg13g2_fill_2 FILLER_77_650 ();
 sg13g2_fill_1 FILLER_77_652 ();
 sg13g2_fill_8 FILLER_77_658 ();
 sg13g2_fill_1 FILLER_77_666 ();
 sg13g2_fill_8 FILLER_77_714 ();
 sg13g2_fill_2 FILLER_77_722 ();
 sg13g2_fill_8 FILLER_77_732 ();
 sg13g2_fill_4 FILLER_77_740 ();
 sg13g2_fill_2 FILLER_77_744 ();
 sg13g2_fill_1 FILLER_77_746 ();
 sg13g2_fill_8 FILLER_77_773 ();
 sg13g2_fill_2 FILLER_77_781 ();
 sg13g2_fill_2 FILLER_77_791 ();
 sg13g2_fill_1 FILLER_77_799 ();
 sg13g2_fill_8 FILLER_77_808 ();
 sg13g2_fill_4 FILLER_77_816 ();
 sg13g2_fill_2 FILLER_77_820 ();
 sg13g2_fill_1 FILLER_77_822 ();
 sg13g2_fill_8 FILLER_77_840 ();
 sg13g2_fill_8 FILLER_77_848 ();
 sg13g2_fill_2 FILLER_77_856 ();
 sg13g2_fill_4 FILLER_77_898 ();
 sg13g2_fill_2 FILLER_77_902 ();
 sg13g2_fill_8 FILLER_77_949 ();
 sg13g2_fill_8 FILLER_77_957 ();
 sg13g2_fill_8 FILLER_77_965 ();
 sg13g2_fill_8 FILLER_77_973 ();
 sg13g2_fill_8 FILLER_77_981 ();
 sg13g2_fill_8 FILLER_77_989 ();
 sg13g2_fill_8 FILLER_77_997 ();
 sg13g2_fill_8 FILLER_77_1005 ();
 sg13g2_fill_8 FILLER_77_1013 ();
 sg13g2_fill_8 FILLER_77_1021 ();
 sg13g2_fill_8 FILLER_77_1029 ();
 sg13g2_fill_8 FILLER_77_1037 ();
 sg13g2_fill_8 FILLER_77_1045 ();
 sg13g2_fill_8 FILLER_77_1053 ();
 sg13g2_fill_8 FILLER_77_1061 ();
 sg13g2_fill_8 FILLER_77_1069 ();
 sg13g2_fill_8 FILLER_77_1077 ();
 sg13g2_fill_8 FILLER_77_1085 ();
 sg13g2_fill_8 FILLER_77_1093 ();
 sg13g2_fill_8 FILLER_77_1101 ();
 sg13g2_fill_8 FILLER_77_1109 ();
 sg13g2_fill_8 FILLER_77_1117 ();
 sg13g2_fill_8 FILLER_77_1125 ();
 sg13g2_fill_8 FILLER_77_1133 ();
 sg13g2_fill_8 FILLER_77_1141 ();
 sg13g2_fill_8 FILLER_77_1149 ();
 sg13g2_fill_8 FILLER_77_1157 ();
 sg13g2_fill_1 FILLER_77_1165 ();
 sg13g2_fill_8 FILLER_78_0 ();
 sg13g2_fill_4 FILLER_78_8 ();
 sg13g2_fill_2 FILLER_78_12 ();
 sg13g2_fill_1 FILLER_78_23 ();
 sg13g2_fill_2 FILLER_78_50 ();
 sg13g2_fill_1 FILLER_78_52 ();
 sg13g2_fill_2 FILLER_78_69 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_fill_4 FILLER_78_76 ();
 sg13g2_fill_8 FILLER_78_101 ();
 sg13g2_fill_4 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_113 ();
 sg13g2_fill_1 FILLER_78_115 ();
 sg13g2_fill_4 FILLER_78_147 ();
 sg13g2_fill_2 FILLER_78_177 ();
 sg13g2_fill_8 FILLER_78_223 ();
 sg13g2_fill_8 FILLER_78_231 ();
 sg13g2_fill_8 FILLER_78_239 ();
 sg13g2_fill_4 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_251 ();
 sg13g2_fill_8 FILLER_78_261 ();
 sg13g2_fill_2 FILLER_78_269 ();
 sg13g2_fill_2 FILLER_78_297 ();
 sg13g2_fill_1 FILLER_78_299 ();
 sg13g2_fill_4 FILLER_78_315 ();
 sg13g2_fill_1 FILLER_78_329 ();
 sg13g2_fill_4 FILLER_78_335 ();
 sg13g2_fill_4 FILLER_78_344 ();
 sg13g2_fill_1 FILLER_78_348 ();
 sg13g2_fill_1 FILLER_78_364 ();
 sg13g2_fill_8 FILLER_78_386 ();
 sg13g2_fill_8 FILLER_78_394 ();
 sg13g2_fill_4 FILLER_78_402 ();
 sg13g2_fill_1 FILLER_78_406 ();
 sg13g2_fill_8 FILLER_78_415 ();
 sg13g2_fill_4 FILLER_78_423 ();
 sg13g2_fill_2 FILLER_78_427 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_fill_4 FILLER_78_436 ();
 sg13g2_fill_1 FILLER_78_440 ();
 sg13g2_fill_4 FILLER_78_447 ();
 sg13g2_fill_2 FILLER_78_451 ();
 sg13g2_fill_2 FILLER_78_472 ();
 sg13g2_fill_1 FILLER_78_474 ();
 sg13g2_fill_4 FILLER_78_485 ();
 sg13g2_fill_2 FILLER_78_489 ();
 sg13g2_fill_2 FILLER_78_496 ();
 sg13g2_fill_1 FILLER_78_498 ();
 sg13g2_fill_4 FILLER_78_515 ();
 sg13g2_fill_4 FILLER_78_562 ();
 sg13g2_fill_2 FILLER_78_589 ();
 sg13g2_fill_1 FILLER_78_601 ();
 sg13g2_fill_8 FILLER_78_608 ();
 sg13g2_fill_4 FILLER_78_616 ();
 sg13g2_fill_8 FILLER_78_625 ();
 sg13g2_fill_8 FILLER_78_633 ();
 sg13g2_fill_8 FILLER_78_641 ();
 sg13g2_fill_4 FILLER_78_649 ();
 sg13g2_fill_8 FILLER_78_672 ();
 sg13g2_fill_2 FILLER_78_680 ();
 sg13g2_fill_4 FILLER_78_709 ();
 sg13g2_fill_1 FILLER_78_723 ();
 sg13g2_fill_1 FILLER_78_754 ();
 sg13g2_fill_2 FILLER_78_802 ();
 sg13g2_fill_8 FILLER_78_834 ();
 sg13g2_fill_8 FILLER_78_842 ();
 sg13g2_fill_1 FILLER_78_850 ();
 sg13g2_fill_8 FILLER_78_897 ();
 sg13g2_fill_8 FILLER_78_905 ();
 sg13g2_fill_8 FILLER_78_913 ();
 sg13g2_fill_4 FILLER_78_921 ();
 sg13g2_fill_1 FILLER_78_930 ();
 sg13g2_fill_8 FILLER_78_964 ();
 sg13g2_fill_8 FILLER_78_972 ();
 sg13g2_fill_8 FILLER_78_980 ();
 sg13g2_fill_8 FILLER_78_988 ();
 sg13g2_fill_8 FILLER_78_1032 ();
 sg13g2_fill_8 FILLER_78_1040 ();
 sg13g2_fill_8 FILLER_78_1048 ();
 sg13g2_fill_8 FILLER_78_1056 ();
 sg13g2_fill_8 FILLER_78_1064 ();
 sg13g2_fill_8 FILLER_78_1072 ();
 sg13g2_fill_8 FILLER_78_1080 ();
 sg13g2_fill_8 FILLER_78_1088 ();
 sg13g2_fill_8 FILLER_78_1096 ();
 sg13g2_fill_8 FILLER_78_1104 ();
 sg13g2_fill_8 FILLER_78_1112 ();
 sg13g2_fill_8 FILLER_78_1120 ();
 sg13g2_fill_8 FILLER_78_1128 ();
 sg13g2_fill_8 FILLER_78_1136 ();
 sg13g2_fill_8 FILLER_78_1144 ();
 sg13g2_fill_8 FILLER_78_1152 ();
 sg13g2_fill_4 FILLER_78_1160 ();
 sg13g2_fill_2 FILLER_78_1164 ();
 sg13g2_fill_8 FILLER_79_0 ();
 sg13g2_fill_4 FILLER_79_8 ();
 sg13g2_fill_1 FILLER_79_12 ();
 sg13g2_fill_8 FILLER_79_21 ();
 sg13g2_fill_4 FILLER_79_29 ();
 sg13g2_fill_1 FILLER_79_33 ();
 sg13g2_fill_2 FILLER_79_64 ();
 sg13g2_fill_1 FILLER_79_66 ();
 sg13g2_fill_2 FILLER_79_72 ();
 sg13g2_fill_1 FILLER_79_74 ();
 sg13g2_fill_8 FILLER_79_107 ();
 sg13g2_fill_1 FILLER_79_115 ();
 sg13g2_fill_2 FILLER_79_122 ();
 sg13g2_fill_1 FILLER_79_124 ();
 sg13g2_fill_2 FILLER_79_151 ();
 sg13g2_fill_2 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_213 ();
 sg13g2_fill_4 FILLER_79_235 ();
 sg13g2_fill_2 FILLER_79_239 ();
 sg13g2_fill_4 FILLER_79_272 ();
 sg13g2_fill_1 FILLER_79_276 ();
 sg13g2_fill_1 FILLER_79_308 ();
 sg13g2_fill_2 FILLER_79_312 ();
 sg13g2_fill_1 FILLER_79_314 ();
 sg13g2_fill_4 FILLER_79_400 ();
 sg13g2_fill_2 FILLER_79_404 ();
 sg13g2_fill_1 FILLER_79_426 ();
 sg13g2_fill_2 FILLER_79_432 ();
 sg13g2_fill_2 FILLER_79_478 ();
 sg13g2_fill_1 FILLER_79_480 ();
 sg13g2_fill_2 FILLER_79_495 ();
 sg13g2_fill_1 FILLER_79_497 ();
 sg13g2_fill_4 FILLER_79_520 ();
 sg13g2_fill_2 FILLER_79_524 ();
 sg13g2_fill_1 FILLER_79_526 ();
 sg13g2_fill_1 FILLER_79_537 ();
 sg13g2_fill_8 FILLER_79_546 ();
 sg13g2_fill_2 FILLER_79_588 ();
 sg13g2_fill_8 FILLER_79_603 ();
 sg13g2_fill_2 FILLER_79_611 ();
 sg13g2_fill_1 FILLER_79_613 ();
 sg13g2_fill_1 FILLER_79_650 ();
 sg13g2_fill_8 FILLER_79_666 ();
 sg13g2_fill_4 FILLER_79_674 ();
 sg13g2_fill_2 FILLER_79_678 ();
 sg13g2_fill_1 FILLER_79_680 ();
 sg13g2_fill_1 FILLER_79_705 ();
 sg13g2_fill_8 FILLER_79_740 ();
 sg13g2_fill_2 FILLER_79_748 ();
 sg13g2_fill_8 FILLER_79_762 ();
 sg13g2_fill_8 FILLER_79_770 ();
 sg13g2_fill_8 FILLER_79_778 ();
 sg13g2_fill_1 FILLER_79_800 ();
 sg13g2_fill_4 FILLER_79_831 ();
 sg13g2_fill_1 FILLER_79_835 ();
 sg13g2_fill_2 FILLER_79_841 ();
 sg13g2_fill_1 FILLER_79_843 ();
 sg13g2_fill_8 FILLER_79_905 ();
 sg13g2_fill_4 FILLER_79_913 ();
 sg13g2_fill_2 FILLER_79_935 ();
 sg13g2_fill_4 FILLER_79_945 ();
 sg13g2_fill_2 FILLER_79_959 ();
 sg13g2_fill_4 FILLER_79_966 ();
 sg13g2_fill_2 FILLER_79_970 ();
 sg13g2_fill_8 FILLER_79_998 ();
 sg13g2_fill_8 FILLER_79_1032 ();
 sg13g2_fill_8 FILLER_79_1040 ();
 sg13g2_fill_8 FILLER_79_1048 ();
 sg13g2_fill_8 FILLER_79_1056 ();
 sg13g2_fill_8 FILLER_79_1064 ();
 sg13g2_fill_8 FILLER_79_1072 ();
 sg13g2_fill_8 FILLER_79_1080 ();
 sg13g2_fill_8 FILLER_79_1088 ();
 sg13g2_fill_8 FILLER_79_1096 ();
 sg13g2_fill_8 FILLER_79_1104 ();
 sg13g2_fill_8 FILLER_79_1112 ();
 sg13g2_fill_8 FILLER_79_1120 ();
 sg13g2_fill_8 FILLER_79_1128 ();
 sg13g2_fill_8 FILLER_79_1136 ();
 sg13g2_fill_8 FILLER_79_1144 ();
 sg13g2_fill_8 FILLER_79_1152 ();
 sg13g2_fill_4 FILLER_79_1160 ();
 sg13g2_fill_2 FILLER_79_1164 ();
 sg13g2_fill_4 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_4 ();
 sg13g2_fill_4 FILLER_80_32 ();
 sg13g2_fill_1 FILLER_80_36 ();
 sg13g2_fill_4 FILLER_80_68 ();
 sg13g2_fill_2 FILLER_80_72 ();
 sg13g2_fill_2 FILLER_80_102 ();
 sg13g2_fill_1 FILLER_80_104 ();
 sg13g2_fill_1 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_129 ();
 sg13g2_fill_4 FILLER_80_156 ();
 sg13g2_fill_2 FILLER_80_160 ();
 sg13g2_fill_1 FILLER_80_162 ();
 sg13g2_fill_4 FILLER_80_174 ();
 sg13g2_fill_1 FILLER_80_178 ();
 sg13g2_fill_4 FILLER_80_200 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_8 FILLER_80_231 ();
 sg13g2_fill_4 FILLER_80_239 ();
 sg13g2_fill_4 FILLER_80_248 ();
 sg13g2_fill_2 FILLER_80_252 ();
 sg13g2_fill_1 FILLER_80_254 ();
 sg13g2_fill_8 FILLER_80_273 ();
 sg13g2_fill_1 FILLER_80_281 ();
 sg13g2_fill_1 FILLER_80_308 ();
 sg13g2_fill_8 FILLER_80_334 ();
 sg13g2_fill_4 FILLER_80_342 ();
 sg13g2_fill_2 FILLER_80_346 ();
 sg13g2_fill_4 FILLER_80_363 ();
 sg13g2_fill_1 FILLER_80_367 ();
 sg13g2_fill_2 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_383 ();
 sg13g2_fill_2 FILLER_80_393 ();
 sg13g2_fill_8 FILLER_80_405 ();
 sg13g2_fill_4 FILLER_80_413 ();
 sg13g2_fill_2 FILLER_80_422 ();
 sg13g2_fill_2 FILLER_80_436 ();
 sg13g2_fill_2 FILLER_80_442 ();
 sg13g2_fill_2 FILLER_80_452 ();
 sg13g2_fill_1 FILLER_80_454 ();
 sg13g2_fill_8 FILLER_80_459 ();
 sg13g2_fill_4 FILLER_80_467 ();
 sg13g2_fill_2 FILLER_80_471 ();
 sg13g2_fill_1 FILLER_80_473 ();
 sg13g2_fill_8 FILLER_80_484 ();
 sg13g2_fill_4 FILLER_80_492 ();
 sg13g2_fill_1 FILLER_80_496 ();
 sg13g2_fill_1 FILLER_80_513 ();
 sg13g2_fill_4 FILLER_80_538 ();
 sg13g2_fill_2 FILLER_80_542 ();
 sg13g2_fill_1 FILLER_80_577 ();
 sg13g2_fill_8 FILLER_80_585 ();
 sg13g2_fill_8 FILLER_80_593 ();
 sg13g2_fill_8 FILLER_80_601 ();
 sg13g2_fill_8 FILLER_80_609 ();
 sg13g2_fill_2 FILLER_80_617 ();
 sg13g2_fill_1 FILLER_80_619 ();
 sg13g2_fill_8 FILLER_80_633 ();
 sg13g2_fill_8 FILLER_80_641 ();
 sg13g2_fill_4 FILLER_80_660 ();
 sg13g2_fill_8 FILLER_80_670 ();
 sg13g2_fill_2 FILLER_80_678 ();
 sg13g2_fill_8 FILLER_80_706 ();
 sg13g2_fill_8 FILLER_80_714 ();
 sg13g2_fill_1 FILLER_80_722 ();
 sg13g2_fill_1 FILLER_80_735 ();
 sg13g2_fill_8 FILLER_80_752 ();
 sg13g2_fill_8 FILLER_80_760 ();
 sg13g2_fill_8 FILLER_80_768 ();
 sg13g2_fill_8 FILLER_80_776 ();
 sg13g2_fill_4 FILLER_80_784 ();
 sg13g2_fill_1 FILLER_80_788 ();
 sg13g2_fill_8 FILLER_80_818 ();
 sg13g2_fill_8 FILLER_80_834 ();
 sg13g2_fill_8 FILLER_80_842 ();
 sg13g2_fill_1 FILLER_80_850 ();
 sg13g2_fill_1 FILLER_80_856 ();
 sg13g2_fill_2 FILLER_80_861 ();
 sg13g2_fill_1 FILLER_80_867 ();
 sg13g2_fill_2 FILLER_80_876 ();
 sg13g2_fill_2 FILLER_80_921 ();
 sg13g2_fill_1 FILLER_80_923 ();
 sg13g2_fill_1 FILLER_80_936 ();
 sg13g2_fill_2 FILLER_80_967 ();
 sg13g2_fill_8 FILLER_80_1042 ();
 sg13g2_fill_8 FILLER_80_1050 ();
 sg13g2_fill_8 FILLER_80_1058 ();
 sg13g2_fill_8 FILLER_80_1066 ();
 sg13g2_fill_8 FILLER_80_1074 ();
 sg13g2_fill_8 FILLER_80_1082 ();
 sg13g2_fill_8 FILLER_80_1090 ();
 sg13g2_fill_8 FILLER_80_1098 ();
 sg13g2_fill_8 FILLER_80_1106 ();
 sg13g2_fill_8 FILLER_80_1114 ();
 sg13g2_fill_8 FILLER_80_1122 ();
 sg13g2_fill_8 FILLER_80_1130 ();
 sg13g2_fill_8 FILLER_80_1138 ();
 sg13g2_fill_8 FILLER_80_1146 ();
 sg13g2_fill_8 FILLER_80_1154 ();
 sg13g2_fill_4 FILLER_80_1162 ();
 sg13g2_fill_4 FILLER_81_0 ();
 sg13g2_fill_2 FILLER_81_4 ();
 sg13g2_fill_8 FILLER_81_27 ();
 sg13g2_fill_8 FILLER_81_35 ();
 sg13g2_fill_4 FILLER_81_43 ();
 sg13g2_fill_1 FILLER_81_47 ();
 sg13g2_fill_4 FILLER_81_53 ();
 sg13g2_fill_2 FILLER_81_57 ();
 sg13g2_fill_1 FILLER_81_59 ();
 sg13g2_fill_8 FILLER_81_107 ();
 sg13g2_fill_4 FILLER_81_115 ();
 sg13g2_fill_2 FILLER_81_119 ();
 sg13g2_fill_1 FILLER_81_129 ();
 sg13g2_fill_4 FILLER_81_143 ();
 sg13g2_fill_2 FILLER_81_147 ();
 sg13g2_fill_1 FILLER_81_149 ();
 sg13g2_fill_8 FILLER_81_153 ();
 sg13g2_fill_8 FILLER_81_161 ();
 sg13g2_fill_8 FILLER_81_169 ();
 sg13g2_fill_8 FILLER_81_177 ();
 sg13g2_fill_2 FILLER_81_185 ();
 sg13g2_fill_4 FILLER_81_192 ();
 sg13g2_fill_4 FILLER_81_233 ();
 sg13g2_fill_2 FILLER_81_237 ();
 sg13g2_fill_1 FILLER_81_239 ();
 sg13g2_fill_8 FILLER_81_269 ();
 sg13g2_fill_8 FILLER_81_277 ();
 sg13g2_fill_4 FILLER_81_285 ();
 sg13g2_fill_2 FILLER_81_289 ();
 sg13g2_fill_1 FILLER_81_316 ();
 sg13g2_fill_2 FILLER_81_323 ();
 sg13g2_fill_1 FILLER_81_356 ();
 sg13g2_fill_8 FILLER_81_363 ();
 sg13g2_fill_8 FILLER_81_371 ();
 sg13g2_fill_1 FILLER_81_379 ();
 sg13g2_fill_8 FILLER_81_385 ();
 sg13g2_fill_2 FILLER_81_393 ();
 sg13g2_fill_8 FILLER_81_400 ();
 sg13g2_fill_4 FILLER_81_421 ();
 sg13g2_fill_2 FILLER_81_425 ();
 sg13g2_fill_1 FILLER_81_427 ();
 sg13g2_fill_8 FILLER_81_442 ();
 sg13g2_fill_8 FILLER_81_450 ();
 sg13g2_fill_4 FILLER_81_458 ();
 sg13g2_fill_1 FILLER_81_462 ();
 sg13g2_fill_8 FILLER_81_467 ();
 sg13g2_fill_8 FILLER_81_489 ();
 sg13g2_fill_4 FILLER_81_497 ();
 sg13g2_fill_2 FILLER_81_501 ();
 sg13g2_fill_1 FILLER_81_503 ();
 sg13g2_fill_8 FILLER_81_508 ();
 sg13g2_fill_2 FILLER_81_516 ();
 sg13g2_fill_1 FILLER_81_518 ();
 sg13g2_fill_8 FILLER_81_525 ();
 sg13g2_fill_8 FILLER_81_533 ();
 sg13g2_fill_4 FILLER_81_541 ();
 sg13g2_fill_1 FILLER_81_545 ();
 sg13g2_fill_4 FILLER_81_572 ();
 sg13g2_fill_8 FILLER_81_676 ();
 sg13g2_fill_2 FILLER_81_684 ();
 sg13g2_fill_4 FILLER_81_712 ();
 sg13g2_fill_2 FILLER_81_716 ();
 sg13g2_fill_1 FILLER_81_749 ();
 sg13g2_fill_8 FILLER_81_814 ();
 sg13g2_fill_8 FILLER_81_822 ();
 sg13g2_fill_4 FILLER_81_834 ();
 sg13g2_fill_4 FILLER_81_846 ();
 sg13g2_fill_2 FILLER_81_850 ();
 sg13g2_fill_1 FILLER_81_852 ();
 sg13g2_fill_2 FILLER_81_883 ();
 sg13g2_fill_1 FILLER_81_885 ();
 sg13g2_fill_4 FILLER_81_892 ();
 sg13g2_fill_2 FILLER_81_896 ();
 sg13g2_fill_4 FILLER_81_960 ();
 sg13g2_fill_2 FILLER_81_964 ();
 sg13g2_fill_1 FILLER_81_966 ();
 sg13g2_fill_8 FILLER_81_995 ();
 sg13g2_fill_2 FILLER_81_1003 ();
 sg13g2_fill_1 FILLER_81_1005 ();
 sg13g2_fill_8 FILLER_81_1016 ();
 sg13g2_fill_8 FILLER_81_1024 ();
 sg13g2_fill_8 FILLER_81_1032 ();
 sg13g2_fill_8 FILLER_81_1040 ();
 sg13g2_fill_8 FILLER_81_1048 ();
 sg13g2_fill_8 FILLER_81_1056 ();
 sg13g2_fill_8 FILLER_81_1064 ();
 sg13g2_fill_8 FILLER_81_1072 ();
 sg13g2_fill_8 FILLER_81_1080 ();
 sg13g2_fill_8 FILLER_81_1088 ();
 sg13g2_fill_8 FILLER_81_1096 ();
 sg13g2_fill_8 FILLER_81_1104 ();
 sg13g2_fill_8 FILLER_81_1112 ();
 sg13g2_fill_8 FILLER_81_1120 ();
 sg13g2_fill_8 FILLER_81_1128 ();
 sg13g2_fill_8 FILLER_81_1136 ();
 sg13g2_fill_8 FILLER_81_1144 ();
 sg13g2_fill_8 FILLER_81_1152 ();
 sg13g2_fill_4 FILLER_81_1160 ();
 sg13g2_fill_2 FILLER_81_1164 ();
 sg13g2_fill_8 FILLER_82_0 ();
 sg13g2_fill_1 FILLER_82_8 ();
 sg13g2_fill_8 FILLER_82_35 ();
 sg13g2_fill_8 FILLER_82_43 ();
 sg13g2_fill_8 FILLER_82_51 ();
 sg13g2_fill_4 FILLER_82_59 ();
 sg13g2_fill_2 FILLER_82_63 ();
 sg13g2_fill_1 FILLER_82_65 ();
 sg13g2_fill_2 FILLER_82_71 ();
 sg13g2_fill_2 FILLER_82_76 ();
 sg13g2_fill_1 FILLER_82_78 ();
 sg13g2_fill_8 FILLER_82_105 ();
 sg13g2_fill_1 FILLER_82_113 ();
 sg13g2_fill_1 FILLER_82_139 ();
 sg13g2_fill_1 FILLER_82_166 ();
 sg13g2_fill_8 FILLER_82_193 ();
 sg13g2_fill_2 FILLER_82_201 ();
 sg13g2_fill_1 FILLER_82_203 ();
 sg13g2_fill_8 FILLER_82_207 ();
 sg13g2_fill_8 FILLER_82_215 ();
 sg13g2_fill_8 FILLER_82_223 ();
 sg13g2_fill_8 FILLER_82_231 ();
 sg13g2_fill_2 FILLER_82_239 ();
 sg13g2_fill_1 FILLER_82_241 ();
 sg13g2_fill_8 FILLER_82_250 ();
 sg13g2_fill_8 FILLER_82_258 ();
 sg13g2_fill_8 FILLER_82_266 ();
 sg13g2_fill_8 FILLER_82_274 ();
 sg13g2_fill_2 FILLER_82_282 ();
 sg13g2_fill_1 FILLER_82_310 ();
 sg13g2_fill_1 FILLER_82_342 ();
 sg13g2_fill_2 FILLER_82_348 ();
 sg13g2_fill_1 FILLER_82_350 ();
 sg13g2_fill_8 FILLER_82_377 ();
 sg13g2_fill_8 FILLER_82_385 ();
 sg13g2_fill_1 FILLER_82_393 ();
 sg13g2_fill_1 FILLER_82_403 ();
 sg13g2_fill_4 FILLER_82_410 ();
 sg13g2_fill_1 FILLER_82_414 ();
 sg13g2_fill_8 FILLER_82_447 ();
 sg13g2_fill_2 FILLER_82_455 ();
 sg13g2_fill_1 FILLER_82_457 ();
 sg13g2_fill_8 FILLER_82_488 ();
 sg13g2_fill_2 FILLER_82_496 ();
 sg13g2_fill_1 FILLER_82_498 ();
 sg13g2_fill_8 FILLER_82_513 ();
 sg13g2_fill_8 FILLER_82_521 ();
 sg13g2_fill_8 FILLER_82_529 ();
 sg13g2_fill_8 FILLER_82_537 ();
 sg13g2_fill_8 FILLER_82_545 ();
 sg13g2_fill_2 FILLER_82_553 ();
 sg13g2_fill_1 FILLER_82_555 ();
 sg13g2_fill_4 FILLER_82_563 ();
 sg13g2_fill_2 FILLER_82_567 ();
 sg13g2_fill_1 FILLER_82_569 ();
 sg13g2_fill_8 FILLER_82_575 ();
 sg13g2_fill_4 FILLER_82_583 ();
 sg13g2_fill_2 FILLER_82_612 ();
 sg13g2_fill_1 FILLER_82_614 ();
 sg13g2_fill_8 FILLER_82_641 ();
 sg13g2_fill_4 FILLER_82_654 ();
 sg13g2_fill_1 FILLER_82_658 ();
 sg13g2_fill_8 FILLER_82_664 ();
 sg13g2_fill_8 FILLER_82_672 ();
 sg13g2_fill_8 FILLER_82_680 ();
 sg13g2_fill_8 FILLER_82_688 ();
 sg13g2_fill_8 FILLER_82_696 ();
 sg13g2_fill_4 FILLER_82_704 ();
 sg13g2_fill_1 FILLER_82_708 ();
 sg13g2_fill_1 FILLER_82_770 ();
 sg13g2_fill_8 FILLER_82_801 ();
 sg13g2_fill_8 FILLER_82_809 ();
 sg13g2_fill_8 FILLER_82_817 ();
 sg13g2_fill_2 FILLER_82_825 ();
 sg13g2_fill_1 FILLER_82_831 ();
 sg13g2_fill_1 FILLER_82_837 ();
 sg13g2_fill_8 FILLER_82_854 ();
 sg13g2_fill_4 FILLER_82_862 ();
 sg13g2_fill_1 FILLER_82_866 ();
 sg13g2_fill_8 FILLER_82_871 ();
 sg13g2_fill_8 FILLER_82_879 ();
 sg13g2_fill_8 FILLER_82_955 ();
 sg13g2_fill_8 FILLER_82_963 ();
 sg13g2_fill_8 FILLER_82_971 ();
 sg13g2_fill_8 FILLER_82_979 ();
 sg13g2_fill_8 FILLER_82_987 ();
 sg13g2_fill_8 FILLER_82_995 ();
 sg13g2_fill_8 FILLER_82_1039 ();
 sg13g2_fill_8 FILLER_82_1047 ();
 sg13g2_fill_8 FILLER_82_1055 ();
 sg13g2_fill_8 FILLER_82_1063 ();
 sg13g2_fill_8 FILLER_82_1071 ();
 sg13g2_fill_8 FILLER_82_1079 ();
 sg13g2_fill_8 FILLER_82_1087 ();
 sg13g2_fill_8 FILLER_82_1095 ();
 sg13g2_fill_8 FILLER_82_1103 ();
 sg13g2_fill_8 FILLER_82_1111 ();
 sg13g2_fill_8 FILLER_82_1119 ();
 sg13g2_fill_8 FILLER_82_1127 ();
 sg13g2_fill_8 FILLER_82_1135 ();
 sg13g2_fill_8 FILLER_82_1143 ();
 sg13g2_fill_8 FILLER_82_1151 ();
 sg13g2_fill_4 FILLER_82_1159 ();
 sg13g2_fill_2 FILLER_82_1163 ();
 sg13g2_fill_1 FILLER_82_1165 ();
 sg13g2_fill_8 FILLER_83_0 ();
 sg13g2_fill_8 FILLER_83_8 ();
 sg13g2_fill_4 FILLER_83_16 ();
 sg13g2_fill_2 FILLER_83_20 ();
 sg13g2_fill_8 FILLER_83_30 ();
 sg13g2_fill_8 FILLER_83_38 ();
 sg13g2_fill_2 FILLER_83_46 ();
 sg13g2_fill_1 FILLER_83_48 ();
 sg13g2_fill_2 FILLER_83_57 ();
 sg13g2_fill_1 FILLER_83_85 ();
 sg13g2_fill_8 FILLER_83_91 ();
 sg13g2_fill_4 FILLER_83_99 ();
 sg13g2_fill_2 FILLER_83_103 ();
 sg13g2_fill_1 FILLER_83_105 ();
 sg13g2_fill_4 FILLER_83_114 ();
 sg13g2_fill_8 FILLER_83_170 ();
 sg13g2_fill_2 FILLER_83_178 ();
 sg13g2_fill_8 FILLER_83_185 ();
 sg13g2_fill_8 FILLER_83_193 ();
 sg13g2_fill_8 FILLER_83_201 ();
 sg13g2_fill_4 FILLER_83_209 ();
 sg13g2_fill_1 FILLER_83_213 ();
 sg13g2_fill_4 FILLER_83_219 ();
 sg13g2_fill_1 FILLER_83_223 ();
 sg13g2_fill_8 FILLER_83_235 ();
 sg13g2_fill_8 FILLER_83_243 ();
 sg13g2_fill_8 FILLER_83_251 ();
 sg13g2_fill_8 FILLER_83_259 ();
 sg13g2_fill_2 FILLER_83_267 ();
 sg13g2_fill_8 FILLER_83_277 ();
 sg13g2_fill_8 FILLER_83_285 ();
 sg13g2_fill_8 FILLER_83_293 ();
 sg13g2_fill_8 FILLER_83_301 ();
 sg13g2_fill_2 FILLER_83_341 ();
 sg13g2_fill_2 FILLER_83_349 ();
 sg13g2_fill_1 FILLER_83_351 ();
 sg13g2_fill_1 FILLER_83_428 ();
 sg13g2_fill_8 FILLER_83_455 ();
 sg13g2_fill_8 FILLER_83_463 ();
 sg13g2_fill_4 FILLER_83_471 ();
 sg13g2_fill_2 FILLER_83_475 ();
 sg13g2_fill_1 FILLER_83_477 ();
 sg13g2_fill_8 FILLER_83_507 ();
 sg13g2_fill_4 FILLER_83_540 ();
 sg13g2_fill_1 FILLER_83_544 ();
 sg13g2_fill_8 FILLER_83_578 ();
 sg13g2_fill_4 FILLER_83_586 ();
 sg13g2_fill_2 FILLER_83_590 ();
 sg13g2_fill_1 FILLER_83_592 ();
 sg13g2_fill_4 FILLER_83_625 ();
 sg13g2_fill_1 FILLER_83_629 ();
 sg13g2_fill_4 FILLER_83_656 ();
 sg13g2_fill_8 FILLER_83_691 ();
 sg13g2_fill_8 FILLER_83_699 ();
 sg13g2_fill_1 FILLER_83_707 ();
 sg13g2_fill_8 FILLER_83_754 ();
 sg13g2_fill_8 FILLER_83_773 ();
 sg13g2_fill_8 FILLER_83_781 ();
 sg13g2_fill_4 FILLER_83_789 ();
 sg13g2_fill_1 FILLER_83_793 ();
 sg13g2_fill_8 FILLER_83_807 ();
 sg13g2_fill_4 FILLER_83_815 ();
 sg13g2_fill_1 FILLER_83_819 ();
 sg13g2_fill_2 FILLER_83_825 ();
 sg13g2_fill_1 FILLER_83_827 ();
 sg13g2_fill_8 FILLER_83_854 ();
 sg13g2_fill_8 FILLER_83_862 ();
 sg13g2_fill_4 FILLER_83_870 ();
 sg13g2_fill_8 FILLER_83_879 ();
 sg13g2_fill_1 FILLER_83_887 ();
 sg13g2_fill_4 FILLER_83_894 ();
 sg13g2_fill_2 FILLER_83_898 ();
 sg13g2_fill_1 FILLER_83_900 ();
 sg13g2_fill_2 FILLER_83_946 ();
 sg13g2_fill_4 FILLER_83_974 ();
 sg13g2_fill_2 FILLER_83_978 ();
 sg13g2_fill_1 FILLER_83_980 ();
 sg13g2_fill_4 FILLER_83_1007 ();
 sg13g2_fill_2 FILLER_83_1011 ();
 sg13g2_fill_8 FILLER_83_1050 ();
 sg13g2_fill_8 FILLER_83_1058 ();
 sg13g2_fill_8 FILLER_83_1066 ();
 sg13g2_fill_8 FILLER_83_1074 ();
 sg13g2_fill_8 FILLER_83_1082 ();
 sg13g2_fill_8 FILLER_83_1090 ();
 sg13g2_fill_8 FILLER_83_1098 ();
 sg13g2_fill_8 FILLER_83_1106 ();
 sg13g2_fill_8 FILLER_83_1114 ();
 sg13g2_fill_8 FILLER_83_1122 ();
 sg13g2_fill_8 FILLER_83_1130 ();
 sg13g2_fill_8 FILLER_83_1138 ();
 sg13g2_fill_8 FILLER_83_1146 ();
 sg13g2_fill_8 FILLER_83_1154 ();
 sg13g2_fill_4 FILLER_83_1162 ();
 sg13g2_fill_4 FILLER_84_0 ();
 sg13g2_fill_1 FILLER_84_4 ();
 sg13g2_fill_2 FILLER_84_20 ();
 sg13g2_fill_8 FILLER_84_27 ();
 sg13g2_fill_8 FILLER_84_35 ();
 sg13g2_fill_8 FILLER_84_43 ();
 sg13g2_fill_1 FILLER_84_51 ();
 sg13g2_fill_8 FILLER_84_56 ();
 sg13g2_fill_1 FILLER_84_64 ();
 sg13g2_fill_4 FILLER_84_70 ();
 sg13g2_fill_2 FILLER_84_99 ();
 sg13g2_fill_2 FILLER_84_131 ();
 sg13g2_fill_1 FILLER_84_133 ();
 sg13g2_fill_1 FILLER_84_139 ();
 sg13g2_fill_2 FILLER_84_145 ();
 sg13g2_fill_8 FILLER_84_150 ();
 sg13g2_fill_8 FILLER_84_158 ();
 sg13g2_fill_8 FILLER_84_166 ();
 sg13g2_fill_8 FILLER_84_182 ();
 sg13g2_fill_8 FILLER_84_190 ();
 sg13g2_fill_8 FILLER_84_198 ();
 sg13g2_fill_4 FILLER_84_206 ();
 sg13g2_fill_2 FILLER_84_240 ();
 sg13g2_fill_8 FILLER_84_272 ();
 sg13g2_fill_4 FILLER_84_280 ();
 sg13g2_fill_2 FILLER_84_284 ();
 sg13g2_fill_1 FILLER_84_286 ();
 sg13g2_fill_8 FILLER_84_300 ();
 sg13g2_fill_4 FILLER_84_308 ();
 sg13g2_fill_4 FILLER_84_337 ();
 sg13g2_fill_1 FILLER_84_341 ();
 sg13g2_fill_8 FILLER_84_367 ();
 sg13g2_fill_8 FILLER_84_375 ();
 sg13g2_fill_1 FILLER_84_400 ();
 sg13g2_fill_8 FILLER_84_442 ();
 sg13g2_fill_2 FILLER_84_450 ();
 sg13g2_fill_8 FILLER_84_492 ();
 sg13g2_fill_8 FILLER_84_500 ();
 sg13g2_fill_8 FILLER_84_508 ();
 sg13g2_fill_8 FILLER_84_542 ();
 sg13g2_fill_2 FILLER_84_550 ();
 sg13g2_fill_8 FILLER_84_578 ();
 sg13g2_fill_8 FILLER_84_586 ();
 sg13g2_fill_1 FILLER_84_594 ();
 sg13g2_fill_4 FILLER_84_602 ();
 sg13g2_fill_2 FILLER_84_606 ();
 sg13g2_fill_1 FILLER_84_608 ();
 sg13g2_fill_8 FILLER_84_615 ();
 sg13g2_fill_8 FILLER_84_623 ();
 sg13g2_fill_4 FILLER_84_631 ();
 sg13g2_fill_8 FILLER_84_666 ();
 sg13g2_fill_4 FILLER_84_674 ();
 sg13g2_fill_2 FILLER_84_678 ();
 sg13g2_fill_8 FILLER_84_710 ();
 sg13g2_fill_4 FILLER_84_718 ();
 sg13g2_fill_2 FILLER_84_726 ();
 sg13g2_fill_1 FILLER_84_728 ();
 sg13g2_fill_2 FILLER_84_735 ();
 sg13g2_fill_8 FILLER_84_741 ();
 sg13g2_fill_8 FILLER_84_749 ();
 sg13g2_fill_8 FILLER_84_778 ();
 sg13g2_fill_8 FILLER_84_786 ();
 sg13g2_fill_4 FILLER_84_794 ();
 sg13g2_fill_2 FILLER_84_798 ();
 sg13g2_fill_1 FILLER_84_815 ();
 sg13g2_fill_1 FILLER_84_846 ();
 sg13g2_fill_1 FILLER_84_855 ();
 sg13g2_fill_8 FILLER_84_886 ();
 sg13g2_fill_8 FILLER_84_894 ();
 sg13g2_fill_2 FILLER_84_902 ();
 sg13g2_fill_1 FILLER_84_904 ();
 sg13g2_fill_2 FILLER_84_919 ();
 sg13g2_fill_4 FILLER_84_931 ();
 sg13g2_fill_2 FILLER_84_935 ();
 sg13g2_fill_4 FILLER_84_973 ();
 sg13g2_fill_8 FILLER_84_1024 ();
 sg13g2_fill_8 FILLER_84_1032 ();
 sg13g2_fill_8 FILLER_84_1040 ();
 sg13g2_fill_8 FILLER_84_1048 ();
 sg13g2_fill_8 FILLER_84_1056 ();
 sg13g2_fill_8 FILLER_84_1064 ();
 sg13g2_fill_8 FILLER_84_1072 ();
 sg13g2_fill_8 FILLER_84_1080 ();
 sg13g2_fill_8 FILLER_84_1088 ();
 sg13g2_fill_8 FILLER_84_1096 ();
 sg13g2_fill_8 FILLER_84_1104 ();
 sg13g2_fill_8 FILLER_84_1112 ();
 sg13g2_fill_8 FILLER_84_1120 ();
 sg13g2_fill_8 FILLER_84_1128 ();
 sg13g2_fill_8 FILLER_84_1136 ();
 sg13g2_fill_8 FILLER_84_1144 ();
 sg13g2_fill_8 FILLER_84_1152 ();
 sg13g2_fill_4 FILLER_84_1160 ();
 sg13g2_fill_2 FILLER_84_1164 ();
 sg13g2_fill_2 FILLER_85_0 ();
 sg13g2_fill_1 FILLER_85_2 ();
 sg13g2_fill_4 FILLER_85_18 ();
 sg13g2_fill_2 FILLER_85_27 ();
 sg13g2_fill_2 FILLER_85_37 ();
 sg13g2_fill_1 FILLER_85_39 ();
 sg13g2_fill_8 FILLER_85_65 ();
 sg13g2_fill_8 FILLER_85_73 ();
 sg13g2_fill_4 FILLER_85_81 ();
 sg13g2_fill_2 FILLER_85_85 ();
 sg13g2_fill_4 FILLER_85_100 ();
 sg13g2_fill_2 FILLER_85_104 ();
 sg13g2_fill_8 FILLER_85_111 ();
 sg13g2_fill_8 FILLER_85_119 ();
 sg13g2_fill_8 FILLER_85_127 ();
 sg13g2_fill_8 FILLER_85_135 ();
 sg13g2_fill_8 FILLER_85_143 ();
 sg13g2_fill_8 FILLER_85_151 ();
 sg13g2_fill_8 FILLER_85_159 ();
 sg13g2_fill_8 FILLER_85_167 ();
 sg13g2_fill_1 FILLER_85_175 ();
 sg13g2_fill_4 FILLER_85_216 ();
 sg13g2_fill_2 FILLER_85_220 ();
 sg13g2_fill_8 FILLER_85_266 ();
 sg13g2_fill_2 FILLER_85_274 ();
 sg13g2_fill_1 FILLER_85_276 ();
 sg13g2_fill_1 FILLER_85_352 ();
 sg13g2_fill_8 FILLER_85_358 ();
 sg13g2_fill_8 FILLER_85_366 ();
 sg13g2_fill_4 FILLER_85_374 ();
 sg13g2_fill_4 FILLER_85_386 ();
 sg13g2_fill_2 FILLER_85_390 ();
 sg13g2_fill_1 FILLER_85_392 ();
 sg13g2_fill_1 FILLER_85_408 ();
 sg13g2_fill_4 FILLER_85_431 ();
 sg13g2_fill_1 FILLER_85_435 ();
 sg13g2_fill_8 FILLER_85_450 ();
 sg13g2_fill_8 FILLER_85_458 ();
 sg13g2_fill_2 FILLER_85_466 ();
 sg13g2_fill_8 FILLER_85_478 ();
 sg13g2_fill_4 FILLER_85_486 ();
 sg13g2_fill_1 FILLER_85_490 ();
 sg13g2_fill_8 FILLER_85_504 ();
 sg13g2_fill_4 FILLER_85_512 ();
 sg13g2_fill_8 FILLER_85_532 ();
 sg13g2_fill_8 FILLER_85_540 ();
 sg13g2_fill_8 FILLER_85_548 ();
 sg13g2_fill_8 FILLER_85_556 ();
 sg13g2_fill_4 FILLER_85_564 ();
 sg13g2_fill_2 FILLER_85_568 ();
 sg13g2_fill_1 FILLER_85_614 ();
 sg13g2_fill_8 FILLER_85_629 ();
 sg13g2_fill_4 FILLER_85_637 ();
 sg13g2_fill_1 FILLER_85_641 ();
 sg13g2_fill_4 FILLER_85_647 ();
 sg13g2_fill_4 FILLER_85_656 ();
 sg13g2_fill_1 FILLER_85_660 ();
 sg13g2_fill_8 FILLER_85_666 ();
 sg13g2_fill_2 FILLER_85_674 ();
 sg13g2_fill_8 FILLER_85_701 ();
 sg13g2_fill_4 FILLER_85_709 ();
 sg13g2_fill_8 FILLER_85_751 ();
 sg13g2_fill_2 FILLER_85_759 ();
 sg13g2_fill_1 FILLER_85_761 ();
 sg13g2_fill_8 FILLER_85_777 ();
 sg13g2_fill_8 FILLER_85_785 ();
 sg13g2_fill_4 FILLER_85_793 ();
 sg13g2_fill_2 FILLER_85_797 ();
 sg13g2_fill_1 FILLER_85_799 ();
 sg13g2_fill_2 FILLER_85_810 ();
 sg13g2_fill_2 FILLER_85_837 ();
 sg13g2_fill_8 FILLER_85_887 ();
 sg13g2_fill_8 FILLER_85_895 ();
 sg13g2_fill_8 FILLER_85_903 ();
 sg13g2_fill_8 FILLER_85_911 ();
 sg13g2_fill_8 FILLER_85_919 ();
 sg13g2_fill_8 FILLER_85_927 ();
 sg13g2_fill_8 FILLER_85_935 ();
 sg13g2_fill_2 FILLER_85_943 ();
 sg13g2_fill_1 FILLER_85_945 ();
 sg13g2_fill_2 FILLER_85_956 ();
 sg13g2_fill_1 FILLER_85_977 ();
 sg13g2_fill_8 FILLER_85_998 ();
 sg13g2_fill_8 FILLER_85_1006 ();
 sg13g2_fill_8 FILLER_85_1014 ();
 sg13g2_fill_8 FILLER_85_1022 ();
 sg13g2_fill_8 FILLER_85_1030 ();
 sg13g2_fill_8 FILLER_85_1038 ();
 sg13g2_fill_8 FILLER_85_1046 ();
 sg13g2_fill_8 FILLER_85_1054 ();
 sg13g2_fill_8 FILLER_85_1062 ();
 sg13g2_fill_8 FILLER_85_1070 ();
 sg13g2_fill_8 FILLER_85_1078 ();
 sg13g2_fill_8 FILLER_85_1086 ();
 sg13g2_fill_8 FILLER_85_1094 ();
 sg13g2_fill_8 FILLER_85_1102 ();
 sg13g2_fill_8 FILLER_85_1110 ();
 sg13g2_fill_8 FILLER_85_1118 ();
 sg13g2_fill_8 FILLER_85_1126 ();
 sg13g2_fill_8 FILLER_85_1134 ();
 sg13g2_fill_8 FILLER_85_1142 ();
 sg13g2_fill_8 FILLER_85_1150 ();
 sg13g2_fill_8 FILLER_85_1158 ();
 sg13g2_fill_8 FILLER_86_0 ();
 sg13g2_fill_2 FILLER_86_8 ();
 sg13g2_fill_2 FILLER_86_37 ();
 sg13g2_fill_8 FILLER_86_59 ();
 sg13g2_fill_4 FILLER_86_67 ();
 sg13g2_fill_2 FILLER_86_71 ();
 sg13g2_fill_1 FILLER_86_73 ();
 sg13g2_fill_1 FILLER_86_102 ();
 sg13g2_fill_2 FILLER_86_111 ();
 sg13g2_fill_4 FILLER_86_128 ();
 sg13g2_fill_2 FILLER_86_132 ();
 sg13g2_fill_1 FILLER_86_134 ();
 sg13g2_fill_4 FILLER_86_150 ();
 sg13g2_fill_2 FILLER_86_154 ();
 sg13g2_fill_2 FILLER_86_161 ();
 sg13g2_fill_1 FILLER_86_163 ();
 sg13g2_fill_2 FILLER_86_174 ();
 sg13g2_fill_4 FILLER_86_250 ();
 sg13g2_fill_2 FILLER_86_254 ();
 sg13g2_fill_1 FILLER_86_256 ();
 sg13g2_fill_2 FILLER_86_288 ();
 sg13g2_fill_1 FILLER_86_290 ();
 sg13g2_fill_2 FILLER_86_296 ();
 sg13g2_fill_1 FILLER_86_303 ();
 sg13g2_fill_2 FILLER_86_324 ();
 sg13g2_fill_4 FILLER_86_343 ();
 sg13g2_fill_4 FILLER_86_361 ();
 sg13g2_fill_2 FILLER_86_365 ();
 sg13g2_fill_1 FILLER_86_407 ();
 sg13g2_fill_1 FILLER_86_419 ();
 sg13g2_fill_1 FILLER_86_433 ();
 sg13g2_fill_2 FILLER_86_438 ();
 sg13g2_fill_8 FILLER_86_464 ();
 sg13g2_fill_8 FILLER_86_472 ();
 sg13g2_fill_4 FILLER_86_480 ();
 sg13g2_fill_1 FILLER_86_484 ();
 sg13g2_fill_1 FILLER_86_501 ();
 sg13g2_fill_1 FILLER_86_538 ();
 sg13g2_fill_8 FILLER_86_544 ();
 sg13g2_fill_4 FILLER_86_552 ();
 sg13g2_fill_1 FILLER_86_556 ();
 sg13g2_fill_1 FILLER_86_571 ();
 sg13g2_fill_4 FILLER_86_609 ();
 sg13g2_fill_1 FILLER_86_613 ();
 sg13g2_fill_2 FILLER_86_644 ();
 sg13g2_fill_1 FILLER_86_651 ();
 sg13g2_fill_8 FILLER_86_657 ();
 sg13g2_fill_8 FILLER_86_665 ();
 sg13g2_fill_8 FILLER_86_673 ();
 sg13g2_fill_4 FILLER_86_681 ();
 sg13g2_fill_1 FILLER_86_685 ();
 sg13g2_fill_2 FILLER_86_713 ();
 sg13g2_fill_2 FILLER_86_726 ();
 sg13g2_fill_8 FILLER_86_742 ();
 sg13g2_fill_1 FILLER_86_755 ();
 sg13g2_fill_4 FILLER_86_761 ();
 sg13g2_fill_1 FILLER_86_765 ();
 sg13g2_fill_4 FILLER_86_806 ();
 sg13g2_fill_2 FILLER_86_810 ();
 sg13g2_fill_1 FILLER_86_812 ();
 sg13g2_fill_8 FILLER_86_858 ();
 sg13g2_fill_4 FILLER_86_866 ();
 sg13g2_fill_2 FILLER_86_870 ();
 sg13g2_fill_1 FILLER_86_872 ();
 sg13g2_fill_4 FILLER_86_881 ();
 sg13g2_fill_2 FILLER_86_885 ();
 sg13g2_fill_8 FILLER_86_899 ();
 sg13g2_fill_2 FILLER_86_907 ();
 sg13g2_fill_8 FILLER_86_917 ();
 sg13g2_fill_8 FILLER_86_925 ();
 sg13g2_fill_8 FILLER_86_933 ();
 sg13g2_fill_4 FILLER_86_951 ();
 sg13g2_fill_2 FILLER_86_955 ();
 sg13g2_fill_1 FILLER_86_957 ();
 sg13g2_fill_8 FILLER_86_983 ();
 sg13g2_fill_8 FILLER_86_991 ();
 sg13g2_fill_4 FILLER_86_999 ();
 sg13g2_fill_1 FILLER_86_1003 ();
 sg13g2_fill_8 FILLER_86_1038 ();
 sg13g2_fill_8 FILLER_86_1046 ();
 sg13g2_fill_8 FILLER_86_1054 ();
 sg13g2_fill_8 FILLER_86_1062 ();
 sg13g2_fill_8 FILLER_86_1070 ();
 sg13g2_fill_8 FILLER_86_1078 ();
 sg13g2_fill_8 FILLER_86_1086 ();
 sg13g2_fill_8 FILLER_86_1094 ();
 sg13g2_fill_8 FILLER_86_1102 ();
 sg13g2_fill_8 FILLER_86_1110 ();
 sg13g2_fill_8 FILLER_86_1118 ();
 sg13g2_fill_8 FILLER_86_1126 ();
 sg13g2_fill_8 FILLER_86_1134 ();
 sg13g2_fill_8 FILLER_86_1142 ();
 sg13g2_fill_8 FILLER_86_1150 ();
 sg13g2_fill_8 FILLER_86_1158 ();
 sg13g2_fill_8 FILLER_87_0 ();
 sg13g2_fill_8 FILLER_87_23 ();
 sg13g2_fill_4 FILLER_87_48 ();
 sg13g2_fill_2 FILLER_87_52 ();
 sg13g2_fill_8 FILLER_87_62 ();
 sg13g2_fill_8 FILLER_87_70 ();
 sg13g2_fill_4 FILLER_87_103 ();
 sg13g2_fill_1 FILLER_87_107 ();
 sg13g2_fill_4 FILLER_87_138 ();
 sg13g2_fill_2 FILLER_87_172 ();
 sg13g2_fill_8 FILLER_87_204 ();
 sg13g2_fill_4 FILLER_87_212 ();
 sg13g2_fill_2 FILLER_87_216 ();
 sg13g2_fill_1 FILLER_87_218 ();
 sg13g2_fill_8 FILLER_87_224 ();
 sg13g2_fill_4 FILLER_87_232 ();
 sg13g2_fill_4 FILLER_87_245 ();
 sg13g2_fill_2 FILLER_87_249 ();
 sg13g2_fill_2 FILLER_87_256 ();
 sg13g2_fill_4 FILLER_87_271 ();
 sg13g2_fill_2 FILLER_87_275 ();
 sg13g2_fill_4 FILLER_87_286 ();
 sg13g2_fill_4 FILLER_87_298 ();
 sg13g2_fill_2 FILLER_87_344 ();
 sg13g2_fill_2 FILLER_87_376 ();
 sg13g2_fill_1 FILLER_87_378 ();
 sg13g2_fill_1 FILLER_87_409 ();
 sg13g2_fill_2 FILLER_87_429 ();
 sg13g2_fill_2 FILLER_87_461 ();
 sg13g2_fill_1 FILLER_87_463 ();
 sg13g2_fill_4 FILLER_87_508 ();
 sg13g2_fill_1 FILLER_87_512 ();
 sg13g2_fill_2 FILLER_87_539 ();
 sg13g2_fill_1 FILLER_87_541 ();
 sg13g2_fill_2 FILLER_87_580 ();
 sg13g2_fill_1 FILLER_87_582 ();
 sg13g2_fill_8 FILLER_87_680 ();
 sg13g2_fill_2 FILLER_87_688 ();
 sg13g2_fill_2 FILLER_87_709 ();
 sg13g2_fill_1 FILLER_87_737 ();
 sg13g2_fill_8 FILLER_87_743 ();
 sg13g2_fill_8 FILLER_87_751 ();
 sg13g2_fill_8 FILLER_87_759 ();
 sg13g2_fill_8 FILLER_87_767 ();
 sg13g2_fill_8 FILLER_87_775 ();
 sg13g2_fill_8 FILLER_87_783 ();
 sg13g2_fill_2 FILLER_87_791 ();
 sg13g2_fill_8 FILLER_87_815 ();
 sg13g2_fill_1 FILLER_87_823 ();
 sg13g2_fill_1 FILLER_87_833 ();
 sg13g2_fill_8 FILLER_87_853 ();
 sg13g2_fill_8 FILLER_87_861 ();
 sg13g2_fill_4 FILLER_87_869 ();
 sg13g2_fill_2 FILLER_87_873 ();
 sg13g2_fill_4 FILLER_87_905 ();
 sg13g2_fill_8 FILLER_87_956 ();
 sg13g2_fill_8 FILLER_87_964 ();
 sg13g2_fill_4 FILLER_87_972 ();
 sg13g2_fill_1 FILLER_87_976 ();
 sg13g2_fill_8 FILLER_87_987 ();
 sg13g2_fill_4 FILLER_87_995 ();
 sg13g2_fill_2 FILLER_87_999 ();
 sg13g2_fill_1 FILLER_87_1001 ();
 sg13g2_fill_8 FILLER_87_1038 ();
 sg13g2_fill_8 FILLER_87_1046 ();
 sg13g2_fill_8 FILLER_87_1054 ();
 sg13g2_fill_8 FILLER_87_1062 ();
 sg13g2_fill_8 FILLER_87_1070 ();
 sg13g2_fill_8 FILLER_87_1078 ();
 sg13g2_fill_8 FILLER_87_1086 ();
 sg13g2_fill_8 FILLER_87_1094 ();
 sg13g2_fill_8 FILLER_87_1102 ();
 sg13g2_fill_8 FILLER_87_1110 ();
 sg13g2_fill_8 FILLER_87_1118 ();
 sg13g2_fill_8 FILLER_87_1126 ();
 sg13g2_fill_8 FILLER_87_1134 ();
 sg13g2_fill_8 FILLER_87_1142 ();
 sg13g2_fill_8 FILLER_87_1150 ();
 sg13g2_fill_8 FILLER_87_1158 ();
 sg13g2_fill_8 FILLER_88_0 ();
 sg13g2_fill_4 FILLER_88_18 ();
 sg13g2_fill_8 FILLER_88_27 ();
 sg13g2_fill_8 FILLER_88_35 ();
 sg13g2_fill_8 FILLER_88_43 ();
 sg13g2_fill_4 FILLER_88_51 ();
 sg13g2_fill_1 FILLER_88_55 ();
 sg13g2_fill_8 FILLER_88_68 ();
 sg13g2_fill_4 FILLER_88_76 ();
 sg13g2_fill_2 FILLER_88_80 ();
 sg13g2_fill_2 FILLER_88_87 ();
 sg13g2_fill_1 FILLER_88_89 ();
 sg13g2_fill_4 FILLER_88_100 ();
 sg13g2_fill_2 FILLER_88_104 ();
 sg13g2_fill_1 FILLER_88_106 ();
 sg13g2_fill_8 FILLER_88_112 ();
 sg13g2_fill_2 FILLER_88_125 ();
 sg13g2_fill_2 FILLER_88_136 ();
 sg13g2_fill_4 FILLER_88_148 ();
 sg13g2_fill_2 FILLER_88_152 ();
 sg13g2_fill_2 FILLER_88_159 ();
 sg13g2_fill_1 FILLER_88_161 ();
 sg13g2_fill_2 FILLER_88_172 ();
 sg13g2_fill_8 FILLER_88_204 ();
 sg13g2_fill_1 FILLER_88_212 ();
 sg13g2_fill_2 FILLER_88_218 ();
 sg13g2_fill_1 FILLER_88_225 ();
 sg13g2_fill_1 FILLER_88_236 ();
 sg13g2_fill_2 FILLER_88_247 ();
 sg13g2_fill_2 FILLER_88_274 ();
 sg13g2_fill_2 FILLER_88_288 ();
 sg13g2_fill_1 FILLER_88_290 ();
 sg13g2_fill_4 FILLER_88_296 ();
 sg13g2_fill_2 FILLER_88_300 ();
 sg13g2_fill_2 FILLER_88_307 ();
 sg13g2_fill_2 FILLER_88_319 ();
 sg13g2_fill_1 FILLER_88_329 ();
 sg13g2_fill_8 FILLER_88_335 ();
 sg13g2_fill_4 FILLER_88_343 ();
 sg13g2_fill_4 FILLER_88_384 ();
 sg13g2_fill_1 FILLER_88_388 ();
 sg13g2_fill_2 FILLER_88_411 ();
 sg13g2_fill_2 FILLER_88_432 ();
 sg13g2_fill_8 FILLER_88_438 ();
 sg13g2_fill_4 FILLER_88_446 ();
 sg13g2_fill_2 FILLER_88_450 ();
 sg13g2_fill_8 FILLER_88_461 ();
 sg13g2_fill_8 FILLER_88_469 ();
 sg13g2_fill_1 FILLER_88_477 ();
 sg13g2_fill_8 FILLER_88_494 ();
 sg13g2_fill_8 FILLER_88_502 ();
 sg13g2_fill_2 FILLER_88_510 ();
 sg13g2_fill_1 FILLER_88_512 ();
 sg13g2_fill_8 FILLER_88_539 ();
 sg13g2_fill_8 FILLER_88_547 ();
 sg13g2_fill_8 FILLER_88_571 ();
 sg13g2_fill_8 FILLER_88_579 ();
 sg13g2_fill_8 FILLER_88_587 ();
 sg13g2_fill_4 FILLER_88_595 ();
 sg13g2_fill_1 FILLER_88_599 ();
 sg13g2_fill_8 FILLER_88_606 ();
 sg13g2_fill_8 FILLER_88_674 ();
 sg13g2_fill_4 FILLER_88_682 ();
 sg13g2_fill_1 FILLER_88_686 ();
 sg13g2_fill_2 FILLER_88_699 ();
 sg13g2_fill_8 FILLER_88_714 ();
 sg13g2_fill_2 FILLER_88_722 ();
 sg13g2_fill_2 FILLER_88_737 ();
 sg13g2_fill_8 FILLER_88_752 ();
 sg13g2_fill_1 FILLER_88_760 ();
 sg13g2_fill_8 FILLER_88_796 ();
 sg13g2_fill_8 FILLER_88_804 ();
 sg13g2_fill_8 FILLER_88_812 ();
 sg13g2_fill_2 FILLER_88_820 ();
 sg13g2_fill_1 FILLER_88_822 ();
 sg13g2_fill_4 FILLER_88_833 ();
 sg13g2_fill_1 FILLER_88_837 ();
 sg13g2_fill_8 FILLER_88_852 ();
 sg13g2_fill_8 FILLER_88_860 ();
 sg13g2_fill_2 FILLER_88_868 ();
 sg13g2_fill_4 FILLER_88_895 ();
 sg13g2_fill_8 FILLER_88_969 ();
 sg13g2_fill_2 FILLER_88_977 ();
 sg13g2_fill_4 FILLER_88_1005 ();
 sg13g2_fill_8 FILLER_88_1019 ();
 sg13g2_fill_1 FILLER_88_1027 ();
 sg13g2_fill_8 FILLER_88_1039 ();
 sg13g2_fill_8 FILLER_88_1047 ();
 sg13g2_fill_8 FILLER_88_1055 ();
 sg13g2_fill_8 FILLER_88_1063 ();
 sg13g2_fill_8 FILLER_88_1071 ();
 sg13g2_fill_8 FILLER_88_1079 ();
 sg13g2_fill_8 FILLER_88_1087 ();
 sg13g2_fill_8 FILLER_88_1095 ();
 sg13g2_fill_8 FILLER_88_1103 ();
 sg13g2_fill_8 FILLER_88_1111 ();
 sg13g2_fill_8 FILLER_88_1119 ();
 sg13g2_fill_8 FILLER_88_1127 ();
 sg13g2_fill_8 FILLER_88_1135 ();
 sg13g2_fill_8 FILLER_88_1143 ();
 sg13g2_fill_8 FILLER_88_1151 ();
 sg13g2_fill_4 FILLER_88_1159 ();
 sg13g2_fill_2 FILLER_88_1163 ();
 sg13g2_fill_1 FILLER_88_1165 ();
 sg13g2_fill_8 FILLER_89_0 ();
 sg13g2_fill_1 FILLER_89_23 ();
 sg13g2_fill_8 FILLER_89_29 ();
 sg13g2_fill_8 FILLER_89_37 ();
 sg13g2_fill_2 FILLER_89_45 ();
 sg13g2_fill_2 FILLER_89_61 ();
 sg13g2_fill_4 FILLER_89_67 ();
 sg13g2_fill_2 FILLER_89_71 ();
 sg13g2_fill_1 FILLER_89_73 ();
 sg13g2_fill_2 FILLER_89_89 ();
 sg13g2_fill_8 FILLER_89_101 ();
 sg13g2_fill_8 FILLER_89_109 ();
 sg13g2_fill_8 FILLER_89_117 ();
 sg13g2_fill_8 FILLER_89_125 ();
 sg13g2_fill_4 FILLER_89_133 ();
 sg13g2_fill_1 FILLER_89_137 ();
 sg13g2_fill_8 FILLER_89_142 ();
 sg13g2_fill_8 FILLER_89_150 ();
 sg13g2_fill_8 FILLER_89_158 ();
 sg13g2_fill_8 FILLER_89_166 ();
 sg13g2_fill_4 FILLER_89_174 ();
 sg13g2_fill_2 FILLER_89_178 ();
 sg13g2_fill_1 FILLER_89_180 ();
 sg13g2_fill_8 FILLER_89_186 ();
 sg13g2_fill_4 FILLER_89_194 ();
 sg13g2_fill_2 FILLER_89_198 ();
 sg13g2_fill_2 FILLER_89_280 ();
 sg13g2_fill_1 FILLER_89_282 ();
 sg13g2_fill_2 FILLER_89_313 ();
 sg13g2_fill_1 FILLER_89_315 ();
 sg13g2_fill_8 FILLER_89_343 ();
 sg13g2_fill_8 FILLER_89_351 ();
 sg13g2_fill_8 FILLER_89_359 ();
 sg13g2_fill_4 FILLER_89_367 ();
 sg13g2_fill_8 FILLER_89_384 ();
 sg13g2_fill_4 FILLER_89_392 ();
 sg13g2_fill_1 FILLER_89_396 ();
 sg13g2_fill_4 FILLER_89_406 ();
 sg13g2_fill_1 FILLER_89_410 ();
 sg13g2_fill_8 FILLER_89_426 ();
 sg13g2_fill_8 FILLER_89_434 ();
 sg13g2_fill_8 FILLER_89_442 ();
 sg13g2_fill_8 FILLER_89_460 ();
 sg13g2_fill_8 FILLER_89_472 ();
 sg13g2_fill_2 FILLER_89_489 ();
 sg13g2_fill_1 FILLER_89_491 ();
 sg13g2_fill_8 FILLER_89_497 ();
 sg13g2_fill_8 FILLER_89_505 ();
 sg13g2_fill_4 FILLER_89_513 ();
 sg13g2_fill_8 FILLER_89_524 ();
 sg13g2_fill_8 FILLER_89_532 ();
 sg13g2_fill_4 FILLER_89_540 ();
 sg13g2_fill_2 FILLER_89_544 ();
 sg13g2_fill_1 FILLER_89_546 ();
 sg13g2_fill_8 FILLER_89_573 ();
 sg13g2_fill_4 FILLER_89_581 ();
 sg13g2_fill_1 FILLER_89_585 ();
 sg13g2_fill_8 FILLER_89_637 ();
 sg13g2_fill_1 FILLER_89_645 ();
 sg13g2_fill_1 FILLER_89_651 ();
 sg13g2_fill_4 FILLER_89_662 ();
 sg13g2_fill_1 FILLER_89_666 ();
 sg13g2_fill_2 FILLER_89_676 ();
 sg13g2_fill_1 FILLER_89_678 ();
 sg13g2_fill_8 FILLER_89_704 ();
 sg13g2_fill_1 FILLER_89_712 ();
 sg13g2_fill_2 FILLER_89_725 ();
 sg13g2_fill_8 FILLER_89_786 ();
 sg13g2_fill_8 FILLER_89_794 ();
 sg13g2_fill_4 FILLER_89_802 ();
 sg13g2_fill_2 FILLER_89_806 ();
 sg13g2_fill_8 FILLER_89_813 ();
 sg13g2_fill_4 FILLER_89_821 ();
 sg13g2_fill_1 FILLER_89_825 ();
 sg13g2_fill_2 FILLER_89_831 ();
 sg13g2_fill_1 FILLER_89_833 ();
 sg13g2_fill_1 FILLER_89_847 ();
 sg13g2_fill_8 FILLER_89_860 ();
 sg13g2_fill_8 FILLER_89_868 ();
 sg13g2_fill_4 FILLER_89_876 ();
 sg13g2_fill_2 FILLER_89_880 ();
 sg13g2_fill_1 FILLER_89_882 ();
 sg13g2_fill_8 FILLER_89_901 ();
 sg13g2_fill_8 FILLER_89_919 ();
 sg13g2_fill_8 FILLER_89_927 ();
 sg13g2_fill_8 FILLER_89_935 ();
 sg13g2_fill_1 FILLER_89_980 ();
 sg13g2_fill_8 FILLER_89_1018 ();
 sg13g2_fill_8 FILLER_89_1026 ();
 sg13g2_fill_8 FILLER_89_1034 ();
 sg13g2_fill_8 FILLER_89_1042 ();
 sg13g2_fill_8 FILLER_89_1050 ();
 sg13g2_fill_8 FILLER_89_1058 ();
 sg13g2_fill_8 FILLER_89_1066 ();
 sg13g2_fill_8 FILLER_89_1074 ();
 sg13g2_fill_8 FILLER_89_1082 ();
 sg13g2_fill_8 FILLER_89_1090 ();
 sg13g2_fill_8 FILLER_89_1098 ();
 sg13g2_fill_8 FILLER_89_1106 ();
 sg13g2_fill_8 FILLER_89_1114 ();
 sg13g2_fill_8 FILLER_89_1122 ();
 sg13g2_fill_8 FILLER_89_1130 ();
 sg13g2_fill_8 FILLER_89_1138 ();
 sg13g2_fill_8 FILLER_89_1146 ();
 sg13g2_fill_8 FILLER_89_1154 ();
 sg13g2_fill_4 FILLER_89_1162 ();
 sg13g2_fill_4 FILLER_90_0 ();
 sg13g2_fill_2 FILLER_90_4 ();
 sg13g2_fill_1 FILLER_90_6 ();
 sg13g2_fill_1 FILLER_90_12 ();
 sg13g2_fill_2 FILLER_90_31 ();
 sg13g2_fill_8 FILLER_90_65 ();
 sg13g2_fill_1 FILLER_90_73 ();
 sg13g2_fill_2 FILLER_90_99 ();
 sg13g2_fill_1 FILLER_90_101 ();
 sg13g2_fill_1 FILLER_90_107 ();
 sg13g2_fill_2 FILLER_90_118 ();
 sg13g2_fill_1 FILLER_90_120 ();
 sg13g2_fill_2 FILLER_90_131 ();
 sg13g2_fill_2 FILLER_90_143 ();
 sg13g2_fill_8 FILLER_90_150 ();
 sg13g2_fill_2 FILLER_90_158 ();
 sg13g2_fill_4 FILLER_90_170 ();
 sg13g2_fill_2 FILLER_90_174 ();
 sg13g2_fill_1 FILLER_90_176 ();
 sg13g2_fill_8 FILLER_90_185 ();
 sg13g2_fill_8 FILLER_90_193 ();
 sg13g2_fill_4 FILLER_90_201 ();
 sg13g2_fill_2 FILLER_90_243 ();
 sg13g2_fill_1 FILLER_90_245 ();
 sg13g2_fill_8 FILLER_90_285 ();
 sg13g2_fill_8 FILLER_90_293 ();
 sg13g2_fill_8 FILLER_90_301 ();
 sg13g2_fill_2 FILLER_90_309 ();
 sg13g2_fill_1 FILLER_90_311 ();
 sg13g2_fill_2 FILLER_90_320 ();
 sg13g2_fill_1 FILLER_90_322 ();
 sg13g2_fill_4 FILLER_90_332 ();
 sg13g2_fill_4 FILLER_90_343 ();
 sg13g2_fill_1 FILLER_90_347 ();
 sg13g2_fill_8 FILLER_90_385 ();
 sg13g2_fill_4 FILLER_90_393 ();
 sg13g2_fill_1 FILLER_90_397 ();
 sg13g2_fill_2 FILLER_90_408 ();
 sg13g2_fill_8 FILLER_90_429 ();
 sg13g2_fill_4 FILLER_90_437 ();
 sg13g2_fill_2 FILLER_90_441 ();
 sg13g2_fill_4 FILLER_90_452 ();
 sg13g2_fill_2 FILLER_90_456 ();
 sg13g2_fill_1 FILLER_90_458 ();
 sg13g2_fill_4 FILLER_90_469 ();
 sg13g2_fill_2 FILLER_90_473 ();
 sg13g2_fill_4 FILLER_90_480 ();
 sg13g2_fill_8 FILLER_90_508 ();
 sg13g2_fill_4 FILLER_90_516 ();
 sg13g2_fill_1 FILLER_90_520 ();
 sg13g2_fill_4 FILLER_90_530 ();
 sg13g2_fill_4 FILLER_90_547 ();
 sg13g2_fill_1 FILLER_90_551 ();
 sg13g2_fill_4 FILLER_90_564 ();
 sg13g2_fill_1 FILLER_90_568 ();
 sg13g2_fill_8 FILLER_90_595 ();
 sg13g2_fill_1 FILLER_90_609 ();
 sg13g2_fill_8 FILLER_90_636 ();
 sg13g2_fill_8 FILLER_90_659 ();
 sg13g2_fill_8 FILLER_90_667 ();
 sg13g2_fill_8 FILLER_90_675 ();
 sg13g2_fill_4 FILLER_90_683 ();
 sg13g2_fill_1 FILLER_90_687 ();
 sg13g2_fill_1 FILLER_90_697 ();
 sg13g2_fill_4 FILLER_90_703 ();
 sg13g2_fill_2 FILLER_90_707 ();
 sg13g2_fill_2 FILLER_90_717 ();
 sg13g2_fill_2 FILLER_90_737 ();
 sg13g2_fill_1 FILLER_90_739 ();
 sg13g2_fill_8 FILLER_90_770 ();
 sg13g2_fill_8 FILLER_90_778 ();
 sg13g2_fill_8 FILLER_90_786 ();
 sg13g2_fill_8 FILLER_90_794 ();
 sg13g2_fill_2 FILLER_90_802 ();
 sg13g2_fill_8 FILLER_90_819 ();
 sg13g2_fill_2 FILLER_90_846 ();
 sg13g2_fill_8 FILLER_90_862 ();
 sg13g2_fill_8 FILLER_90_870 ();
 sg13g2_fill_8 FILLER_90_878 ();
 sg13g2_fill_8 FILLER_90_886 ();
 sg13g2_fill_8 FILLER_90_894 ();
 sg13g2_fill_8 FILLER_90_902 ();
 sg13g2_fill_8 FILLER_90_910 ();
 sg13g2_fill_8 FILLER_90_918 ();
 sg13g2_fill_8 FILLER_90_926 ();
 sg13g2_fill_8 FILLER_90_934 ();
 sg13g2_fill_8 FILLER_90_942 ();
 sg13g2_fill_8 FILLER_90_950 ();
 sg13g2_fill_8 FILLER_90_958 ();
 sg13g2_fill_8 FILLER_90_966 ();
 sg13g2_fill_1 FILLER_90_974 ();
 sg13g2_fill_8 FILLER_90_985 ();
 sg13g2_fill_1 FILLER_90_993 ();
 sg13g2_fill_8 FILLER_90_1019 ();
 sg13g2_fill_8 FILLER_90_1027 ();
 sg13g2_fill_8 FILLER_90_1035 ();
 sg13g2_fill_8 FILLER_90_1043 ();
 sg13g2_fill_8 FILLER_90_1051 ();
 sg13g2_fill_8 FILLER_90_1059 ();
 sg13g2_fill_8 FILLER_90_1067 ();
 sg13g2_fill_8 FILLER_90_1075 ();
 sg13g2_fill_8 FILLER_90_1083 ();
 sg13g2_fill_8 FILLER_90_1091 ();
 sg13g2_fill_8 FILLER_90_1099 ();
 sg13g2_fill_8 FILLER_90_1107 ();
 sg13g2_fill_8 FILLER_90_1115 ();
 sg13g2_fill_8 FILLER_90_1123 ();
 sg13g2_fill_8 FILLER_90_1131 ();
 sg13g2_fill_8 FILLER_90_1139 ();
 sg13g2_fill_8 FILLER_90_1147 ();
 sg13g2_fill_8 FILLER_90_1155 ();
 sg13g2_fill_2 FILLER_90_1163 ();
 sg13g2_fill_1 FILLER_90_1165 ();
 sg13g2_fill_4 FILLER_91_0 ();
 sg13g2_fill_1 FILLER_91_4 ();
 sg13g2_fill_2 FILLER_91_23 ();
 sg13g2_fill_1 FILLER_91_25 ();
 sg13g2_fill_2 FILLER_91_31 ();
 sg13g2_fill_4 FILLER_91_53 ();
 sg13g2_fill_2 FILLER_91_57 ();
 sg13g2_fill_4 FILLER_91_65 ();
 sg13g2_fill_1 FILLER_91_69 ();
 sg13g2_fill_2 FILLER_91_85 ();
 sg13g2_fill_2 FILLER_91_120 ();
 sg13g2_fill_2 FILLER_91_155 ();
 sg13g2_fill_1 FILLER_91_157 ();
 sg13g2_fill_2 FILLER_91_198 ();
 sg13g2_fill_8 FILLER_91_215 ();
 sg13g2_fill_4 FILLER_91_223 ();
 sg13g2_fill_2 FILLER_91_227 ();
 sg13g2_fill_1 FILLER_91_229 ();
 sg13g2_fill_1 FILLER_91_237 ();
 sg13g2_fill_1 FILLER_91_278 ();
 sg13g2_fill_8 FILLER_91_296 ();
 sg13g2_fill_2 FILLER_91_338 ();
 sg13g2_fill_4 FILLER_91_370 ();
 sg13g2_fill_2 FILLER_91_374 ();
 sg13g2_fill_8 FILLER_91_428 ();
 sg13g2_fill_2 FILLER_91_462 ();
 sg13g2_fill_4 FILLER_91_542 ();
 sg13g2_fill_1 FILLER_91_546 ();
 sg13g2_fill_1 FILLER_91_560 ();
 sg13g2_fill_4 FILLER_91_605 ();
 sg13g2_fill_1 FILLER_91_609 ();
 sg13g2_fill_2 FILLER_91_636 ();
 sg13g2_fill_1 FILLER_91_638 ();
 sg13g2_fill_4 FILLER_91_649 ();
 sg13g2_fill_2 FILLER_91_653 ();
 sg13g2_fill_8 FILLER_91_661 ();
 sg13g2_fill_4 FILLER_91_669 ();
 sg13g2_fill_1 FILLER_91_673 ();
 sg13g2_fill_2 FILLER_91_682 ();
 sg13g2_fill_8 FILLER_91_710 ();
 sg13g2_fill_4 FILLER_91_718 ();
 sg13g2_fill_8 FILLER_91_752 ();
 sg13g2_fill_8 FILLER_91_760 ();
 sg13g2_fill_8 FILLER_91_768 ();
 sg13g2_fill_8 FILLER_91_776 ();
 sg13g2_fill_4 FILLER_91_784 ();
 sg13g2_fill_2 FILLER_91_788 ();
 sg13g2_fill_4 FILLER_91_820 ();
 sg13g2_fill_2 FILLER_91_824 ();
 sg13g2_fill_1 FILLER_91_826 ();
 sg13g2_fill_4 FILLER_91_832 ();
 sg13g2_fill_2 FILLER_91_836 ();
 sg13g2_fill_1 FILLER_91_838 ();
 sg13g2_fill_8 FILLER_91_848 ();
 sg13g2_fill_8 FILLER_91_856 ();
 sg13g2_fill_8 FILLER_91_864 ();
 sg13g2_fill_8 FILLER_91_872 ();
 sg13g2_fill_8 FILLER_91_880 ();
 sg13g2_fill_8 FILLER_91_888 ();
 sg13g2_fill_8 FILLER_91_896 ();
 sg13g2_fill_4 FILLER_91_904 ();
 sg13g2_fill_2 FILLER_91_908 ();
 sg13g2_fill_1 FILLER_91_910 ();
 sg13g2_fill_4 FILLER_91_937 ();
 sg13g2_fill_2 FILLER_91_941 ();
 sg13g2_fill_8 FILLER_91_961 ();
 sg13g2_fill_8 FILLER_91_969 ();
 sg13g2_fill_4 FILLER_91_977 ();
 sg13g2_fill_1 FILLER_91_981 ();
 sg13g2_fill_1 FILLER_91_992 ();
 sg13g2_fill_8 FILLER_91_1019 ();
 sg13g2_fill_8 FILLER_91_1027 ();
 sg13g2_fill_8 FILLER_91_1035 ();
 sg13g2_fill_8 FILLER_91_1043 ();
 sg13g2_fill_8 FILLER_91_1051 ();
 sg13g2_fill_8 FILLER_91_1059 ();
 sg13g2_fill_8 FILLER_91_1067 ();
 sg13g2_fill_8 FILLER_91_1075 ();
 sg13g2_fill_8 FILLER_91_1083 ();
 sg13g2_fill_8 FILLER_91_1091 ();
 sg13g2_fill_8 FILLER_91_1099 ();
 sg13g2_fill_8 FILLER_91_1107 ();
 sg13g2_fill_8 FILLER_91_1115 ();
 sg13g2_fill_8 FILLER_91_1123 ();
 sg13g2_fill_8 FILLER_91_1131 ();
 sg13g2_fill_8 FILLER_91_1139 ();
 sg13g2_fill_8 FILLER_91_1147 ();
 sg13g2_fill_8 FILLER_91_1155 ();
 sg13g2_fill_2 FILLER_91_1163 ();
 sg13g2_fill_1 FILLER_91_1165 ();
 sg13g2_fill_8 FILLER_92_0 ();
 sg13g2_fill_4 FILLER_92_8 ();
 sg13g2_fill_4 FILLER_92_32 ();
 sg13g2_fill_2 FILLER_92_36 ();
 sg13g2_fill_8 FILLER_92_63 ();
 sg13g2_fill_4 FILLER_92_71 ();
 sg13g2_fill_2 FILLER_92_75 ();
 sg13g2_fill_8 FILLER_92_82 ();
 sg13g2_fill_1 FILLER_92_90 ();
 sg13g2_fill_1 FILLER_92_111 ();
 sg13g2_fill_4 FILLER_92_138 ();
 sg13g2_fill_2 FILLER_92_152 ();
 sg13g2_fill_1 FILLER_92_154 ();
 sg13g2_fill_4 FILLER_92_200 ();
 sg13g2_fill_2 FILLER_92_204 ();
 sg13g2_fill_1 FILLER_92_206 ();
 sg13g2_fill_1 FILLER_92_232 ();
 sg13g2_fill_8 FILLER_92_268 ();
 sg13g2_fill_8 FILLER_92_276 ();
 sg13g2_fill_4 FILLER_92_284 ();
 sg13g2_fill_4 FILLER_92_318 ();
 sg13g2_fill_2 FILLER_92_322 ();
 sg13g2_fill_8 FILLER_92_387 ();
 sg13g2_fill_4 FILLER_92_395 ();
 sg13g2_fill_1 FILLER_92_399 ();
 sg13g2_fill_4 FILLER_92_437 ();
 sg13g2_fill_2 FILLER_92_441 ();
 sg13g2_fill_1 FILLER_92_443 ();
 sg13g2_fill_1 FILLER_92_451 ();
 sg13g2_fill_8 FILLER_92_488 ();
 sg13g2_fill_1 FILLER_92_496 ();
 sg13g2_fill_4 FILLER_92_507 ();
 sg13g2_fill_1 FILLER_92_511 ();
 sg13g2_fill_8 FILLER_92_538 ();
 sg13g2_fill_4 FILLER_92_546 ();
 sg13g2_fill_2 FILLER_92_550 ();
 sg13g2_fill_1 FILLER_92_552 ();
 sg13g2_fill_8 FILLER_92_611 ();
 sg13g2_fill_8 FILLER_92_619 ();
 sg13g2_fill_2 FILLER_92_627 ();
 sg13g2_fill_8 FILLER_92_634 ();
 sg13g2_fill_2 FILLER_92_642 ();
 sg13g2_fill_1 FILLER_92_644 ();
 sg13g2_fill_8 FILLER_92_674 ();
 sg13g2_fill_8 FILLER_92_682 ();
 sg13g2_fill_2 FILLER_92_695 ();
 sg13g2_fill_4 FILLER_92_709 ();
 sg13g2_fill_8 FILLER_92_718 ();
 sg13g2_fill_1 FILLER_92_726 ();
 sg13g2_fill_1 FILLER_92_732 ();
 sg13g2_fill_8 FILLER_92_763 ();
 sg13g2_fill_8 FILLER_92_771 ();
 sg13g2_fill_8 FILLER_92_779 ();
 sg13g2_fill_2 FILLER_92_787 ();
 sg13g2_fill_1 FILLER_92_789 ();
 sg13g2_fill_1 FILLER_92_810 ();
 sg13g2_fill_1 FILLER_92_834 ();
 sg13g2_fill_8 FILLER_92_855 ();
 sg13g2_fill_8 FILLER_92_863 ();
 sg13g2_fill_8 FILLER_92_871 ();
 sg13g2_fill_8 FILLER_92_879 ();
 sg13g2_fill_8 FILLER_92_887 ();
 sg13g2_fill_4 FILLER_92_895 ();
 sg13g2_fill_2 FILLER_92_899 ();
 sg13g2_fill_4 FILLER_92_948 ();
 sg13g2_fill_2 FILLER_92_952 ();
 sg13g2_fill_4 FILLER_92_980 ();
 sg13g2_fill_2 FILLER_92_984 ();
 sg13g2_fill_1 FILLER_92_986 ();
 sg13g2_fill_8 FILLER_92_1024 ();
 sg13g2_fill_8 FILLER_92_1032 ();
 sg13g2_fill_8 FILLER_92_1040 ();
 sg13g2_fill_8 FILLER_92_1048 ();
 sg13g2_fill_8 FILLER_92_1056 ();
 sg13g2_fill_8 FILLER_92_1064 ();
 sg13g2_fill_8 FILLER_92_1072 ();
 sg13g2_fill_8 FILLER_92_1080 ();
 sg13g2_fill_8 FILLER_92_1088 ();
 sg13g2_fill_8 FILLER_92_1096 ();
 sg13g2_fill_8 FILLER_92_1104 ();
 sg13g2_fill_8 FILLER_92_1112 ();
 sg13g2_fill_8 FILLER_92_1120 ();
 sg13g2_fill_8 FILLER_92_1128 ();
 sg13g2_fill_8 FILLER_92_1136 ();
 sg13g2_fill_8 FILLER_92_1144 ();
 sg13g2_fill_8 FILLER_92_1152 ();
 sg13g2_fill_4 FILLER_92_1160 ();
 sg13g2_fill_2 FILLER_92_1164 ();
 sg13g2_fill_8 FILLER_93_0 ();
 sg13g2_fill_8 FILLER_93_8 ();
 sg13g2_fill_8 FILLER_93_16 ();
 sg13g2_fill_8 FILLER_93_24 ();
 sg13g2_fill_8 FILLER_93_32 ();
 sg13g2_fill_8 FILLER_93_40 ();
 sg13g2_fill_4 FILLER_93_48 ();
 sg13g2_fill_2 FILLER_93_52 ();
 sg13g2_fill_8 FILLER_93_79 ();
 sg13g2_fill_8 FILLER_93_87 ();
 sg13g2_fill_8 FILLER_93_95 ();
 sg13g2_fill_8 FILLER_93_103 ();
 sg13g2_fill_8 FILLER_93_116 ();
 sg13g2_fill_4 FILLER_93_124 ();
 sg13g2_fill_2 FILLER_93_128 ();
 sg13g2_fill_8 FILLER_93_155 ();
 sg13g2_fill_4 FILLER_93_163 ();
 sg13g2_fill_1 FILLER_93_167 ();
 sg13g2_fill_4 FILLER_93_198 ();
 sg13g2_fill_2 FILLER_93_202 ();
 sg13g2_fill_4 FILLER_93_279 ();
 sg13g2_fill_4 FILLER_93_313 ();
 sg13g2_fill_2 FILLER_93_317 ();
 sg13g2_fill_2 FILLER_93_358 ();
 sg13g2_fill_8 FILLER_93_368 ();
 sg13g2_fill_2 FILLER_93_376 ();
 sg13g2_fill_8 FILLER_93_440 ();
 sg13g2_fill_8 FILLER_93_448 ();
 sg13g2_fill_2 FILLER_93_456 ();
 sg13g2_fill_4 FILLER_93_475 ();
 sg13g2_fill_2 FILLER_93_479 ();
 sg13g2_fill_4 FILLER_93_485 ();
 sg13g2_fill_2 FILLER_93_489 ();
 sg13g2_fill_1 FILLER_93_491 ();
 sg13g2_fill_8 FILLER_93_498 ();
 sg13g2_fill_8 FILLER_93_506 ();
 sg13g2_fill_4 FILLER_93_514 ();
 sg13g2_fill_2 FILLER_93_518 ();
 sg13g2_fill_1 FILLER_93_520 ();
 sg13g2_fill_8 FILLER_93_597 ();
 sg13g2_fill_4 FILLER_93_605 ();
 sg13g2_fill_4 FILLER_93_622 ();
 sg13g2_fill_1 FILLER_93_626 ();
 sg13g2_fill_8 FILLER_93_630 ();
 sg13g2_fill_2 FILLER_93_699 ();
 sg13g2_fill_1 FILLER_93_701 ();
 sg13g2_fill_8 FILLER_93_762 ();
 sg13g2_fill_8 FILLER_93_770 ();
 sg13g2_fill_8 FILLER_93_778 ();
 sg13g2_fill_8 FILLER_93_786 ();
 sg13g2_fill_1 FILLER_93_794 ();
 sg13g2_fill_2 FILLER_93_832 ();
 sg13g2_fill_1 FILLER_93_834 ();
 sg13g2_fill_8 FILLER_93_861 ();
 sg13g2_fill_8 FILLER_93_869 ();
 sg13g2_fill_8 FILLER_93_877 ();
 sg13g2_fill_8 FILLER_93_885 ();
 sg13g2_fill_8 FILLER_93_893 ();
 sg13g2_fill_8 FILLER_93_901 ();
 sg13g2_fill_2 FILLER_93_919 ();
 sg13g2_fill_1 FILLER_93_921 ();
 sg13g2_fill_8 FILLER_93_930 ();
 sg13g2_fill_8 FILLER_93_938 ();
 sg13g2_fill_2 FILLER_93_946 ();
 sg13g2_fill_4 FILLER_93_984 ();
 sg13g2_fill_1 FILLER_93_988 ();
 sg13g2_fill_8 FILLER_93_999 ();
 sg13g2_fill_8 FILLER_93_1007 ();
 sg13g2_fill_8 FILLER_93_1015 ();
 sg13g2_fill_8 FILLER_93_1023 ();
 sg13g2_fill_8 FILLER_93_1031 ();
 sg13g2_fill_8 FILLER_93_1039 ();
 sg13g2_fill_8 FILLER_93_1047 ();
 sg13g2_fill_8 FILLER_93_1055 ();
 sg13g2_fill_8 FILLER_93_1063 ();
 sg13g2_fill_8 FILLER_93_1071 ();
 sg13g2_fill_8 FILLER_93_1079 ();
 sg13g2_fill_8 FILLER_93_1087 ();
 sg13g2_fill_8 FILLER_93_1095 ();
 sg13g2_fill_8 FILLER_93_1103 ();
 sg13g2_fill_8 FILLER_93_1111 ();
 sg13g2_fill_8 FILLER_93_1119 ();
 sg13g2_fill_8 FILLER_93_1127 ();
 sg13g2_fill_8 FILLER_93_1135 ();
 sg13g2_fill_8 FILLER_93_1143 ();
 sg13g2_fill_8 FILLER_93_1151 ();
 sg13g2_fill_4 FILLER_93_1159 ();
 sg13g2_fill_2 FILLER_93_1163 ();
 sg13g2_fill_1 FILLER_93_1165 ();
 sg13g2_fill_8 FILLER_94_0 ();
 sg13g2_fill_8 FILLER_94_8 ();
 sg13g2_fill_8 FILLER_94_16 ();
 sg13g2_fill_8 FILLER_94_24 ();
 sg13g2_fill_8 FILLER_94_32 ();
 sg13g2_fill_8 FILLER_94_40 ();
 sg13g2_fill_8 FILLER_94_48 ();
 sg13g2_fill_8 FILLER_94_56 ();
 sg13g2_fill_8 FILLER_94_64 ();
 sg13g2_fill_8 FILLER_94_72 ();
 sg13g2_fill_8 FILLER_94_80 ();
 sg13g2_fill_8 FILLER_94_88 ();
 sg13g2_fill_8 FILLER_94_96 ();
 sg13g2_fill_8 FILLER_94_104 ();
 sg13g2_fill_8 FILLER_94_112 ();
 sg13g2_fill_8 FILLER_94_120 ();
 sg13g2_fill_8 FILLER_94_128 ();
 sg13g2_fill_8 FILLER_94_136 ();
 sg13g2_fill_8 FILLER_94_144 ();
 sg13g2_fill_8 FILLER_94_152 ();
 sg13g2_fill_8 FILLER_94_160 ();
 sg13g2_fill_8 FILLER_94_168 ();
 sg13g2_fill_8 FILLER_94_176 ();
 sg13g2_fill_8 FILLER_94_184 ();
 sg13g2_fill_2 FILLER_94_192 ();
 sg13g2_fill_4 FILLER_94_234 ();
 sg13g2_fill_2 FILLER_94_238 ();
 sg13g2_fill_1 FILLER_94_240 ();
 sg13g2_fill_8 FILLER_94_281 ();
 sg13g2_fill_1 FILLER_94_319 ();
 sg13g2_fill_4 FILLER_94_357 ();
 sg13g2_fill_1 FILLER_94_361 ();
 sg13g2_fill_8 FILLER_94_370 ();
 sg13g2_fill_4 FILLER_94_408 ();
 sg13g2_fill_2 FILLER_94_435 ();
 sg13g2_fill_8 FILLER_94_446 ();
 sg13g2_fill_8 FILLER_94_462 ();
 sg13g2_fill_2 FILLER_94_470 ();
 sg13g2_fill_1 FILLER_94_472 ();
 sg13g2_fill_4 FILLER_94_502 ();
 sg13g2_fill_8 FILLER_94_516 ();
 sg13g2_fill_8 FILLER_94_524 ();
 sg13g2_fill_4 FILLER_94_532 ();
 sg13g2_fill_1 FILLER_94_536 ();
 sg13g2_fill_4 FILLER_94_543 ();
 sg13g2_fill_1 FILLER_94_547 ();
 sg13g2_fill_8 FILLER_94_579 ();
 sg13g2_fill_8 FILLER_94_587 ();
 sg13g2_fill_2 FILLER_94_595 ();
 sg13g2_fill_1 FILLER_94_622 ();
 sg13g2_fill_4 FILLER_94_640 ();
 sg13g2_fill_8 FILLER_94_677 ();
 sg13g2_fill_4 FILLER_94_685 ();
 sg13g2_fill_1 FILLER_94_689 ();
 sg13g2_fill_1 FILLER_94_695 ();
 sg13g2_fill_8 FILLER_94_726 ();
 sg13g2_fill_8 FILLER_94_734 ();
 sg13g2_fill_8 FILLER_94_742 ();
 sg13g2_fill_8 FILLER_94_750 ();
 sg13g2_fill_8 FILLER_94_758 ();
 sg13g2_fill_8 FILLER_94_766 ();
 sg13g2_fill_8 FILLER_94_774 ();
 sg13g2_fill_8 FILLER_94_782 ();
 sg13g2_fill_8 FILLER_94_790 ();
 sg13g2_fill_8 FILLER_94_798 ();
 sg13g2_fill_8 FILLER_94_806 ();
 sg13g2_fill_4 FILLER_94_814 ();
 sg13g2_fill_2 FILLER_94_844 ();
 sg13g2_fill_8 FILLER_94_860 ();
 sg13g2_fill_8 FILLER_94_868 ();
 sg13g2_fill_8 FILLER_94_876 ();
 sg13g2_fill_8 FILLER_94_884 ();
 sg13g2_fill_8 FILLER_94_892 ();
 sg13g2_fill_8 FILLER_94_900 ();
 sg13g2_fill_8 FILLER_94_908 ();
 sg13g2_fill_8 FILLER_94_916 ();
 sg13g2_fill_4 FILLER_94_924 ();
 sg13g2_fill_2 FILLER_94_928 ();
 sg13g2_fill_1 FILLER_94_930 ();
 sg13g2_fill_4 FILLER_94_971 ();
 sg13g2_fill_2 FILLER_94_975 ();
 sg13g2_fill_8 FILLER_94_988 ();
 sg13g2_fill_8 FILLER_94_996 ();
 sg13g2_fill_8 FILLER_94_1004 ();
 sg13g2_fill_8 FILLER_94_1012 ();
 sg13g2_fill_8 FILLER_94_1020 ();
 sg13g2_fill_8 FILLER_94_1028 ();
 sg13g2_fill_8 FILLER_94_1036 ();
 sg13g2_fill_8 FILLER_94_1044 ();
 sg13g2_fill_8 FILLER_94_1052 ();
 sg13g2_fill_8 FILLER_94_1060 ();
 sg13g2_fill_8 FILLER_94_1068 ();
 sg13g2_fill_8 FILLER_94_1076 ();
 sg13g2_fill_8 FILLER_94_1084 ();
 sg13g2_fill_8 FILLER_94_1092 ();
 sg13g2_fill_8 FILLER_94_1100 ();
 sg13g2_fill_8 FILLER_94_1108 ();
 sg13g2_fill_8 FILLER_94_1116 ();
 sg13g2_fill_8 FILLER_94_1124 ();
 sg13g2_fill_8 FILLER_94_1132 ();
 sg13g2_fill_8 FILLER_94_1140 ();
 sg13g2_fill_8 FILLER_94_1148 ();
 sg13g2_fill_8 FILLER_94_1156 ();
 sg13g2_fill_2 FILLER_94_1164 ();
 sg13g2_fill_8 FILLER_95_0 ();
 sg13g2_fill_8 FILLER_95_8 ();
 sg13g2_fill_8 FILLER_95_16 ();
 sg13g2_fill_8 FILLER_95_24 ();
 sg13g2_fill_8 FILLER_95_32 ();
 sg13g2_fill_8 FILLER_95_40 ();
 sg13g2_fill_8 FILLER_95_48 ();
 sg13g2_fill_8 FILLER_95_56 ();
 sg13g2_fill_8 FILLER_95_64 ();
 sg13g2_fill_8 FILLER_95_72 ();
 sg13g2_fill_8 FILLER_95_80 ();
 sg13g2_fill_8 FILLER_95_88 ();
 sg13g2_fill_8 FILLER_95_96 ();
 sg13g2_fill_8 FILLER_95_104 ();
 sg13g2_fill_8 FILLER_95_112 ();
 sg13g2_fill_8 FILLER_95_120 ();
 sg13g2_fill_8 FILLER_95_128 ();
 sg13g2_fill_8 FILLER_95_136 ();
 sg13g2_fill_8 FILLER_95_144 ();
 sg13g2_fill_8 FILLER_95_152 ();
 sg13g2_fill_8 FILLER_95_160 ();
 sg13g2_fill_8 FILLER_95_168 ();
 sg13g2_fill_8 FILLER_95_176 ();
 sg13g2_fill_8 FILLER_95_184 ();
 sg13g2_fill_8 FILLER_95_192 ();
 sg13g2_fill_8 FILLER_95_200 ();
 sg13g2_fill_8 FILLER_95_208 ();
 sg13g2_fill_8 FILLER_95_216 ();
 sg13g2_fill_8 FILLER_95_224 ();
 sg13g2_fill_4 FILLER_95_232 ();
 sg13g2_fill_2 FILLER_95_236 ();
 sg13g2_fill_1 FILLER_95_238 ();
 sg13g2_fill_1 FILLER_95_269 ();
 sg13g2_fill_8 FILLER_95_300 ();
 sg13g2_fill_8 FILLER_95_308 ();
 sg13g2_fill_2 FILLER_95_316 ();
 sg13g2_fill_1 FILLER_95_318 ();
 sg13g2_fill_8 FILLER_95_381 ();
 sg13g2_fill_8 FILLER_95_389 ();
 sg13g2_fill_8 FILLER_95_397 ();
 sg13g2_fill_4 FILLER_95_405 ();
 sg13g2_fill_1 FILLER_95_409 ();
 sg13g2_fill_2 FILLER_95_471 ();
 sg13g2_fill_1 FILLER_95_473 ();
 sg13g2_fill_2 FILLER_95_483 ();
 sg13g2_fill_1 FILLER_95_485 ();
 sg13g2_fill_8 FILLER_95_504 ();
 sg13g2_fill_8 FILLER_95_512 ();
 sg13g2_fill_8 FILLER_95_520 ();
 sg13g2_fill_2 FILLER_95_528 ();
 sg13g2_fill_1 FILLER_95_530 ();
 sg13g2_fill_8 FILLER_95_566 ();
 sg13g2_fill_1 FILLER_95_574 ();
 sg13g2_fill_2 FILLER_95_601 ();
 sg13g2_fill_2 FILLER_95_617 ();
 sg13g2_fill_1 FILLER_95_650 ();
 sg13g2_fill_8 FILLER_95_676 ();
 sg13g2_fill_8 FILLER_95_684 ();
 sg13g2_fill_8 FILLER_95_692 ();
 sg13g2_fill_8 FILLER_95_700 ();
 sg13g2_fill_8 FILLER_95_708 ();
 sg13g2_fill_8 FILLER_95_716 ();
 sg13g2_fill_8 FILLER_95_724 ();
 sg13g2_fill_8 FILLER_95_732 ();
 sg13g2_fill_8 FILLER_95_740 ();
 sg13g2_fill_8 FILLER_95_748 ();
 sg13g2_fill_8 FILLER_95_756 ();
 sg13g2_fill_8 FILLER_95_764 ();
 sg13g2_fill_8 FILLER_95_772 ();
 sg13g2_fill_8 FILLER_95_780 ();
 sg13g2_fill_8 FILLER_95_788 ();
 sg13g2_fill_8 FILLER_95_796 ();
 sg13g2_fill_8 FILLER_95_804 ();
 sg13g2_fill_8 FILLER_95_812 ();
 sg13g2_fill_8 FILLER_95_820 ();
 sg13g2_fill_8 FILLER_95_828 ();
 sg13g2_fill_8 FILLER_95_836 ();
 sg13g2_fill_8 FILLER_95_844 ();
 sg13g2_fill_8 FILLER_95_852 ();
 sg13g2_fill_8 FILLER_95_860 ();
 sg13g2_fill_8 FILLER_95_868 ();
 sg13g2_fill_8 FILLER_95_876 ();
 sg13g2_fill_8 FILLER_95_884 ();
 sg13g2_fill_8 FILLER_95_892 ();
 sg13g2_fill_8 FILLER_95_900 ();
 sg13g2_fill_4 FILLER_95_908 ();
 sg13g2_fill_2 FILLER_95_912 ();
 sg13g2_fill_1 FILLER_95_914 ();
 sg13g2_fill_4 FILLER_95_941 ();
 sg13g2_fill_2 FILLER_95_945 ();
 sg13g2_fill_8 FILLER_95_973 ();
 sg13g2_fill_4 FILLER_95_981 ();
 sg13g2_fill_8 FILLER_95_1011 ();
 sg13g2_fill_8 FILLER_95_1019 ();
 sg13g2_fill_8 FILLER_95_1027 ();
 sg13g2_fill_8 FILLER_95_1035 ();
 sg13g2_fill_8 FILLER_95_1043 ();
 sg13g2_fill_8 FILLER_95_1051 ();
 sg13g2_fill_8 FILLER_95_1059 ();
 sg13g2_fill_8 FILLER_95_1067 ();
 sg13g2_fill_8 FILLER_95_1075 ();
 sg13g2_fill_8 FILLER_95_1083 ();
 sg13g2_fill_8 FILLER_95_1091 ();
 sg13g2_fill_8 FILLER_95_1099 ();
 sg13g2_fill_8 FILLER_95_1107 ();
 sg13g2_fill_8 FILLER_95_1115 ();
 sg13g2_fill_8 FILLER_95_1123 ();
 sg13g2_fill_8 FILLER_95_1131 ();
 sg13g2_fill_8 FILLER_95_1139 ();
 sg13g2_fill_8 FILLER_95_1147 ();
 sg13g2_fill_8 FILLER_95_1155 ();
 sg13g2_fill_2 FILLER_95_1163 ();
 sg13g2_fill_1 FILLER_95_1165 ();
 sg13g2_fill_8 FILLER_96_0 ();
 sg13g2_fill_8 FILLER_96_8 ();
 sg13g2_fill_8 FILLER_96_16 ();
 sg13g2_fill_8 FILLER_96_24 ();
 sg13g2_fill_8 FILLER_96_32 ();
 sg13g2_fill_8 FILLER_96_40 ();
 sg13g2_fill_8 FILLER_96_48 ();
 sg13g2_fill_8 FILLER_96_56 ();
 sg13g2_fill_8 FILLER_96_64 ();
 sg13g2_fill_8 FILLER_96_72 ();
 sg13g2_fill_8 FILLER_96_80 ();
 sg13g2_fill_8 FILLER_96_88 ();
 sg13g2_fill_8 FILLER_96_96 ();
 sg13g2_fill_8 FILLER_96_104 ();
 sg13g2_fill_8 FILLER_96_112 ();
 sg13g2_fill_8 FILLER_96_120 ();
 sg13g2_fill_8 FILLER_96_128 ();
 sg13g2_fill_8 FILLER_96_136 ();
 sg13g2_fill_8 FILLER_96_144 ();
 sg13g2_fill_8 FILLER_96_152 ();
 sg13g2_fill_8 FILLER_96_160 ();
 sg13g2_fill_8 FILLER_96_168 ();
 sg13g2_fill_8 FILLER_96_176 ();
 sg13g2_fill_8 FILLER_96_184 ();
 sg13g2_fill_8 FILLER_96_192 ();
 sg13g2_fill_8 FILLER_96_200 ();
 sg13g2_fill_8 FILLER_96_208 ();
 sg13g2_fill_8 FILLER_96_216 ();
 sg13g2_fill_8 FILLER_96_224 ();
 sg13g2_fill_8 FILLER_96_232 ();
 sg13g2_fill_8 FILLER_96_240 ();
 sg13g2_fill_8 FILLER_96_248 ();
 sg13g2_fill_8 FILLER_96_256 ();
 sg13g2_fill_8 FILLER_96_264 ();
 sg13g2_fill_8 FILLER_96_272 ();
 sg13g2_fill_8 FILLER_96_280 ();
 sg13g2_fill_8 FILLER_96_288 ();
 sg13g2_fill_8 FILLER_96_296 ();
 sg13g2_fill_8 FILLER_96_304 ();
 sg13g2_fill_8 FILLER_96_312 ();
 sg13g2_fill_8 FILLER_96_320 ();
 sg13g2_fill_8 FILLER_96_328 ();
 sg13g2_fill_8 FILLER_96_336 ();
 sg13g2_fill_8 FILLER_96_344 ();
 sg13g2_fill_8 FILLER_96_352 ();
 sg13g2_fill_8 FILLER_96_360 ();
 sg13g2_fill_8 FILLER_96_368 ();
 sg13g2_fill_8 FILLER_96_376 ();
 sg13g2_fill_4 FILLER_96_384 ();
 sg13g2_fill_2 FILLER_96_388 ();
 sg13g2_fill_1 FILLER_96_390 ();
 sg13g2_fill_8 FILLER_96_399 ();
 sg13g2_fill_8 FILLER_96_407 ();
 sg13g2_fill_4 FILLER_96_415 ();
 sg13g2_fill_8 FILLER_96_445 ();
 sg13g2_fill_1 FILLER_96_453 ();
 sg13g2_fill_2 FILLER_96_513 ();
 sg13g2_fill_2 FILLER_96_520 ();
 sg13g2_fill_2 FILLER_96_548 ();
 sg13g2_fill_8 FILLER_96_648 ();
 sg13g2_fill_8 FILLER_96_656 ();
 sg13g2_fill_8 FILLER_96_664 ();
 sg13g2_fill_8 FILLER_96_672 ();
 sg13g2_fill_8 FILLER_96_680 ();
 sg13g2_fill_8 FILLER_96_688 ();
 sg13g2_fill_8 FILLER_96_696 ();
 sg13g2_fill_8 FILLER_96_704 ();
 sg13g2_fill_8 FILLER_96_712 ();
 sg13g2_fill_8 FILLER_96_720 ();
 sg13g2_fill_8 FILLER_96_728 ();
 sg13g2_fill_8 FILLER_96_736 ();
 sg13g2_fill_8 FILLER_96_744 ();
 sg13g2_fill_8 FILLER_96_752 ();
 sg13g2_fill_8 FILLER_96_760 ();
 sg13g2_fill_8 FILLER_96_768 ();
 sg13g2_fill_8 FILLER_96_776 ();
 sg13g2_fill_8 FILLER_96_784 ();
 sg13g2_fill_8 FILLER_96_792 ();
 sg13g2_fill_8 FILLER_96_800 ();
 sg13g2_fill_8 FILLER_96_808 ();
 sg13g2_fill_8 FILLER_96_816 ();
 sg13g2_fill_8 FILLER_96_824 ();
 sg13g2_fill_8 FILLER_96_832 ();
 sg13g2_fill_8 FILLER_96_840 ();
 sg13g2_fill_8 FILLER_96_848 ();
 sg13g2_fill_8 FILLER_96_856 ();
 sg13g2_fill_8 FILLER_96_864 ();
 sg13g2_fill_8 FILLER_96_872 ();
 sg13g2_fill_8 FILLER_96_880 ();
 sg13g2_fill_8 FILLER_96_888 ();
 sg13g2_fill_8 FILLER_96_896 ();
 sg13g2_fill_1 FILLER_96_904 ();
 sg13g2_fill_4 FILLER_96_941 ();
 sg13g2_fill_2 FILLER_96_945 ();
 sg13g2_fill_1 FILLER_96_973 ();
 sg13g2_fill_8 FILLER_96_1021 ();
 sg13g2_fill_8 FILLER_96_1029 ();
 sg13g2_fill_8 FILLER_96_1037 ();
 sg13g2_fill_8 FILLER_96_1045 ();
 sg13g2_fill_8 FILLER_96_1053 ();
 sg13g2_fill_8 FILLER_96_1061 ();
 sg13g2_fill_8 FILLER_96_1069 ();
 sg13g2_fill_8 FILLER_96_1077 ();
 sg13g2_fill_8 FILLER_96_1085 ();
 sg13g2_fill_8 FILLER_96_1093 ();
 sg13g2_fill_8 FILLER_96_1101 ();
 sg13g2_fill_8 FILLER_96_1109 ();
 sg13g2_fill_8 FILLER_96_1117 ();
 sg13g2_fill_8 FILLER_96_1125 ();
 sg13g2_fill_8 FILLER_96_1133 ();
 sg13g2_fill_8 FILLER_96_1141 ();
 sg13g2_fill_8 FILLER_96_1149 ();
 sg13g2_fill_8 FILLER_96_1157 ();
 sg13g2_fill_1 FILLER_96_1165 ();
 sg13g2_fill_8 FILLER_97_0 ();
 sg13g2_fill_8 FILLER_97_8 ();
 sg13g2_fill_8 FILLER_97_16 ();
 sg13g2_fill_8 FILLER_97_24 ();
 sg13g2_fill_8 FILLER_97_32 ();
 sg13g2_fill_8 FILLER_97_40 ();
 sg13g2_fill_8 FILLER_97_48 ();
 sg13g2_fill_8 FILLER_97_56 ();
 sg13g2_fill_8 FILLER_97_64 ();
 sg13g2_fill_8 FILLER_97_72 ();
 sg13g2_fill_8 FILLER_97_80 ();
 sg13g2_fill_8 FILLER_97_88 ();
 sg13g2_fill_8 FILLER_97_96 ();
 sg13g2_fill_8 FILLER_97_104 ();
 sg13g2_fill_8 FILLER_97_112 ();
 sg13g2_fill_8 FILLER_97_120 ();
 sg13g2_fill_8 FILLER_97_128 ();
 sg13g2_fill_8 FILLER_97_136 ();
 sg13g2_fill_8 FILLER_97_144 ();
 sg13g2_fill_8 FILLER_97_152 ();
 sg13g2_fill_8 FILLER_97_160 ();
 sg13g2_fill_8 FILLER_97_168 ();
 sg13g2_fill_8 FILLER_97_176 ();
 sg13g2_fill_8 FILLER_97_184 ();
 sg13g2_fill_8 FILLER_97_192 ();
 sg13g2_fill_8 FILLER_97_200 ();
 sg13g2_fill_8 FILLER_97_208 ();
 sg13g2_fill_8 FILLER_97_216 ();
 sg13g2_fill_8 FILLER_97_224 ();
 sg13g2_fill_8 FILLER_97_232 ();
 sg13g2_fill_8 FILLER_97_240 ();
 sg13g2_fill_8 FILLER_97_248 ();
 sg13g2_fill_8 FILLER_97_256 ();
 sg13g2_fill_8 FILLER_97_264 ();
 sg13g2_fill_8 FILLER_97_272 ();
 sg13g2_fill_8 FILLER_97_280 ();
 sg13g2_fill_8 FILLER_97_288 ();
 sg13g2_fill_8 FILLER_97_296 ();
 sg13g2_fill_8 FILLER_97_304 ();
 sg13g2_fill_8 FILLER_97_312 ();
 sg13g2_fill_8 FILLER_97_320 ();
 sg13g2_fill_8 FILLER_97_328 ();
 sg13g2_fill_8 FILLER_97_336 ();
 sg13g2_fill_8 FILLER_97_344 ();
 sg13g2_fill_8 FILLER_97_352 ();
 sg13g2_fill_8 FILLER_97_360 ();
 sg13g2_fill_8 FILLER_97_368 ();
 sg13g2_fill_8 FILLER_97_376 ();
 sg13g2_fill_4 FILLER_97_384 ();
 sg13g2_fill_1 FILLER_97_388 ();
 sg13g2_fill_8 FILLER_97_413 ();
 sg13g2_fill_8 FILLER_97_421 ();
 sg13g2_fill_2 FILLER_97_429 ();
 sg13g2_fill_8 FILLER_97_438 ();
 sg13g2_fill_8 FILLER_97_446 ();
 sg13g2_fill_8 FILLER_97_454 ();
 sg13g2_fill_4 FILLER_97_469 ();
 sg13g2_fill_2 FILLER_97_482 ();
 sg13g2_fill_1 FILLER_97_484 ();
 sg13g2_fill_1 FILLER_97_563 ();
 sg13g2_fill_1 FILLER_97_570 ();
 sg13g2_fill_8 FILLER_97_597 ();
 sg13g2_fill_4 FILLER_97_605 ();
 sg13g2_fill_2 FILLER_97_609 ();
 sg13g2_fill_2 FILLER_97_621 ();
 sg13g2_fill_1 FILLER_97_623 ();
 sg13g2_fill_8 FILLER_97_627 ();
 sg13g2_fill_8 FILLER_97_635 ();
 sg13g2_fill_8 FILLER_97_643 ();
 sg13g2_fill_8 FILLER_97_651 ();
 sg13g2_fill_8 FILLER_97_659 ();
 sg13g2_fill_8 FILLER_97_667 ();
 sg13g2_fill_8 FILLER_97_675 ();
 sg13g2_fill_8 FILLER_97_683 ();
 sg13g2_fill_8 FILLER_97_691 ();
 sg13g2_fill_8 FILLER_97_699 ();
 sg13g2_fill_8 FILLER_97_707 ();
 sg13g2_fill_8 FILLER_97_715 ();
 sg13g2_fill_8 FILLER_97_723 ();
 sg13g2_fill_8 FILLER_97_731 ();
 sg13g2_fill_8 FILLER_97_739 ();
 sg13g2_fill_8 FILLER_97_747 ();
 sg13g2_fill_8 FILLER_97_755 ();
 sg13g2_fill_8 FILLER_97_763 ();
 sg13g2_fill_8 FILLER_97_771 ();
 sg13g2_fill_8 FILLER_97_779 ();
 sg13g2_fill_8 FILLER_97_787 ();
 sg13g2_fill_8 FILLER_97_795 ();
 sg13g2_fill_8 FILLER_97_803 ();
 sg13g2_fill_8 FILLER_97_811 ();
 sg13g2_fill_8 FILLER_97_819 ();
 sg13g2_fill_8 FILLER_97_827 ();
 sg13g2_fill_8 FILLER_97_835 ();
 sg13g2_fill_8 FILLER_97_843 ();
 sg13g2_fill_8 FILLER_97_851 ();
 sg13g2_fill_8 FILLER_97_859 ();
 sg13g2_fill_8 FILLER_97_867 ();
 sg13g2_fill_8 FILLER_97_875 ();
 sg13g2_fill_8 FILLER_97_883 ();
 sg13g2_fill_8 FILLER_97_891 ();
 sg13g2_fill_8 FILLER_97_899 ();
 sg13g2_fill_4 FILLER_97_907 ();
 sg13g2_fill_2 FILLER_97_911 ();
 sg13g2_fill_8 FILLER_97_923 ();
 sg13g2_fill_2 FILLER_97_931 ();
 sg13g2_fill_1 FILLER_97_933 ();
 sg13g2_fill_8 FILLER_97_955 ();
 sg13g2_fill_4 FILLER_97_963 ();
 sg13g2_fill_2 FILLER_97_978 ();
 sg13g2_fill_8 FILLER_97_990 ();
 sg13g2_fill_8 FILLER_97_998 ();
 sg13g2_fill_8 FILLER_97_1006 ();
 sg13g2_fill_8 FILLER_97_1014 ();
 sg13g2_fill_8 FILLER_97_1022 ();
 sg13g2_fill_8 FILLER_97_1030 ();
 sg13g2_fill_8 FILLER_97_1038 ();
 sg13g2_fill_8 FILLER_97_1046 ();
 sg13g2_fill_8 FILLER_97_1054 ();
 sg13g2_fill_8 FILLER_97_1062 ();
 sg13g2_fill_8 FILLER_97_1070 ();
 sg13g2_fill_8 FILLER_97_1078 ();
 sg13g2_fill_8 FILLER_97_1086 ();
 sg13g2_fill_8 FILLER_97_1094 ();
 sg13g2_fill_8 FILLER_97_1102 ();
 sg13g2_fill_8 FILLER_97_1110 ();
 sg13g2_fill_8 FILLER_97_1118 ();
 sg13g2_fill_8 FILLER_97_1126 ();
 sg13g2_fill_8 FILLER_97_1134 ();
 sg13g2_fill_8 FILLER_97_1142 ();
 sg13g2_fill_8 FILLER_97_1150 ();
 sg13g2_fill_8 FILLER_97_1158 ();
 sg13g2_fill_8 FILLER_98_0 ();
 sg13g2_fill_8 FILLER_98_8 ();
 sg13g2_fill_8 FILLER_98_16 ();
 sg13g2_fill_8 FILLER_98_24 ();
 sg13g2_fill_8 FILLER_98_32 ();
 sg13g2_fill_8 FILLER_98_40 ();
 sg13g2_fill_8 FILLER_98_48 ();
 sg13g2_fill_8 FILLER_98_56 ();
 sg13g2_fill_8 FILLER_98_64 ();
 sg13g2_fill_8 FILLER_98_72 ();
 sg13g2_fill_8 FILLER_98_80 ();
 sg13g2_fill_8 FILLER_98_88 ();
 sg13g2_fill_8 FILLER_98_96 ();
 sg13g2_fill_8 FILLER_98_104 ();
 sg13g2_fill_8 FILLER_98_112 ();
 sg13g2_fill_8 FILLER_98_120 ();
 sg13g2_fill_8 FILLER_98_128 ();
 sg13g2_fill_8 FILLER_98_136 ();
 sg13g2_fill_8 FILLER_98_144 ();
 sg13g2_fill_8 FILLER_98_152 ();
 sg13g2_fill_8 FILLER_98_160 ();
 sg13g2_fill_8 FILLER_98_168 ();
 sg13g2_fill_8 FILLER_98_176 ();
 sg13g2_fill_8 FILLER_98_184 ();
 sg13g2_fill_8 FILLER_98_192 ();
 sg13g2_fill_8 FILLER_98_200 ();
 sg13g2_fill_8 FILLER_98_208 ();
 sg13g2_fill_8 FILLER_98_216 ();
 sg13g2_fill_8 FILLER_98_224 ();
 sg13g2_fill_8 FILLER_98_232 ();
 sg13g2_fill_8 FILLER_98_240 ();
 sg13g2_fill_8 FILLER_98_248 ();
 sg13g2_fill_8 FILLER_98_256 ();
 sg13g2_fill_8 FILLER_98_264 ();
 sg13g2_fill_8 FILLER_98_272 ();
 sg13g2_fill_8 FILLER_98_280 ();
 sg13g2_fill_8 FILLER_98_288 ();
 sg13g2_fill_8 FILLER_98_296 ();
 sg13g2_fill_8 FILLER_98_304 ();
 sg13g2_fill_8 FILLER_98_312 ();
 sg13g2_fill_8 FILLER_98_320 ();
 sg13g2_fill_8 FILLER_98_328 ();
 sg13g2_fill_8 FILLER_98_336 ();
 sg13g2_fill_8 FILLER_98_344 ();
 sg13g2_fill_8 FILLER_98_352 ();
 sg13g2_fill_8 FILLER_98_360 ();
 sg13g2_fill_8 FILLER_98_368 ();
 sg13g2_fill_8 FILLER_98_376 ();
 sg13g2_fill_8 FILLER_98_384 ();
 sg13g2_fill_8 FILLER_98_392 ();
 sg13g2_fill_8 FILLER_98_400 ();
 sg13g2_fill_8 FILLER_98_408 ();
 sg13g2_fill_8 FILLER_98_416 ();
 sg13g2_fill_8 FILLER_98_424 ();
 sg13g2_fill_8 FILLER_98_432 ();
 sg13g2_fill_8 FILLER_98_440 ();
 sg13g2_fill_8 FILLER_98_448 ();
 sg13g2_fill_8 FILLER_98_456 ();
 sg13g2_fill_8 FILLER_98_464 ();
 sg13g2_fill_8 FILLER_98_472 ();
 sg13g2_fill_8 FILLER_98_480 ();
 sg13g2_fill_8 FILLER_98_488 ();
 sg13g2_fill_8 FILLER_98_496 ();
 sg13g2_fill_1 FILLER_98_504 ();
 sg13g2_fill_8 FILLER_98_511 ();
 sg13g2_fill_4 FILLER_98_519 ();
 sg13g2_fill_2 FILLER_98_529 ();
 sg13g2_fill_1 FILLER_98_531 ();
 sg13g2_fill_8 FILLER_98_555 ();
 sg13g2_fill_8 FILLER_98_563 ();
 sg13g2_fill_8 FILLER_98_571 ();
 sg13g2_fill_8 FILLER_98_579 ();
 sg13g2_fill_8 FILLER_98_587 ();
 sg13g2_fill_8 FILLER_98_595 ();
 sg13g2_fill_8 FILLER_98_603 ();
 sg13g2_fill_8 FILLER_98_611 ();
 sg13g2_fill_8 FILLER_98_619 ();
 sg13g2_fill_8 FILLER_98_627 ();
 sg13g2_fill_8 FILLER_98_635 ();
 sg13g2_fill_8 FILLER_98_643 ();
 sg13g2_fill_8 FILLER_98_651 ();
 sg13g2_fill_8 FILLER_98_659 ();
 sg13g2_fill_8 FILLER_98_667 ();
 sg13g2_fill_8 FILLER_98_675 ();
 sg13g2_fill_8 FILLER_98_683 ();
 sg13g2_fill_8 FILLER_98_691 ();
 sg13g2_fill_8 FILLER_98_699 ();
 sg13g2_fill_8 FILLER_98_707 ();
 sg13g2_fill_8 FILLER_98_715 ();
 sg13g2_fill_8 FILLER_98_723 ();
 sg13g2_fill_8 FILLER_98_731 ();
 sg13g2_fill_8 FILLER_98_739 ();
 sg13g2_fill_8 FILLER_98_747 ();
 sg13g2_fill_8 FILLER_98_755 ();
 sg13g2_fill_8 FILLER_98_763 ();
 sg13g2_fill_8 FILLER_98_771 ();
 sg13g2_fill_8 FILLER_98_779 ();
 sg13g2_fill_8 FILLER_98_787 ();
 sg13g2_fill_8 FILLER_98_795 ();
 sg13g2_fill_8 FILLER_98_803 ();
 sg13g2_fill_8 FILLER_98_811 ();
 sg13g2_fill_8 FILLER_98_819 ();
 sg13g2_fill_8 FILLER_98_827 ();
 sg13g2_fill_8 FILLER_98_835 ();
 sg13g2_fill_8 FILLER_98_843 ();
 sg13g2_fill_8 FILLER_98_851 ();
 sg13g2_fill_8 FILLER_98_859 ();
 sg13g2_fill_8 FILLER_98_867 ();
 sg13g2_fill_8 FILLER_98_875 ();
 sg13g2_fill_8 FILLER_98_883 ();
 sg13g2_fill_8 FILLER_98_891 ();
 sg13g2_fill_8 FILLER_98_899 ();
 sg13g2_fill_8 FILLER_98_907 ();
 sg13g2_fill_8 FILLER_98_915 ();
 sg13g2_fill_8 FILLER_98_923 ();
 sg13g2_fill_8 FILLER_98_931 ();
 sg13g2_fill_8 FILLER_98_939 ();
 sg13g2_fill_8 FILLER_98_947 ();
 sg13g2_fill_8 FILLER_98_955 ();
 sg13g2_fill_8 FILLER_98_963 ();
 sg13g2_fill_8 FILLER_98_971 ();
 sg13g2_fill_8 FILLER_98_979 ();
 sg13g2_fill_8 FILLER_98_987 ();
 sg13g2_fill_8 FILLER_98_995 ();
 sg13g2_fill_8 FILLER_98_1003 ();
 sg13g2_fill_8 FILLER_98_1011 ();
 sg13g2_fill_8 FILLER_98_1019 ();
 sg13g2_fill_8 FILLER_98_1027 ();
 sg13g2_fill_8 FILLER_98_1035 ();
 sg13g2_fill_8 FILLER_98_1043 ();
 sg13g2_fill_8 FILLER_98_1051 ();
 sg13g2_fill_8 FILLER_98_1059 ();
 sg13g2_fill_8 FILLER_98_1067 ();
 sg13g2_fill_8 FILLER_98_1075 ();
 sg13g2_fill_8 FILLER_98_1083 ();
 sg13g2_fill_8 FILLER_98_1091 ();
 sg13g2_fill_8 FILLER_98_1099 ();
 sg13g2_fill_8 FILLER_98_1107 ();
 sg13g2_fill_8 FILLER_98_1115 ();
 sg13g2_fill_8 FILLER_98_1123 ();
 sg13g2_fill_8 FILLER_98_1131 ();
 sg13g2_fill_8 FILLER_98_1139 ();
 sg13g2_fill_8 FILLER_98_1147 ();
 sg13g2_fill_8 FILLER_98_1155 ();
 sg13g2_fill_2 FILLER_98_1163 ();
 sg13g2_fill_1 FILLER_98_1165 ();
 sg13g2_fill_8 FILLER_99_0 ();
 sg13g2_fill_8 FILLER_99_8 ();
 sg13g2_fill_8 FILLER_99_16 ();
 sg13g2_fill_8 FILLER_99_24 ();
 sg13g2_fill_8 FILLER_99_32 ();
 sg13g2_fill_8 FILLER_99_40 ();
 sg13g2_fill_8 FILLER_99_48 ();
 sg13g2_fill_8 FILLER_99_56 ();
 sg13g2_fill_8 FILLER_99_64 ();
 sg13g2_fill_8 FILLER_99_72 ();
 sg13g2_fill_8 FILLER_99_80 ();
 sg13g2_fill_8 FILLER_99_88 ();
 sg13g2_fill_8 FILLER_99_96 ();
 sg13g2_fill_8 FILLER_99_104 ();
 sg13g2_fill_8 FILLER_99_112 ();
 sg13g2_fill_8 FILLER_99_120 ();
 sg13g2_fill_8 FILLER_99_128 ();
 sg13g2_fill_8 FILLER_99_136 ();
 sg13g2_fill_8 FILLER_99_144 ();
 sg13g2_fill_8 FILLER_99_152 ();
 sg13g2_fill_8 FILLER_99_160 ();
 sg13g2_fill_8 FILLER_99_168 ();
 sg13g2_fill_8 FILLER_99_176 ();
 sg13g2_fill_8 FILLER_99_184 ();
 sg13g2_fill_8 FILLER_99_192 ();
 sg13g2_fill_8 FILLER_99_200 ();
 sg13g2_fill_8 FILLER_99_208 ();
 sg13g2_fill_8 FILLER_99_216 ();
 sg13g2_fill_8 FILLER_99_224 ();
 sg13g2_fill_8 FILLER_99_232 ();
 sg13g2_fill_8 FILLER_99_240 ();
 sg13g2_fill_8 FILLER_99_248 ();
 sg13g2_fill_8 FILLER_99_256 ();
 sg13g2_fill_8 FILLER_99_264 ();
 sg13g2_fill_8 FILLER_99_272 ();
 sg13g2_fill_8 FILLER_99_280 ();
 sg13g2_fill_8 FILLER_99_288 ();
 sg13g2_fill_8 FILLER_99_296 ();
 sg13g2_fill_8 FILLER_99_304 ();
 sg13g2_fill_8 FILLER_99_312 ();
 sg13g2_fill_8 FILLER_99_320 ();
 sg13g2_fill_8 FILLER_99_328 ();
 sg13g2_fill_8 FILLER_99_336 ();
 sg13g2_fill_8 FILLER_99_344 ();
 sg13g2_fill_8 FILLER_99_352 ();
 sg13g2_fill_8 FILLER_99_360 ();
 sg13g2_fill_8 FILLER_99_368 ();
 sg13g2_fill_8 FILLER_99_376 ();
 sg13g2_fill_8 FILLER_99_384 ();
 sg13g2_fill_8 FILLER_99_392 ();
 sg13g2_fill_8 FILLER_99_400 ();
 sg13g2_fill_8 FILLER_99_408 ();
 sg13g2_fill_8 FILLER_99_416 ();
 sg13g2_fill_8 FILLER_99_424 ();
 sg13g2_fill_8 FILLER_99_432 ();
 sg13g2_fill_8 FILLER_99_440 ();
 sg13g2_fill_8 FILLER_99_448 ();
 sg13g2_fill_8 FILLER_99_456 ();
 sg13g2_fill_8 FILLER_99_464 ();
 sg13g2_fill_8 FILLER_99_472 ();
 sg13g2_fill_8 FILLER_99_480 ();
 sg13g2_fill_8 FILLER_99_488 ();
 sg13g2_fill_8 FILLER_99_496 ();
 sg13g2_fill_8 FILLER_99_504 ();
 sg13g2_fill_8 FILLER_99_512 ();
 sg13g2_fill_4 FILLER_99_520 ();
 sg13g2_fill_2 FILLER_99_524 ();
 sg13g2_fill_1 FILLER_99_526 ();
 sg13g2_fill_8 FILLER_99_532 ();
 sg13g2_fill_8 FILLER_99_540 ();
 sg13g2_fill_8 FILLER_99_548 ();
 sg13g2_fill_8 FILLER_99_556 ();
 sg13g2_fill_8 FILLER_99_564 ();
 sg13g2_fill_8 FILLER_99_572 ();
 sg13g2_fill_8 FILLER_99_580 ();
 sg13g2_fill_8 FILLER_99_588 ();
 sg13g2_fill_8 FILLER_99_596 ();
 sg13g2_fill_8 FILLER_99_604 ();
 sg13g2_fill_8 FILLER_99_612 ();
 sg13g2_fill_8 FILLER_99_620 ();
 sg13g2_fill_8 FILLER_99_628 ();
 sg13g2_fill_8 FILLER_99_636 ();
 sg13g2_fill_8 FILLER_99_644 ();
 sg13g2_fill_8 FILLER_99_652 ();
 sg13g2_fill_8 FILLER_99_660 ();
 sg13g2_fill_8 FILLER_99_668 ();
 sg13g2_fill_8 FILLER_99_676 ();
 sg13g2_fill_8 FILLER_99_684 ();
 sg13g2_fill_8 FILLER_99_692 ();
 sg13g2_fill_8 FILLER_99_700 ();
 sg13g2_fill_8 FILLER_99_708 ();
 sg13g2_fill_8 FILLER_99_716 ();
 sg13g2_fill_8 FILLER_99_724 ();
 sg13g2_fill_8 FILLER_99_732 ();
 sg13g2_fill_8 FILLER_99_740 ();
 sg13g2_fill_8 FILLER_99_748 ();
 sg13g2_fill_8 FILLER_99_756 ();
 sg13g2_fill_8 FILLER_99_764 ();
 sg13g2_fill_8 FILLER_99_772 ();
 sg13g2_fill_8 FILLER_99_780 ();
 sg13g2_fill_8 FILLER_99_788 ();
 sg13g2_fill_8 FILLER_99_796 ();
 sg13g2_fill_8 FILLER_99_804 ();
 sg13g2_fill_8 FILLER_99_812 ();
 sg13g2_fill_8 FILLER_99_820 ();
 sg13g2_fill_8 FILLER_99_828 ();
 sg13g2_fill_8 FILLER_99_836 ();
 sg13g2_fill_8 FILLER_99_844 ();
 sg13g2_fill_8 FILLER_99_852 ();
 sg13g2_fill_8 FILLER_99_860 ();
 sg13g2_fill_8 FILLER_99_868 ();
 sg13g2_fill_8 FILLER_99_876 ();
 sg13g2_fill_8 FILLER_99_884 ();
 sg13g2_fill_8 FILLER_99_892 ();
 sg13g2_fill_8 FILLER_99_900 ();
 sg13g2_fill_8 FILLER_99_908 ();
 sg13g2_fill_8 FILLER_99_916 ();
 sg13g2_fill_8 FILLER_99_924 ();
 sg13g2_fill_8 FILLER_99_932 ();
 sg13g2_fill_8 FILLER_99_940 ();
 sg13g2_fill_8 FILLER_99_948 ();
 sg13g2_fill_8 FILLER_99_956 ();
 sg13g2_fill_8 FILLER_99_964 ();
 sg13g2_fill_8 FILLER_99_972 ();
 sg13g2_fill_8 FILLER_99_980 ();
 sg13g2_fill_8 FILLER_99_988 ();
 sg13g2_fill_8 FILLER_99_996 ();
 sg13g2_fill_8 FILLER_99_1004 ();
 sg13g2_fill_8 FILLER_99_1012 ();
 sg13g2_fill_8 FILLER_99_1020 ();
 sg13g2_fill_8 FILLER_99_1028 ();
 sg13g2_fill_8 FILLER_99_1036 ();
 sg13g2_fill_8 FILLER_99_1044 ();
 sg13g2_fill_8 FILLER_99_1052 ();
 sg13g2_fill_8 FILLER_99_1060 ();
 sg13g2_fill_8 FILLER_99_1068 ();
 sg13g2_fill_8 FILLER_99_1076 ();
 sg13g2_fill_8 FILLER_99_1084 ();
 sg13g2_fill_8 FILLER_99_1092 ();
 sg13g2_fill_8 FILLER_99_1100 ();
 sg13g2_fill_8 FILLER_99_1108 ();
 sg13g2_fill_8 FILLER_99_1116 ();
 sg13g2_fill_8 FILLER_99_1124 ();
 sg13g2_fill_8 FILLER_99_1132 ();
 sg13g2_fill_8 FILLER_99_1140 ();
 sg13g2_fill_8 FILLER_99_1148 ();
 sg13g2_fill_8 FILLER_99_1156 ();
 sg13g2_fill_2 FILLER_99_1164 ();
 sg13g2_fill_8 FILLER_100_0 ();
 sg13g2_fill_8 FILLER_100_8 ();
 sg13g2_fill_8 FILLER_100_16 ();
 sg13g2_fill_8 FILLER_100_24 ();
 sg13g2_fill_8 FILLER_100_32 ();
 sg13g2_fill_8 FILLER_100_40 ();
 sg13g2_fill_8 FILLER_100_48 ();
 sg13g2_fill_8 FILLER_100_56 ();
 sg13g2_fill_8 FILLER_100_64 ();
 sg13g2_fill_8 FILLER_100_72 ();
 sg13g2_fill_8 FILLER_100_80 ();
 sg13g2_fill_8 FILLER_100_88 ();
 sg13g2_fill_8 FILLER_100_96 ();
 sg13g2_fill_8 FILLER_100_104 ();
 sg13g2_fill_8 FILLER_100_112 ();
 sg13g2_fill_8 FILLER_100_120 ();
 sg13g2_fill_8 FILLER_100_128 ();
 sg13g2_fill_8 FILLER_100_136 ();
 sg13g2_fill_8 FILLER_100_144 ();
 sg13g2_fill_8 FILLER_100_152 ();
 sg13g2_fill_8 FILLER_100_160 ();
 sg13g2_fill_8 FILLER_100_168 ();
 sg13g2_fill_8 FILLER_100_176 ();
 sg13g2_fill_8 FILLER_100_184 ();
 sg13g2_fill_8 FILLER_100_192 ();
 sg13g2_fill_8 FILLER_100_200 ();
 sg13g2_fill_8 FILLER_100_208 ();
 sg13g2_fill_8 FILLER_100_216 ();
 sg13g2_fill_8 FILLER_100_224 ();
 sg13g2_fill_8 FILLER_100_232 ();
 sg13g2_fill_8 FILLER_100_240 ();
 sg13g2_fill_8 FILLER_100_248 ();
 sg13g2_fill_8 FILLER_100_256 ();
 sg13g2_fill_8 FILLER_100_264 ();
 sg13g2_fill_8 FILLER_100_272 ();
 sg13g2_fill_8 FILLER_100_280 ();
 sg13g2_fill_8 FILLER_100_288 ();
 sg13g2_fill_8 FILLER_100_296 ();
 sg13g2_fill_8 FILLER_100_304 ();
 sg13g2_fill_8 FILLER_100_312 ();
 sg13g2_fill_8 FILLER_100_320 ();
 sg13g2_fill_8 FILLER_100_328 ();
 sg13g2_fill_8 FILLER_100_336 ();
 sg13g2_fill_8 FILLER_100_344 ();
 sg13g2_fill_8 FILLER_100_352 ();
 sg13g2_fill_8 FILLER_100_360 ();
 sg13g2_fill_8 FILLER_100_368 ();
 sg13g2_fill_8 FILLER_100_376 ();
 sg13g2_fill_8 FILLER_100_384 ();
 sg13g2_fill_8 FILLER_100_392 ();
 sg13g2_fill_8 FILLER_100_400 ();
 sg13g2_fill_8 FILLER_100_408 ();
 sg13g2_fill_8 FILLER_100_416 ();
 sg13g2_fill_8 FILLER_100_424 ();
 sg13g2_fill_8 FILLER_100_432 ();
 sg13g2_fill_8 FILLER_100_440 ();
 sg13g2_fill_8 FILLER_100_448 ();
 sg13g2_fill_8 FILLER_100_456 ();
 sg13g2_fill_8 FILLER_100_464 ();
 sg13g2_fill_8 FILLER_100_472 ();
 sg13g2_fill_8 FILLER_100_480 ();
 sg13g2_fill_8 FILLER_100_488 ();
 sg13g2_fill_8 FILLER_100_496 ();
 sg13g2_fill_8 FILLER_100_504 ();
 sg13g2_fill_8 FILLER_100_512 ();
 sg13g2_fill_8 FILLER_100_520 ();
 sg13g2_fill_8 FILLER_100_528 ();
 sg13g2_fill_8 FILLER_100_536 ();
 sg13g2_fill_8 FILLER_100_544 ();
 sg13g2_fill_8 FILLER_100_552 ();
 sg13g2_fill_8 FILLER_100_560 ();
 sg13g2_fill_8 FILLER_100_568 ();
 sg13g2_fill_8 FILLER_100_576 ();
 sg13g2_fill_8 FILLER_100_584 ();
 sg13g2_fill_8 FILLER_100_592 ();
 sg13g2_fill_8 FILLER_100_600 ();
 sg13g2_fill_8 FILLER_100_608 ();
 sg13g2_fill_8 FILLER_100_616 ();
 sg13g2_fill_8 FILLER_100_624 ();
 sg13g2_fill_8 FILLER_100_632 ();
 sg13g2_fill_8 FILLER_100_640 ();
 sg13g2_fill_8 FILLER_100_648 ();
 sg13g2_fill_8 FILLER_100_656 ();
 sg13g2_fill_8 FILLER_100_664 ();
 sg13g2_fill_8 FILLER_100_672 ();
 sg13g2_fill_8 FILLER_100_680 ();
 sg13g2_fill_8 FILLER_100_688 ();
 sg13g2_fill_8 FILLER_100_696 ();
 sg13g2_fill_8 FILLER_100_704 ();
 sg13g2_fill_8 FILLER_100_712 ();
 sg13g2_fill_8 FILLER_100_720 ();
 sg13g2_fill_8 FILLER_100_728 ();
 sg13g2_fill_8 FILLER_100_736 ();
 sg13g2_fill_8 FILLER_100_744 ();
 sg13g2_fill_8 FILLER_100_752 ();
 sg13g2_fill_8 FILLER_100_760 ();
 sg13g2_fill_8 FILLER_100_768 ();
 sg13g2_fill_8 FILLER_100_776 ();
 sg13g2_fill_8 FILLER_100_784 ();
 sg13g2_fill_8 FILLER_100_792 ();
 sg13g2_fill_8 FILLER_100_800 ();
 sg13g2_fill_8 FILLER_100_808 ();
 sg13g2_fill_8 FILLER_100_816 ();
 sg13g2_fill_8 FILLER_100_824 ();
 sg13g2_fill_8 FILLER_100_832 ();
 sg13g2_fill_8 FILLER_100_840 ();
 sg13g2_fill_8 FILLER_100_848 ();
 sg13g2_fill_8 FILLER_100_856 ();
 sg13g2_fill_8 FILLER_100_864 ();
 sg13g2_fill_8 FILLER_100_872 ();
 sg13g2_fill_8 FILLER_100_880 ();
 sg13g2_fill_8 FILLER_100_888 ();
 sg13g2_fill_8 FILLER_100_896 ();
 sg13g2_fill_8 FILLER_100_904 ();
 sg13g2_fill_8 FILLER_100_912 ();
 sg13g2_fill_8 FILLER_100_920 ();
 sg13g2_fill_8 FILLER_100_928 ();
 sg13g2_fill_8 FILLER_100_936 ();
 sg13g2_fill_8 FILLER_100_944 ();
 sg13g2_fill_8 FILLER_100_952 ();
 sg13g2_fill_8 FILLER_100_960 ();
 sg13g2_fill_8 FILLER_100_968 ();
 sg13g2_fill_8 FILLER_100_976 ();
 sg13g2_fill_8 FILLER_100_984 ();
 sg13g2_fill_8 FILLER_100_992 ();
 sg13g2_fill_8 FILLER_100_1000 ();
 sg13g2_fill_8 FILLER_100_1008 ();
 sg13g2_fill_8 FILLER_100_1016 ();
 sg13g2_fill_8 FILLER_100_1024 ();
 sg13g2_fill_8 FILLER_100_1032 ();
 sg13g2_fill_8 FILLER_100_1040 ();
 sg13g2_fill_8 FILLER_100_1048 ();
 sg13g2_fill_8 FILLER_100_1056 ();
 sg13g2_fill_8 FILLER_100_1064 ();
 sg13g2_fill_8 FILLER_100_1072 ();
 sg13g2_fill_8 FILLER_100_1080 ();
 sg13g2_fill_8 FILLER_100_1088 ();
 sg13g2_fill_8 FILLER_100_1096 ();
 sg13g2_fill_8 FILLER_100_1104 ();
 sg13g2_fill_8 FILLER_100_1112 ();
 sg13g2_fill_8 FILLER_100_1120 ();
 sg13g2_fill_8 FILLER_100_1128 ();
 sg13g2_fill_8 FILLER_100_1136 ();
 sg13g2_fill_8 FILLER_100_1144 ();
 sg13g2_fill_8 FILLER_100_1152 ();
 sg13g2_fill_4 FILLER_100_1160 ();
 sg13g2_fill_2 FILLER_100_1164 ();
 sg13g2_fill_8 FILLER_101_0 ();
 sg13g2_fill_8 FILLER_101_8 ();
 sg13g2_fill_8 FILLER_101_16 ();
 sg13g2_fill_8 FILLER_101_24 ();
 sg13g2_fill_8 FILLER_101_32 ();
 sg13g2_fill_8 FILLER_101_40 ();
 sg13g2_fill_8 FILLER_101_48 ();
 sg13g2_fill_8 FILLER_101_56 ();
 sg13g2_fill_8 FILLER_101_64 ();
 sg13g2_fill_8 FILLER_101_72 ();
 sg13g2_fill_8 FILLER_101_80 ();
 sg13g2_fill_8 FILLER_101_88 ();
 sg13g2_fill_8 FILLER_101_96 ();
 sg13g2_fill_8 FILLER_101_104 ();
 sg13g2_fill_8 FILLER_101_112 ();
 sg13g2_fill_8 FILLER_101_120 ();
 sg13g2_fill_8 FILLER_101_128 ();
 sg13g2_fill_8 FILLER_101_136 ();
 sg13g2_fill_8 FILLER_101_144 ();
 sg13g2_fill_8 FILLER_101_152 ();
 sg13g2_fill_8 FILLER_101_160 ();
 sg13g2_fill_8 FILLER_101_168 ();
 sg13g2_fill_8 FILLER_101_176 ();
 sg13g2_fill_8 FILLER_101_184 ();
 sg13g2_fill_8 FILLER_101_192 ();
 sg13g2_fill_8 FILLER_101_200 ();
 sg13g2_fill_8 FILLER_101_208 ();
 sg13g2_fill_8 FILLER_101_216 ();
 sg13g2_fill_8 FILLER_101_224 ();
 sg13g2_fill_8 FILLER_101_232 ();
 sg13g2_fill_8 FILLER_101_240 ();
 sg13g2_fill_8 FILLER_101_248 ();
 sg13g2_fill_8 FILLER_101_256 ();
 sg13g2_fill_8 FILLER_101_264 ();
 sg13g2_fill_8 FILLER_101_272 ();
 sg13g2_fill_8 FILLER_101_280 ();
 sg13g2_fill_8 FILLER_101_288 ();
 sg13g2_fill_8 FILLER_101_296 ();
 sg13g2_fill_8 FILLER_101_304 ();
 sg13g2_fill_8 FILLER_101_312 ();
 sg13g2_fill_8 FILLER_101_320 ();
 sg13g2_fill_8 FILLER_101_328 ();
 sg13g2_fill_8 FILLER_101_336 ();
 sg13g2_fill_8 FILLER_101_344 ();
 sg13g2_fill_8 FILLER_101_352 ();
 sg13g2_fill_8 FILLER_101_360 ();
 sg13g2_fill_8 FILLER_101_368 ();
 sg13g2_fill_8 FILLER_101_376 ();
 sg13g2_fill_8 FILLER_101_384 ();
 sg13g2_fill_8 FILLER_101_392 ();
 sg13g2_fill_8 FILLER_101_400 ();
 sg13g2_fill_8 FILLER_101_408 ();
 sg13g2_fill_8 FILLER_101_416 ();
 sg13g2_fill_8 FILLER_101_424 ();
 sg13g2_fill_8 FILLER_101_432 ();
 sg13g2_fill_8 FILLER_101_440 ();
 sg13g2_fill_8 FILLER_101_448 ();
 sg13g2_fill_8 FILLER_101_456 ();
 sg13g2_fill_8 FILLER_101_464 ();
 sg13g2_fill_8 FILLER_101_472 ();
 sg13g2_fill_8 FILLER_101_480 ();
 sg13g2_fill_8 FILLER_101_488 ();
 sg13g2_fill_8 FILLER_101_496 ();
 sg13g2_fill_8 FILLER_101_504 ();
 sg13g2_fill_8 FILLER_101_512 ();
 sg13g2_fill_8 FILLER_101_520 ();
 sg13g2_fill_8 FILLER_101_528 ();
 sg13g2_fill_8 FILLER_101_536 ();
 sg13g2_fill_8 FILLER_101_544 ();
 sg13g2_fill_8 FILLER_101_552 ();
 sg13g2_fill_8 FILLER_101_560 ();
 sg13g2_fill_8 FILLER_101_568 ();
 sg13g2_fill_8 FILLER_101_576 ();
 sg13g2_fill_8 FILLER_101_584 ();
 sg13g2_fill_8 FILLER_101_592 ();
 sg13g2_fill_8 FILLER_101_600 ();
 sg13g2_fill_8 FILLER_101_608 ();
 sg13g2_fill_8 FILLER_101_616 ();
 sg13g2_fill_8 FILLER_101_624 ();
 sg13g2_fill_8 FILLER_101_632 ();
 sg13g2_fill_8 FILLER_101_640 ();
 sg13g2_fill_8 FILLER_101_648 ();
 sg13g2_fill_8 FILLER_101_656 ();
 sg13g2_fill_8 FILLER_101_664 ();
 sg13g2_fill_8 FILLER_101_672 ();
 sg13g2_fill_8 FILLER_101_680 ();
 sg13g2_fill_8 FILLER_101_688 ();
 sg13g2_fill_8 FILLER_101_696 ();
 sg13g2_fill_8 FILLER_101_704 ();
 sg13g2_fill_8 FILLER_101_712 ();
 sg13g2_fill_8 FILLER_101_720 ();
 sg13g2_fill_8 FILLER_101_728 ();
 sg13g2_fill_8 FILLER_101_736 ();
 sg13g2_fill_8 FILLER_101_744 ();
 sg13g2_fill_8 FILLER_101_752 ();
 sg13g2_fill_8 FILLER_101_760 ();
 sg13g2_fill_8 FILLER_101_768 ();
 sg13g2_fill_8 FILLER_101_776 ();
 sg13g2_fill_8 FILLER_101_784 ();
 sg13g2_fill_8 FILLER_101_792 ();
 sg13g2_fill_8 FILLER_101_800 ();
 sg13g2_fill_8 FILLER_101_808 ();
 sg13g2_fill_8 FILLER_101_816 ();
 sg13g2_fill_8 FILLER_101_824 ();
 sg13g2_fill_8 FILLER_101_832 ();
 sg13g2_fill_8 FILLER_101_840 ();
 sg13g2_fill_8 FILLER_101_848 ();
 sg13g2_fill_8 FILLER_101_856 ();
 sg13g2_fill_8 FILLER_101_864 ();
 sg13g2_fill_8 FILLER_101_872 ();
 sg13g2_fill_8 FILLER_101_880 ();
 sg13g2_fill_8 FILLER_101_888 ();
 sg13g2_fill_8 FILLER_101_896 ();
 sg13g2_fill_8 FILLER_101_904 ();
 sg13g2_fill_8 FILLER_101_912 ();
 sg13g2_fill_8 FILLER_101_920 ();
 sg13g2_fill_8 FILLER_101_928 ();
 sg13g2_fill_8 FILLER_101_936 ();
 sg13g2_fill_8 FILLER_101_944 ();
 sg13g2_fill_8 FILLER_101_952 ();
 sg13g2_fill_8 FILLER_101_960 ();
 sg13g2_fill_8 FILLER_101_968 ();
 sg13g2_fill_8 FILLER_101_976 ();
 sg13g2_fill_8 FILLER_101_984 ();
 sg13g2_fill_8 FILLER_101_992 ();
 sg13g2_fill_8 FILLER_101_1000 ();
 sg13g2_fill_8 FILLER_101_1008 ();
 sg13g2_fill_8 FILLER_101_1016 ();
 sg13g2_fill_8 FILLER_101_1024 ();
 sg13g2_fill_8 FILLER_101_1032 ();
 sg13g2_fill_8 FILLER_101_1040 ();
 sg13g2_fill_8 FILLER_101_1048 ();
 sg13g2_fill_8 FILLER_101_1056 ();
 sg13g2_fill_8 FILLER_101_1064 ();
 sg13g2_fill_8 FILLER_101_1072 ();
 sg13g2_fill_8 FILLER_101_1080 ();
 sg13g2_fill_8 FILLER_101_1088 ();
 sg13g2_fill_8 FILLER_101_1096 ();
 sg13g2_fill_8 FILLER_101_1104 ();
 sg13g2_fill_8 FILLER_101_1112 ();
 sg13g2_fill_8 FILLER_101_1120 ();
 sg13g2_fill_8 FILLER_101_1128 ();
 sg13g2_fill_8 FILLER_101_1136 ();
 sg13g2_fill_8 FILLER_101_1144 ();
 sg13g2_fill_8 FILLER_101_1152 ();
 sg13g2_fill_4 FILLER_101_1160 ();
 sg13g2_fill_2 FILLER_101_1164 ();
 sg13g2_fill_8 FILLER_102_0 ();
 sg13g2_fill_8 FILLER_102_8 ();
 sg13g2_fill_8 FILLER_102_16 ();
 sg13g2_fill_8 FILLER_102_24 ();
 sg13g2_fill_8 FILLER_102_32 ();
 sg13g2_fill_8 FILLER_102_40 ();
 sg13g2_fill_8 FILLER_102_48 ();
 sg13g2_fill_8 FILLER_102_56 ();
 sg13g2_fill_8 FILLER_102_64 ();
 sg13g2_fill_8 FILLER_102_72 ();
 sg13g2_fill_8 FILLER_102_80 ();
 sg13g2_fill_8 FILLER_102_88 ();
 sg13g2_fill_8 FILLER_102_96 ();
 sg13g2_fill_8 FILLER_102_104 ();
 sg13g2_fill_8 FILLER_102_112 ();
 sg13g2_fill_8 FILLER_102_120 ();
 sg13g2_fill_8 FILLER_102_128 ();
 sg13g2_fill_8 FILLER_102_136 ();
 sg13g2_fill_8 FILLER_102_144 ();
 sg13g2_fill_8 FILLER_102_152 ();
 sg13g2_fill_8 FILLER_102_160 ();
 sg13g2_fill_8 FILLER_102_168 ();
 sg13g2_fill_8 FILLER_102_176 ();
 sg13g2_fill_8 FILLER_102_184 ();
 sg13g2_fill_8 FILLER_102_192 ();
 sg13g2_fill_8 FILLER_102_200 ();
 sg13g2_fill_8 FILLER_102_208 ();
 sg13g2_fill_8 FILLER_102_216 ();
 sg13g2_fill_8 FILLER_102_224 ();
 sg13g2_fill_8 FILLER_102_232 ();
 sg13g2_fill_8 FILLER_102_240 ();
 sg13g2_fill_8 FILLER_102_248 ();
 sg13g2_fill_8 FILLER_102_256 ();
 sg13g2_fill_8 FILLER_102_264 ();
 sg13g2_fill_8 FILLER_102_272 ();
 sg13g2_fill_8 FILLER_102_280 ();
 sg13g2_fill_8 FILLER_102_288 ();
 sg13g2_fill_8 FILLER_102_296 ();
 sg13g2_fill_8 FILLER_102_304 ();
 sg13g2_fill_8 FILLER_102_312 ();
 sg13g2_fill_8 FILLER_102_320 ();
 sg13g2_fill_8 FILLER_102_328 ();
 sg13g2_fill_8 FILLER_102_336 ();
 sg13g2_fill_8 FILLER_102_344 ();
 sg13g2_fill_8 FILLER_102_352 ();
 sg13g2_fill_8 FILLER_102_360 ();
 sg13g2_fill_8 FILLER_102_368 ();
 sg13g2_fill_8 FILLER_102_376 ();
 sg13g2_fill_8 FILLER_102_384 ();
 sg13g2_fill_8 FILLER_102_392 ();
 sg13g2_fill_8 FILLER_102_400 ();
 sg13g2_fill_8 FILLER_102_408 ();
 sg13g2_fill_8 FILLER_102_416 ();
 sg13g2_fill_8 FILLER_102_424 ();
 sg13g2_fill_8 FILLER_102_432 ();
 sg13g2_fill_8 FILLER_102_440 ();
 sg13g2_fill_8 FILLER_102_448 ();
 sg13g2_fill_8 FILLER_102_456 ();
 sg13g2_fill_8 FILLER_102_464 ();
 sg13g2_fill_8 FILLER_102_472 ();
 sg13g2_fill_8 FILLER_102_480 ();
 sg13g2_fill_8 FILLER_102_488 ();
 sg13g2_fill_8 FILLER_102_496 ();
 sg13g2_fill_8 FILLER_102_504 ();
 sg13g2_fill_8 FILLER_102_512 ();
 sg13g2_fill_8 FILLER_102_520 ();
 sg13g2_fill_8 FILLER_102_528 ();
 sg13g2_fill_8 FILLER_102_536 ();
 sg13g2_fill_8 FILLER_102_544 ();
 sg13g2_fill_8 FILLER_102_552 ();
 sg13g2_fill_8 FILLER_102_560 ();
 sg13g2_fill_8 FILLER_102_568 ();
 sg13g2_fill_8 FILLER_102_576 ();
 sg13g2_fill_8 FILLER_102_584 ();
 sg13g2_fill_8 FILLER_102_592 ();
 sg13g2_fill_8 FILLER_102_600 ();
 sg13g2_fill_8 FILLER_102_608 ();
 sg13g2_fill_8 FILLER_102_616 ();
 sg13g2_fill_8 FILLER_102_624 ();
 sg13g2_fill_8 FILLER_102_632 ();
 sg13g2_fill_8 FILLER_102_640 ();
 sg13g2_fill_8 FILLER_102_648 ();
 sg13g2_fill_8 FILLER_102_656 ();
 sg13g2_fill_8 FILLER_102_664 ();
 sg13g2_fill_8 FILLER_102_672 ();
 sg13g2_fill_8 FILLER_102_680 ();
 sg13g2_fill_8 FILLER_102_688 ();
 sg13g2_fill_8 FILLER_102_696 ();
 sg13g2_fill_8 FILLER_102_704 ();
 sg13g2_fill_8 FILLER_102_712 ();
 sg13g2_fill_8 FILLER_102_720 ();
 sg13g2_fill_8 FILLER_102_728 ();
 sg13g2_fill_8 FILLER_102_736 ();
 sg13g2_fill_8 FILLER_102_744 ();
 sg13g2_fill_8 FILLER_102_752 ();
 sg13g2_fill_8 FILLER_102_760 ();
 sg13g2_fill_8 FILLER_102_768 ();
 sg13g2_fill_8 FILLER_102_776 ();
 sg13g2_fill_8 FILLER_102_784 ();
 sg13g2_fill_8 FILLER_102_792 ();
 sg13g2_fill_8 FILLER_102_800 ();
 sg13g2_fill_8 FILLER_102_808 ();
 sg13g2_fill_8 FILLER_102_816 ();
 sg13g2_fill_8 FILLER_102_824 ();
 sg13g2_fill_8 FILLER_102_832 ();
 sg13g2_fill_8 FILLER_102_840 ();
 sg13g2_fill_8 FILLER_102_848 ();
 sg13g2_fill_8 FILLER_102_856 ();
 sg13g2_fill_8 FILLER_102_864 ();
 sg13g2_fill_8 FILLER_102_872 ();
 sg13g2_fill_8 FILLER_102_880 ();
 sg13g2_fill_8 FILLER_102_888 ();
 sg13g2_fill_8 FILLER_102_896 ();
 sg13g2_fill_8 FILLER_102_904 ();
 sg13g2_fill_8 FILLER_102_912 ();
 sg13g2_fill_8 FILLER_102_920 ();
 sg13g2_fill_8 FILLER_102_928 ();
 sg13g2_fill_8 FILLER_102_936 ();
 sg13g2_fill_8 FILLER_102_944 ();
 sg13g2_fill_8 FILLER_102_952 ();
 sg13g2_fill_8 FILLER_102_960 ();
 sg13g2_fill_8 FILLER_102_968 ();
 sg13g2_fill_8 FILLER_102_976 ();
 sg13g2_fill_8 FILLER_102_984 ();
 sg13g2_fill_8 FILLER_102_992 ();
 sg13g2_fill_8 FILLER_102_1000 ();
 sg13g2_fill_8 FILLER_102_1008 ();
 sg13g2_fill_8 FILLER_102_1016 ();
 sg13g2_fill_8 FILLER_102_1024 ();
 sg13g2_fill_8 FILLER_102_1032 ();
 sg13g2_fill_8 FILLER_102_1040 ();
 sg13g2_fill_8 FILLER_102_1048 ();
 sg13g2_fill_8 FILLER_102_1056 ();
 sg13g2_fill_8 FILLER_102_1064 ();
 sg13g2_fill_8 FILLER_102_1072 ();
 sg13g2_fill_8 FILLER_102_1080 ();
 sg13g2_fill_8 FILLER_102_1088 ();
 sg13g2_fill_8 FILLER_102_1096 ();
 sg13g2_fill_8 FILLER_102_1104 ();
 sg13g2_fill_8 FILLER_102_1112 ();
 sg13g2_fill_8 FILLER_102_1120 ();
 sg13g2_fill_8 FILLER_102_1128 ();
 sg13g2_fill_8 FILLER_102_1136 ();
 sg13g2_fill_8 FILLER_102_1144 ();
 sg13g2_fill_8 FILLER_102_1152 ();
 sg13g2_fill_4 FILLER_102_1160 ();
 sg13g2_fill_2 FILLER_102_1164 ();
 sg13g2_fill_8 FILLER_103_0 ();
 sg13g2_fill_8 FILLER_103_8 ();
 sg13g2_fill_8 FILLER_103_16 ();
 sg13g2_fill_8 FILLER_103_24 ();
 sg13g2_fill_8 FILLER_103_32 ();
 sg13g2_fill_8 FILLER_103_40 ();
 sg13g2_fill_8 FILLER_103_48 ();
 sg13g2_fill_8 FILLER_103_56 ();
 sg13g2_fill_8 FILLER_103_64 ();
 sg13g2_fill_8 FILLER_103_72 ();
 sg13g2_fill_8 FILLER_103_80 ();
 sg13g2_fill_8 FILLER_103_88 ();
 sg13g2_fill_8 FILLER_103_96 ();
 sg13g2_fill_8 FILLER_103_104 ();
 sg13g2_fill_8 FILLER_103_112 ();
 sg13g2_fill_8 FILLER_103_120 ();
 sg13g2_fill_8 FILLER_103_128 ();
 sg13g2_fill_8 FILLER_103_136 ();
 sg13g2_fill_8 FILLER_103_144 ();
 sg13g2_fill_8 FILLER_103_152 ();
 sg13g2_fill_8 FILLER_103_160 ();
 sg13g2_fill_8 FILLER_103_168 ();
 sg13g2_fill_8 FILLER_103_176 ();
 sg13g2_fill_8 FILLER_103_184 ();
 sg13g2_fill_8 FILLER_103_192 ();
 sg13g2_fill_8 FILLER_103_200 ();
 sg13g2_fill_8 FILLER_103_208 ();
 sg13g2_fill_8 FILLER_103_216 ();
 sg13g2_fill_8 FILLER_103_224 ();
 sg13g2_fill_8 FILLER_103_232 ();
 sg13g2_fill_8 FILLER_103_240 ();
 sg13g2_fill_8 FILLER_103_248 ();
 sg13g2_fill_8 FILLER_103_256 ();
 sg13g2_fill_8 FILLER_103_264 ();
 sg13g2_fill_8 FILLER_103_272 ();
 sg13g2_fill_8 FILLER_103_280 ();
 sg13g2_fill_8 FILLER_103_288 ();
 sg13g2_fill_8 FILLER_103_296 ();
 sg13g2_fill_8 FILLER_103_304 ();
 sg13g2_fill_8 FILLER_103_312 ();
 sg13g2_fill_8 FILLER_103_320 ();
 sg13g2_fill_8 FILLER_103_328 ();
 sg13g2_fill_8 FILLER_103_336 ();
 sg13g2_fill_8 FILLER_103_344 ();
 sg13g2_fill_8 FILLER_103_352 ();
 sg13g2_fill_8 FILLER_103_360 ();
 sg13g2_fill_8 FILLER_103_368 ();
 sg13g2_fill_8 FILLER_103_376 ();
 sg13g2_fill_8 FILLER_103_384 ();
 sg13g2_fill_8 FILLER_103_392 ();
 sg13g2_fill_8 FILLER_103_400 ();
 sg13g2_fill_8 FILLER_103_408 ();
 sg13g2_fill_8 FILLER_103_416 ();
 sg13g2_fill_8 FILLER_103_424 ();
 sg13g2_fill_8 FILLER_103_432 ();
 sg13g2_fill_8 FILLER_103_440 ();
 sg13g2_fill_8 FILLER_103_448 ();
 sg13g2_fill_8 FILLER_103_456 ();
 sg13g2_fill_8 FILLER_103_464 ();
 sg13g2_fill_8 FILLER_103_472 ();
 sg13g2_fill_8 FILLER_103_480 ();
 sg13g2_fill_8 FILLER_103_488 ();
 sg13g2_fill_8 FILLER_103_496 ();
 sg13g2_fill_8 FILLER_103_504 ();
 sg13g2_fill_8 FILLER_103_512 ();
 sg13g2_fill_8 FILLER_103_520 ();
 sg13g2_fill_8 FILLER_103_528 ();
 sg13g2_fill_8 FILLER_103_536 ();
 sg13g2_fill_8 FILLER_103_544 ();
 sg13g2_fill_8 FILLER_103_552 ();
 sg13g2_fill_8 FILLER_103_560 ();
 sg13g2_fill_8 FILLER_103_568 ();
 sg13g2_fill_8 FILLER_103_576 ();
 sg13g2_fill_8 FILLER_103_584 ();
 sg13g2_fill_8 FILLER_103_592 ();
 sg13g2_fill_8 FILLER_103_600 ();
 sg13g2_fill_8 FILLER_103_608 ();
 sg13g2_fill_8 FILLER_103_616 ();
 sg13g2_fill_8 FILLER_103_624 ();
 sg13g2_fill_8 FILLER_103_632 ();
 sg13g2_fill_8 FILLER_103_640 ();
 sg13g2_fill_8 FILLER_103_648 ();
 sg13g2_fill_8 FILLER_103_656 ();
 sg13g2_fill_8 FILLER_103_664 ();
 sg13g2_fill_8 FILLER_103_672 ();
 sg13g2_fill_8 FILLER_103_680 ();
 sg13g2_fill_8 FILLER_103_688 ();
 sg13g2_fill_8 FILLER_103_696 ();
 sg13g2_fill_8 FILLER_103_704 ();
 sg13g2_fill_8 FILLER_103_712 ();
 sg13g2_fill_8 FILLER_103_720 ();
 sg13g2_fill_8 FILLER_103_728 ();
 sg13g2_fill_8 FILLER_103_736 ();
 sg13g2_fill_8 FILLER_103_744 ();
 sg13g2_fill_8 FILLER_103_752 ();
 sg13g2_fill_8 FILLER_103_760 ();
 sg13g2_fill_8 FILLER_103_768 ();
 sg13g2_fill_8 FILLER_103_776 ();
 sg13g2_fill_8 FILLER_103_784 ();
 sg13g2_fill_8 FILLER_103_792 ();
 sg13g2_fill_8 FILLER_103_800 ();
 sg13g2_fill_8 FILLER_103_808 ();
 sg13g2_fill_8 FILLER_103_816 ();
 sg13g2_fill_8 FILLER_103_824 ();
 sg13g2_fill_8 FILLER_103_832 ();
 sg13g2_fill_8 FILLER_103_840 ();
 sg13g2_fill_8 FILLER_103_848 ();
 sg13g2_fill_8 FILLER_103_856 ();
 sg13g2_fill_8 FILLER_103_864 ();
 sg13g2_fill_8 FILLER_103_872 ();
 sg13g2_fill_8 FILLER_103_880 ();
 sg13g2_fill_8 FILLER_103_888 ();
 sg13g2_fill_8 FILLER_103_896 ();
 sg13g2_fill_8 FILLER_103_904 ();
 sg13g2_fill_8 FILLER_103_912 ();
 sg13g2_fill_8 FILLER_103_920 ();
 sg13g2_fill_8 FILLER_103_928 ();
 sg13g2_fill_8 FILLER_103_936 ();
 sg13g2_fill_8 FILLER_103_944 ();
 sg13g2_fill_8 FILLER_103_952 ();
 sg13g2_fill_8 FILLER_103_960 ();
 sg13g2_fill_8 FILLER_103_968 ();
 sg13g2_fill_8 FILLER_103_976 ();
 sg13g2_fill_8 FILLER_103_984 ();
 sg13g2_fill_8 FILLER_103_992 ();
 sg13g2_fill_8 FILLER_103_1000 ();
 sg13g2_fill_8 FILLER_103_1008 ();
 sg13g2_fill_8 FILLER_103_1016 ();
 sg13g2_fill_8 FILLER_103_1024 ();
 sg13g2_fill_8 FILLER_103_1032 ();
 sg13g2_fill_8 FILLER_103_1040 ();
 sg13g2_fill_8 FILLER_103_1048 ();
 sg13g2_fill_8 FILLER_103_1056 ();
 sg13g2_fill_8 FILLER_103_1064 ();
 sg13g2_fill_8 FILLER_103_1072 ();
 sg13g2_fill_8 FILLER_103_1080 ();
 sg13g2_fill_8 FILLER_103_1088 ();
 sg13g2_fill_8 FILLER_103_1096 ();
 sg13g2_fill_8 FILLER_103_1104 ();
 sg13g2_fill_8 FILLER_103_1112 ();
 sg13g2_fill_8 FILLER_103_1120 ();
 sg13g2_fill_8 FILLER_103_1128 ();
 sg13g2_fill_8 FILLER_103_1136 ();
 sg13g2_fill_8 FILLER_103_1144 ();
 sg13g2_fill_8 FILLER_103_1152 ();
 sg13g2_fill_4 FILLER_103_1160 ();
 sg13g2_fill_2 FILLER_103_1164 ();
 sg13g2_fill_8 FILLER_104_0 ();
 sg13g2_fill_8 FILLER_104_8 ();
 sg13g2_fill_8 FILLER_104_16 ();
 sg13g2_fill_8 FILLER_104_24 ();
 sg13g2_fill_8 FILLER_104_32 ();
 sg13g2_fill_8 FILLER_104_40 ();
 sg13g2_fill_8 FILLER_104_48 ();
 sg13g2_fill_8 FILLER_104_56 ();
 sg13g2_fill_8 FILLER_104_64 ();
 sg13g2_fill_8 FILLER_104_72 ();
 sg13g2_fill_8 FILLER_104_80 ();
 sg13g2_fill_8 FILLER_104_88 ();
 sg13g2_fill_8 FILLER_104_96 ();
 sg13g2_fill_8 FILLER_104_104 ();
 sg13g2_fill_8 FILLER_104_112 ();
 sg13g2_fill_8 FILLER_104_120 ();
 sg13g2_fill_8 FILLER_104_128 ();
 sg13g2_fill_8 FILLER_104_136 ();
 sg13g2_fill_8 FILLER_104_144 ();
 sg13g2_fill_8 FILLER_104_152 ();
 sg13g2_fill_8 FILLER_104_160 ();
 sg13g2_fill_8 FILLER_104_168 ();
 sg13g2_fill_8 FILLER_104_176 ();
 sg13g2_fill_8 FILLER_104_184 ();
 sg13g2_fill_8 FILLER_104_192 ();
 sg13g2_fill_8 FILLER_104_200 ();
 sg13g2_fill_8 FILLER_104_208 ();
 sg13g2_fill_8 FILLER_104_216 ();
 sg13g2_fill_8 FILLER_104_224 ();
 sg13g2_fill_8 FILLER_104_232 ();
 sg13g2_fill_8 FILLER_104_240 ();
 sg13g2_fill_8 FILLER_104_248 ();
 sg13g2_fill_8 FILLER_104_256 ();
 sg13g2_fill_8 FILLER_104_264 ();
 sg13g2_fill_8 FILLER_104_272 ();
 sg13g2_fill_8 FILLER_104_280 ();
 sg13g2_fill_8 FILLER_104_288 ();
 sg13g2_fill_8 FILLER_104_296 ();
 sg13g2_fill_8 FILLER_104_304 ();
 sg13g2_fill_8 FILLER_104_312 ();
 sg13g2_fill_8 FILLER_104_320 ();
 sg13g2_fill_8 FILLER_104_328 ();
 sg13g2_fill_8 FILLER_104_336 ();
 sg13g2_fill_8 FILLER_104_344 ();
 sg13g2_fill_8 FILLER_104_352 ();
 sg13g2_fill_8 FILLER_104_360 ();
 sg13g2_fill_8 FILLER_104_368 ();
 sg13g2_fill_8 FILLER_104_376 ();
 sg13g2_fill_8 FILLER_104_384 ();
 sg13g2_fill_8 FILLER_104_392 ();
 sg13g2_fill_8 FILLER_104_400 ();
 sg13g2_fill_8 FILLER_104_408 ();
 sg13g2_fill_8 FILLER_104_416 ();
 sg13g2_fill_8 FILLER_104_424 ();
 sg13g2_fill_8 FILLER_104_432 ();
 sg13g2_fill_8 FILLER_104_440 ();
 sg13g2_fill_8 FILLER_104_448 ();
 sg13g2_fill_8 FILLER_104_456 ();
 sg13g2_fill_8 FILLER_104_464 ();
 sg13g2_fill_8 FILLER_104_472 ();
 sg13g2_fill_8 FILLER_104_480 ();
 sg13g2_fill_8 FILLER_104_488 ();
 sg13g2_fill_8 FILLER_104_496 ();
 sg13g2_fill_8 FILLER_104_504 ();
 sg13g2_fill_8 FILLER_104_512 ();
 sg13g2_fill_8 FILLER_104_520 ();
 sg13g2_fill_8 FILLER_104_528 ();
 sg13g2_fill_8 FILLER_104_536 ();
 sg13g2_fill_8 FILLER_104_544 ();
 sg13g2_fill_8 FILLER_104_552 ();
 sg13g2_fill_8 FILLER_104_560 ();
 sg13g2_fill_8 FILLER_104_568 ();
 sg13g2_fill_8 FILLER_104_576 ();
 sg13g2_fill_8 FILLER_104_584 ();
 sg13g2_fill_8 FILLER_104_592 ();
 sg13g2_fill_8 FILLER_104_600 ();
 sg13g2_fill_8 FILLER_104_608 ();
 sg13g2_fill_8 FILLER_104_616 ();
 sg13g2_fill_8 FILLER_104_624 ();
 sg13g2_fill_8 FILLER_104_632 ();
 sg13g2_fill_8 FILLER_104_640 ();
 sg13g2_fill_8 FILLER_104_648 ();
 sg13g2_fill_8 FILLER_104_656 ();
 sg13g2_fill_8 FILLER_104_664 ();
 sg13g2_fill_8 FILLER_104_672 ();
 sg13g2_fill_8 FILLER_104_680 ();
 sg13g2_fill_8 FILLER_104_688 ();
 sg13g2_fill_8 FILLER_104_696 ();
 sg13g2_fill_8 FILLER_104_704 ();
 sg13g2_fill_8 FILLER_104_712 ();
 sg13g2_fill_8 FILLER_104_720 ();
 sg13g2_fill_8 FILLER_104_728 ();
 sg13g2_fill_8 FILLER_104_736 ();
 sg13g2_fill_8 FILLER_104_744 ();
 sg13g2_fill_8 FILLER_104_752 ();
 sg13g2_fill_8 FILLER_104_760 ();
 sg13g2_fill_8 FILLER_104_768 ();
 sg13g2_fill_8 FILLER_104_776 ();
 sg13g2_fill_8 FILLER_104_784 ();
 sg13g2_fill_8 FILLER_104_792 ();
 sg13g2_fill_8 FILLER_104_800 ();
 sg13g2_fill_8 FILLER_104_808 ();
 sg13g2_fill_8 FILLER_104_816 ();
 sg13g2_fill_8 FILLER_104_824 ();
 sg13g2_fill_8 FILLER_104_832 ();
 sg13g2_fill_8 FILLER_104_840 ();
 sg13g2_fill_8 FILLER_104_848 ();
 sg13g2_fill_8 FILLER_104_856 ();
 sg13g2_fill_8 FILLER_104_864 ();
 sg13g2_fill_8 FILLER_104_872 ();
 sg13g2_fill_8 FILLER_104_880 ();
 sg13g2_fill_8 FILLER_104_888 ();
 sg13g2_fill_8 FILLER_104_896 ();
 sg13g2_fill_8 FILLER_104_904 ();
 sg13g2_fill_8 FILLER_104_912 ();
 sg13g2_fill_8 FILLER_104_920 ();
 sg13g2_fill_8 FILLER_104_928 ();
 sg13g2_fill_8 FILLER_104_936 ();
 sg13g2_fill_8 FILLER_104_944 ();
 sg13g2_fill_8 FILLER_104_952 ();
 sg13g2_fill_8 FILLER_104_960 ();
 sg13g2_fill_8 FILLER_104_968 ();
 sg13g2_fill_8 FILLER_104_976 ();
 sg13g2_fill_8 FILLER_104_984 ();
 sg13g2_fill_8 FILLER_104_992 ();
 sg13g2_fill_8 FILLER_104_1000 ();
 sg13g2_fill_8 FILLER_104_1008 ();
 sg13g2_fill_8 FILLER_104_1016 ();
 sg13g2_fill_8 FILLER_104_1024 ();
 sg13g2_fill_8 FILLER_104_1032 ();
 sg13g2_fill_8 FILLER_104_1040 ();
 sg13g2_fill_8 FILLER_104_1048 ();
 sg13g2_fill_8 FILLER_104_1056 ();
 sg13g2_fill_8 FILLER_104_1064 ();
 sg13g2_fill_8 FILLER_104_1072 ();
 sg13g2_fill_8 FILLER_104_1080 ();
 sg13g2_fill_8 FILLER_104_1088 ();
 sg13g2_fill_8 FILLER_104_1096 ();
 sg13g2_fill_8 FILLER_104_1104 ();
 sg13g2_fill_8 FILLER_104_1112 ();
 sg13g2_fill_8 FILLER_104_1120 ();
 sg13g2_fill_8 FILLER_104_1128 ();
 sg13g2_fill_8 FILLER_104_1136 ();
 sg13g2_fill_8 FILLER_104_1144 ();
 sg13g2_fill_8 FILLER_104_1152 ();
 sg13g2_fill_4 FILLER_104_1160 ();
 sg13g2_fill_2 FILLER_104_1164 ();
 sg13g2_fill_8 FILLER_105_0 ();
 sg13g2_fill_8 FILLER_105_8 ();
 sg13g2_fill_8 FILLER_105_16 ();
 sg13g2_fill_8 FILLER_105_24 ();
 sg13g2_fill_8 FILLER_105_32 ();
 sg13g2_fill_8 FILLER_105_40 ();
 sg13g2_fill_8 FILLER_105_48 ();
 sg13g2_fill_8 FILLER_105_56 ();
 sg13g2_fill_8 FILLER_105_64 ();
 sg13g2_fill_8 FILLER_105_72 ();
 sg13g2_fill_8 FILLER_105_80 ();
 sg13g2_fill_8 FILLER_105_88 ();
 sg13g2_fill_8 FILLER_105_96 ();
 sg13g2_fill_8 FILLER_105_104 ();
 sg13g2_fill_8 FILLER_105_112 ();
 sg13g2_fill_8 FILLER_105_120 ();
 sg13g2_fill_8 FILLER_105_128 ();
 sg13g2_fill_8 FILLER_105_136 ();
 sg13g2_fill_8 FILLER_105_144 ();
 sg13g2_fill_8 FILLER_105_152 ();
 sg13g2_fill_8 FILLER_105_160 ();
 sg13g2_fill_8 FILLER_105_168 ();
 sg13g2_fill_8 FILLER_105_176 ();
 sg13g2_fill_8 FILLER_105_184 ();
 sg13g2_fill_8 FILLER_105_192 ();
 sg13g2_fill_8 FILLER_105_200 ();
 sg13g2_fill_8 FILLER_105_208 ();
 sg13g2_fill_8 FILLER_105_216 ();
 sg13g2_fill_8 FILLER_105_224 ();
 sg13g2_fill_8 FILLER_105_232 ();
 sg13g2_fill_8 FILLER_105_240 ();
 sg13g2_fill_8 FILLER_105_248 ();
 sg13g2_fill_8 FILLER_105_256 ();
 sg13g2_fill_8 FILLER_105_264 ();
 sg13g2_fill_8 FILLER_105_272 ();
 sg13g2_fill_8 FILLER_105_280 ();
 sg13g2_fill_8 FILLER_105_288 ();
 sg13g2_fill_8 FILLER_105_296 ();
 sg13g2_fill_8 FILLER_105_304 ();
 sg13g2_fill_8 FILLER_105_312 ();
 sg13g2_fill_8 FILLER_105_320 ();
 sg13g2_fill_8 FILLER_105_328 ();
 sg13g2_fill_8 FILLER_105_336 ();
 sg13g2_fill_8 FILLER_105_344 ();
 sg13g2_fill_8 FILLER_105_352 ();
 sg13g2_fill_8 FILLER_105_360 ();
 sg13g2_fill_8 FILLER_105_368 ();
 sg13g2_fill_8 FILLER_105_376 ();
 sg13g2_fill_8 FILLER_105_384 ();
 sg13g2_fill_8 FILLER_105_392 ();
 sg13g2_fill_8 FILLER_105_400 ();
 sg13g2_fill_8 FILLER_105_408 ();
 sg13g2_fill_8 FILLER_105_416 ();
 sg13g2_fill_8 FILLER_105_424 ();
 sg13g2_fill_8 FILLER_105_432 ();
 sg13g2_fill_8 FILLER_105_440 ();
 sg13g2_fill_8 FILLER_105_448 ();
 sg13g2_fill_8 FILLER_105_456 ();
 sg13g2_fill_8 FILLER_105_464 ();
 sg13g2_fill_8 FILLER_105_472 ();
 sg13g2_fill_8 FILLER_105_480 ();
 sg13g2_fill_8 FILLER_105_488 ();
 sg13g2_fill_8 FILLER_105_496 ();
 sg13g2_fill_8 FILLER_105_504 ();
 sg13g2_fill_8 FILLER_105_512 ();
 sg13g2_fill_8 FILLER_105_520 ();
 sg13g2_fill_8 FILLER_105_528 ();
 sg13g2_fill_8 FILLER_105_536 ();
 sg13g2_fill_8 FILLER_105_544 ();
 sg13g2_fill_8 FILLER_105_552 ();
 sg13g2_fill_8 FILLER_105_560 ();
 sg13g2_fill_8 FILLER_105_568 ();
 sg13g2_fill_8 FILLER_105_576 ();
 sg13g2_fill_8 FILLER_105_584 ();
 sg13g2_fill_8 FILLER_105_592 ();
 sg13g2_fill_8 FILLER_105_600 ();
 sg13g2_fill_8 FILLER_105_608 ();
 sg13g2_fill_8 FILLER_105_616 ();
 sg13g2_fill_8 FILLER_105_624 ();
 sg13g2_fill_8 FILLER_105_632 ();
 sg13g2_fill_8 FILLER_105_640 ();
 sg13g2_fill_8 FILLER_105_648 ();
 sg13g2_fill_8 FILLER_105_656 ();
 sg13g2_fill_8 FILLER_105_664 ();
 sg13g2_fill_8 FILLER_105_672 ();
 sg13g2_fill_8 FILLER_105_680 ();
 sg13g2_fill_8 FILLER_105_688 ();
 sg13g2_fill_8 FILLER_105_696 ();
 sg13g2_fill_8 FILLER_105_704 ();
 sg13g2_fill_8 FILLER_105_712 ();
 sg13g2_fill_8 FILLER_105_720 ();
 sg13g2_fill_8 FILLER_105_728 ();
 sg13g2_fill_8 FILLER_105_736 ();
 sg13g2_fill_8 FILLER_105_744 ();
 sg13g2_fill_8 FILLER_105_752 ();
 sg13g2_fill_8 FILLER_105_760 ();
 sg13g2_fill_8 FILLER_105_768 ();
 sg13g2_fill_8 FILLER_105_776 ();
 sg13g2_fill_8 FILLER_105_784 ();
 sg13g2_fill_8 FILLER_105_792 ();
 sg13g2_fill_8 FILLER_105_800 ();
 sg13g2_fill_8 FILLER_105_808 ();
 sg13g2_fill_8 FILLER_105_816 ();
 sg13g2_fill_8 FILLER_105_824 ();
 sg13g2_fill_8 FILLER_105_832 ();
 sg13g2_fill_8 FILLER_105_840 ();
 sg13g2_fill_8 FILLER_105_848 ();
 sg13g2_fill_8 FILLER_105_856 ();
 sg13g2_fill_8 FILLER_105_864 ();
 sg13g2_fill_8 FILLER_105_872 ();
 sg13g2_fill_8 FILLER_105_880 ();
 sg13g2_fill_8 FILLER_105_888 ();
 sg13g2_fill_8 FILLER_105_896 ();
 sg13g2_fill_8 FILLER_105_904 ();
 sg13g2_fill_8 FILLER_105_912 ();
 sg13g2_fill_8 FILLER_105_920 ();
 sg13g2_fill_8 FILLER_105_928 ();
 sg13g2_fill_8 FILLER_105_936 ();
 sg13g2_fill_8 FILLER_105_944 ();
 sg13g2_fill_8 FILLER_105_952 ();
 sg13g2_fill_8 FILLER_105_960 ();
 sg13g2_fill_8 FILLER_105_968 ();
 sg13g2_fill_8 FILLER_105_976 ();
 sg13g2_fill_8 FILLER_105_984 ();
 sg13g2_fill_8 FILLER_105_992 ();
 sg13g2_fill_8 FILLER_105_1000 ();
 sg13g2_fill_8 FILLER_105_1008 ();
 sg13g2_fill_8 FILLER_105_1016 ();
 sg13g2_fill_8 FILLER_105_1024 ();
 sg13g2_fill_8 FILLER_105_1032 ();
 sg13g2_fill_8 FILLER_105_1040 ();
 sg13g2_fill_8 FILLER_105_1048 ();
 sg13g2_fill_8 FILLER_105_1056 ();
 sg13g2_fill_8 FILLER_105_1064 ();
 sg13g2_fill_8 FILLER_105_1072 ();
 sg13g2_fill_8 FILLER_105_1080 ();
 sg13g2_fill_8 FILLER_105_1088 ();
 sg13g2_fill_8 FILLER_105_1096 ();
 sg13g2_fill_8 FILLER_105_1104 ();
 sg13g2_fill_8 FILLER_105_1112 ();
 sg13g2_fill_8 FILLER_105_1120 ();
 sg13g2_fill_8 FILLER_105_1128 ();
 sg13g2_fill_8 FILLER_105_1136 ();
 sg13g2_fill_8 FILLER_105_1144 ();
 sg13g2_fill_8 FILLER_105_1152 ();
 sg13g2_fill_4 FILLER_105_1160 ();
 sg13g2_fill_2 FILLER_105_1164 ();
 sg13g2_fill_8 FILLER_106_0 ();
 sg13g2_fill_8 FILLER_106_8 ();
 sg13g2_fill_8 FILLER_106_16 ();
 sg13g2_fill_8 FILLER_106_24 ();
 sg13g2_fill_8 FILLER_106_32 ();
 sg13g2_fill_8 FILLER_106_40 ();
 sg13g2_fill_8 FILLER_106_48 ();
 sg13g2_fill_8 FILLER_106_56 ();
 sg13g2_fill_8 FILLER_106_64 ();
 sg13g2_fill_8 FILLER_106_72 ();
 sg13g2_fill_8 FILLER_106_80 ();
 sg13g2_fill_8 FILLER_106_88 ();
 sg13g2_fill_8 FILLER_106_96 ();
 sg13g2_fill_8 FILLER_106_104 ();
 sg13g2_fill_8 FILLER_106_112 ();
 sg13g2_fill_8 FILLER_106_120 ();
 sg13g2_fill_8 FILLER_106_128 ();
 sg13g2_fill_8 FILLER_106_136 ();
 sg13g2_fill_8 FILLER_106_144 ();
 sg13g2_fill_8 FILLER_106_152 ();
 sg13g2_fill_8 FILLER_106_160 ();
 sg13g2_fill_8 FILLER_106_168 ();
 sg13g2_fill_8 FILLER_106_176 ();
 sg13g2_fill_8 FILLER_106_184 ();
 sg13g2_fill_8 FILLER_106_192 ();
 sg13g2_fill_8 FILLER_106_200 ();
 sg13g2_fill_8 FILLER_106_208 ();
 sg13g2_fill_8 FILLER_106_216 ();
 sg13g2_fill_8 FILLER_106_224 ();
 sg13g2_fill_8 FILLER_106_232 ();
 sg13g2_fill_8 FILLER_106_240 ();
 sg13g2_fill_8 FILLER_106_248 ();
 sg13g2_fill_8 FILLER_106_256 ();
 sg13g2_fill_8 FILLER_106_264 ();
 sg13g2_fill_8 FILLER_106_272 ();
 sg13g2_fill_8 FILLER_106_280 ();
 sg13g2_fill_8 FILLER_106_288 ();
 sg13g2_fill_8 FILLER_106_296 ();
 sg13g2_fill_8 FILLER_106_304 ();
 sg13g2_fill_8 FILLER_106_312 ();
 sg13g2_fill_8 FILLER_106_320 ();
 sg13g2_fill_8 FILLER_106_328 ();
 sg13g2_fill_8 FILLER_106_336 ();
 sg13g2_fill_8 FILLER_106_344 ();
 sg13g2_fill_8 FILLER_106_352 ();
 sg13g2_fill_8 FILLER_106_360 ();
 sg13g2_fill_8 FILLER_106_368 ();
 sg13g2_fill_8 FILLER_106_376 ();
 sg13g2_fill_8 FILLER_106_384 ();
 sg13g2_fill_8 FILLER_106_392 ();
 sg13g2_fill_8 FILLER_106_400 ();
 sg13g2_fill_8 FILLER_106_408 ();
 sg13g2_fill_8 FILLER_106_416 ();
 sg13g2_fill_8 FILLER_106_424 ();
 sg13g2_fill_8 FILLER_106_432 ();
 sg13g2_fill_8 FILLER_106_440 ();
 sg13g2_fill_8 FILLER_106_448 ();
 sg13g2_fill_8 FILLER_106_456 ();
 sg13g2_fill_8 FILLER_106_464 ();
 sg13g2_fill_8 FILLER_106_472 ();
 sg13g2_fill_8 FILLER_106_480 ();
 sg13g2_fill_8 FILLER_106_488 ();
 sg13g2_fill_8 FILLER_106_496 ();
 sg13g2_fill_8 FILLER_106_504 ();
 sg13g2_fill_8 FILLER_106_512 ();
 sg13g2_fill_8 FILLER_106_520 ();
 sg13g2_fill_8 FILLER_106_528 ();
 sg13g2_fill_8 FILLER_106_536 ();
 sg13g2_fill_8 FILLER_106_544 ();
 sg13g2_fill_8 FILLER_106_552 ();
 sg13g2_fill_8 FILLER_106_560 ();
 sg13g2_fill_8 FILLER_106_568 ();
 sg13g2_fill_8 FILLER_106_576 ();
 sg13g2_fill_8 FILLER_106_584 ();
 sg13g2_fill_8 FILLER_106_592 ();
 sg13g2_fill_8 FILLER_106_600 ();
 sg13g2_fill_8 FILLER_106_608 ();
 sg13g2_fill_8 FILLER_106_616 ();
 sg13g2_fill_8 FILLER_106_624 ();
 sg13g2_fill_8 FILLER_106_632 ();
 sg13g2_fill_8 FILLER_106_640 ();
 sg13g2_fill_8 FILLER_106_648 ();
 sg13g2_fill_8 FILLER_106_656 ();
 sg13g2_fill_8 FILLER_106_664 ();
 sg13g2_fill_8 FILLER_106_672 ();
 sg13g2_fill_8 FILLER_106_680 ();
 sg13g2_fill_8 FILLER_106_688 ();
 sg13g2_fill_8 FILLER_106_696 ();
 sg13g2_fill_8 FILLER_106_704 ();
 sg13g2_fill_8 FILLER_106_712 ();
 sg13g2_fill_8 FILLER_106_720 ();
 sg13g2_fill_8 FILLER_106_728 ();
 sg13g2_fill_8 FILLER_106_736 ();
 sg13g2_fill_8 FILLER_106_744 ();
 sg13g2_fill_8 FILLER_106_752 ();
 sg13g2_fill_8 FILLER_106_760 ();
 sg13g2_fill_8 FILLER_106_768 ();
 sg13g2_fill_8 FILLER_106_776 ();
 sg13g2_fill_8 FILLER_106_784 ();
 sg13g2_fill_8 FILLER_106_792 ();
 sg13g2_fill_8 FILLER_106_800 ();
 sg13g2_fill_8 FILLER_106_808 ();
 sg13g2_fill_8 FILLER_106_816 ();
 sg13g2_fill_8 FILLER_106_824 ();
 sg13g2_fill_8 FILLER_106_832 ();
 sg13g2_fill_8 FILLER_106_840 ();
 sg13g2_fill_8 FILLER_106_848 ();
 sg13g2_fill_8 FILLER_106_856 ();
 sg13g2_fill_8 FILLER_106_864 ();
 sg13g2_fill_8 FILLER_106_872 ();
 sg13g2_fill_8 FILLER_106_880 ();
 sg13g2_fill_8 FILLER_106_888 ();
 sg13g2_fill_8 FILLER_106_896 ();
 sg13g2_fill_8 FILLER_106_904 ();
 sg13g2_fill_8 FILLER_106_912 ();
 sg13g2_fill_8 FILLER_106_920 ();
 sg13g2_fill_8 FILLER_106_928 ();
 sg13g2_fill_8 FILLER_106_936 ();
 sg13g2_fill_8 FILLER_106_944 ();
 sg13g2_fill_8 FILLER_106_952 ();
 sg13g2_fill_8 FILLER_106_960 ();
 sg13g2_fill_8 FILLER_106_968 ();
 sg13g2_fill_8 FILLER_106_976 ();
 sg13g2_fill_8 FILLER_106_984 ();
 sg13g2_fill_8 FILLER_106_992 ();
 sg13g2_fill_8 FILLER_106_1000 ();
 sg13g2_fill_8 FILLER_106_1008 ();
 sg13g2_fill_8 FILLER_106_1016 ();
 sg13g2_fill_8 FILLER_106_1024 ();
 sg13g2_fill_8 FILLER_106_1032 ();
 sg13g2_fill_8 FILLER_106_1040 ();
 sg13g2_fill_8 FILLER_106_1048 ();
 sg13g2_fill_8 FILLER_106_1056 ();
 sg13g2_fill_8 FILLER_106_1064 ();
 sg13g2_fill_8 FILLER_106_1072 ();
 sg13g2_fill_8 FILLER_106_1080 ();
 sg13g2_fill_8 FILLER_106_1088 ();
 sg13g2_fill_8 FILLER_106_1096 ();
 sg13g2_fill_8 FILLER_106_1104 ();
 sg13g2_fill_8 FILLER_106_1112 ();
 sg13g2_fill_8 FILLER_106_1120 ();
 sg13g2_fill_8 FILLER_106_1128 ();
 sg13g2_fill_8 FILLER_106_1136 ();
 sg13g2_fill_8 FILLER_106_1144 ();
 sg13g2_fill_8 FILLER_106_1152 ();
 sg13g2_fill_4 FILLER_106_1160 ();
 sg13g2_fill_2 FILLER_106_1164 ();
 sg13g2_fill_8 FILLER_107_0 ();
 sg13g2_fill_8 FILLER_107_8 ();
 sg13g2_fill_8 FILLER_107_16 ();
 sg13g2_fill_8 FILLER_107_24 ();
 sg13g2_fill_8 FILLER_107_32 ();
 sg13g2_fill_8 FILLER_107_40 ();
 sg13g2_fill_8 FILLER_107_48 ();
 sg13g2_fill_8 FILLER_107_56 ();
 sg13g2_fill_8 FILLER_107_64 ();
 sg13g2_fill_8 FILLER_107_72 ();
 sg13g2_fill_8 FILLER_107_80 ();
 sg13g2_fill_8 FILLER_107_88 ();
 sg13g2_fill_8 FILLER_107_96 ();
 sg13g2_fill_8 FILLER_107_104 ();
 sg13g2_fill_8 FILLER_107_112 ();
 sg13g2_fill_8 FILLER_107_120 ();
 sg13g2_fill_8 FILLER_107_128 ();
 sg13g2_fill_8 FILLER_107_136 ();
 sg13g2_fill_8 FILLER_107_144 ();
 sg13g2_fill_8 FILLER_107_152 ();
 sg13g2_fill_8 FILLER_107_160 ();
 sg13g2_fill_8 FILLER_107_168 ();
 sg13g2_fill_8 FILLER_107_176 ();
 sg13g2_fill_8 FILLER_107_184 ();
 sg13g2_fill_8 FILLER_107_192 ();
 sg13g2_fill_8 FILLER_107_200 ();
 sg13g2_fill_8 FILLER_107_208 ();
 sg13g2_fill_8 FILLER_107_216 ();
 sg13g2_fill_8 FILLER_107_224 ();
 sg13g2_fill_8 FILLER_107_232 ();
 sg13g2_fill_8 FILLER_107_240 ();
 sg13g2_fill_8 FILLER_107_248 ();
 sg13g2_fill_8 FILLER_107_256 ();
 sg13g2_fill_8 FILLER_107_264 ();
 sg13g2_fill_8 FILLER_107_272 ();
 sg13g2_fill_8 FILLER_107_280 ();
 sg13g2_fill_8 FILLER_107_288 ();
 sg13g2_fill_8 FILLER_107_296 ();
 sg13g2_fill_8 FILLER_107_304 ();
 sg13g2_fill_8 FILLER_107_312 ();
 sg13g2_fill_8 FILLER_107_320 ();
 sg13g2_fill_8 FILLER_107_328 ();
 sg13g2_fill_8 FILLER_107_336 ();
 sg13g2_fill_8 FILLER_107_344 ();
 sg13g2_fill_8 FILLER_107_352 ();
 sg13g2_fill_8 FILLER_107_360 ();
 sg13g2_fill_8 FILLER_107_368 ();
 sg13g2_fill_8 FILLER_107_376 ();
 sg13g2_fill_8 FILLER_107_384 ();
 sg13g2_fill_8 FILLER_107_392 ();
 sg13g2_fill_8 FILLER_107_400 ();
 sg13g2_fill_8 FILLER_107_408 ();
 sg13g2_fill_8 FILLER_107_416 ();
 sg13g2_fill_8 FILLER_107_424 ();
 sg13g2_fill_8 FILLER_107_432 ();
 sg13g2_fill_8 FILLER_107_440 ();
 sg13g2_fill_8 FILLER_107_448 ();
 sg13g2_fill_8 FILLER_107_456 ();
 sg13g2_fill_8 FILLER_107_464 ();
 sg13g2_fill_8 FILLER_107_472 ();
 sg13g2_fill_8 FILLER_107_480 ();
 sg13g2_fill_8 FILLER_107_488 ();
 sg13g2_fill_8 FILLER_107_496 ();
 sg13g2_fill_8 FILLER_107_504 ();
 sg13g2_fill_8 FILLER_107_512 ();
 sg13g2_fill_8 FILLER_107_520 ();
 sg13g2_fill_8 FILLER_107_528 ();
 sg13g2_fill_8 FILLER_107_536 ();
 sg13g2_fill_8 FILLER_107_544 ();
 sg13g2_fill_8 FILLER_107_552 ();
 sg13g2_fill_8 FILLER_107_560 ();
 sg13g2_fill_8 FILLER_107_568 ();
 sg13g2_fill_8 FILLER_107_576 ();
 sg13g2_fill_8 FILLER_107_584 ();
 sg13g2_fill_8 FILLER_107_592 ();
 sg13g2_fill_8 FILLER_107_600 ();
 sg13g2_fill_8 FILLER_107_608 ();
 sg13g2_fill_8 FILLER_107_616 ();
 sg13g2_fill_8 FILLER_107_624 ();
 sg13g2_fill_8 FILLER_107_632 ();
 sg13g2_fill_8 FILLER_107_640 ();
 sg13g2_fill_8 FILLER_107_648 ();
 sg13g2_fill_8 FILLER_107_656 ();
 sg13g2_fill_8 FILLER_107_664 ();
 sg13g2_fill_8 FILLER_107_672 ();
 sg13g2_fill_8 FILLER_107_680 ();
 sg13g2_fill_8 FILLER_107_688 ();
 sg13g2_fill_8 FILLER_107_696 ();
 sg13g2_fill_8 FILLER_107_704 ();
 sg13g2_fill_8 FILLER_107_712 ();
 sg13g2_fill_8 FILLER_107_720 ();
 sg13g2_fill_8 FILLER_107_728 ();
 sg13g2_fill_8 FILLER_107_736 ();
 sg13g2_fill_8 FILLER_107_744 ();
 sg13g2_fill_8 FILLER_107_752 ();
 sg13g2_fill_8 FILLER_107_760 ();
 sg13g2_fill_8 FILLER_107_768 ();
 sg13g2_fill_8 FILLER_107_776 ();
 sg13g2_fill_8 FILLER_107_784 ();
 sg13g2_fill_8 FILLER_107_792 ();
 sg13g2_fill_8 FILLER_107_800 ();
 sg13g2_fill_8 FILLER_107_808 ();
 sg13g2_fill_8 FILLER_107_816 ();
 sg13g2_fill_8 FILLER_107_824 ();
 sg13g2_fill_8 FILLER_107_832 ();
 sg13g2_fill_8 FILLER_107_840 ();
 sg13g2_fill_8 FILLER_107_848 ();
 sg13g2_fill_8 FILLER_107_856 ();
 sg13g2_fill_8 FILLER_107_864 ();
 sg13g2_fill_8 FILLER_107_872 ();
 sg13g2_fill_8 FILLER_107_880 ();
 sg13g2_fill_8 FILLER_107_888 ();
 sg13g2_fill_8 FILLER_107_896 ();
 sg13g2_fill_8 FILLER_107_904 ();
 sg13g2_fill_8 FILLER_107_912 ();
 sg13g2_fill_8 FILLER_107_920 ();
 sg13g2_fill_8 FILLER_107_928 ();
 sg13g2_fill_8 FILLER_107_936 ();
 sg13g2_fill_8 FILLER_107_944 ();
 sg13g2_fill_8 FILLER_107_952 ();
 sg13g2_fill_8 FILLER_107_960 ();
 sg13g2_fill_8 FILLER_107_968 ();
 sg13g2_fill_8 FILLER_107_976 ();
 sg13g2_fill_8 FILLER_107_984 ();
 sg13g2_fill_8 FILLER_107_992 ();
 sg13g2_fill_8 FILLER_107_1000 ();
 sg13g2_fill_8 FILLER_107_1008 ();
 sg13g2_fill_8 FILLER_107_1016 ();
 sg13g2_fill_8 FILLER_107_1024 ();
 sg13g2_fill_8 FILLER_107_1032 ();
 sg13g2_fill_8 FILLER_107_1040 ();
 sg13g2_fill_8 FILLER_107_1048 ();
 sg13g2_fill_8 FILLER_107_1056 ();
 sg13g2_fill_8 FILLER_107_1064 ();
 sg13g2_fill_8 FILLER_107_1072 ();
 sg13g2_fill_8 FILLER_107_1080 ();
 sg13g2_fill_8 FILLER_107_1088 ();
 sg13g2_fill_8 FILLER_107_1096 ();
 sg13g2_fill_8 FILLER_107_1104 ();
 sg13g2_fill_8 FILLER_107_1112 ();
 sg13g2_fill_8 FILLER_107_1120 ();
 sg13g2_fill_8 FILLER_107_1128 ();
 sg13g2_fill_8 FILLER_107_1136 ();
 sg13g2_fill_8 FILLER_107_1144 ();
 sg13g2_fill_8 FILLER_107_1152 ();
 sg13g2_fill_4 FILLER_107_1160 ();
 sg13g2_fill_2 FILLER_107_1164 ();
 sg13g2_fill_8 FILLER_108_0 ();
 sg13g2_fill_8 FILLER_108_8 ();
 sg13g2_fill_8 FILLER_108_16 ();
 sg13g2_fill_8 FILLER_108_24 ();
 sg13g2_fill_8 FILLER_108_32 ();
 sg13g2_fill_8 FILLER_108_40 ();
 sg13g2_fill_8 FILLER_108_48 ();
 sg13g2_fill_8 FILLER_108_56 ();
 sg13g2_fill_8 FILLER_108_64 ();
 sg13g2_fill_8 FILLER_108_72 ();
 sg13g2_fill_8 FILLER_108_80 ();
 sg13g2_fill_8 FILLER_108_88 ();
 sg13g2_fill_8 FILLER_108_96 ();
 sg13g2_fill_8 FILLER_108_104 ();
 sg13g2_fill_8 FILLER_108_112 ();
 sg13g2_fill_8 FILLER_108_120 ();
 sg13g2_fill_8 FILLER_108_128 ();
 sg13g2_fill_8 FILLER_108_136 ();
 sg13g2_fill_8 FILLER_108_144 ();
 sg13g2_fill_8 FILLER_108_152 ();
 sg13g2_fill_8 FILLER_108_160 ();
 sg13g2_fill_8 FILLER_108_168 ();
 sg13g2_fill_8 FILLER_108_176 ();
 sg13g2_fill_8 FILLER_108_184 ();
 sg13g2_fill_8 FILLER_108_192 ();
 sg13g2_fill_8 FILLER_108_200 ();
 sg13g2_fill_8 FILLER_108_208 ();
 sg13g2_fill_8 FILLER_108_216 ();
 sg13g2_fill_8 FILLER_108_224 ();
 sg13g2_fill_8 FILLER_108_232 ();
 sg13g2_fill_8 FILLER_108_240 ();
 sg13g2_fill_8 FILLER_108_248 ();
 sg13g2_fill_8 FILLER_108_256 ();
 sg13g2_fill_8 FILLER_108_264 ();
 sg13g2_fill_8 FILLER_108_272 ();
 sg13g2_fill_8 FILLER_108_280 ();
 sg13g2_fill_8 FILLER_108_288 ();
 sg13g2_fill_8 FILLER_108_296 ();
 sg13g2_fill_8 FILLER_108_304 ();
 sg13g2_fill_8 FILLER_108_312 ();
 sg13g2_fill_8 FILLER_108_320 ();
 sg13g2_fill_8 FILLER_108_328 ();
 sg13g2_fill_8 FILLER_108_336 ();
 sg13g2_fill_8 FILLER_108_344 ();
 sg13g2_fill_8 FILLER_108_352 ();
 sg13g2_fill_8 FILLER_108_360 ();
 sg13g2_fill_8 FILLER_108_368 ();
 sg13g2_fill_8 FILLER_108_376 ();
 sg13g2_fill_8 FILLER_108_384 ();
 sg13g2_fill_8 FILLER_108_392 ();
 sg13g2_fill_8 FILLER_108_400 ();
 sg13g2_fill_8 FILLER_108_408 ();
 sg13g2_fill_8 FILLER_108_416 ();
 sg13g2_fill_8 FILLER_108_424 ();
 sg13g2_fill_8 FILLER_108_432 ();
 sg13g2_fill_8 FILLER_108_440 ();
 sg13g2_fill_8 FILLER_108_448 ();
 sg13g2_fill_8 FILLER_108_456 ();
 sg13g2_fill_8 FILLER_108_464 ();
 sg13g2_fill_8 FILLER_108_472 ();
 sg13g2_fill_8 FILLER_108_480 ();
 sg13g2_fill_8 FILLER_108_488 ();
 sg13g2_fill_8 FILLER_108_496 ();
 sg13g2_fill_8 FILLER_108_504 ();
 sg13g2_fill_8 FILLER_108_512 ();
 sg13g2_fill_8 FILLER_108_520 ();
 sg13g2_fill_8 FILLER_108_528 ();
 sg13g2_fill_8 FILLER_108_536 ();
 sg13g2_fill_8 FILLER_108_544 ();
 sg13g2_fill_8 FILLER_108_552 ();
 sg13g2_fill_8 FILLER_108_560 ();
 sg13g2_fill_8 FILLER_108_568 ();
 sg13g2_fill_8 FILLER_108_576 ();
 sg13g2_fill_8 FILLER_108_584 ();
 sg13g2_fill_8 FILLER_108_592 ();
 sg13g2_fill_8 FILLER_108_600 ();
 sg13g2_fill_8 FILLER_108_608 ();
 sg13g2_fill_8 FILLER_108_616 ();
 sg13g2_fill_8 FILLER_108_624 ();
 sg13g2_fill_8 FILLER_108_632 ();
 sg13g2_fill_8 FILLER_108_640 ();
 sg13g2_fill_8 FILLER_108_648 ();
 sg13g2_fill_8 FILLER_108_656 ();
 sg13g2_fill_8 FILLER_108_664 ();
 sg13g2_fill_8 FILLER_108_672 ();
 sg13g2_fill_8 FILLER_108_680 ();
 sg13g2_fill_8 FILLER_108_688 ();
 sg13g2_fill_8 FILLER_108_696 ();
 sg13g2_fill_8 FILLER_108_704 ();
 sg13g2_fill_8 FILLER_108_712 ();
 sg13g2_fill_8 FILLER_108_720 ();
 sg13g2_fill_8 FILLER_108_728 ();
 sg13g2_fill_8 FILLER_108_736 ();
 sg13g2_fill_8 FILLER_108_744 ();
 sg13g2_fill_8 FILLER_108_752 ();
 sg13g2_fill_8 FILLER_108_760 ();
 sg13g2_fill_8 FILLER_108_768 ();
 sg13g2_fill_8 FILLER_108_776 ();
 sg13g2_fill_8 FILLER_108_784 ();
 sg13g2_fill_8 FILLER_108_792 ();
 sg13g2_fill_8 FILLER_108_800 ();
 sg13g2_fill_8 FILLER_108_808 ();
 sg13g2_fill_8 FILLER_108_816 ();
 sg13g2_fill_8 FILLER_108_824 ();
 sg13g2_fill_8 FILLER_108_832 ();
 sg13g2_fill_8 FILLER_108_840 ();
 sg13g2_fill_8 FILLER_108_848 ();
 sg13g2_fill_8 FILLER_108_856 ();
 sg13g2_fill_8 FILLER_108_864 ();
 sg13g2_fill_8 FILLER_108_872 ();
 sg13g2_fill_8 FILLER_108_880 ();
 sg13g2_fill_8 FILLER_108_888 ();
 sg13g2_fill_8 FILLER_108_896 ();
 sg13g2_fill_8 FILLER_108_904 ();
 sg13g2_fill_8 FILLER_108_912 ();
 sg13g2_fill_8 FILLER_108_920 ();
 sg13g2_fill_8 FILLER_108_928 ();
 sg13g2_fill_8 FILLER_108_936 ();
 sg13g2_fill_8 FILLER_108_944 ();
 sg13g2_fill_8 FILLER_108_952 ();
 sg13g2_fill_8 FILLER_108_960 ();
 sg13g2_fill_8 FILLER_108_968 ();
 sg13g2_fill_8 FILLER_108_976 ();
 sg13g2_fill_8 FILLER_108_984 ();
 sg13g2_fill_8 FILLER_108_992 ();
 sg13g2_fill_8 FILLER_108_1000 ();
 sg13g2_fill_8 FILLER_108_1008 ();
 sg13g2_fill_8 FILLER_108_1016 ();
 sg13g2_fill_8 FILLER_108_1024 ();
 sg13g2_fill_8 FILLER_108_1032 ();
 sg13g2_fill_8 FILLER_108_1040 ();
 sg13g2_fill_8 FILLER_108_1048 ();
 sg13g2_fill_8 FILLER_108_1056 ();
 sg13g2_fill_8 FILLER_108_1064 ();
 sg13g2_fill_8 FILLER_108_1072 ();
 sg13g2_fill_8 FILLER_108_1080 ();
 sg13g2_fill_8 FILLER_108_1088 ();
 sg13g2_fill_8 FILLER_108_1096 ();
 sg13g2_fill_8 FILLER_108_1104 ();
 sg13g2_fill_8 FILLER_108_1112 ();
 sg13g2_fill_8 FILLER_108_1120 ();
 sg13g2_fill_8 FILLER_108_1128 ();
 sg13g2_fill_8 FILLER_108_1136 ();
 sg13g2_fill_8 FILLER_108_1144 ();
 sg13g2_fill_8 FILLER_108_1152 ();
 sg13g2_fill_4 FILLER_108_1160 ();
 sg13g2_fill_2 FILLER_108_1164 ();
 sg13g2_fill_8 FILLER_109_0 ();
 sg13g2_fill_8 FILLER_109_8 ();
 sg13g2_fill_8 FILLER_109_16 ();
 sg13g2_fill_8 FILLER_109_24 ();
 sg13g2_fill_8 FILLER_109_32 ();
 sg13g2_fill_8 FILLER_109_40 ();
 sg13g2_fill_8 FILLER_109_48 ();
 sg13g2_fill_8 FILLER_109_56 ();
 sg13g2_fill_8 FILLER_109_64 ();
 sg13g2_fill_8 FILLER_109_72 ();
 sg13g2_fill_8 FILLER_109_80 ();
 sg13g2_fill_8 FILLER_109_88 ();
 sg13g2_fill_8 FILLER_109_96 ();
 sg13g2_fill_8 FILLER_109_104 ();
 sg13g2_fill_8 FILLER_109_112 ();
 sg13g2_fill_8 FILLER_109_120 ();
 sg13g2_fill_8 FILLER_109_128 ();
 sg13g2_fill_8 FILLER_109_136 ();
 sg13g2_fill_8 FILLER_109_144 ();
 sg13g2_fill_8 FILLER_109_152 ();
 sg13g2_fill_8 FILLER_109_160 ();
 sg13g2_fill_8 FILLER_109_168 ();
 sg13g2_fill_8 FILLER_109_176 ();
 sg13g2_fill_8 FILLER_109_184 ();
 sg13g2_fill_8 FILLER_109_192 ();
 sg13g2_fill_8 FILLER_109_200 ();
 sg13g2_fill_8 FILLER_109_208 ();
 sg13g2_fill_8 FILLER_109_216 ();
 sg13g2_fill_8 FILLER_109_224 ();
 sg13g2_fill_8 FILLER_109_232 ();
 sg13g2_fill_8 FILLER_109_240 ();
 sg13g2_fill_8 FILLER_109_248 ();
 sg13g2_fill_8 FILLER_109_256 ();
 sg13g2_fill_8 FILLER_109_264 ();
 sg13g2_fill_8 FILLER_109_272 ();
 sg13g2_fill_8 FILLER_109_280 ();
 sg13g2_fill_8 FILLER_109_288 ();
 sg13g2_fill_8 FILLER_109_296 ();
 sg13g2_fill_8 FILLER_109_304 ();
 sg13g2_fill_8 FILLER_109_312 ();
 sg13g2_fill_8 FILLER_109_320 ();
 sg13g2_fill_8 FILLER_109_328 ();
 sg13g2_fill_8 FILLER_109_336 ();
 sg13g2_fill_8 FILLER_109_344 ();
 sg13g2_fill_8 FILLER_109_352 ();
 sg13g2_fill_8 FILLER_109_360 ();
 sg13g2_fill_8 FILLER_109_368 ();
 sg13g2_fill_8 FILLER_109_376 ();
 sg13g2_fill_8 FILLER_109_384 ();
 sg13g2_fill_8 FILLER_109_392 ();
 sg13g2_fill_8 FILLER_109_400 ();
 sg13g2_fill_8 FILLER_109_408 ();
 sg13g2_fill_8 FILLER_109_416 ();
 sg13g2_fill_8 FILLER_109_424 ();
 sg13g2_fill_8 FILLER_109_432 ();
 sg13g2_fill_8 FILLER_109_440 ();
 sg13g2_fill_8 FILLER_109_448 ();
 sg13g2_fill_8 FILLER_109_456 ();
 sg13g2_fill_8 FILLER_109_464 ();
 sg13g2_fill_8 FILLER_109_472 ();
 sg13g2_fill_8 FILLER_109_480 ();
 sg13g2_fill_8 FILLER_109_488 ();
 sg13g2_fill_8 FILLER_109_496 ();
 sg13g2_fill_8 FILLER_109_504 ();
 sg13g2_fill_8 FILLER_109_512 ();
 sg13g2_fill_8 FILLER_109_520 ();
 sg13g2_fill_8 FILLER_109_528 ();
 sg13g2_fill_8 FILLER_109_536 ();
 sg13g2_fill_8 FILLER_109_544 ();
 sg13g2_fill_8 FILLER_109_552 ();
 sg13g2_fill_8 FILLER_109_560 ();
 sg13g2_fill_8 FILLER_109_568 ();
 sg13g2_fill_8 FILLER_109_576 ();
 sg13g2_fill_8 FILLER_109_584 ();
 sg13g2_fill_8 FILLER_109_592 ();
 sg13g2_fill_8 FILLER_109_600 ();
 sg13g2_fill_8 FILLER_109_608 ();
 sg13g2_fill_8 FILLER_109_616 ();
 sg13g2_fill_8 FILLER_109_624 ();
 sg13g2_fill_8 FILLER_109_632 ();
 sg13g2_fill_8 FILLER_109_640 ();
 sg13g2_fill_8 FILLER_109_648 ();
 sg13g2_fill_8 FILLER_109_656 ();
 sg13g2_fill_8 FILLER_109_664 ();
 sg13g2_fill_8 FILLER_109_672 ();
 sg13g2_fill_8 FILLER_109_680 ();
 sg13g2_fill_8 FILLER_109_688 ();
 sg13g2_fill_8 FILLER_109_696 ();
 sg13g2_fill_8 FILLER_109_704 ();
 sg13g2_fill_8 FILLER_109_712 ();
 sg13g2_fill_8 FILLER_109_720 ();
 sg13g2_fill_8 FILLER_109_728 ();
 sg13g2_fill_8 FILLER_109_736 ();
 sg13g2_fill_8 FILLER_109_744 ();
 sg13g2_fill_8 FILLER_109_752 ();
 sg13g2_fill_8 FILLER_109_760 ();
 sg13g2_fill_8 FILLER_109_768 ();
 sg13g2_fill_8 FILLER_109_776 ();
 sg13g2_fill_8 FILLER_109_784 ();
 sg13g2_fill_8 FILLER_109_792 ();
 sg13g2_fill_8 FILLER_109_800 ();
 sg13g2_fill_8 FILLER_109_808 ();
 sg13g2_fill_8 FILLER_109_816 ();
 sg13g2_fill_8 FILLER_109_824 ();
 sg13g2_fill_8 FILLER_109_832 ();
 sg13g2_fill_8 FILLER_109_840 ();
 sg13g2_fill_8 FILLER_109_848 ();
 sg13g2_fill_8 FILLER_109_856 ();
 sg13g2_fill_8 FILLER_109_864 ();
 sg13g2_fill_8 FILLER_109_872 ();
 sg13g2_fill_8 FILLER_109_880 ();
 sg13g2_fill_8 FILLER_109_888 ();
 sg13g2_fill_8 FILLER_109_896 ();
 sg13g2_fill_8 FILLER_109_904 ();
 sg13g2_fill_8 FILLER_109_912 ();
 sg13g2_fill_8 FILLER_109_920 ();
 sg13g2_fill_8 FILLER_109_928 ();
 sg13g2_fill_8 FILLER_109_936 ();
 sg13g2_fill_8 FILLER_109_944 ();
 sg13g2_fill_8 FILLER_109_952 ();
 sg13g2_fill_8 FILLER_109_960 ();
 sg13g2_fill_8 FILLER_109_968 ();
 sg13g2_fill_8 FILLER_109_976 ();
 sg13g2_fill_8 FILLER_109_984 ();
 sg13g2_fill_8 FILLER_109_992 ();
 sg13g2_fill_8 FILLER_109_1000 ();
 sg13g2_fill_8 FILLER_109_1008 ();
 sg13g2_fill_8 FILLER_109_1016 ();
 sg13g2_fill_8 FILLER_109_1024 ();
 sg13g2_fill_8 FILLER_109_1032 ();
 sg13g2_fill_8 FILLER_109_1040 ();
 sg13g2_fill_8 FILLER_109_1048 ();
 sg13g2_fill_8 FILLER_109_1056 ();
 sg13g2_fill_8 FILLER_109_1064 ();
 sg13g2_fill_8 FILLER_109_1072 ();
 sg13g2_fill_8 FILLER_109_1080 ();
 sg13g2_fill_8 FILLER_109_1088 ();
 sg13g2_fill_8 FILLER_109_1096 ();
 sg13g2_fill_8 FILLER_109_1104 ();
 sg13g2_fill_8 FILLER_109_1112 ();
 sg13g2_fill_8 FILLER_109_1120 ();
 sg13g2_fill_8 FILLER_109_1128 ();
 sg13g2_fill_8 FILLER_109_1136 ();
 sg13g2_fill_8 FILLER_109_1144 ();
 sg13g2_fill_8 FILLER_109_1152 ();
 sg13g2_fill_4 FILLER_109_1160 ();
 sg13g2_fill_2 FILLER_109_1164 ();
 sg13g2_fill_8 FILLER_110_0 ();
 sg13g2_fill_8 FILLER_110_8 ();
 sg13g2_fill_8 FILLER_110_16 ();
 sg13g2_fill_8 FILLER_110_24 ();
 sg13g2_fill_8 FILLER_110_32 ();
 sg13g2_fill_8 FILLER_110_40 ();
 sg13g2_fill_8 FILLER_110_48 ();
 sg13g2_fill_8 FILLER_110_56 ();
 sg13g2_fill_8 FILLER_110_64 ();
 sg13g2_fill_8 FILLER_110_72 ();
 sg13g2_fill_8 FILLER_110_80 ();
 sg13g2_fill_8 FILLER_110_88 ();
 sg13g2_fill_8 FILLER_110_96 ();
 sg13g2_fill_8 FILLER_110_104 ();
 sg13g2_fill_8 FILLER_110_112 ();
 sg13g2_fill_8 FILLER_110_120 ();
 sg13g2_fill_8 FILLER_110_128 ();
 sg13g2_fill_8 FILLER_110_136 ();
 sg13g2_fill_8 FILLER_110_144 ();
 sg13g2_fill_8 FILLER_110_152 ();
 sg13g2_fill_8 FILLER_110_160 ();
 sg13g2_fill_8 FILLER_110_168 ();
 sg13g2_fill_8 FILLER_110_176 ();
 sg13g2_fill_8 FILLER_110_184 ();
 sg13g2_fill_8 FILLER_110_192 ();
 sg13g2_fill_8 FILLER_110_200 ();
 sg13g2_fill_8 FILLER_110_208 ();
 sg13g2_fill_8 FILLER_110_216 ();
 sg13g2_fill_8 FILLER_110_224 ();
 sg13g2_fill_8 FILLER_110_232 ();
 sg13g2_fill_8 FILLER_110_240 ();
 sg13g2_fill_8 FILLER_110_248 ();
 sg13g2_fill_8 FILLER_110_256 ();
 sg13g2_fill_8 FILLER_110_264 ();
 sg13g2_fill_8 FILLER_110_272 ();
 sg13g2_fill_8 FILLER_110_280 ();
 sg13g2_fill_8 FILLER_110_288 ();
 sg13g2_fill_8 FILLER_110_296 ();
 sg13g2_fill_8 FILLER_110_304 ();
 sg13g2_fill_8 FILLER_110_312 ();
 sg13g2_fill_8 FILLER_110_320 ();
 sg13g2_fill_8 FILLER_110_328 ();
 sg13g2_fill_8 FILLER_110_336 ();
 sg13g2_fill_8 FILLER_110_344 ();
 sg13g2_fill_8 FILLER_110_352 ();
 sg13g2_fill_8 FILLER_110_360 ();
 sg13g2_fill_8 FILLER_110_368 ();
 sg13g2_fill_8 FILLER_110_376 ();
 sg13g2_fill_8 FILLER_110_384 ();
 sg13g2_fill_8 FILLER_110_392 ();
 sg13g2_fill_8 FILLER_110_400 ();
 sg13g2_fill_8 FILLER_110_408 ();
 sg13g2_fill_8 FILLER_110_416 ();
 sg13g2_fill_8 FILLER_110_424 ();
 sg13g2_fill_8 FILLER_110_432 ();
 sg13g2_fill_8 FILLER_110_440 ();
 sg13g2_fill_8 FILLER_110_448 ();
 sg13g2_fill_8 FILLER_110_456 ();
 sg13g2_fill_8 FILLER_110_464 ();
 sg13g2_fill_8 FILLER_110_472 ();
 sg13g2_fill_8 FILLER_110_480 ();
 sg13g2_fill_8 FILLER_110_488 ();
 sg13g2_fill_8 FILLER_110_496 ();
 sg13g2_fill_8 FILLER_110_504 ();
 sg13g2_fill_8 FILLER_110_512 ();
 sg13g2_fill_8 FILLER_110_520 ();
 sg13g2_fill_8 FILLER_110_528 ();
 sg13g2_fill_8 FILLER_110_536 ();
 sg13g2_fill_8 FILLER_110_544 ();
 sg13g2_fill_8 FILLER_110_552 ();
 sg13g2_fill_8 FILLER_110_560 ();
 sg13g2_fill_8 FILLER_110_568 ();
 sg13g2_fill_8 FILLER_110_576 ();
 sg13g2_fill_8 FILLER_110_584 ();
 sg13g2_fill_8 FILLER_110_592 ();
 sg13g2_fill_8 FILLER_110_600 ();
 sg13g2_fill_8 FILLER_110_608 ();
 sg13g2_fill_8 FILLER_110_616 ();
 sg13g2_fill_8 FILLER_110_624 ();
 sg13g2_fill_8 FILLER_110_632 ();
 sg13g2_fill_8 FILLER_110_640 ();
 sg13g2_fill_8 FILLER_110_648 ();
 sg13g2_fill_8 FILLER_110_656 ();
 sg13g2_fill_8 FILLER_110_664 ();
 sg13g2_fill_8 FILLER_110_672 ();
 sg13g2_fill_8 FILLER_110_680 ();
 sg13g2_fill_8 FILLER_110_688 ();
 sg13g2_fill_8 FILLER_110_696 ();
 sg13g2_fill_8 FILLER_110_704 ();
 sg13g2_fill_8 FILLER_110_712 ();
 sg13g2_fill_8 FILLER_110_720 ();
 sg13g2_fill_8 FILLER_110_728 ();
 sg13g2_fill_8 FILLER_110_736 ();
 sg13g2_fill_8 FILLER_110_744 ();
 sg13g2_fill_8 FILLER_110_752 ();
 sg13g2_fill_8 FILLER_110_760 ();
 sg13g2_fill_8 FILLER_110_768 ();
 sg13g2_fill_8 FILLER_110_776 ();
 sg13g2_fill_8 FILLER_110_784 ();
 sg13g2_fill_8 FILLER_110_792 ();
 sg13g2_fill_8 FILLER_110_800 ();
 sg13g2_fill_8 FILLER_110_808 ();
 sg13g2_fill_8 FILLER_110_816 ();
 sg13g2_fill_8 FILLER_110_824 ();
 sg13g2_fill_8 FILLER_110_832 ();
 sg13g2_fill_8 FILLER_110_840 ();
 sg13g2_fill_8 FILLER_110_848 ();
 sg13g2_fill_8 FILLER_110_856 ();
 sg13g2_fill_8 FILLER_110_864 ();
 sg13g2_fill_8 FILLER_110_872 ();
 sg13g2_fill_8 FILLER_110_880 ();
 sg13g2_fill_8 FILLER_110_888 ();
 sg13g2_fill_8 FILLER_110_896 ();
 sg13g2_fill_8 FILLER_110_904 ();
 sg13g2_fill_8 FILLER_110_912 ();
 sg13g2_fill_8 FILLER_110_920 ();
 sg13g2_fill_8 FILLER_110_928 ();
 sg13g2_fill_8 FILLER_110_936 ();
 sg13g2_fill_8 FILLER_110_944 ();
 sg13g2_fill_8 FILLER_110_952 ();
 sg13g2_fill_8 FILLER_110_960 ();
 sg13g2_fill_8 FILLER_110_968 ();
 sg13g2_fill_8 FILLER_110_976 ();
 sg13g2_fill_8 FILLER_110_984 ();
 sg13g2_fill_8 FILLER_110_992 ();
 sg13g2_fill_8 FILLER_110_1000 ();
 sg13g2_fill_8 FILLER_110_1008 ();
 sg13g2_fill_8 FILLER_110_1016 ();
 sg13g2_fill_8 FILLER_110_1024 ();
 sg13g2_fill_8 FILLER_110_1032 ();
 sg13g2_fill_8 FILLER_110_1040 ();
 sg13g2_fill_8 FILLER_110_1048 ();
 sg13g2_fill_8 FILLER_110_1056 ();
 sg13g2_fill_8 FILLER_110_1064 ();
 sg13g2_fill_8 FILLER_110_1072 ();
 sg13g2_fill_8 FILLER_110_1080 ();
 sg13g2_fill_8 FILLER_110_1088 ();
 sg13g2_fill_8 FILLER_110_1096 ();
 sg13g2_fill_8 FILLER_110_1104 ();
 sg13g2_fill_8 FILLER_110_1112 ();
 sg13g2_fill_8 FILLER_110_1120 ();
 sg13g2_fill_8 FILLER_110_1128 ();
 sg13g2_fill_8 FILLER_110_1136 ();
 sg13g2_fill_8 FILLER_110_1144 ();
 sg13g2_fill_8 FILLER_110_1152 ();
 sg13g2_fill_4 FILLER_110_1160 ();
 sg13g2_fill_2 FILLER_110_1164 ();
 sg13g2_fill_8 FILLER_111_0 ();
 sg13g2_fill_8 FILLER_111_8 ();
 sg13g2_fill_8 FILLER_111_16 ();
 sg13g2_fill_8 FILLER_111_24 ();
 sg13g2_fill_8 FILLER_111_32 ();
 sg13g2_fill_8 FILLER_111_40 ();
 sg13g2_fill_8 FILLER_111_48 ();
 sg13g2_fill_8 FILLER_111_56 ();
 sg13g2_fill_8 FILLER_111_64 ();
 sg13g2_fill_8 FILLER_111_72 ();
 sg13g2_fill_8 FILLER_111_80 ();
 sg13g2_fill_8 FILLER_111_88 ();
 sg13g2_fill_8 FILLER_111_96 ();
 sg13g2_fill_8 FILLER_111_104 ();
 sg13g2_fill_8 FILLER_111_112 ();
 sg13g2_fill_8 FILLER_111_120 ();
 sg13g2_fill_8 FILLER_111_128 ();
 sg13g2_fill_8 FILLER_111_136 ();
 sg13g2_fill_8 FILLER_111_144 ();
 sg13g2_fill_8 FILLER_111_152 ();
 sg13g2_fill_8 FILLER_111_160 ();
 sg13g2_fill_8 FILLER_111_168 ();
 sg13g2_fill_8 FILLER_111_176 ();
 sg13g2_fill_8 FILLER_111_184 ();
 sg13g2_fill_8 FILLER_111_192 ();
 sg13g2_fill_8 FILLER_111_200 ();
 sg13g2_fill_8 FILLER_111_208 ();
 sg13g2_fill_8 FILLER_111_216 ();
 sg13g2_fill_8 FILLER_111_224 ();
 sg13g2_fill_8 FILLER_111_232 ();
 sg13g2_fill_8 FILLER_111_240 ();
 sg13g2_fill_8 FILLER_111_248 ();
 sg13g2_fill_8 FILLER_111_256 ();
 sg13g2_fill_8 FILLER_111_264 ();
 sg13g2_fill_8 FILLER_111_272 ();
 sg13g2_fill_8 FILLER_111_280 ();
 sg13g2_fill_8 FILLER_111_288 ();
 sg13g2_fill_8 FILLER_111_296 ();
 sg13g2_fill_8 FILLER_111_304 ();
 sg13g2_fill_8 FILLER_111_312 ();
 sg13g2_fill_8 FILLER_111_320 ();
 sg13g2_fill_8 FILLER_111_328 ();
 sg13g2_fill_8 FILLER_111_336 ();
 sg13g2_fill_8 FILLER_111_344 ();
 sg13g2_fill_8 FILLER_111_352 ();
 sg13g2_fill_8 FILLER_111_360 ();
 sg13g2_fill_8 FILLER_111_368 ();
 sg13g2_fill_8 FILLER_111_376 ();
 sg13g2_fill_8 FILLER_111_384 ();
 sg13g2_fill_8 FILLER_111_392 ();
 sg13g2_fill_8 FILLER_111_400 ();
 sg13g2_fill_8 FILLER_111_408 ();
 sg13g2_fill_8 FILLER_111_416 ();
 sg13g2_fill_8 FILLER_111_424 ();
 sg13g2_fill_8 FILLER_111_432 ();
 sg13g2_fill_8 FILLER_111_440 ();
 sg13g2_fill_8 FILLER_111_448 ();
 sg13g2_fill_8 FILLER_111_456 ();
 sg13g2_fill_8 FILLER_111_464 ();
 sg13g2_fill_8 FILLER_111_472 ();
 sg13g2_fill_8 FILLER_111_480 ();
 sg13g2_fill_8 FILLER_111_488 ();
 sg13g2_fill_8 FILLER_111_496 ();
 sg13g2_fill_8 FILLER_111_504 ();
 sg13g2_fill_8 FILLER_111_512 ();
 sg13g2_fill_8 FILLER_111_520 ();
 sg13g2_fill_8 FILLER_111_528 ();
 sg13g2_fill_8 FILLER_111_536 ();
 sg13g2_fill_8 FILLER_111_544 ();
 sg13g2_fill_8 FILLER_111_552 ();
 sg13g2_fill_8 FILLER_111_560 ();
 sg13g2_fill_8 FILLER_111_568 ();
 sg13g2_fill_8 FILLER_111_576 ();
 sg13g2_fill_8 FILLER_111_584 ();
 sg13g2_fill_8 FILLER_111_592 ();
 sg13g2_fill_8 FILLER_111_600 ();
 sg13g2_fill_8 FILLER_111_608 ();
 sg13g2_fill_8 FILLER_111_616 ();
 sg13g2_fill_8 FILLER_111_624 ();
 sg13g2_fill_8 FILLER_111_632 ();
 sg13g2_fill_8 FILLER_111_640 ();
 sg13g2_fill_8 FILLER_111_648 ();
 sg13g2_fill_8 FILLER_111_656 ();
 sg13g2_fill_8 FILLER_111_664 ();
 sg13g2_fill_8 FILLER_111_672 ();
 sg13g2_fill_8 FILLER_111_680 ();
 sg13g2_fill_8 FILLER_111_688 ();
 sg13g2_fill_8 FILLER_111_696 ();
 sg13g2_fill_8 FILLER_111_704 ();
 sg13g2_fill_8 FILLER_111_712 ();
 sg13g2_fill_8 FILLER_111_720 ();
 sg13g2_fill_8 FILLER_111_728 ();
 sg13g2_fill_8 FILLER_111_736 ();
 sg13g2_fill_8 FILLER_111_744 ();
 sg13g2_fill_8 FILLER_111_752 ();
 sg13g2_fill_8 FILLER_111_760 ();
 sg13g2_fill_8 FILLER_111_768 ();
 sg13g2_fill_8 FILLER_111_776 ();
 sg13g2_fill_8 FILLER_111_784 ();
 sg13g2_fill_8 FILLER_111_792 ();
 sg13g2_fill_8 FILLER_111_800 ();
 sg13g2_fill_8 FILLER_111_808 ();
 sg13g2_fill_8 FILLER_111_816 ();
 sg13g2_fill_8 FILLER_111_824 ();
 sg13g2_fill_8 FILLER_111_832 ();
 sg13g2_fill_8 FILLER_111_840 ();
 sg13g2_fill_8 FILLER_111_848 ();
 sg13g2_fill_8 FILLER_111_856 ();
 sg13g2_fill_8 FILLER_111_864 ();
 sg13g2_fill_8 FILLER_111_872 ();
 sg13g2_fill_8 FILLER_111_880 ();
 sg13g2_fill_8 FILLER_111_888 ();
 sg13g2_fill_8 FILLER_111_896 ();
 sg13g2_fill_8 FILLER_111_904 ();
 sg13g2_fill_8 FILLER_111_912 ();
 sg13g2_fill_8 FILLER_111_920 ();
 sg13g2_fill_8 FILLER_111_928 ();
 sg13g2_fill_8 FILLER_111_936 ();
 sg13g2_fill_8 FILLER_111_944 ();
 sg13g2_fill_8 FILLER_111_952 ();
 sg13g2_fill_8 FILLER_111_960 ();
 sg13g2_fill_8 FILLER_111_968 ();
 sg13g2_fill_8 FILLER_111_976 ();
 sg13g2_fill_8 FILLER_111_984 ();
 sg13g2_fill_8 FILLER_111_992 ();
 sg13g2_fill_8 FILLER_111_1000 ();
 sg13g2_fill_8 FILLER_111_1008 ();
 sg13g2_fill_8 FILLER_111_1016 ();
 sg13g2_fill_8 FILLER_111_1024 ();
 sg13g2_fill_8 FILLER_111_1032 ();
 sg13g2_fill_8 FILLER_111_1040 ();
 sg13g2_fill_8 FILLER_111_1048 ();
 sg13g2_fill_8 FILLER_111_1056 ();
 sg13g2_fill_8 FILLER_111_1064 ();
 sg13g2_fill_8 FILLER_111_1072 ();
 sg13g2_fill_8 FILLER_111_1080 ();
 sg13g2_fill_8 FILLER_111_1088 ();
 sg13g2_fill_8 FILLER_111_1096 ();
 sg13g2_fill_8 FILLER_111_1104 ();
 sg13g2_fill_8 FILLER_111_1112 ();
 sg13g2_fill_8 FILLER_111_1120 ();
 sg13g2_fill_8 FILLER_111_1128 ();
 sg13g2_fill_8 FILLER_111_1136 ();
 sg13g2_fill_8 FILLER_111_1144 ();
 sg13g2_fill_8 FILLER_111_1152 ();
 sg13g2_fill_4 FILLER_111_1160 ();
 sg13g2_fill_2 FILLER_111_1164 ();
 sg13g2_fill_8 FILLER_112_0 ();
 sg13g2_fill_8 FILLER_112_8 ();
 sg13g2_fill_8 FILLER_112_16 ();
 sg13g2_fill_8 FILLER_112_24 ();
 sg13g2_fill_8 FILLER_112_32 ();
 sg13g2_fill_8 FILLER_112_40 ();
 sg13g2_fill_8 FILLER_112_48 ();
 sg13g2_fill_8 FILLER_112_56 ();
 sg13g2_fill_8 FILLER_112_64 ();
 sg13g2_fill_8 FILLER_112_72 ();
 sg13g2_fill_8 FILLER_112_80 ();
 sg13g2_fill_8 FILLER_112_88 ();
 sg13g2_fill_8 FILLER_112_96 ();
 sg13g2_fill_8 FILLER_112_104 ();
 sg13g2_fill_8 FILLER_112_112 ();
 sg13g2_fill_8 FILLER_112_120 ();
 sg13g2_fill_8 FILLER_112_128 ();
 sg13g2_fill_8 FILLER_112_136 ();
 sg13g2_fill_8 FILLER_112_144 ();
 sg13g2_fill_8 FILLER_112_152 ();
 sg13g2_fill_8 FILLER_112_160 ();
 sg13g2_fill_8 FILLER_112_168 ();
 sg13g2_fill_8 FILLER_112_176 ();
 sg13g2_fill_8 FILLER_112_184 ();
 sg13g2_fill_8 FILLER_112_192 ();
 sg13g2_fill_8 FILLER_112_200 ();
 sg13g2_fill_8 FILLER_112_208 ();
 sg13g2_fill_8 FILLER_112_216 ();
 sg13g2_fill_8 FILLER_112_224 ();
 sg13g2_fill_8 FILLER_112_232 ();
 sg13g2_fill_8 FILLER_112_240 ();
 sg13g2_fill_8 FILLER_112_248 ();
 sg13g2_fill_8 FILLER_112_256 ();
 sg13g2_fill_8 FILLER_112_264 ();
 sg13g2_fill_8 FILLER_112_272 ();
 sg13g2_fill_8 FILLER_112_280 ();
 sg13g2_fill_8 FILLER_112_288 ();
 sg13g2_fill_8 FILLER_112_296 ();
 sg13g2_fill_8 FILLER_112_304 ();
 sg13g2_fill_8 FILLER_112_312 ();
 sg13g2_fill_8 FILLER_112_320 ();
 sg13g2_fill_8 FILLER_112_328 ();
 sg13g2_fill_8 FILLER_112_336 ();
 sg13g2_fill_8 FILLER_112_344 ();
 sg13g2_fill_8 FILLER_112_352 ();
 sg13g2_fill_8 FILLER_112_360 ();
 sg13g2_fill_8 FILLER_112_368 ();
 sg13g2_fill_8 FILLER_112_376 ();
 sg13g2_fill_8 FILLER_112_384 ();
 sg13g2_fill_8 FILLER_112_392 ();
 sg13g2_fill_8 FILLER_112_400 ();
 sg13g2_fill_8 FILLER_112_408 ();
 sg13g2_fill_8 FILLER_112_416 ();
 sg13g2_fill_8 FILLER_112_424 ();
 sg13g2_fill_8 FILLER_112_432 ();
 sg13g2_fill_8 FILLER_112_440 ();
 sg13g2_fill_8 FILLER_112_448 ();
 sg13g2_fill_8 FILLER_112_456 ();
 sg13g2_fill_8 FILLER_112_464 ();
 sg13g2_fill_8 FILLER_112_472 ();
 sg13g2_fill_8 FILLER_112_480 ();
 sg13g2_fill_8 FILLER_112_488 ();
 sg13g2_fill_8 FILLER_112_496 ();
 sg13g2_fill_8 FILLER_112_504 ();
 sg13g2_fill_8 FILLER_112_512 ();
 sg13g2_fill_8 FILLER_112_520 ();
 sg13g2_fill_8 FILLER_112_528 ();
 sg13g2_fill_8 FILLER_112_536 ();
 sg13g2_fill_8 FILLER_112_544 ();
 sg13g2_fill_8 FILLER_112_552 ();
 sg13g2_fill_8 FILLER_112_560 ();
 sg13g2_fill_8 FILLER_112_568 ();
 sg13g2_fill_8 FILLER_112_576 ();
 sg13g2_fill_8 FILLER_112_584 ();
 sg13g2_fill_8 FILLER_112_592 ();
 sg13g2_fill_8 FILLER_112_600 ();
 sg13g2_fill_8 FILLER_112_608 ();
 sg13g2_fill_8 FILLER_112_616 ();
 sg13g2_fill_8 FILLER_112_624 ();
 sg13g2_fill_8 FILLER_112_632 ();
 sg13g2_fill_8 FILLER_112_640 ();
 sg13g2_fill_8 FILLER_112_648 ();
 sg13g2_fill_8 FILLER_112_656 ();
 sg13g2_fill_8 FILLER_112_664 ();
 sg13g2_fill_8 FILLER_112_672 ();
 sg13g2_fill_8 FILLER_112_680 ();
 sg13g2_fill_8 FILLER_112_688 ();
 sg13g2_fill_8 FILLER_112_696 ();
 sg13g2_fill_8 FILLER_112_704 ();
 sg13g2_fill_8 FILLER_112_712 ();
 sg13g2_fill_8 FILLER_112_720 ();
 sg13g2_fill_8 FILLER_112_728 ();
 sg13g2_fill_8 FILLER_112_736 ();
 sg13g2_fill_8 FILLER_112_744 ();
 sg13g2_fill_8 FILLER_112_752 ();
 sg13g2_fill_8 FILLER_112_760 ();
 sg13g2_fill_8 FILLER_112_768 ();
 sg13g2_fill_8 FILLER_112_776 ();
 sg13g2_fill_8 FILLER_112_784 ();
 sg13g2_fill_8 FILLER_112_792 ();
 sg13g2_fill_8 FILLER_112_800 ();
 sg13g2_fill_8 FILLER_112_808 ();
 sg13g2_fill_8 FILLER_112_816 ();
 sg13g2_fill_8 FILLER_112_824 ();
 sg13g2_fill_8 FILLER_112_832 ();
 sg13g2_fill_8 FILLER_112_840 ();
 sg13g2_fill_8 FILLER_112_848 ();
 sg13g2_fill_8 FILLER_112_856 ();
 sg13g2_fill_8 FILLER_112_864 ();
 sg13g2_fill_8 FILLER_112_872 ();
 sg13g2_fill_8 FILLER_112_880 ();
 sg13g2_fill_8 FILLER_112_888 ();
 sg13g2_fill_8 FILLER_112_896 ();
 sg13g2_fill_8 FILLER_112_904 ();
 sg13g2_fill_8 FILLER_112_912 ();
 sg13g2_fill_8 FILLER_112_920 ();
 sg13g2_fill_8 FILLER_112_928 ();
 sg13g2_fill_8 FILLER_112_936 ();
 sg13g2_fill_8 FILLER_112_944 ();
 sg13g2_fill_8 FILLER_112_952 ();
 sg13g2_fill_8 FILLER_112_960 ();
 sg13g2_fill_8 FILLER_112_968 ();
 sg13g2_fill_8 FILLER_112_976 ();
 sg13g2_fill_8 FILLER_112_984 ();
 sg13g2_fill_8 FILLER_112_992 ();
 sg13g2_fill_8 FILLER_112_1000 ();
 sg13g2_fill_8 FILLER_112_1008 ();
 sg13g2_fill_8 FILLER_112_1016 ();
 sg13g2_fill_8 FILLER_112_1024 ();
 sg13g2_fill_8 FILLER_112_1032 ();
 sg13g2_fill_8 FILLER_112_1040 ();
 sg13g2_fill_8 FILLER_112_1048 ();
 sg13g2_fill_8 FILLER_112_1056 ();
 sg13g2_fill_8 FILLER_112_1064 ();
 sg13g2_fill_8 FILLER_112_1072 ();
 sg13g2_fill_8 FILLER_112_1080 ();
 sg13g2_fill_8 FILLER_112_1088 ();
 sg13g2_fill_8 FILLER_112_1096 ();
 sg13g2_fill_8 FILLER_112_1104 ();
 sg13g2_fill_8 FILLER_112_1112 ();
 sg13g2_fill_8 FILLER_112_1120 ();
 sg13g2_fill_8 FILLER_112_1128 ();
 sg13g2_fill_8 FILLER_112_1136 ();
 sg13g2_fill_8 FILLER_112_1144 ();
 sg13g2_fill_8 FILLER_112_1152 ();
 sg13g2_fill_4 FILLER_112_1160 ();
 sg13g2_fill_2 FILLER_112_1164 ();
 sg13g2_fill_8 FILLER_113_0 ();
 sg13g2_fill_8 FILLER_113_8 ();
 sg13g2_fill_8 FILLER_113_16 ();
 sg13g2_fill_8 FILLER_113_24 ();
 sg13g2_fill_8 FILLER_113_32 ();
 sg13g2_fill_8 FILLER_113_40 ();
 sg13g2_fill_8 FILLER_113_48 ();
 sg13g2_fill_8 FILLER_113_56 ();
 sg13g2_fill_8 FILLER_113_64 ();
 sg13g2_fill_8 FILLER_113_72 ();
 sg13g2_fill_8 FILLER_113_80 ();
 sg13g2_fill_8 FILLER_113_88 ();
 sg13g2_fill_8 FILLER_113_96 ();
 sg13g2_fill_8 FILLER_113_104 ();
 sg13g2_fill_8 FILLER_113_112 ();
 sg13g2_fill_8 FILLER_113_120 ();
 sg13g2_fill_8 FILLER_113_128 ();
 sg13g2_fill_8 FILLER_113_136 ();
 sg13g2_fill_8 FILLER_113_144 ();
 sg13g2_fill_8 FILLER_113_152 ();
 sg13g2_fill_8 FILLER_113_160 ();
 sg13g2_fill_8 FILLER_113_168 ();
 sg13g2_fill_8 FILLER_113_176 ();
 sg13g2_fill_8 FILLER_113_184 ();
 sg13g2_fill_8 FILLER_113_192 ();
 sg13g2_fill_8 FILLER_113_200 ();
 sg13g2_fill_8 FILLER_113_208 ();
 sg13g2_fill_8 FILLER_113_216 ();
 sg13g2_fill_8 FILLER_113_224 ();
 sg13g2_fill_8 FILLER_113_232 ();
 sg13g2_fill_8 FILLER_113_240 ();
 sg13g2_fill_8 FILLER_113_248 ();
 sg13g2_fill_8 FILLER_113_256 ();
 sg13g2_fill_8 FILLER_113_264 ();
 sg13g2_fill_8 FILLER_113_272 ();
 sg13g2_fill_8 FILLER_113_280 ();
 sg13g2_fill_8 FILLER_113_288 ();
 sg13g2_fill_8 FILLER_113_296 ();
 sg13g2_fill_8 FILLER_113_304 ();
 sg13g2_fill_8 FILLER_113_312 ();
 sg13g2_fill_8 FILLER_113_320 ();
 sg13g2_fill_8 FILLER_113_328 ();
 sg13g2_fill_8 FILLER_113_336 ();
 sg13g2_fill_8 FILLER_113_344 ();
 sg13g2_fill_8 FILLER_113_352 ();
 sg13g2_fill_8 FILLER_113_360 ();
 sg13g2_fill_8 FILLER_113_368 ();
 sg13g2_fill_8 FILLER_113_376 ();
 sg13g2_fill_8 FILLER_113_384 ();
 sg13g2_fill_8 FILLER_113_392 ();
 sg13g2_fill_8 FILLER_113_400 ();
 sg13g2_fill_8 FILLER_113_408 ();
 sg13g2_fill_8 FILLER_113_416 ();
 sg13g2_fill_8 FILLER_113_424 ();
 sg13g2_fill_8 FILLER_113_432 ();
 sg13g2_fill_8 FILLER_113_440 ();
 sg13g2_fill_8 FILLER_113_448 ();
 sg13g2_fill_8 FILLER_113_456 ();
 sg13g2_fill_8 FILLER_113_464 ();
 sg13g2_fill_8 FILLER_113_472 ();
 sg13g2_fill_8 FILLER_113_480 ();
 sg13g2_fill_8 FILLER_113_488 ();
 sg13g2_fill_8 FILLER_113_496 ();
 sg13g2_fill_8 FILLER_113_504 ();
 sg13g2_fill_8 FILLER_113_512 ();
 sg13g2_fill_8 FILLER_113_520 ();
 sg13g2_fill_8 FILLER_113_528 ();
 sg13g2_fill_8 FILLER_113_536 ();
 sg13g2_fill_8 FILLER_113_544 ();
 sg13g2_fill_8 FILLER_113_552 ();
 sg13g2_fill_8 FILLER_113_560 ();
 sg13g2_fill_8 FILLER_113_568 ();
 sg13g2_fill_8 FILLER_113_576 ();
 sg13g2_fill_8 FILLER_113_584 ();
 sg13g2_fill_8 FILLER_113_592 ();
 sg13g2_fill_8 FILLER_113_600 ();
 sg13g2_fill_8 FILLER_113_608 ();
 sg13g2_fill_8 FILLER_113_616 ();
 sg13g2_fill_8 FILLER_113_624 ();
 sg13g2_fill_8 FILLER_113_632 ();
 sg13g2_fill_8 FILLER_113_640 ();
 sg13g2_fill_8 FILLER_113_648 ();
 sg13g2_fill_8 FILLER_113_656 ();
 sg13g2_fill_8 FILLER_113_664 ();
 sg13g2_fill_8 FILLER_113_672 ();
 sg13g2_fill_8 FILLER_113_680 ();
 sg13g2_fill_8 FILLER_113_688 ();
 sg13g2_fill_8 FILLER_113_696 ();
 sg13g2_fill_8 FILLER_113_704 ();
 sg13g2_fill_8 FILLER_113_712 ();
 sg13g2_fill_8 FILLER_113_720 ();
 sg13g2_fill_8 FILLER_113_728 ();
 sg13g2_fill_8 FILLER_113_736 ();
 sg13g2_fill_8 FILLER_113_744 ();
 sg13g2_fill_8 FILLER_113_752 ();
 sg13g2_fill_8 FILLER_113_760 ();
 sg13g2_fill_8 FILLER_113_768 ();
 sg13g2_fill_8 FILLER_113_776 ();
 sg13g2_fill_8 FILLER_113_784 ();
 sg13g2_fill_8 FILLER_113_792 ();
 sg13g2_fill_8 FILLER_113_800 ();
 sg13g2_fill_8 FILLER_113_808 ();
 sg13g2_fill_8 FILLER_113_816 ();
 sg13g2_fill_8 FILLER_113_824 ();
 sg13g2_fill_8 FILLER_113_832 ();
 sg13g2_fill_8 FILLER_113_840 ();
 sg13g2_fill_8 FILLER_113_848 ();
 sg13g2_fill_8 FILLER_113_856 ();
 sg13g2_fill_8 FILLER_113_864 ();
 sg13g2_fill_8 FILLER_113_872 ();
 sg13g2_fill_8 FILLER_113_880 ();
 sg13g2_fill_8 FILLER_113_888 ();
 sg13g2_fill_8 FILLER_113_896 ();
 sg13g2_fill_8 FILLER_113_904 ();
 sg13g2_fill_8 FILLER_113_912 ();
 sg13g2_fill_8 FILLER_113_920 ();
 sg13g2_fill_8 FILLER_113_928 ();
 sg13g2_fill_8 FILLER_113_936 ();
 sg13g2_fill_8 FILLER_113_944 ();
 sg13g2_fill_8 FILLER_113_952 ();
 sg13g2_fill_8 FILLER_113_960 ();
 sg13g2_fill_8 FILLER_113_968 ();
 sg13g2_fill_8 FILLER_113_976 ();
 sg13g2_fill_8 FILLER_113_984 ();
 sg13g2_fill_8 FILLER_113_992 ();
 sg13g2_fill_8 FILLER_113_1000 ();
 sg13g2_fill_8 FILLER_113_1008 ();
 sg13g2_fill_8 FILLER_113_1016 ();
 sg13g2_fill_8 FILLER_113_1024 ();
 sg13g2_fill_8 FILLER_113_1032 ();
 sg13g2_fill_8 FILLER_113_1040 ();
 sg13g2_fill_8 FILLER_113_1048 ();
 sg13g2_fill_8 FILLER_113_1056 ();
 sg13g2_fill_8 FILLER_113_1064 ();
 sg13g2_fill_8 FILLER_113_1072 ();
 sg13g2_fill_8 FILLER_113_1080 ();
 sg13g2_fill_8 FILLER_113_1088 ();
 sg13g2_fill_8 FILLER_113_1096 ();
 sg13g2_fill_8 FILLER_113_1104 ();
 sg13g2_fill_8 FILLER_113_1112 ();
 sg13g2_fill_8 FILLER_113_1120 ();
 sg13g2_fill_8 FILLER_113_1128 ();
 sg13g2_fill_8 FILLER_113_1136 ();
 sg13g2_fill_8 FILLER_113_1144 ();
 sg13g2_fill_8 FILLER_113_1152 ();
 sg13g2_fill_4 FILLER_113_1160 ();
 sg13g2_fill_2 FILLER_113_1164 ();
 sg13g2_fill_8 FILLER_114_0 ();
 sg13g2_fill_8 FILLER_114_8 ();
 sg13g2_fill_8 FILLER_114_16 ();
 sg13g2_fill_8 FILLER_114_24 ();
 sg13g2_fill_8 FILLER_114_32 ();
 sg13g2_fill_8 FILLER_114_40 ();
 sg13g2_fill_8 FILLER_114_48 ();
 sg13g2_fill_8 FILLER_114_56 ();
 sg13g2_fill_8 FILLER_114_64 ();
 sg13g2_fill_8 FILLER_114_72 ();
 sg13g2_fill_8 FILLER_114_80 ();
 sg13g2_fill_8 FILLER_114_88 ();
 sg13g2_fill_8 FILLER_114_96 ();
 sg13g2_fill_8 FILLER_114_104 ();
 sg13g2_fill_8 FILLER_114_112 ();
 sg13g2_fill_8 FILLER_114_120 ();
 sg13g2_fill_8 FILLER_114_128 ();
 sg13g2_fill_8 FILLER_114_136 ();
 sg13g2_fill_8 FILLER_114_144 ();
 sg13g2_fill_8 FILLER_114_152 ();
 sg13g2_fill_8 FILLER_114_160 ();
 sg13g2_fill_8 FILLER_114_168 ();
 sg13g2_fill_8 FILLER_114_176 ();
 sg13g2_fill_8 FILLER_114_184 ();
 sg13g2_fill_8 FILLER_114_192 ();
 sg13g2_fill_8 FILLER_114_200 ();
 sg13g2_fill_8 FILLER_114_208 ();
 sg13g2_fill_8 FILLER_114_216 ();
 sg13g2_fill_8 FILLER_114_224 ();
 sg13g2_fill_8 FILLER_114_232 ();
 sg13g2_fill_8 FILLER_114_240 ();
 sg13g2_fill_8 FILLER_114_248 ();
 sg13g2_fill_8 FILLER_114_256 ();
 sg13g2_fill_8 FILLER_114_264 ();
 sg13g2_fill_8 FILLER_114_272 ();
 sg13g2_fill_8 FILLER_114_280 ();
 sg13g2_fill_8 FILLER_114_288 ();
 sg13g2_fill_8 FILLER_114_296 ();
 sg13g2_fill_8 FILLER_114_304 ();
 sg13g2_fill_8 FILLER_114_312 ();
 sg13g2_fill_8 FILLER_114_320 ();
 sg13g2_fill_8 FILLER_114_328 ();
 sg13g2_fill_8 FILLER_114_336 ();
 sg13g2_fill_8 FILLER_114_344 ();
 sg13g2_fill_8 FILLER_114_352 ();
 sg13g2_fill_8 FILLER_114_360 ();
 sg13g2_fill_8 FILLER_114_368 ();
 sg13g2_fill_8 FILLER_114_376 ();
 sg13g2_fill_8 FILLER_114_384 ();
 sg13g2_fill_8 FILLER_114_392 ();
 sg13g2_fill_8 FILLER_114_400 ();
 sg13g2_fill_8 FILLER_114_408 ();
 sg13g2_fill_8 FILLER_114_416 ();
 sg13g2_fill_8 FILLER_114_424 ();
 sg13g2_fill_8 FILLER_114_432 ();
 sg13g2_fill_8 FILLER_114_440 ();
 sg13g2_fill_8 FILLER_114_448 ();
 sg13g2_fill_8 FILLER_114_456 ();
 sg13g2_fill_8 FILLER_114_464 ();
 sg13g2_fill_8 FILLER_114_472 ();
 sg13g2_fill_8 FILLER_114_480 ();
 sg13g2_fill_8 FILLER_114_488 ();
 sg13g2_fill_8 FILLER_114_496 ();
 sg13g2_fill_8 FILLER_114_504 ();
 sg13g2_fill_8 FILLER_114_512 ();
 sg13g2_fill_8 FILLER_114_520 ();
 sg13g2_fill_8 FILLER_114_528 ();
 sg13g2_fill_8 FILLER_114_536 ();
 sg13g2_fill_8 FILLER_114_544 ();
 sg13g2_fill_8 FILLER_114_552 ();
 sg13g2_fill_8 FILLER_114_560 ();
 sg13g2_fill_8 FILLER_114_568 ();
 sg13g2_fill_8 FILLER_114_576 ();
 sg13g2_fill_8 FILLER_114_584 ();
 sg13g2_fill_8 FILLER_114_592 ();
 sg13g2_fill_8 FILLER_114_600 ();
 sg13g2_fill_8 FILLER_114_608 ();
 sg13g2_fill_8 FILLER_114_616 ();
 sg13g2_fill_8 FILLER_114_624 ();
 sg13g2_fill_8 FILLER_114_632 ();
 sg13g2_fill_8 FILLER_114_640 ();
 sg13g2_fill_8 FILLER_114_648 ();
 sg13g2_fill_8 FILLER_114_656 ();
 sg13g2_fill_8 FILLER_114_664 ();
 sg13g2_fill_8 FILLER_114_672 ();
 sg13g2_fill_8 FILLER_114_680 ();
 sg13g2_fill_8 FILLER_114_688 ();
 sg13g2_fill_8 FILLER_114_696 ();
 sg13g2_fill_8 FILLER_114_704 ();
 sg13g2_fill_8 FILLER_114_712 ();
 sg13g2_fill_8 FILLER_114_720 ();
 sg13g2_fill_8 FILLER_114_728 ();
 sg13g2_fill_8 FILLER_114_736 ();
 sg13g2_fill_8 FILLER_114_744 ();
 sg13g2_fill_8 FILLER_114_752 ();
 sg13g2_fill_8 FILLER_114_760 ();
 sg13g2_fill_8 FILLER_114_768 ();
 sg13g2_fill_8 FILLER_114_776 ();
 sg13g2_fill_8 FILLER_114_784 ();
 sg13g2_fill_8 FILLER_114_792 ();
 sg13g2_fill_8 FILLER_114_800 ();
 sg13g2_fill_8 FILLER_114_808 ();
 sg13g2_fill_8 FILLER_114_816 ();
 sg13g2_fill_8 FILLER_114_824 ();
 sg13g2_fill_8 FILLER_114_832 ();
 sg13g2_fill_8 FILLER_114_840 ();
 sg13g2_fill_8 FILLER_114_848 ();
 sg13g2_fill_8 FILLER_114_856 ();
 sg13g2_fill_8 FILLER_114_864 ();
 sg13g2_fill_8 FILLER_114_872 ();
 sg13g2_fill_8 FILLER_114_880 ();
 sg13g2_fill_8 FILLER_114_888 ();
 sg13g2_fill_8 FILLER_114_896 ();
 sg13g2_fill_8 FILLER_114_904 ();
 sg13g2_fill_8 FILLER_114_912 ();
 sg13g2_fill_8 FILLER_114_920 ();
 sg13g2_fill_8 FILLER_114_928 ();
 sg13g2_fill_8 FILLER_114_936 ();
 sg13g2_fill_8 FILLER_114_944 ();
 sg13g2_fill_8 FILLER_114_952 ();
 sg13g2_fill_8 FILLER_114_960 ();
 sg13g2_fill_8 FILLER_114_968 ();
 sg13g2_fill_8 FILLER_114_976 ();
 sg13g2_fill_8 FILLER_114_984 ();
 sg13g2_fill_8 FILLER_114_992 ();
 sg13g2_fill_8 FILLER_114_1000 ();
 sg13g2_fill_8 FILLER_114_1008 ();
 sg13g2_fill_8 FILLER_114_1016 ();
 sg13g2_fill_8 FILLER_114_1024 ();
 sg13g2_fill_8 FILLER_114_1032 ();
 sg13g2_fill_8 FILLER_114_1040 ();
 sg13g2_fill_8 FILLER_114_1048 ();
 sg13g2_fill_8 FILLER_114_1056 ();
 sg13g2_fill_8 FILLER_114_1064 ();
 sg13g2_fill_8 FILLER_114_1072 ();
 sg13g2_fill_8 FILLER_114_1080 ();
 sg13g2_fill_8 FILLER_114_1088 ();
 sg13g2_fill_8 FILLER_114_1096 ();
 sg13g2_fill_8 FILLER_114_1104 ();
 sg13g2_fill_8 FILLER_114_1112 ();
 sg13g2_fill_8 FILLER_114_1120 ();
 sg13g2_fill_8 FILLER_114_1128 ();
 sg13g2_fill_8 FILLER_114_1136 ();
 sg13g2_fill_8 FILLER_114_1144 ();
 sg13g2_fill_8 FILLER_114_1152 ();
 sg13g2_fill_4 FILLER_114_1160 ();
 sg13g2_fill_2 FILLER_114_1164 ();
 sg13g2_fill_8 FILLER_115_0 ();
 sg13g2_fill_8 FILLER_115_8 ();
 sg13g2_fill_8 FILLER_115_16 ();
 sg13g2_fill_8 FILLER_115_24 ();
 sg13g2_fill_8 FILLER_115_32 ();
 sg13g2_fill_8 FILLER_115_40 ();
 sg13g2_fill_8 FILLER_115_48 ();
 sg13g2_fill_8 FILLER_115_56 ();
 sg13g2_fill_8 FILLER_115_64 ();
 sg13g2_fill_8 FILLER_115_72 ();
 sg13g2_fill_8 FILLER_115_80 ();
 sg13g2_fill_8 FILLER_115_88 ();
 sg13g2_fill_8 FILLER_115_96 ();
 sg13g2_fill_8 FILLER_115_104 ();
 sg13g2_fill_8 FILLER_115_112 ();
 sg13g2_fill_8 FILLER_115_120 ();
 sg13g2_fill_8 FILLER_115_128 ();
 sg13g2_fill_8 FILLER_115_136 ();
 sg13g2_fill_8 FILLER_115_144 ();
 sg13g2_fill_8 FILLER_115_152 ();
 sg13g2_fill_8 FILLER_115_160 ();
 sg13g2_fill_8 FILLER_115_168 ();
 sg13g2_fill_8 FILLER_115_176 ();
 sg13g2_fill_8 FILLER_115_184 ();
 sg13g2_fill_8 FILLER_115_192 ();
 sg13g2_fill_8 FILLER_115_200 ();
 sg13g2_fill_8 FILLER_115_208 ();
 sg13g2_fill_8 FILLER_115_216 ();
 sg13g2_fill_8 FILLER_115_224 ();
 sg13g2_fill_8 FILLER_115_232 ();
 sg13g2_fill_8 FILLER_115_240 ();
 sg13g2_fill_8 FILLER_115_248 ();
 sg13g2_fill_8 FILLER_115_256 ();
 sg13g2_fill_8 FILLER_115_264 ();
 sg13g2_fill_8 FILLER_115_272 ();
 sg13g2_fill_8 FILLER_115_280 ();
 sg13g2_fill_8 FILLER_115_288 ();
 sg13g2_fill_8 FILLER_115_296 ();
 sg13g2_fill_8 FILLER_115_304 ();
 sg13g2_fill_8 FILLER_115_312 ();
 sg13g2_fill_8 FILLER_115_320 ();
 sg13g2_fill_8 FILLER_115_328 ();
 sg13g2_fill_8 FILLER_115_336 ();
 sg13g2_fill_8 FILLER_115_344 ();
 sg13g2_fill_8 FILLER_115_352 ();
 sg13g2_fill_8 FILLER_115_360 ();
 sg13g2_fill_8 FILLER_115_368 ();
 sg13g2_fill_8 FILLER_115_376 ();
 sg13g2_fill_8 FILLER_115_384 ();
 sg13g2_fill_8 FILLER_115_392 ();
 sg13g2_fill_8 FILLER_115_400 ();
 sg13g2_fill_8 FILLER_115_408 ();
 sg13g2_fill_8 FILLER_115_416 ();
 sg13g2_fill_8 FILLER_115_424 ();
 sg13g2_fill_8 FILLER_115_432 ();
 sg13g2_fill_8 FILLER_115_440 ();
 sg13g2_fill_8 FILLER_115_448 ();
 sg13g2_fill_8 FILLER_115_456 ();
 sg13g2_fill_8 FILLER_115_464 ();
 sg13g2_fill_8 FILLER_115_472 ();
 sg13g2_fill_8 FILLER_115_480 ();
 sg13g2_fill_8 FILLER_115_488 ();
 sg13g2_fill_8 FILLER_115_496 ();
 sg13g2_fill_8 FILLER_115_504 ();
 sg13g2_fill_8 FILLER_115_512 ();
 sg13g2_fill_8 FILLER_115_520 ();
 sg13g2_fill_8 FILLER_115_528 ();
 sg13g2_fill_8 FILLER_115_536 ();
 sg13g2_fill_8 FILLER_115_544 ();
 sg13g2_fill_8 FILLER_115_552 ();
 sg13g2_fill_8 FILLER_115_560 ();
 sg13g2_fill_8 FILLER_115_568 ();
 sg13g2_fill_8 FILLER_115_576 ();
 sg13g2_fill_8 FILLER_115_584 ();
 sg13g2_fill_8 FILLER_115_592 ();
 sg13g2_fill_8 FILLER_115_600 ();
 sg13g2_fill_8 FILLER_115_608 ();
 sg13g2_fill_8 FILLER_115_616 ();
 sg13g2_fill_8 FILLER_115_624 ();
 sg13g2_fill_8 FILLER_115_632 ();
 sg13g2_fill_8 FILLER_115_640 ();
 sg13g2_fill_8 FILLER_115_648 ();
 sg13g2_fill_8 FILLER_115_656 ();
 sg13g2_fill_8 FILLER_115_664 ();
 sg13g2_fill_8 FILLER_115_672 ();
 sg13g2_fill_8 FILLER_115_680 ();
 sg13g2_fill_8 FILLER_115_688 ();
 sg13g2_fill_8 FILLER_115_696 ();
 sg13g2_fill_8 FILLER_115_704 ();
 sg13g2_fill_8 FILLER_115_712 ();
 sg13g2_fill_8 FILLER_115_720 ();
 sg13g2_fill_8 FILLER_115_728 ();
 sg13g2_fill_8 FILLER_115_736 ();
 sg13g2_fill_8 FILLER_115_744 ();
 sg13g2_fill_8 FILLER_115_752 ();
 sg13g2_fill_8 FILLER_115_760 ();
 sg13g2_fill_8 FILLER_115_768 ();
 sg13g2_fill_8 FILLER_115_776 ();
 sg13g2_fill_8 FILLER_115_784 ();
 sg13g2_fill_8 FILLER_115_792 ();
 sg13g2_fill_8 FILLER_115_800 ();
 sg13g2_fill_8 FILLER_115_808 ();
 sg13g2_fill_8 FILLER_115_816 ();
 sg13g2_fill_8 FILLER_115_824 ();
 sg13g2_fill_8 FILLER_115_832 ();
 sg13g2_fill_8 FILLER_115_840 ();
 sg13g2_fill_8 FILLER_115_848 ();
 sg13g2_fill_8 FILLER_115_856 ();
 sg13g2_fill_8 FILLER_115_864 ();
 sg13g2_fill_8 FILLER_115_872 ();
 sg13g2_fill_8 FILLER_115_880 ();
 sg13g2_fill_8 FILLER_115_888 ();
 sg13g2_fill_8 FILLER_115_896 ();
 sg13g2_fill_8 FILLER_115_904 ();
 sg13g2_fill_8 FILLER_115_912 ();
 sg13g2_fill_8 FILLER_115_920 ();
 sg13g2_fill_8 FILLER_115_928 ();
 sg13g2_fill_8 FILLER_115_936 ();
 sg13g2_fill_8 FILLER_115_944 ();
 sg13g2_fill_8 FILLER_115_952 ();
 sg13g2_fill_8 FILLER_115_960 ();
 sg13g2_fill_8 FILLER_115_968 ();
 sg13g2_fill_8 FILLER_115_976 ();
 sg13g2_fill_8 FILLER_115_984 ();
 sg13g2_fill_8 FILLER_115_992 ();
 sg13g2_fill_8 FILLER_115_1000 ();
 sg13g2_fill_8 FILLER_115_1008 ();
 sg13g2_fill_8 FILLER_115_1016 ();
 sg13g2_fill_8 FILLER_115_1024 ();
 sg13g2_fill_8 FILLER_115_1032 ();
 sg13g2_fill_8 FILLER_115_1040 ();
 sg13g2_fill_8 FILLER_115_1048 ();
 sg13g2_fill_8 FILLER_115_1056 ();
 sg13g2_fill_8 FILLER_115_1064 ();
 sg13g2_fill_8 FILLER_115_1072 ();
 sg13g2_fill_8 FILLER_115_1080 ();
 sg13g2_fill_8 FILLER_115_1088 ();
 sg13g2_fill_8 FILLER_115_1096 ();
 sg13g2_fill_8 FILLER_115_1104 ();
 sg13g2_fill_8 FILLER_115_1112 ();
 sg13g2_fill_8 FILLER_115_1120 ();
 sg13g2_fill_8 FILLER_115_1128 ();
 sg13g2_fill_8 FILLER_115_1136 ();
 sg13g2_fill_8 FILLER_115_1144 ();
 sg13g2_fill_8 FILLER_115_1152 ();
 sg13g2_fill_4 FILLER_115_1160 ();
 sg13g2_fill_2 FILLER_115_1164 ();
 sg13g2_fill_8 FILLER_116_0 ();
 sg13g2_fill_8 FILLER_116_8 ();
 sg13g2_fill_8 FILLER_116_16 ();
 sg13g2_fill_8 FILLER_116_24 ();
 sg13g2_fill_8 FILLER_116_32 ();
 sg13g2_fill_8 FILLER_116_40 ();
 sg13g2_fill_8 FILLER_116_48 ();
 sg13g2_fill_8 FILLER_116_56 ();
 sg13g2_fill_8 FILLER_116_64 ();
 sg13g2_fill_8 FILLER_116_72 ();
 sg13g2_fill_8 FILLER_116_80 ();
 sg13g2_fill_8 FILLER_116_88 ();
 sg13g2_fill_8 FILLER_116_96 ();
 sg13g2_fill_8 FILLER_116_104 ();
 sg13g2_fill_8 FILLER_116_112 ();
 sg13g2_fill_8 FILLER_116_120 ();
 sg13g2_fill_8 FILLER_116_128 ();
 sg13g2_fill_8 FILLER_116_136 ();
 sg13g2_fill_8 FILLER_116_144 ();
 sg13g2_fill_8 FILLER_116_152 ();
 sg13g2_fill_8 FILLER_116_160 ();
 sg13g2_fill_8 FILLER_116_168 ();
 sg13g2_fill_8 FILLER_116_176 ();
 sg13g2_fill_8 FILLER_116_184 ();
 sg13g2_fill_8 FILLER_116_192 ();
 sg13g2_fill_8 FILLER_116_200 ();
 sg13g2_fill_8 FILLER_116_208 ();
 sg13g2_fill_8 FILLER_116_216 ();
 sg13g2_fill_8 FILLER_116_224 ();
 sg13g2_fill_8 FILLER_116_232 ();
 sg13g2_fill_8 FILLER_116_240 ();
 sg13g2_fill_8 FILLER_116_248 ();
 sg13g2_fill_8 FILLER_116_256 ();
 sg13g2_fill_8 FILLER_116_264 ();
 sg13g2_fill_8 FILLER_116_272 ();
 sg13g2_fill_8 FILLER_116_280 ();
 sg13g2_fill_8 FILLER_116_288 ();
 sg13g2_fill_8 FILLER_116_296 ();
 sg13g2_fill_8 FILLER_116_304 ();
 sg13g2_fill_8 FILLER_116_312 ();
 sg13g2_fill_8 FILLER_116_320 ();
 sg13g2_fill_8 FILLER_116_328 ();
 sg13g2_fill_8 FILLER_116_336 ();
 sg13g2_fill_8 FILLER_116_344 ();
 sg13g2_fill_8 FILLER_116_352 ();
 sg13g2_fill_8 FILLER_116_360 ();
 sg13g2_fill_8 FILLER_116_368 ();
 sg13g2_fill_8 FILLER_116_376 ();
 sg13g2_fill_8 FILLER_116_384 ();
 sg13g2_fill_8 FILLER_116_392 ();
 sg13g2_fill_8 FILLER_116_400 ();
 sg13g2_fill_8 FILLER_116_408 ();
 sg13g2_fill_8 FILLER_116_416 ();
 sg13g2_fill_8 FILLER_116_424 ();
 sg13g2_fill_8 FILLER_116_432 ();
 sg13g2_fill_8 FILLER_116_440 ();
 sg13g2_fill_8 FILLER_116_448 ();
 sg13g2_fill_8 FILLER_116_456 ();
 sg13g2_fill_8 FILLER_116_464 ();
 sg13g2_fill_8 FILLER_116_472 ();
 sg13g2_fill_8 FILLER_116_480 ();
 sg13g2_fill_8 FILLER_116_488 ();
 sg13g2_fill_8 FILLER_116_496 ();
 sg13g2_fill_8 FILLER_116_504 ();
 sg13g2_fill_8 FILLER_116_512 ();
 sg13g2_fill_8 FILLER_116_520 ();
 sg13g2_fill_8 FILLER_116_528 ();
 sg13g2_fill_8 FILLER_116_536 ();
 sg13g2_fill_8 FILLER_116_544 ();
 sg13g2_fill_8 FILLER_116_552 ();
 sg13g2_fill_8 FILLER_116_560 ();
 sg13g2_fill_8 FILLER_116_568 ();
 sg13g2_fill_8 FILLER_116_576 ();
 sg13g2_fill_8 FILLER_116_584 ();
 sg13g2_fill_8 FILLER_116_592 ();
 sg13g2_fill_8 FILLER_116_600 ();
 sg13g2_fill_8 FILLER_116_608 ();
 sg13g2_fill_8 FILLER_116_616 ();
 sg13g2_fill_8 FILLER_116_624 ();
 sg13g2_fill_8 FILLER_116_632 ();
 sg13g2_fill_8 FILLER_116_640 ();
 sg13g2_fill_8 FILLER_116_648 ();
 sg13g2_fill_8 FILLER_116_656 ();
 sg13g2_fill_8 FILLER_116_664 ();
 sg13g2_fill_8 FILLER_116_672 ();
 sg13g2_fill_8 FILLER_116_680 ();
 sg13g2_fill_8 FILLER_116_688 ();
 sg13g2_fill_8 FILLER_116_696 ();
 sg13g2_fill_8 FILLER_116_704 ();
 sg13g2_fill_8 FILLER_116_712 ();
 sg13g2_fill_8 FILLER_116_720 ();
 sg13g2_fill_8 FILLER_116_728 ();
 sg13g2_fill_8 FILLER_116_736 ();
 sg13g2_fill_8 FILLER_116_744 ();
 sg13g2_fill_8 FILLER_116_752 ();
 sg13g2_fill_8 FILLER_116_760 ();
 sg13g2_fill_8 FILLER_116_768 ();
 sg13g2_fill_8 FILLER_116_776 ();
 sg13g2_fill_8 FILLER_116_784 ();
 sg13g2_fill_8 FILLER_116_792 ();
 sg13g2_fill_8 FILLER_116_800 ();
 sg13g2_fill_8 FILLER_116_808 ();
 sg13g2_fill_8 FILLER_116_816 ();
 sg13g2_fill_8 FILLER_116_824 ();
 sg13g2_fill_8 FILLER_116_832 ();
 sg13g2_fill_8 FILLER_116_840 ();
 sg13g2_fill_8 FILLER_116_848 ();
 sg13g2_fill_8 FILLER_116_856 ();
 sg13g2_fill_8 FILLER_116_864 ();
 sg13g2_fill_8 FILLER_116_872 ();
 sg13g2_fill_8 FILLER_116_880 ();
 sg13g2_fill_8 FILLER_116_888 ();
 sg13g2_fill_8 FILLER_116_896 ();
 sg13g2_fill_8 FILLER_116_904 ();
 sg13g2_fill_8 FILLER_116_912 ();
 sg13g2_fill_8 FILLER_116_920 ();
 sg13g2_fill_8 FILLER_116_928 ();
 sg13g2_fill_8 FILLER_116_936 ();
 sg13g2_fill_8 FILLER_116_944 ();
 sg13g2_fill_8 FILLER_116_952 ();
 sg13g2_fill_8 FILLER_116_960 ();
 sg13g2_fill_8 FILLER_116_968 ();
 sg13g2_fill_8 FILLER_116_976 ();
 sg13g2_fill_8 FILLER_116_984 ();
 sg13g2_fill_8 FILLER_116_992 ();
 sg13g2_fill_8 FILLER_116_1000 ();
 sg13g2_fill_8 FILLER_116_1008 ();
 sg13g2_fill_8 FILLER_116_1016 ();
 sg13g2_fill_8 FILLER_116_1024 ();
 sg13g2_fill_8 FILLER_116_1032 ();
 sg13g2_fill_8 FILLER_116_1040 ();
 sg13g2_fill_8 FILLER_116_1048 ();
 sg13g2_fill_8 FILLER_116_1056 ();
 sg13g2_fill_8 FILLER_116_1064 ();
 sg13g2_fill_8 FILLER_116_1072 ();
 sg13g2_fill_8 FILLER_116_1080 ();
 sg13g2_fill_8 FILLER_116_1088 ();
 sg13g2_fill_8 FILLER_116_1096 ();
 sg13g2_fill_8 FILLER_116_1104 ();
 sg13g2_fill_8 FILLER_116_1112 ();
 sg13g2_fill_8 FILLER_116_1120 ();
 sg13g2_fill_8 FILLER_116_1128 ();
 sg13g2_fill_8 FILLER_116_1136 ();
 sg13g2_fill_8 FILLER_116_1144 ();
 sg13g2_fill_8 FILLER_116_1152 ();
 sg13g2_fill_4 FILLER_116_1160 ();
 sg13g2_fill_2 FILLER_116_1164 ();
 sg13g2_fill_8 FILLER_117_0 ();
 sg13g2_fill_8 FILLER_117_8 ();
 sg13g2_fill_8 FILLER_117_16 ();
 sg13g2_fill_8 FILLER_117_24 ();
 sg13g2_fill_8 FILLER_117_32 ();
 sg13g2_fill_8 FILLER_117_40 ();
 sg13g2_fill_8 FILLER_117_48 ();
 sg13g2_fill_8 FILLER_117_56 ();
 sg13g2_fill_8 FILLER_117_64 ();
 sg13g2_fill_8 FILLER_117_72 ();
 sg13g2_fill_8 FILLER_117_80 ();
 sg13g2_fill_8 FILLER_117_88 ();
 sg13g2_fill_8 FILLER_117_96 ();
 sg13g2_fill_8 FILLER_117_104 ();
 sg13g2_fill_8 FILLER_117_112 ();
 sg13g2_fill_8 FILLER_117_120 ();
 sg13g2_fill_8 FILLER_117_128 ();
 sg13g2_fill_8 FILLER_117_136 ();
 sg13g2_fill_8 FILLER_117_144 ();
 sg13g2_fill_8 FILLER_117_152 ();
 sg13g2_fill_8 FILLER_117_160 ();
 sg13g2_fill_8 FILLER_117_168 ();
 sg13g2_fill_8 FILLER_117_176 ();
 sg13g2_fill_8 FILLER_117_184 ();
 sg13g2_fill_8 FILLER_117_192 ();
 sg13g2_fill_8 FILLER_117_200 ();
 sg13g2_fill_8 FILLER_117_208 ();
 sg13g2_fill_8 FILLER_117_216 ();
 sg13g2_fill_8 FILLER_117_224 ();
 sg13g2_fill_8 FILLER_117_232 ();
 sg13g2_fill_8 FILLER_117_240 ();
 sg13g2_fill_8 FILLER_117_248 ();
 sg13g2_fill_8 FILLER_117_256 ();
 sg13g2_fill_8 FILLER_117_264 ();
 sg13g2_fill_8 FILLER_117_272 ();
 sg13g2_fill_8 FILLER_117_280 ();
 sg13g2_fill_8 FILLER_117_288 ();
 sg13g2_fill_8 FILLER_117_296 ();
 sg13g2_fill_8 FILLER_117_304 ();
 sg13g2_fill_8 FILLER_117_312 ();
 sg13g2_fill_8 FILLER_117_320 ();
 sg13g2_fill_8 FILLER_117_328 ();
 sg13g2_fill_8 FILLER_117_336 ();
 sg13g2_fill_8 FILLER_117_344 ();
 sg13g2_fill_8 FILLER_117_352 ();
 sg13g2_fill_8 FILLER_117_360 ();
 sg13g2_fill_8 FILLER_117_368 ();
 sg13g2_fill_8 FILLER_117_376 ();
 sg13g2_fill_8 FILLER_117_384 ();
 sg13g2_fill_8 FILLER_117_392 ();
 sg13g2_fill_8 FILLER_117_400 ();
 sg13g2_fill_8 FILLER_117_408 ();
 sg13g2_fill_8 FILLER_117_416 ();
 sg13g2_fill_8 FILLER_117_424 ();
 sg13g2_fill_8 FILLER_117_432 ();
 sg13g2_fill_8 FILLER_117_440 ();
 sg13g2_fill_8 FILLER_117_448 ();
 sg13g2_fill_8 FILLER_117_456 ();
 sg13g2_fill_8 FILLER_117_464 ();
 sg13g2_fill_8 FILLER_117_472 ();
 sg13g2_fill_8 FILLER_117_480 ();
 sg13g2_fill_8 FILLER_117_488 ();
 sg13g2_fill_8 FILLER_117_496 ();
 sg13g2_fill_8 FILLER_117_504 ();
 sg13g2_fill_8 FILLER_117_512 ();
 sg13g2_fill_8 FILLER_117_520 ();
 sg13g2_fill_8 FILLER_117_528 ();
 sg13g2_fill_8 FILLER_117_536 ();
 sg13g2_fill_8 FILLER_117_544 ();
 sg13g2_fill_8 FILLER_117_552 ();
 sg13g2_fill_8 FILLER_117_560 ();
 sg13g2_fill_8 FILLER_117_568 ();
 sg13g2_fill_8 FILLER_117_576 ();
 sg13g2_fill_8 FILLER_117_584 ();
 sg13g2_fill_8 FILLER_117_592 ();
 sg13g2_fill_8 FILLER_117_600 ();
 sg13g2_fill_8 FILLER_117_608 ();
 sg13g2_fill_8 FILLER_117_616 ();
 sg13g2_fill_8 FILLER_117_624 ();
 sg13g2_fill_8 FILLER_117_632 ();
 sg13g2_fill_8 FILLER_117_640 ();
 sg13g2_fill_8 FILLER_117_648 ();
 sg13g2_fill_8 FILLER_117_656 ();
 sg13g2_fill_8 FILLER_117_664 ();
 sg13g2_fill_8 FILLER_117_672 ();
 sg13g2_fill_8 FILLER_117_680 ();
 sg13g2_fill_8 FILLER_117_688 ();
 sg13g2_fill_8 FILLER_117_696 ();
 sg13g2_fill_8 FILLER_117_704 ();
 sg13g2_fill_8 FILLER_117_712 ();
 sg13g2_fill_8 FILLER_117_720 ();
 sg13g2_fill_8 FILLER_117_728 ();
 sg13g2_fill_8 FILLER_117_736 ();
 sg13g2_fill_8 FILLER_117_744 ();
 sg13g2_fill_8 FILLER_117_752 ();
 sg13g2_fill_8 FILLER_117_760 ();
 sg13g2_fill_8 FILLER_117_768 ();
 sg13g2_fill_8 FILLER_117_776 ();
 sg13g2_fill_8 FILLER_117_784 ();
 sg13g2_fill_8 FILLER_117_792 ();
 sg13g2_fill_8 FILLER_117_800 ();
 sg13g2_fill_8 FILLER_117_808 ();
 sg13g2_fill_8 FILLER_117_816 ();
 sg13g2_fill_8 FILLER_117_824 ();
 sg13g2_fill_8 FILLER_117_832 ();
 sg13g2_fill_8 FILLER_117_840 ();
 sg13g2_fill_8 FILLER_117_848 ();
 sg13g2_fill_8 FILLER_117_856 ();
 sg13g2_fill_8 FILLER_117_864 ();
 sg13g2_fill_8 FILLER_117_872 ();
 sg13g2_fill_8 FILLER_117_880 ();
 sg13g2_fill_8 FILLER_117_888 ();
 sg13g2_fill_8 FILLER_117_896 ();
 sg13g2_fill_8 FILLER_117_904 ();
 sg13g2_fill_8 FILLER_117_912 ();
 sg13g2_fill_8 FILLER_117_920 ();
 sg13g2_fill_8 FILLER_117_928 ();
 sg13g2_fill_8 FILLER_117_936 ();
 sg13g2_fill_8 FILLER_117_944 ();
 sg13g2_fill_8 FILLER_117_952 ();
 sg13g2_fill_8 FILLER_117_960 ();
 sg13g2_fill_8 FILLER_117_968 ();
 sg13g2_fill_8 FILLER_117_976 ();
 sg13g2_fill_8 FILLER_117_984 ();
 sg13g2_fill_8 FILLER_117_992 ();
 sg13g2_fill_8 FILLER_117_1000 ();
 sg13g2_fill_8 FILLER_117_1008 ();
 sg13g2_fill_8 FILLER_117_1016 ();
 sg13g2_fill_8 FILLER_117_1024 ();
 sg13g2_fill_8 FILLER_117_1032 ();
 sg13g2_fill_8 FILLER_117_1040 ();
 sg13g2_fill_8 FILLER_117_1048 ();
 sg13g2_fill_8 FILLER_117_1056 ();
 sg13g2_fill_8 FILLER_117_1064 ();
 sg13g2_fill_8 FILLER_117_1072 ();
 sg13g2_fill_8 FILLER_117_1080 ();
 sg13g2_fill_8 FILLER_117_1088 ();
 sg13g2_fill_8 FILLER_117_1096 ();
 sg13g2_fill_8 FILLER_117_1104 ();
 sg13g2_fill_8 FILLER_117_1112 ();
 sg13g2_fill_8 FILLER_117_1120 ();
 sg13g2_fill_8 FILLER_117_1128 ();
 sg13g2_fill_8 FILLER_117_1136 ();
 sg13g2_fill_8 FILLER_117_1144 ();
 sg13g2_fill_8 FILLER_117_1152 ();
 sg13g2_fill_4 FILLER_117_1160 ();
 sg13g2_fill_2 FILLER_117_1164 ();
 sg13g2_fill_8 FILLER_118_0 ();
 sg13g2_fill_4 FILLER_118_8 ();
 sg13g2_fill_2 FILLER_118_12 ();
 sg13g2_fill_8 FILLER_118_22 ();
 sg13g2_fill_8 FILLER_118_30 ();
 sg13g2_fill_8 FILLER_118_38 ();
 sg13g2_fill_8 FILLER_118_46 ();
 sg13g2_fill_8 FILLER_118_54 ();
 sg13g2_fill_8 FILLER_118_62 ();
 sg13g2_fill_8 FILLER_118_70 ();
 sg13g2_fill_8 FILLER_118_78 ();
 sg13g2_fill_8 FILLER_118_86 ();
 sg13g2_fill_8 FILLER_118_94 ();
 sg13g2_fill_8 FILLER_118_102 ();
 sg13g2_fill_8 FILLER_118_110 ();
 sg13g2_fill_8 FILLER_118_118 ();
 sg13g2_fill_8 FILLER_118_126 ();
 sg13g2_fill_8 FILLER_118_134 ();
 sg13g2_fill_8 FILLER_118_142 ();
 sg13g2_fill_8 FILLER_118_150 ();
 sg13g2_fill_8 FILLER_118_158 ();
 sg13g2_fill_8 FILLER_118_166 ();
 sg13g2_fill_8 FILLER_118_174 ();
 sg13g2_fill_8 FILLER_118_182 ();
 sg13g2_fill_8 FILLER_118_190 ();
 sg13g2_fill_8 FILLER_118_198 ();
 sg13g2_fill_8 FILLER_118_206 ();
 sg13g2_fill_8 FILLER_118_214 ();
 sg13g2_fill_8 FILLER_118_222 ();
 sg13g2_fill_8 FILLER_118_230 ();
 sg13g2_fill_8 FILLER_118_238 ();
 sg13g2_fill_8 FILLER_118_246 ();
 sg13g2_fill_8 FILLER_118_254 ();
 sg13g2_fill_8 FILLER_118_262 ();
 sg13g2_fill_8 FILLER_118_270 ();
 sg13g2_fill_8 FILLER_118_278 ();
 sg13g2_fill_8 FILLER_118_286 ();
 sg13g2_fill_8 FILLER_118_294 ();
 sg13g2_fill_8 FILLER_118_302 ();
 sg13g2_fill_8 FILLER_118_310 ();
 sg13g2_fill_8 FILLER_118_318 ();
 sg13g2_fill_8 FILLER_118_326 ();
 sg13g2_fill_8 FILLER_118_334 ();
 sg13g2_fill_8 FILLER_118_342 ();
 sg13g2_fill_8 FILLER_118_350 ();
 sg13g2_fill_8 FILLER_118_358 ();
 sg13g2_fill_8 FILLER_118_366 ();
 sg13g2_fill_8 FILLER_118_374 ();
 sg13g2_fill_8 FILLER_118_382 ();
 sg13g2_fill_8 FILLER_118_390 ();
 sg13g2_fill_8 FILLER_118_398 ();
 sg13g2_fill_8 FILLER_118_406 ();
 sg13g2_fill_8 FILLER_118_414 ();
 sg13g2_fill_8 FILLER_118_422 ();
 sg13g2_fill_8 FILLER_118_430 ();
 sg13g2_fill_8 FILLER_118_438 ();
 sg13g2_fill_8 FILLER_118_446 ();
 sg13g2_fill_8 FILLER_118_454 ();
 sg13g2_fill_8 FILLER_118_462 ();
 sg13g2_fill_8 FILLER_118_470 ();
 sg13g2_fill_8 FILLER_118_478 ();
 sg13g2_fill_8 FILLER_118_486 ();
 sg13g2_fill_8 FILLER_118_494 ();
 sg13g2_fill_8 FILLER_118_502 ();
 sg13g2_fill_8 FILLER_118_510 ();
 sg13g2_fill_8 FILLER_118_518 ();
 sg13g2_fill_8 FILLER_118_526 ();
 sg13g2_fill_8 FILLER_118_534 ();
 sg13g2_fill_8 FILLER_118_542 ();
 sg13g2_fill_8 FILLER_118_550 ();
 sg13g2_fill_8 FILLER_118_558 ();
 sg13g2_fill_8 FILLER_118_566 ();
 sg13g2_fill_8 FILLER_118_574 ();
 sg13g2_fill_8 FILLER_118_582 ();
 sg13g2_fill_8 FILLER_118_590 ();
 sg13g2_fill_8 FILLER_118_598 ();
 sg13g2_fill_8 FILLER_118_606 ();
 sg13g2_fill_8 FILLER_118_614 ();
 sg13g2_fill_8 FILLER_118_622 ();
 sg13g2_fill_8 FILLER_118_630 ();
 sg13g2_fill_8 FILLER_118_638 ();
 sg13g2_fill_8 FILLER_118_646 ();
 sg13g2_fill_8 FILLER_118_654 ();
 sg13g2_fill_8 FILLER_118_662 ();
 sg13g2_fill_8 FILLER_118_670 ();
 sg13g2_fill_8 FILLER_118_678 ();
 sg13g2_fill_8 FILLER_118_686 ();
 sg13g2_fill_8 FILLER_118_694 ();
 sg13g2_fill_8 FILLER_118_702 ();
 sg13g2_fill_8 FILLER_118_710 ();
 sg13g2_fill_8 FILLER_118_718 ();
 sg13g2_fill_8 FILLER_118_726 ();
 sg13g2_fill_8 FILLER_118_734 ();
 sg13g2_fill_8 FILLER_118_742 ();
 sg13g2_fill_8 FILLER_118_750 ();
 sg13g2_fill_8 FILLER_118_758 ();
 sg13g2_fill_8 FILLER_118_766 ();
 sg13g2_fill_8 FILLER_118_774 ();
 sg13g2_fill_8 FILLER_118_782 ();
 sg13g2_fill_8 FILLER_118_790 ();
 sg13g2_fill_8 FILLER_118_798 ();
 sg13g2_fill_8 FILLER_118_806 ();
 sg13g2_fill_8 FILLER_118_814 ();
 sg13g2_fill_8 FILLER_118_822 ();
 sg13g2_fill_8 FILLER_118_830 ();
 sg13g2_fill_8 FILLER_118_838 ();
 sg13g2_fill_8 FILLER_118_846 ();
 sg13g2_fill_8 FILLER_118_854 ();
 sg13g2_fill_8 FILLER_118_862 ();
 sg13g2_fill_8 FILLER_118_870 ();
 sg13g2_fill_8 FILLER_118_878 ();
 sg13g2_fill_8 FILLER_118_886 ();
 sg13g2_fill_8 FILLER_118_894 ();
 sg13g2_fill_8 FILLER_118_902 ();
 sg13g2_fill_8 FILLER_118_910 ();
 sg13g2_fill_8 FILLER_118_918 ();
 sg13g2_fill_8 FILLER_118_926 ();
 sg13g2_fill_8 FILLER_118_934 ();
 sg13g2_fill_8 FILLER_118_942 ();
 sg13g2_fill_8 FILLER_118_950 ();
 sg13g2_fill_8 FILLER_118_958 ();
 sg13g2_fill_8 FILLER_118_966 ();
 sg13g2_fill_8 FILLER_118_974 ();
 sg13g2_fill_8 FILLER_118_982 ();
 sg13g2_fill_8 FILLER_118_990 ();
 sg13g2_fill_8 FILLER_118_998 ();
 sg13g2_fill_8 FILLER_118_1006 ();
 sg13g2_fill_8 FILLER_118_1014 ();
 sg13g2_fill_8 FILLER_118_1022 ();
 sg13g2_fill_8 FILLER_118_1030 ();
 sg13g2_fill_8 FILLER_118_1038 ();
 sg13g2_fill_8 FILLER_118_1046 ();
 sg13g2_fill_8 FILLER_118_1054 ();
 sg13g2_fill_8 FILLER_118_1062 ();
 sg13g2_fill_8 FILLER_118_1070 ();
 sg13g2_fill_8 FILLER_118_1078 ();
 sg13g2_fill_8 FILLER_118_1086 ();
 sg13g2_fill_8 FILLER_118_1094 ();
 sg13g2_fill_8 FILLER_118_1102 ();
 sg13g2_fill_8 FILLER_118_1110 ();
 sg13g2_fill_8 FILLER_118_1118 ();
 sg13g2_fill_8 FILLER_118_1126 ();
 sg13g2_fill_8 FILLER_118_1134 ();
 sg13g2_fill_8 FILLER_118_1142 ();
 sg13g2_fill_8 FILLER_118_1150 ();
 sg13g2_fill_8 FILLER_118_1158 ();
 sg13g2_fill_8 FILLER_119_0 ();
 sg13g2_fill_8 FILLER_119_8 ();
 sg13g2_fill_8 FILLER_119_16 ();
 sg13g2_fill_8 FILLER_119_24 ();
 sg13g2_fill_8 FILLER_119_32 ();
 sg13g2_fill_8 FILLER_119_40 ();
 sg13g2_fill_8 FILLER_119_48 ();
 sg13g2_fill_8 FILLER_119_56 ();
 sg13g2_fill_8 FILLER_119_64 ();
 sg13g2_fill_8 FILLER_119_72 ();
 sg13g2_fill_8 FILLER_119_80 ();
 sg13g2_fill_8 FILLER_119_88 ();
 sg13g2_fill_8 FILLER_119_96 ();
 sg13g2_fill_8 FILLER_119_104 ();
 sg13g2_fill_8 FILLER_119_112 ();
 sg13g2_fill_8 FILLER_119_120 ();
 sg13g2_fill_8 FILLER_119_128 ();
 sg13g2_fill_8 FILLER_119_136 ();
 sg13g2_fill_8 FILLER_119_144 ();
 sg13g2_fill_8 FILLER_119_152 ();
 sg13g2_fill_8 FILLER_119_160 ();
 sg13g2_fill_8 FILLER_119_168 ();
 sg13g2_fill_8 FILLER_119_176 ();
 sg13g2_fill_8 FILLER_119_184 ();
 sg13g2_fill_8 FILLER_119_192 ();
 sg13g2_fill_8 FILLER_119_200 ();
 sg13g2_fill_8 FILLER_119_208 ();
 sg13g2_fill_8 FILLER_119_216 ();
 sg13g2_fill_8 FILLER_119_224 ();
 sg13g2_fill_8 FILLER_119_232 ();
 sg13g2_fill_8 FILLER_119_240 ();
 sg13g2_fill_8 FILLER_119_248 ();
 sg13g2_fill_8 FILLER_119_256 ();
 sg13g2_fill_8 FILLER_119_264 ();
 sg13g2_fill_8 FILLER_119_272 ();
 sg13g2_fill_8 FILLER_119_280 ();
 sg13g2_fill_8 FILLER_119_288 ();
 sg13g2_fill_8 FILLER_119_296 ();
 sg13g2_fill_8 FILLER_119_304 ();
 sg13g2_fill_8 FILLER_119_312 ();
 sg13g2_fill_8 FILLER_119_320 ();
 sg13g2_fill_8 FILLER_119_328 ();
 sg13g2_fill_8 FILLER_119_336 ();
 sg13g2_fill_8 FILLER_119_344 ();
 sg13g2_fill_8 FILLER_119_352 ();
 sg13g2_fill_8 FILLER_119_360 ();
 sg13g2_fill_8 FILLER_119_368 ();
 sg13g2_fill_8 FILLER_119_376 ();
 sg13g2_fill_8 FILLER_119_384 ();
 sg13g2_fill_8 FILLER_119_392 ();
 sg13g2_fill_8 FILLER_119_400 ();
 sg13g2_fill_8 FILLER_119_408 ();
 sg13g2_fill_8 FILLER_119_416 ();
 sg13g2_fill_8 FILLER_119_424 ();
 sg13g2_fill_8 FILLER_119_432 ();
 sg13g2_fill_8 FILLER_119_440 ();
 sg13g2_fill_8 FILLER_119_448 ();
 sg13g2_fill_8 FILLER_119_456 ();
 sg13g2_fill_8 FILLER_119_464 ();
 sg13g2_fill_8 FILLER_119_472 ();
 sg13g2_fill_8 FILLER_119_480 ();
 sg13g2_fill_8 FILLER_119_488 ();
 sg13g2_fill_8 FILLER_119_496 ();
 sg13g2_fill_8 FILLER_119_504 ();
 sg13g2_fill_8 FILLER_119_512 ();
 sg13g2_fill_8 FILLER_119_520 ();
 sg13g2_fill_8 FILLER_119_528 ();
 sg13g2_fill_8 FILLER_119_536 ();
 sg13g2_fill_8 FILLER_119_544 ();
 sg13g2_fill_8 FILLER_119_552 ();
 sg13g2_fill_8 FILLER_119_560 ();
 sg13g2_fill_8 FILLER_119_568 ();
 sg13g2_fill_8 FILLER_119_576 ();
 sg13g2_fill_8 FILLER_119_584 ();
 sg13g2_fill_8 FILLER_119_592 ();
 sg13g2_fill_8 FILLER_119_600 ();
 sg13g2_fill_8 FILLER_119_608 ();
 sg13g2_fill_8 FILLER_119_616 ();
 sg13g2_fill_8 FILLER_119_624 ();
 sg13g2_fill_8 FILLER_119_632 ();
 sg13g2_fill_8 FILLER_119_640 ();
 sg13g2_fill_8 FILLER_119_648 ();
 sg13g2_fill_8 FILLER_119_656 ();
 sg13g2_fill_8 FILLER_119_664 ();
 sg13g2_fill_8 FILLER_119_672 ();
 sg13g2_fill_8 FILLER_119_680 ();
 sg13g2_fill_8 FILLER_119_688 ();
 sg13g2_fill_8 FILLER_119_696 ();
 sg13g2_fill_8 FILLER_119_704 ();
 sg13g2_fill_8 FILLER_119_712 ();
 sg13g2_fill_8 FILLER_119_720 ();
 sg13g2_fill_8 FILLER_119_728 ();
 sg13g2_fill_8 FILLER_119_736 ();
 sg13g2_fill_8 FILLER_119_744 ();
 sg13g2_fill_8 FILLER_119_752 ();
 sg13g2_fill_8 FILLER_119_760 ();
 sg13g2_fill_8 FILLER_119_768 ();
 sg13g2_fill_8 FILLER_119_776 ();
 sg13g2_fill_8 FILLER_119_784 ();
 sg13g2_fill_8 FILLER_119_792 ();
 sg13g2_fill_8 FILLER_119_800 ();
 sg13g2_fill_8 FILLER_119_808 ();
 sg13g2_fill_8 FILLER_119_816 ();
 sg13g2_fill_8 FILLER_119_824 ();
 sg13g2_fill_8 FILLER_119_832 ();
 sg13g2_fill_8 FILLER_119_840 ();
 sg13g2_fill_8 FILLER_119_848 ();
 sg13g2_fill_8 FILLER_119_856 ();
 sg13g2_fill_8 FILLER_119_864 ();
 sg13g2_fill_8 FILLER_119_872 ();
 sg13g2_fill_8 FILLER_119_880 ();
 sg13g2_fill_8 FILLER_119_888 ();
 sg13g2_fill_8 FILLER_119_896 ();
 sg13g2_fill_8 FILLER_119_904 ();
 sg13g2_fill_8 FILLER_119_912 ();
 sg13g2_fill_8 FILLER_119_920 ();
 sg13g2_fill_8 FILLER_119_928 ();
 sg13g2_fill_8 FILLER_119_936 ();
 sg13g2_fill_8 FILLER_119_944 ();
 sg13g2_fill_8 FILLER_119_952 ();
 sg13g2_fill_8 FILLER_119_960 ();
 sg13g2_fill_8 FILLER_119_968 ();
 sg13g2_fill_8 FILLER_119_976 ();
 sg13g2_fill_8 FILLER_119_984 ();
 sg13g2_fill_8 FILLER_119_992 ();
 sg13g2_fill_8 FILLER_119_1000 ();
 sg13g2_fill_8 FILLER_119_1008 ();
 sg13g2_fill_8 FILLER_119_1016 ();
 sg13g2_fill_8 FILLER_119_1024 ();
 sg13g2_fill_8 FILLER_119_1032 ();
 sg13g2_fill_8 FILLER_119_1040 ();
 sg13g2_fill_8 FILLER_119_1048 ();
 sg13g2_fill_8 FILLER_119_1056 ();
 sg13g2_fill_8 FILLER_119_1064 ();
 sg13g2_fill_8 FILLER_119_1072 ();
 sg13g2_fill_8 FILLER_119_1080 ();
 sg13g2_fill_8 FILLER_119_1088 ();
 sg13g2_fill_8 FILLER_119_1096 ();
 sg13g2_fill_8 FILLER_119_1104 ();
 sg13g2_fill_8 FILLER_119_1112 ();
 sg13g2_fill_8 FILLER_119_1120 ();
 sg13g2_fill_8 FILLER_119_1128 ();
 sg13g2_fill_8 FILLER_119_1136 ();
 sg13g2_fill_8 FILLER_119_1144 ();
 sg13g2_fill_8 FILLER_119_1152 ();
 sg13g2_fill_4 FILLER_119_1160 ();
 sg13g2_fill_2 FILLER_119_1164 ();
 sg13g2_fill_8 FILLER_120_0 ();
 sg13g2_fill_8 FILLER_120_8 ();
 sg13g2_fill_8 FILLER_120_16 ();
 sg13g2_fill_8 FILLER_120_24 ();
 sg13g2_fill_8 FILLER_120_32 ();
 sg13g2_fill_8 FILLER_120_40 ();
 sg13g2_fill_8 FILLER_120_48 ();
 sg13g2_fill_8 FILLER_120_56 ();
 sg13g2_fill_8 FILLER_120_64 ();
 sg13g2_fill_8 FILLER_120_72 ();
 sg13g2_fill_8 FILLER_120_80 ();
 sg13g2_fill_8 FILLER_120_88 ();
 sg13g2_fill_8 FILLER_120_96 ();
 sg13g2_fill_8 FILLER_120_104 ();
 sg13g2_fill_8 FILLER_120_112 ();
 sg13g2_fill_8 FILLER_120_120 ();
 sg13g2_fill_8 FILLER_120_128 ();
 sg13g2_fill_8 FILLER_120_136 ();
 sg13g2_fill_8 FILLER_120_144 ();
 sg13g2_fill_8 FILLER_120_152 ();
 sg13g2_fill_8 FILLER_120_160 ();
 sg13g2_fill_8 FILLER_120_168 ();
 sg13g2_fill_8 FILLER_120_176 ();
 sg13g2_fill_8 FILLER_120_184 ();
 sg13g2_fill_8 FILLER_120_192 ();
 sg13g2_fill_8 FILLER_120_200 ();
 sg13g2_fill_8 FILLER_120_208 ();
 sg13g2_fill_8 FILLER_120_216 ();
 sg13g2_fill_8 FILLER_120_224 ();
 sg13g2_fill_8 FILLER_120_232 ();
 sg13g2_fill_8 FILLER_120_240 ();
 sg13g2_fill_8 FILLER_120_248 ();
 sg13g2_fill_8 FILLER_120_256 ();
 sg13g2_fill_8 FILLER_120_264 ();
 sg13g2_fill_8 FILLER_120_272 ();
 sg13g2_fill_8 FILLER_120_280 ();
 sg13g2_fill_8 FILLER_120_288 ();
 sg13g2_fill_8 FILLER_120_296 ();
 sg13g2_fill_8 FILLER_120_304 ();
 sg13g2_fill_8 FILLER_120_312 ();
 sg13g2_fill_8 FILLER_120_320 ();
 sg13g2_fill_8 FILLER_120_328 ();
 sg13g2_fill_8 FILLER_120_336 ();
 sg13g2_fill_8 FILLER_120_344 ();
 sg13g2_fill_8 FILLER_120_352 ();
 sg13g2_fill_8 FILLER_120_360 ();
 sg13g2_fill_8 FILLER_120_368 ();
 sg13g2_fill_8 FILLER_120_376 ();
 sg13g2_fill_8 FILLER_120_384 ();
 sg13g2_fill_8 FILLER_120_392 ();
 sg13g2_fill_8 FILLER_120_400 ();
 sg13g2_fill_8 FILLER_120_408 ();
 sg13g2_fill_8 FILLER_120_416 ();
 sg13g2_fill_8 FILLER_120_424 ();
 sg13g2_fill_8 FILLER_120_432 ();
 sg13g2_fill_8 FILLER_120_440 ();
 sg13g2_fill_8 FILLER_120_448 ();
 sg13g2_fill_8 FILLER_120_456 ();
 sg13g2_fill_8 FILLER_120_464 ();
 sg13g2_fill_8 FILLER_120_472 ();
 sg13g2_fill_8 FILLER_120_480 ();
 sg13g2_fill_8 FILLER_120_488 ();
 sg13g2_fill_8 FILLER_120_496 ();
 sg13g2_fill_8 FILLER_120_504 ();
 sg13g2_fill_8 FILLER_120_512 ();
 sg13g2_fill_8 FILLER_120_520 ();
 sg13g2_fill_8 FILLER_120_528 ();
 sg13g2_fill_8 FILLER_120_536 ();
 sg13g2_fill_8 FILLER_120_544 ();
 sg13g2_fill_8 FILLER_120_552 ();
 sg13g2_fill_8 FILLER_120_560 ();
 sg13g2_fill_8 FILLER_120_568 ();
 sg13g2_fill_8 FILLER_120_576 ();
 sg13g2_fill_8 FILLER_120_584 ();
 sg13g2_fill_8 FILLER_120_592 ();
 sg13g2_fill_8 FILLER_120_600 ();
 sg13g2_fill_8 FILLER_120_608 ();
 sg13g2_fill_8 FILLER_120_616 ();
 sg13g2_fill_8 FILLER_120_624 ();
 sg13g2_fill_8 FILLER_120_632 ();
 sg13g2_fill_8 FILLER_120_640 ();
 sg13g2_fill_8 FILLER_120_648 ();
 sg13g2_fill_8 FILLER_120_656 ();
 sg13g2_fill_8 FILLER_120_664 ();
 sg13g2_fill_8 FILLER_120_672 ();
 sg13g2_fill_8 FILLER_120_680 ();
 sg13g2_fill_8 FILLER_120_688 ();
 sg13g2_fill_8 FILLER_120_696 ();
 sg13g2_fill_8 FILLER_120_704 ();
 sg13g2_fill_8 FILLER_120_712 ();
 sg13g2_fill_8 FILLER_120_720 ();
 sg13g2_fill_8 FILLER_120_728 ();
 sg13g2_fill_8 FILLER_120_736 ();
 sg13g2_fill_8 FILLER_120_744 ();
 sg13g2_fill_8 FILLER_120_752 ();
 sg13g2_fill_8 FILLER_120_760 ();
 sg13g2_fill_8 FILLER_120_768 ();
 sg13g2_fill_8 FILLER_120_776 ();
 sg13g2_fill_8 FILLER_120_784 ();
 sg13g2_fill_8 FILLER_120_792 ();
 sg13g2_fill_8 FILLER_120_800 ();
 sg13g2_fill_8 FILLER_120_808 ();
 sg13g2_fill_8 FILLER_120_816 ();
 sg13g2_fill_8 FILLER_120_824 ();
 sg13g2_fill_8 FILLER_120_832 ();
 sg13g2_fill_8 FILLER_120_840 ();
 sg13g2_fill_8 FILLER_120_848 ();
 sg13g2_fill_8 FILLER_120_856 ();
 sg13g2_fill_8 FILLER_120_864 ();
 sg13g2_fill_8 FILLER_120_872 ();
 sg13g2_fill_8 FILLER_120_880 ();
 sg13g2_fill_8 FILLER_120_888 ();
 sg13g2_fill_8 FILLER_120_896 ();
 sg13g2_fill_8 FILLER_120_904 ();
 sg13g2_fill_8 FILLER_120_912 ();
 sg13g2_fill_8 FILLER_120_920 ();
 sg13g2_fill_8 FILLER_120_928 ();
 sg13g2_fill_8 FILLER_120_936 ();
 sg13g2_fill_8 FILLER_120_944 ();
 sg13g2_fill_8 FILLER_120_952 ();
 sg13g2_fill_8 FILLER_120_960 ();
 sg13g2_fill_8 FILLER_120_968 ();
 sg13g2_fill_8 FILLER_120_976 ();
 sg13g2_fill_8 FILLER_120_984 ();
 sg13g2_fill_8 FILLER_120_992 ();
 sg13g2_fill_8 FILLER_120_1000 ();
 sg13g2_fill_8 FILLER_120_1008 ();
 sg13g2_fill_8 FILLER_120_1016 ();
 sg13g2_fill_8 FILLER_120_1024 ();
 sg13g2_fill_8 FILLER_120_1032 ();
 sg13g2_fill_8 FILLER_120_1040 ();
 sg13g2_fill_8 FILLER_120_1048 ();
 sg13g2_fill_8 FILLER_120_1056 ();
 sg13g2_fill_8 FILLER_120_1064 ();
 sg13g2_fill_8 FILLER_120_1072 ();
 sg13g2_fill_8 FILLER_120_1080 ();
 sg13g2_fill_8 FILLER_120_1088 ();
 sg13g2_fill_8 FILLER_120_1096 ();
 sg13g2_fill_8 FILLER_120_1104 ();
 sg13g2_fill_8 FILLER_120_1112 ();
 sg13g2_fill_8 FILLER_120_1120 ();
 sg13g2_fill_8 FILLER_120_1128 ();
 sg13g2_fill_8 FILLER_120_1136 ();
 sg13g2_fill_8 FILLER_120_1144 ();
 sg13g2_fill_8 FILLER_120_1152 ();
 sg13g2_fill_4 FILLER_120_1160 ();
 sg13g2_fill_2 FILLER_120_1164 ();
 sg13g2_fill_8 FILLER_121_0 ();
 sg13g2_fill_8 FILLER_121_8 ();
 sg13g2_fill_8 FILLER_121_16 ();
 sg13g2_fill_8 FILLER_121_24 ();
 sg13g2_fill_8 FILLER_121_32 ();
 sg13g2_fill_8 FILLER_121_40 ();
 sg13g2_fill_8 FILLER_121_48 ();
 sg13g2_fill_8 FILLER_121_56 ();
 sg13g2_fill_8 FILLER_121_64 ();
 sg13g2_fill_8 FILLER_121_72 ();
 sg13g2_fill_8 FILLER_121_80 ();
 sg13g2_fill_8 FILLER_121_88 ();
 sg13g2_fill_8 FILLER_121_96 ();
 sg13g2_fill_8 FILLER_121_104 ();
 sg13g2_fill_8 FILLER_121_112 ();
 sg13g2_fill_8 FILLER_121_120 ();
 sg13g2_fill_8 FILLER_121_128 ();
 sg13g2_fill_8 FILLER_121_136 ();
 sg13g2_fill_8 FILLER_121_144 ();
 sg13g2_fill_8 FILLER_121_152 ();
 sg13g2_fill_8 FILLER_121_160 ();
 sg13g2_fill_8 FILLER_121_168 ();
 sg13g2_fill_8 FILLER_121_176 ();
 sg13g2_fill_8 FILLER_121_184 ();
 sg13g2_fill_8 FILLER_121_192 ();
 sg13g2_fill_8 FILLER_121_200 ();
 sg13g2_fill_8 FILLER_121_208 ();
 sg13g2_fill_8 FILLER_121_216 ();
 sg13g2_fill_8 FILLER_121_224 ();
 sg13g2_fill_8 FILLER_121_232 ();
 sg13g2_fill_8 FILLER_121_240 ();
 sg13g2_fill_8 FILLER_121_248 ();
 sg13g2_fill_8 FILLER_121_256 ();
 sg13g2_fill_8 FILLER_121_264 ();
 sg13g2_fill_8 FILLER_121_272 ();
 sg13g2_fill_8 FILLER_121_280 ();
 sg13g2_fill_8 FILLER_121_288 ();
 sg13g2_fill_8 FILLER_121_296 ();
 sg13g2_fill_8 FILLER_121_304 ();
 sg13g2_fill_8 FILLER_121_312 ();
 sg13g2_fill_8 FILLER_121_320 ();
 sg13g2_fill_8 FILLER_121_328 ();
 sg13g2_fill_8 FILLER_121_336 ();
 sg13g2_fill_8 FILLER_121_344 ();
 sg13g2_fill_8 FILLER_121_352 ();
 sg13g2_fill_8 FILLER_121_360 ();
 sg13g2_fill_8 FILLER_121_368 ();
 sg13g2_fill_8 FILLER_121_376 ();
 sg13g2_fill_8 FILLER_121_384 ();
 sg13g2_fill_8 FILLER_121_392 ();
 sg13g2_fill_8 FILLER_121_400 ();
 sg13g2_fill_8 FILLER_121_408 ();
 sg13g2_fill_8 FILLER_121_416 ();
 sg13g2_fill_8 FILLER_121_424 ();
 sg13g2_fill_8 FILLER_121_432 ();
 sg13g2_fill_8 FILLER_121_440 ();
 sg13g2_fill_8 FILLER_121_448 ();
 sg13g2_fill_8 FILLER_121_456 ();
 sg13g2_fill_8 FILLER_121_464 ();
 sg13g2_fill_8 FILLER_121_472 ();
 sg13g2_fill_8 FILLER_121_480 ();
 sg13g2_fill_8 FILLER_121_488 ();
 sg13g2_fill_8 FILLER_121_496 ();
 sg13g2_fill_8 FILLER_121_504 ();
 sg13g2_fill_8 FILLER_121_512 ();
 sg13g2_fill_8 FILLER_121_520 ();
 sg13g2_fill_8 FILLER_121_528 ();
 sg13g2_fill_8 FILLER_121_536 ();
 sg13g2_fill_8 FILLER_121_544 ();
 sg13g2_fill_8 FILLER_121_552 ();
 sg13g2_fill_8 FILLER_121_560 ();
 sg13g2_fill_8 FILLER_121_568 ();
 sg13g2_fill_8 FILLER_121_576 ();
 sg13g2_fill_8 FILLER_121_584 ();
 sg13g2_fill_8 FILLER_121_592 ();
 sg13g2_fill_8 FILLER_121_600 ();
 sg13g2_fill_8 FILLER_121_608 ();
 sg13g2_fill_8 FILLER_121_616 ();
 sg13g2_fill_8 FILLER_121_624 ();
 sg13g2_fill_8 FILLER_121_632 ();
 sg13g2_fill_8 FILLER_121_640 ();
 sg13g2_fill_8 FILLER_121_648 ();
 sg13g2_fill_8 FILLER_121_656 ();
 sg13g2_fill_8 FILLER_121_664 ();
 sg13g2_fill_8 FILLER_121_672 ();
 sg13g2_fill_8 FILLER_121_680 ();
 sg13g2_fill_8 FILLER_121_688 ();
 sg13g2_fill_8 FILLER_121_696 ();
 sg13g2_fill_8 FILLER_121_704 ();
 sg13g2_fill_8 FILLER_121_712 ();
 sg13g2_fill_8 FILLER_121_720 ();
 sg13g2_fill_8 FILLER_121_728 ();
 sg13g2_fill_8 FILLER_121_736 ();
 sg13g2_fill_8 FILLER_121_744 ();
 sg13g2_fill_8 FILLER_121_752 ();
 sg13g2_fill_8 FILLER_121_760 ();
 sg13g2_fill_8 FILLER_121_768 ();
 sg13g2_fill_8 FILLER_121_776 ();
 sg13g2_fill_8 FILLER_121_784 ();
 sg13g2_fill_8 FILLER_121_792 ();
 sg13g2_fill_8 FILLER_121_800 ();
 sg13g2_fill_8 FILLER_121_808 ();
 sg13g2_fill_8 FILLER_121_816 ();
 sg13g2_fill_8 FILLER_121_824 ();
 sg13g2_fill_8 FILLER_121_832 ();
 sg13g2_fill_8 FILLER_121_840 ();
 sg13g2_fill_8 FILLER_121_848 ();
 sg13g2_fill_8 FILLER_121_856 ();
 sg13g2_fill_8 FILLER_121_864 ();
 sg13g2_fill_8 FILLER_121_872 ();
 sg13g2_fill_8 FILLER_121_880 ();
 sg13g2_fill_8 FILLER_121_888 ();
 sg13g2_fill_8 FILLER_121_896 ();
 sg13g2_fill_8 FILLER_121_904 ();
 sg13g2_fill_8 FILLER_121_912 ();
 sg13g2_fill_8 FILLER_121_920 ();
 sg13g2_fill_8 FILLER_121_928 ();
 sg13g2_fill_8 FILLER_121_936 ();
 sg13g2_fill_8 FILLER_121_944 ();
 sg13g2_fill_8 FILLER_121_952 ();
 sg13g2_fill_8 FILLER_121_960 ();
 sg13g2_fill_8 FILLER_121_968 ();
 sg13g2_fill_8 FILLER_121_976 ();
 sg13g2_fill_8 FILLER_121_984 ();
 sg13g2_fill_8 FILLER_121_992 ();
 sg13g2_fill_8 FILLER_121_1000 ();
 sg13g2_fill_8 FILLER_121_1008 ();
 sg13g2_fill_8 FILLER_121_1016 ();
 sg13g2_fill_8 FILLER_121_1024 ();
 sg13g2_fill_8 FILLER_121_1032 ();
 sg13g2_fill_8 FILLER_121_1040 ();
 sg13g2_fill_8 FILLER_121_1048 ();
 sg13g2_fill_8 FILLER_121_1056 ();
 sg13g2_fill_8 FILLER_121_1064 ();
 sg13g2_fill_8 FILLER_121_1072 ();
 sg13g2_fill_8 FILLER_121_1080 ();
 sg13g2_fill_8 FILLER_121_1088 ();
 sg13g2_fill_8 FILLER_121_1096 ();
 sg13g2_fill_8 FILLER_121_1104 ();
 sg13g2_fill_8 FILLER_121_1112 ();
 sg13g2_fill_8 FILLER_121_1120 ();
 sg13g2_fill_8 FILLER_121_1128 ();
 sg13g2_fill_8 FILLER_121_1136 ();
 sg13g2_fill_8 FILLER_121_1144 ();
 sg13g2_fill_8 FILLER_121_1152 ();
 sg13g2_fill_4 FILLER_121_1160 ();
 sg13g2_fill_2 FILLER_121_1164 ();
 sg13g2_fill_8 FILLER_122_0 ();
 sg13g2_fill_8 FILLER_122_8 ();
 sg13g2_fill_8 FILLER_122_16 ();
 sg13g2_fill_8 FILLER_122_24 ();
 sg13g2_fill_8 FILLER_122_32 ();
 sg13g2_fill_8 FILLER_122_40 ();
 sg13g2_fill_8 FILLER_122_48 ();
 sg13g2_fill_8 FILLER_122_56 ();
 sg13g2_fill_8 FILLER_122_64 ();
 sg13g2_fill_8 FILLER_122_72 ();
 sg13g2_fill_8 FILLER_122_80 ();
 sg13g2_fill_8 FILLER_122_88 ();
 sg13g2_fill_8 FILLER_122_96 ();
 sg13g2_fill_8 FILLER_122_104 ();
 sg13g2_fill_8 FILLER_122_112 ();
 sg13g2_fill_8 FILLER_122_120 ();
 sg13g2_fill_8 FILLER_122_128 ();
 sg13g2_fill_8 FILLER_122_136 ();
 sg13g2_fill_8 FILLER_122_144 ();
 sg13g2_fill_8 FILLER_122_152 ();
 sg13g2_fill_8 FILLER_122_160 ();
 sg13g2_fill_8 FILLER_122_168 ();
 sg13g2_fill_8 FILLER_122_176 ();
 sg13g2_fill_8 FILLER_122_184 ();
 sg13g2_fill_8 FILLER_122_192 ();
 sg13g2_fill_8 FILLER_122_200 ();
 sg13g2_fill_8 FILLER_122_208 ();
 sg13g2_fill_8 FILLER_122_216 ();
 sg13g2_fill_8 FILLER_122_224 ();
 sg13g2_fill_8 FILLER_122_232 ();
 sg13g2_fill_8 FILLER_122_240 ();
 sg13g2_fill_8 FILLER_122_248 ();
 sg13g2_fill_8 FILLER_122_256 ();
 sg13g2_fill_8 FILLER_122_264 ();
 sg13g2_fill_8 FILLER_122_272 ();
 sg13g2_fill_8 FILLER_122_280 ();
 sg13g2_fill_8 FILLER_122_288 ();
 sg13g2_fill_8 FILLER_122_296 ();
 sg13g2_fill_8 FILLER_122_304 ();
 sg13g2_fill_8 FILLER_122_312 ();
 sg13g2_fill_8 FILLER_122_320 ();
 sg13g2_fill_8 FILLER_122_328 ();
 sg13g2_fill_8 FILLER_122_336 ();
 sg13g2_fill_8 FILLER_122_344 ();
 sg13g2_fill_8 FILLER_122_352 ();
 sg13g2_fill_8 FILLER_122_360 ();
 sg13g2_fill_8 FILLER_122_368 ();
 sg13g2_fill_8 FILLER_122_376 ();
 sg13g2_fill_8 FILLER_122_384 ();
 sg13g2_fill_8 FILLER_122_392 ();
 sg13g2_fill_8 FILLER_122_400 ();
 sg13g2_fill_8 FILLER_122_408 ();
 sg13g2_fill_8 FILLER_122_416 ();
 sg13g2_fill_8 FILLER_122_424 ();
 sg13g2_fill_8 FILLER_122_432 ();
 sg13g2_fill_8 FILLER_122_440 ();
 sg13g2_fill_8 FILLER_122_448 ();
 sg13g2_fill_8 FILLER_122_456 ();
 sg13g2_fill_8 FILLER_122_464 ();
 sg13g2_fill_8 FILLER_122_472 ();
 sg13g2_fill_8 FILLER_122_480 ();
 sg13g2_fill_8 FILLER_122_488 ();
 sg13g2_fill_8 FILLER_122_496 ();
 sg13g2_fill_8 FILLER_122_504 ();
 sg13g2_fill_8 FILLER_122_512 ();
 sg13g2_fill_8 FILLER_122_520 ();
 sg13g2_fill_8 FILLER_122_528 ();
 sg13g2_fill_8 FILLER_122_536 ();
 sg13g2_fill_8 FILLER_122_544 ();
 sg13g2_fill_8 FILLER_122_552 ();
 sg13g2_fill_8 FILLER_122_560 ();
 sg13g2_fill_8 FILLER_122_568 ();
 sg13g2_fill_8 FILLER_122_576 ();
 sg13g2_fill_8 FILLER_122_584 ();
 sg13g2_fill_8 FILLER_122_592 ();
 sg13g2_fill_8 FILLER_122_600 ();
 sg13g2_fill_8 FILLER_122_608 ();
 sg13g2_fill_8 FILLER_122_616 ();
 sg13g2_fill_8 FILLER_122_624 ();
 sg13g2_fill_8 FILLER_122_632 ();
 sg13g2_fill_8 FILLER_122_640 ();
 sg13g2_fill_8 FILLER_122_648 ();
 sg13g2_fill_8 FILLER_122_656 ();
 sg13g2_fill_8 FILLER_122_664 ();
 sg13g2_fill_8 FILLER_122_672 ();
 sg13g2_fill_8 FILLER_122_680 ();
 sg13g2_fill_8 FILLER_122_688 ();
 sg13g2_fill_8 FILLER_122_696 ();
 sg13g2_fill_8 FILLER_122_704 ();
 sg13g2_fill_8 FILLER_122_712 ();
 sg13g2_fill_8 FILLER_122_720 ();
 sg13g2_fill_8 FILLER_122_728 ();
 sg13g2_fill_8 FILLER_122_736 ();
 sg13g2_fill_8 FILLER_122_744 ();
 sg13g2_fill_8 FILLER_122_752 ();
 sg13g2_fill_8 FILLER_122_760 ();
 sg13g2_fill_8 FILLER_122_768 ();
 sg13g2_fill_8 FILLER_122_776 ();
 sg13g2_fill_8 FILLER_122_784 ();
 sg13g2_fill_8 FILLER_122_792 ();
 sg13g2_fill_8 FILLER_122_800 ();
 sg13g2_fill_8 FILLER_122_808 ();
 sg13g2_fill_8 FILLER_122_816 ();
 sg13g2_fill_8 FILLER_122_824 ();
 sg13g2_fill_8 FILLER_122_832 ();
 sg13g2_fill_8 FILLER_122_840 ();
 sg13g2_fill_8 FILLER_122_848 ();
 sg13g2_fill_8 FILLER_122_856 ();
 sg13g2_fill_8 FILLER_122_864 ();
 sg13g2_fill_8 FILLER_122_872 ();
 sg13g2_fill_8 FILLER_122_880 ();
 sg13g2_fill_8 FILLER_122_888 ();
 sg13g2_fill_8 FILLER_122_896 ();
 sg13g2_fill_8 FILLER_122_904 ();
 sg13g2_fill_8 FILLER_122_912 ();
 sg13g2_fill_8 FILLER_122_920 ();
 sg13g2_fill_8 FILLER_122_928 ();
 sg13g2_fill_8 FILLER_122_936 ();
 sg13g2_fill_8 FILLER_122_944 ();
 sg13g2_fill_8 FILLER_122_952 ();
 sg13g2_fill_8 FILLER_122_960 ();
 sg13g2_fill_8 FILLER_122_968 ();
 sg13g2_fill_8 FILLER_122_976 ();
 sg13g2_fill_8 FILLER_122_984 ();
 sg13g2_fill_8 FILLER_122_992 ();
 sg13g2_fill_8 FILLER_122_1000 ();
 sg13g2_fill_8 FILLER_122_1008 ();
 sg13g2_fill_8 FILLER_122_1016 ();
 sg13g2_fill_8 FILLER_122_1024 ();
 sg13g2_fill_8 FILLER_122_1032 ();
 sg13g2_fill_8 FILLER_122_1040 ();
 sg13g2_fill_8 FILLER_122_1048 ();
 sg13g2_fill_8 FILLER_122_1056 ();
 sg13g2_fill_8 FILLER_122_1064 ();
 sg13g2_fill_8 FILLER_122_1072 ();
 sg13g2_fill_8 FILLER_122_1080 ();
 sg13g2_fill_8 FILLER_122_1088 ();
 sg13g2_fill_8 FILLER_122_1096 ();
 sg13g2_fill_8 FILLER_122_1104 ();
 sg13g2_fill_8 FILLER_122_1112 ();
 sg13g2_fill_8 FILLER_122_1120 ();
 sg13g2_fill_8 FILLER_122_1128 ();
 sg13g2_fill_8 FILLER_122_1136 ();
 sg13g2_fill_8 FILLER_122_1144 ();
 sg13g2_fill_8 FILLER_122_1152 ();
 sg13g2_fill_4 FILLER_122_1160 ();
 sg13g2_fill_2 FILLER_122_1164 ();
 sg13g2_fill_8 FILLER_123_0 ();
 sg13g2_fill_8 FILLER_123_8 ();
 sg13g2_fill_8 FILLER_123_16 ();
 sg13g2_fill_8 FILLER_123_24 ();
 sg13g2_fill_8 FILLER_123_32 ();
 sg13g2_fill_8 FILLER_123_40 ();
 sg13g2_fill_8 FILLER_123_48 ();
 sg13g2_fill_8 FILLER_123_56 ();
 sg13g2_fill_8 FILLER_123_64 ();
 sg13g2_fill_8 FILLER_123_72 ();
 sg13g2_fill_8 FILLER_123_80 ();
 sg13g2_fill_8 FILLER_123_88 ();
 sg13g2_fill_8 FILLER_123_96 ();
 sg13g2_fill_8 FILLER_123_104 ();
 sg13g2_fill_8 FILLER_123_112 ();
 sg13g2_fill_8 FILLER_123_120 ();
 sg13g2_fill_8 FILLER_123_128 ();
 sg13g2_fill_8 FILLER_123_136 ();
 sg13g2_fill_8 FILLER_123_144 ();
 sg13g2_fill_8 FILLER_123_152 ();
 sg13g2_fill_8 FILLER_123_160 ();
 sg13g2_fill_8 FILLER_123_168 ();
 sg13g2_fill_8 FILLER_123_176 ();
 sg13g2_fill_8 FILLER_123_184 ();
 sg13g2_fill_8 FILLER_123_192 ();
 sg13g2_fill_8 FILLER_123_200 ();
 sg13g2_fill_8 FILLER_123_208 ();
 sg13g2_fill_8 FILLER_123_216 ();
 sg13g2_fill_8 FILLER_123_224 ();
 sg13g2_fill_8 FILLER_123_232 ();
 sg13g2_fill_8 FILLER_123_240 ();
 sg13g2_fill_8 FILLER_123_248 ();
 sg13g2_fill_8 FILLER_123_256 ();
 sg13g2_fill_8 FILLER_123_264 ();
 sg13g2_fill_8 FILLER_123_272 ();
 sg13g2_fill_8 FILLER_123_280 ();
 sg13g2_fill_8 FILLER_123_288 ();
 sg13g2_fill_8 FILLER_123_296 ();
 sg13g2_fill_8 FILLER_123_304 ();
 sg13g2_fill_8 FILLER_123_312 ();
 sg13g2_fill_8 FILLER_123_320 ();
 sg13g2_fill_8 FILLER_123_328 ();
 sg13g2_fill_8 FILLER_123_336 ();
 sg13g2_fill_8 FILLER_123_344 ();
 sg13g2_fill_8 FILLER_123_352 ();
 sg13g2_fill_8 FILLER_123_360 ();
 sg13g2_fill_8 FILLER_123_368 ();
 sg13g2_fill_8 FILLER_123_376 ();
 sg13g2_fill_8 FILLER_123_384 ();
 sg13g2_fill_8 FILLER_123_392 ();
 sg13g2_fill_8 FILLER_123_400 ();
 sg13g2_fill_8 FILLER_123_408 ();
 sg13g2_fill_8 FILLER_123_416 ();
 sg13g2_fill_8 FILLER_123_424 ();
 sg13g2_fill_8 FILLER_123_432 ();
 sg13g2_fill_8 FILLER_123_440 ();
 sg13g2_fill_8 FILLER_123_448 ();
 sg13g2_fill_8 FILLER_123_456 ();
 sg13g2_fill_8 FILLER_123_464 ();
 sg13g2_fill_8 FILLER_123_472 ();
 sg13g2_fill_8 FILLER_123_480 ();
 sg13g2_fill_8 FILLER_123_488 ();
 sg13g2_fill_8 FILLER_123_496 ();
 sg13g2_fill_8 FILLER_123_504 ();
 sg13g2_fill_8 FILLER_123_512 ();
 sg13g2_fill_8 FILLER_123_520 ();
 sg13g2_fill_8 FILLER_123_528 ();
 sg13g2_fill_8 FILLER_123_536 ();
 sg13g2_fill_8 FILLER_123_544 ();
 sg13g2_fill_8 FILLER_123_552 ();
 sg13g2_fill_8 FILLER_123_560 ();
 sg13g2_fill_8 FILLER_123_568 ();
 sg13g2_fill_8 FILLER_123_576 ();
 sg13g2_fill_8 FILLER_123_584 ();
 sg13g2_fill_8 FILLER_123_592 ();
 sg13g2_fill_8 FILLER_123_600 ();
 sg13g2_fill_8 FILLER_123_608 ();
 sg13g2_fill_8 FILLER_123_616 ();
 sg13g2_fill_8 FILLER_123_624 ();
 sg13g2_fill_8 FILLER_123_632 ();
 sg13g2_fill_8 FILLER_123_640 ();
 sg13g2_fill_8 FILLER_123_648 ();
 sg13g2_fill_8 FILLER_123_656 ();
 sg13g2_fill_8 FILLER_123_664 ();
 sg13g2_fill_8 FILLER_123_672 ();
 sg13g2_fill_8 FILLER_123_680 ();
 sg13g2_fill_8 FILLER_123_688 ();
 sg13g2_fill_8 FILLER_123_696 ();
 sg13g2_fill_8 FILLER_123_704 ();
 sg13g2_fill_8 FILLER_123_712 ();
 sg13g2_fill_8 FILLER_123_720 ();
 sg13g2_fill_8 FILLER_123_728 ();
 sg13g2_fill_8 FILLER_123_736 ();
 sg13g2_fill_8 FILLER_123_744 ();
 sg13g2_fill_8 FILLER_123_752 ();
 sg13g2_fill_8 FILLER_123_760 ();
 sg13g2_fill_8 FILLER_123_768 ();
 sg13g2_fill_8 FILLER_123_776 ();
 sg13g2_fill_8 FILLER_123_784 ();
 sg13g2_fill_8 FILLER_123_792 ();
 sg13g2_fill_8 FILLER_123_800 ();
 sg13g2_fill_8 FILLER_123_808 ();
 sg13g2_fill_8 FILLER_123_816 ();
 sg13g2_fill_8 FILLER_123_824 ();
 sg13g2_fill_8 FILLER_123_832 ();
 sg13g2_fill_8 FILLER_123_840 ();
 sg13g2_fill_8 FILLER_123_848 ();
 sg13g2_fill_8 FILLER_123_856 ();
 sg13g2_fill_8 FILLER_123_864 ();
 sg13g2_fill_8 FILLER_123_872 ();
 sg13g2_fill_8 FILLER_123_880 ();
 sg13g2_fill_8 FILLER_123_888 ();
 sg13g2_fill_8 FILLER_123_896 ();
 sg13g2_fill_8 FILLER_123_904 ();
 sg13g2_fill_8 FILLER_123_912 ();
 sg13g2_fill_8 FILLER_123_920 ();
 sg13g2_fill_8 FILLER_123_928 ();
 sg13g2_fill_8 FILLER_123_936 ();
 sg13g2_fill_8 FILLER_123_944 ();
 sg13g2_fill_8 FILLER_123_952 ();
 sg13g2_fill_8 FILLER_123_960 ();
 sg13g2_fill_8 FILLER_123_968 ();
 sg13g2_fill_8 FILLER_123_976 ();
 sg13g2_fill_8 FILLER_123_984 ();
 sg13g2_fill_8 FILLER_123_992 ();
 sg13g2_fill_8 FILLER_123_1000 ();
 sg13g2_fill_8 FILLER_123_1008 ();
 sg13g2_fill_8 FILLER_123_1016 ();
 sg13g2_fill_8 FILLER_123_1024 ();
 sg13g2_fill_8 FILLER_123_1032 ();
 sg13g2_fill_8 FILLER_123_1040 ();
 sg13g2_fill_8 FILLER_123_1048 ();
 sg13g2_fill_8 FILLER_123_1056 ();
 sg13g2_fill_8 FILLER_123_1064 ();
 sg13g2_fill_8 FILLER_123_1072 ();
 sg13g2_fill_8 FILLER_123_1080 ();
 sg13g2_fill_8 FILLER_123_1088 ();
 sg13g2_fill_8 FILLER_123_1096 ();
 sg13g2_fill_8 FILLER_123_1104 ();
 sg13g2_fill_8 FILLER_123_1112 ();
 sg13g2_fill_8 FILLER_123_1120 ();
 sg13g2_fill_8 FILLER_123_1128 ();
 sg13g2_fill_8 FILLER_123_1136 ();
 sg13g2_fill_8 FILLER_123_1144 ();
 sg13g2_fill_8 FILLER_123_1152 ();
 sg13g2_fill_4 FILLER_123_1160 ();
 sg13g2_fill_2 FILLER_123_1164 ();
 sg13g2_fill_8 FILLER_124_0 ();
 sg13g2_fill_8 FILLER_124_8 ();
 sg13g2_fill_8 FILLER_124_16 ();
 sg13g2_fill_8 FILLER_124_24 ();
 sg13g2_fill_8 FILLER_124_32 ();
 sg13g2_fill_8 FILLER_124_40 ();
 sg13g2_fill_8 FILLER_124_48 ();
 sg13g2_fill_8 FILLER_124_56 ();
 sg13g2_fill_8 FILLER_124_64 ();
 sg13g2_fill_8 FILLER_124_72 ();
 sg13g2_fill_8 FILLER_124_80 ();
 sg13g2_fill_8 FILLER_124_88 ();
 sg13g2_fill_8 FILLER_124_96 ();
 sg13g2_fill_8 FILLER_124_104 ();
 sg13g2_fill_8 FILLER_124_112 ();
 sg13g2_fill_8 FILLER_124_120 ();
 sg13g2_fill_8 FILLER_124_128 ();
 sg13g2_fill_8 FILLER_124_136 ();
 sg13g2_fill_8 FILLER_124_144 ();
 sg13g2_fill_8 FILLER_124_152 ();
 sg13g2_fill_8 FILLER_124_160 ();
 sg13g2_fill_8 FILLER_124_168 ();
 sg13g2_fill_8 FILLER_124_176 ();
 sg13g2_fill_8 FILLER_124_184 ();
 sg13g2_fill_8 FILLER_124_192 ();
 sg13g2_fill_8 FILLER_124_200 ();
 sg13g2_fill_8 FILLER_124_208 ();
 sg13g2_fill_8 FILLER_124_216 ();
 sg13g2_fill_8 FILLER_124_224 ();
 sg13g2_fill_8 FILLER_124_232 ();
 sg13g2_fill_8 FILLER_124_240 ();
 sg13g2_fill_8 FILLER_124_248 ();
 sg13g2_fill_8 FILLER_124_256 ();
 sg13g2_fill_8 FILLER_124_264 ();
 sg13g2_fill_8 FILLER_124_272 ();
 sg13g2_fill_8 FILLER_124_280 ();
 sg13g2_fill_8 FILLER_124_288 ();
 sg13g2_fill_8 FILLER_124_296 ();
 sg13g2_fill_8 FILLER_124_304 ();
 sg13g2_fill_8 FILLER_124_312 ();
 sg13g2_fill_8 FILLER_124_320 ();
 sg13g2_fill_8 FILLER_124_328 ();
 sg13g2_fill_8 FILLER_124_336 ();
 sg13g2_fill_8 FILLER_124_344 ();
 sg13g2_fill_8 FILLER_124_352 ();
 sg13g2_fill_8 FILLER_124_360 ();
 sg13g2_fill_8 FILLER_124_368 ();
 sg13g2_fill_8 FILLER_124_376 ();
 sg13g2_fill_8 FILLER_124_384 ();
 sg13g2_fill_8 FILLER_124_392 ();
 sg13g2_fill_8 FILLER_124_400 ();
 sg13g2_fill_8 FILLER_124_408 ();
 sg13g2_fill_8 FILLER_124_416 ();
 sg13g2_fill_8 FILLER_124_424 ();
 sg13g2_fill_8 FILLER_124_432 ();
 sg13g2_fill_8 FILLER_124_440 ();
 sg13g2_fill_8 FILLER_124_448 ();
 sg13g2_fill_8 FILLER_124_456 ();
 sg13g2_fill_8 FILLER_124_464 ();
 sg13g2_fill_8 FILLER_124_472 ();
 sg13g2_fill_8 FILLER_124_480 ();
 sg13g2_fill_8 FILLER_124_488 ();
 sg13g2_fill_8 FILLER_124_496 ();
 sg13g2_fill_8 FILLER_124_504 ();
 sg13g2_fill_8 FILLER_124_512 ();
 sg13g2_fill_8 FILLER_124_520 ();
 sg13g2_fill_8 FILLER_124_528 ();
 sg13g2_fill_8 FILLER_124_536 ();
 sg13g2_fill_8 FILLER_124_544 ();
 sg13g2_fill_8 FILLER_124_552 ();
 sg13g2_fill_8 FILLER_124_560 ();
 sg13g2_fill_8 FILLER_124_568 ();
 sg13g2_fill_8 FILLER_124_576 ();
 sg13g2_fill_8 FILLER_124_584 ();
 sg13g2_fill_8 FILLER_124_592 ();
 sg13g2_fill_8 FILLER_124_600 ();
 sg13g2_fill_8 FILLER_124_608 ();
 sg13g2_fill_8 FILLER_124_616 ();
 sg13g2_fill_8 FILLER_124_624 ();
 sg13g2_fill_8 FILLER_124_632 ();
 sg13g2_fill_8 FILLER_124_640 ();
 sg13g2_fill_8 FILLER_124_648 ();
 sg13g2_fill_8 FILLER_124_656 ();
 sg13g2_fill_8 FILLER_124_664 ();
 sg13g2_fill_8 FILLER_124_672 ();
 sg13g2_fill_8 FILLER_124_680 ();
 sg13g2_fill_8 FILLER_124_688 ();
 sg13g2_fill_8 FILLER_124_696 ();
 sg13g2_fill_8 FILLER_124_704 ();
 sg13g2_fill_8 FILLER_124_712 ();
 sg13g2_fill_8 FILLER_124_720 ();
 sg13g2_fill_8 FILLER_124_728 ();
 sg13g2_fill_8 FILLER_124_736 ();
 sg13g2_fill_8 FILLER_124_744 ();
 sg13g2_fill_8 FILLER_124_752 ();
 sg13g2_fill_8 FILLER_124_760 ();
 sg13g2_fill_8 FILLER_124_768 ();
 sg13g2_fill_8 FILLER_124_776 ();
 sg13g2_fill_8 FILLER_124_784 ();
 sg13g2_fill_8 FILLER_124_792 ();
 sg13g2_fill_8 FILLER_124_800 ();
 sg13g2_fill_8 FILLER_124_808 ();
 sg13g2_fill_8 FILLER_124_816 ();
 sg13g2_fill_8 FILLER_124_824 ();
 sg13g2_fill_8 FILLER_124_832 ();
 sg13g2_fill_8 FILLER_124_840 ();
 sg13g2_fill_8 FILLER_124_848 ();
 sg13g2_fill_8 FILLER_124_856 ();
 sg13g2_fill_8 FILLER_124_864 ();
 sg13g2_fill_8 FILLER_124_872 ();
 sg13g2_fill_8 FILLER_124_880 ();
 sg13g2_fill_8 FILLER_124_888 ();
 sg13g2_fill_8 FILLER_124_896 ();
 sg13g2_fill_8 FILLER_124_904 ();
 sg13g2_fill_8 FILLER_124_912 ();
 sg13g2_fill_8 FILLER_124_920 ();
 sg13g2_fill_8 FILLER_124_928 ();
 sg13g2_fill_8 FILLER_124_936 ();
 sg13g2_fill_8 FILLER_124_944 ();
 sg13g2_fill_8 FILLER_124_952 ();
 sg13g2_fill_8 FILLER_124_960 ();
 sg13g2_fill_8 FILLER_124_968 ();
 sg13g2_fill_8 FILLER_124_976 ();
 sg13g2_fill_8 FILLER_124_984 ();
 sg13g2_fill_8 FILLER_124_992 ();
 sg13g2_fill_8 FILLER_124_1000 ();
 sg13g2_fill_8 FILLER_124_1008 ();
 sg13g2_fill_8 FILLER_124_1016 ();
 sg13g2_fill_8 FILLER_124_1024 ();
 sg13g2_fill_8 FILLER_124_1032 ();
 sg13g2_fill_8 FILLER_124_1040 ();
 sg13g2_fill_8 FILLER_124_1048 ();
 sg13g2_fill_8 FILLER_124_1056 ();
 sg13g2_fill_8 FILLER_124_1064 ();
 sg13g2_fill_8 FILLER_124_1072 ();
 sg13g2_fill_8 FILLER_124_1080 ();
 sg13g2_fill_8 FILLER_124_1088 ();
 sg13g2_fill_8 FILLER_124_1096 ();
 sg13g2_fill_8 FILLER_124_1104 ();
 sg13g2_fill_8 FILLER_124_1112 ();
 sg13g2_fill_8 FILLER_124_1120 ();
 sg13g2_fill_8 FILLER_124_1128 ();
 sg13g2_fill_8 FILLER_124_1136 ();
 sg13g2_fill_8 FILLER_124_1144 ();
 sg13g2_fill_8 FILLER_124_1152 ();
 sg13g2_fill_4 FILLER_124_1160 ();
 sg13g2_fill_2 FILLER_124_1164 ();
 sg13g2_fill_8 FILLER_125_0 ();
 sg13g2_fill_8 FILLER_125_8 ();
 sg13g2_fill_8 FILLER_125_16 ();
 sg13g2_fill_8 FILLER_125_24 ();
 sg13g2_fill_8 FILLER_125_32 ();
 sg13g2_fill_8 FILLER_125_40 ();
 sg13g2_fill_8 FILLER_125_48 ();
 sg13g2_fill_8 FILLER_125_56 ();
 sg13g2_fill_8 FILLER_125_64 ();
 sg13g2_fill_8 FILLER_125_72 ();
 sg13g2_fill_8 FILLER_125_80 ();
 sg13g2_fill_8 FILLER_125_88 ();
 sg13g2_fill_8 FILLER_125_96 ();
 sg13g2_fill_8 FILLER_125_104 ();
 sg13g2_fill_8 FILLER_125_112 ();
 sg13g2_fill_8 FILLER_125_120 ();
 sg13g2_fill_8 FILLER_125_128 ();
 sg13g2_fill_8 FILLER_125_136 ();
 sg13g2_fill_8 FILLER_125_144 ();
 sg13g2_fill_8 FILLER_125_152 ();
 sg13g2_fill_8 FILLER_125_160 ();
 sg13g2_fill_8 FILLER_125_168 ();
 sg13g2_fill_8 FILLER_125_176 ();
 sg13g2_fill_8 FILLER_125_184 ();
 sg13g2_fill_8 FILLER_125_192 ();
 sg13g2_fill_8 FILLER_125_200 ();
 sg13g2_fill_8 FILLER_125_208 ();
 sg13g2_fill_8 FILLER_125_216 ();
 sg13g2_fill_8 FILLER_125_224 ();
 sg13g2_fill_8 FILLER_125_232 ();
 sg13g2_fill_8 FILLER_125_240 ();
 sg13g2_fill_8 FILLER_125_248 ();
 sg13g2_fill_8 FILLER_125_256 ();
 sg13g2_fill_8 FILLER_125_264 ();
 sg13g2_fill_8 FILLER_125_272 ();
 sg13g2_fill_8 FILLER_125_280 ();
 sg13g2_fill_8 FILLER_125_288 ();
 sg13g2_fill_8 FILLER_125_296 ();
 sg13g2_fill_8 FILLER_125_304 ();
 sg13g2_fill_8 FILLER_125_312 ();
 sg13g2_fill_8 FILLER_125_320 ();
 sg13g2_fill_8 FILLER_125_328 ();
 sg13g2_fill_8 FILLER_125_336 ();
 sg13g2_fill_8 FILLER_125_344 ();
 sg13g2_fill_8 FILLER_125_352 ();
 sg13g2_fill_8 FILLER_125_360 ();
 sg13g2_fill_8 FILLER_125_368 ();
 sg13g2_fill_8 FILLER_125_376 ();
 sg13g2_fill_8 FILLER_125_384 ();
 sg13g2_fill_8 FILLER_125_392 ();
 sg13g2_fill_8 FILLER_125_400 ();
 sg13g2_fill_8 FILLER_125_408 ();
 sg13g2_fill_8 FILLER_125_416 ();
 sg13g2_fill_8 FILLER_125_424 ();
 sg13g2_fill_8 FILLER_125_432 ();
 sg13g2_fill_8 FILLER_125_440 ();
 sg13g2_fill_8 FILLER_125_448 ();
 sg13g2_fill_8 FILLER_125_456 ();
 sg13g2_fill_8 FILLER_125_464 ();
 sg13g2_fill_8 FILLER_125_472 ();
 sg13g2_fill_8 FILLER_125_480 ();
 sg13g2_fill_8 FILLER_125_488 ();
 sg13g2_fill_8 FILLER_125_496 ();
 sg13g2_fill_8 FILLER_125_504 ();
 sg13g2_fill_8 FILLER_125_512 ();
 sg13g2_fill_8 FILLER_125_520 ();
 sg13g2_fill_8 FILLER_125_528 ();
 sg13g2_fill_8 FILLER_125_536 ();
 sg13g2_fill_8 FILLER_125_544 ();
 sg13g2_fill_8 FILLER_125_552 ();
 sg13g2_fill_8 FILLER_125_560 ();
 sg13g2_fill_8 FILLER_125_568 ();
 sg13g2_fill_8 FILLER_125_576 ();
 sg13g2_fill_8 FILLER_125_584 ();
 sg13g2_fill_8 FILLER_125_592 ();
 sg13g2_fill_8 FILLER_125_600 ();
 sg13g2_fill_8 FILLER_125_608 ();
 sg13g2_fill_8 FILLER_125_616 ();
 sg13g2_fill_8 FILLER_125_624 ();
 sg13g2_fill_8 FILLER_125_632 ();
 sg13g2_fill_8 FILLER_125_640 ();
 sg13g2_fill_8 FILLER_125_648 ();
 sg13g2_fill_8 FILLER_125_656 ();
 sg13g2_fill_8 FILLER_125_664 ();
 sg13g2_fill_8 FILLER_125_672 ();
 sg13g2_fill_8 FILLER_125_680 ();
 sg13g2_fill_8 FILLER_125_688 ();
 sg13g2_fill_8 FILLER_125_696 ();
 sg13g2_fill_8 FILLER_125_704 ();
 sg13g2_fill_8 FILLER_125_712 ();
 sg13g2_fill_8 FILLER_125_720 ();
 sg13g2_fill_8 FILLER_125_728 ();
 sg13g2_fill_8 FILLER_125_736 ();
 sg13g2_fill_8 FILLER_125_744 ();
 sg13g2_fill_8 FILLER_125_752 ();
 sg13g2_fill_8 FILLER_125_760 ();
 sg13g2_fill_8 FILLER_125_768 ();
 sg13g2_fill_8 FILLER_125_776 ();
 sg13g2_fill_8 FILLER_125_784 ();
 sg13g2_fill_8 FILLER_125_792 ();
 sg13g2_fill_8 FILLER_125_800 ();
 sg13g2_fill_8 FILLER_125_808 ();
 sg13g2_fill_8 FILLER_125_816 ();
 sg13g2_fill_8 FILLER_125_824 ();
 sg13g2_fill_8 FILLER_125_832 ();
 sg13g2_fill_8 FILLER_125_840 ();
 sg13g2_fill_8 FILLER_125_848 ();
 sg13g2_fill_8 FILLER_125_856 ();
 sg13g2_fill_8 FILLER_125_864 ();
 sg13g2_fill_8 FILLER_125_872 ();
 sg13g2_fill_8 FILLER_125_880 ();
 sg13g2_fill_8 FILLER_125_888 ();
 sg13g2_fill_8 FILLER_125_896 ();
 sg13g2_fill_8 FILLER_125_904 ();
 sg13g2_fill_8 FILLER_125_912 ();
 sg13g2_fill_8 FILLER_125_920 ();
 sg13g2_fill_8 FILLER_125_928 ();
 sg13g2_fill_8 FILLER_125_936 ();
 sg13g2_fill_8 FILLER_125_944 ();
 sg13g2_fill_8 FILLER_125_952 ();
 sg13g2_fill_8 FILLER_125_960 ();
 sg13g2_fill_8 FILLER_125_968 ();
 sg13g2_fill_8 FILLER_125_976 ();
 sg13g2_fill_8 FILLER_125_984 ();
 sg13g2_fill_8 FILLER_125_992 ();
 sg13g2_fill_8 FILLER_125_1000 ();
 sg13g2_fill_8 FILLER_125_1008 ();
 sg13g2_fill_8 FILLER_125_1016 ();
 sg13g2_fill_8 FILLER_125_1024 ();
 sg13g2_fill_8 FILLER_125_1032 ();
 sg13g2_fill_8 FILLER_125_1040 ();
 sg13g2_fill_8 FILLER_125_1048 ();
 sg13g2_fill_8 FILLER_125_1056 ();
 sg13g2_fill_8 FILLER_125_1064 ();
 sg13g2_fill_8 FILLER_125_1072 ();
 sg13g2_fill_8 FILLER_125_1080 ();
 sg13g2_fill_8 FILLER_125_1088 ();
 sg13g2_fill_8 FILLER_125_1096 ();
 sg13g2_fill_8 FILLER_125_1104 ();
 sg13g2_fill_8 FILLER_125_1112 ();
 sg13g2_fill_8 FILLER_125_1120 ();
 sg13g2_fill_8 FILLER_125_1128 ();
 sg13g2_fill_8 FILLER_125_1136 ();
 sg13g2_fill_8 FILLER_125_1144 ();
 sg13g2_fill_8 FILLER_125_1152 ();
 sg13g2_fill_4 FILLER_125_1160 ();
 sg13g2_fill_2 FILLER_125_1164 ();
 sg13g2_fill_8 FILLER_126_0 ();
 sg13g2_fill_8 FILLER_126_8 ();
 sg13g2_fill_8 FILLER_126_16 ();
 sg13g2_fill_8 FILLER_126_24 ();
 sg13g2_fill_8 FILLER_126_32 ();
 sg13g2_fill_8 FILLER_126_40 ();
 sg13g2_fill_8 FILLER_126_48 ();
 sg13g2_fill_8 FILLER_126_56 ();
 sg13g2_fill_8 FILLER_126_64 ();
 sg13g2_fill_8 FILLER_126_72 ();
 sg13g2_fill_8 FILLER_126_80 ();
 sg13g2_fill_8 FILLER_126_88 ();
 sg13g2_fill_8 FILLER_126_96 ();
 sg13g2_fill_8 FILLER_126_104 ();
 sg13g2_fill_8 FILLER_126_112 ();
 sg13g2_fill_8 FILLER_126_120 ();
 sg13g2_fill_8 FILLER_126_128 ();
 sg13g2_fill_8 FILLER_126_136 ();
 sg13g2_fill_8 FILLER_126_144 ();
 sg13g2_fill_8 FILLER_126_152 ();
 sg13g2_fill_8 FILLER_126_160 ();
 sg13g2_fill_8 FILLER_126_168 ();
 sg13g2_fill_8 FILLER_126_176 ();
 sg13g2_fill_8 FILLER_126_184 ();
 sg13g2_fill_8 FILLER_126_192 ();
 sg13g2_fill_8 FILLER_126_200 ();
 sg13g2_fill_8 FILLER_126_208 ();
 sg13g2_fill_8 FILLER_126_216 ();
 sg13g2_fill_8 FILLER_126_224 ();
 sg13g2_fill_8 FILLER_126_232 ();
 sg13g2_fill_8 FILLER_126_240 ();
 sg13g2_fill_8 FILLER_126_248 ();
 sg13g2_fill_8 FILLER_126_256 ();
 sg13g2_fill_8 FILLER_126_264 ();
 sg13g2_fill_8 FILLER_126_272 ();
 sg13g2_fill_8 FILLER_126_280 ();
 sg13g2_fill_8 FILLER_126_288 ();
 sg13g2_fill_8 FILLER_126_296 ();
 sg13g2_fill_8 FILLER_126_304 ();
 sg13g2_fill_8 FILLER_126_312 ();
 sg13g2_fill_8 FILLER_126_320 ();
 sg13g2_fill_8 FILLER_126_328 ();
 sg13g2_fill_8 FILLER_126_336 ();
 sg13g2_fill_8 FILLER_126_344 ();
 sg13g2_fill_8 FILLER_126_352 ();
 sg13g2_fill_8 FILLER_126_360 ();
 sg13g2_fill_8 FILLER_126_368 ();
 sg13g2_fill_8 FILLER_126_376 ();
 sg13g2_fill_8 FILLER_126_384 ();
 sg13g2_fill_8 FILLER_126_392 ();
 sg13g2_fill_8 FILLER_126_400 ();
 sg13g2_fill_8 FILLER_126_408 ();
 sg13g2_fill_8 FILLER_126_416 ();
 sg13g2_fill_8 FILLER_126_424 ();
 sg13g2_fill_8 FILLER_126_432 ();
 sg13g2_fill_8 FILLER_126_440 ();
 sg13g2_fill_8 FILLER_126_448 ();
 sg13g2_fill_8 FILLER_126_456 ();
 sg13g2_fill_8 FILLER_126_464 ();
 sg13g2_fill_8 FILLER_126_472 ();
 sg13g2_fill_8 FILLER_126_480 ();
 sg13g2_fill_8 FILLER_126_488 ();
 sg13g2_fill_8 FILLER_126_496 ();
 sg13g2_fill_8 FILLER_126_504 ();
 sg13g2_fill_8 FILLER_126_512 ();
 sg13g2_fill_8 FILLER_126_520 ();
 sg13g2_fill_8 FILLER_126_528 ();
 sg13g2_fill_8 FILLER_126_536 ();
 sg13g2_fill_8 FILLER_126_544 ();
 sg13g2_fill_8 FILLER_126_552 ();
 sg13g2_fill_8 FILLER_126_560 ();
 sg13g2_fill_8 FILLER_126_568 ();
 sg13g2_fill_8 FILLER_126_576 ();
 sg13g2_fill_8 FILLER_126_584 ();
 sg13g2_fill_8 FILLER_126_592 ();
 sg13g2_fill_8 FILLER_126_600 ();
 sg13g2_fill_8 FILLER_126_608 ();
 sg13g2_fill_8 FILLER_126_616 ();
 sg13g2_fill_8 FILLER_126_624 ();
 sg13g2_fill_8 FILLER_126_632 ();
 sg13g2_fill_8 FILLER_126_640 ();
 sg13g2_fill_8 FILLER_126_648 ();
 sg13g2_fill_8 FILLER_126_656 ();
 sg13g2_fill_8 FILLER_126_664 ();
 sg13g2_fill_8 FILLER_126_672 ();
 sg13g2_fill_8 FILLER_126_680 ();
 sg13g2_fill_8 FILLER_126_688 ();
 sg13g2_fill_8 FILLER_126_696 ();
 sg13g2_fill_8 FILLER_126_704 ();
 sg13g2_fill_8 FILLER_126_712 ();
 sg13g2_fill_8 FILLER_126_720 ();
 sg13g2_fill_8 FILLER_126_728 ();
 sg13g2_fill_8 FILLER_126_736 ();
 sg13g2_fill_8 FILLER_126_744 ();
 sg13g2_fill_8 FILLER_126_752 ();
 sg13g2_fill_8 FILLER_126_760 ();
 sg13g2_fill_8 FILLER_126_768 ();
 sg13g2_fill_8 FILLER_126_776 ();
 sg13g2_fill_8 FILLER_126_784 ();
 sg13g2_fill_8 FILLER_126_792 ();
 sg13g2_fill_8 FILLER_126_800 ();
 sg13g2_fill_8 FILLER_126_808 ();
 sg13g2_fill_8 FILLER_126_816 ();
 sg13g2_fill_8 FILLER_126_824 ();
 sg13g2_fill_8 FILLER_126_832 ();
 sg13g2_fill_8 FILLER_126_840 ();
 sg13g2_fill_8 FILLER_126_848 ();
 sg13g2_fill_8 FILLER_126_856 ();
 sg13g2_fill_8 FILLER_126_864 ();
 sg13g2_fill_8 FILLER_126_872 ();
 sg13g2_fill_8 FILLER_126_880 ();
 sg13g2_fill_8 FILLER_126_888 ();
 sg13g2_fill_8 FILLER_126_896 ();
 sg13g2_fill_8 FILLER_126_904 ();
 sg13g2_fill_8 FILLER_126_912 ();
 sg13g2_fill_8 FILLER_126_920 ();
 sg13g2_fill_8 FILLER_126_928 ();
 sg13g2_fill_8 FILLER_126_936 ();
 sg13g2_fill_8 FILLER_126_944 ();
 sg13g2_fill_8 FILLER_126_952 ();
 sg13g2_fill_8 FILLER_126_960 ();
 sg13g2_fill_8 FILLER_126_968 ();
 sg13g2_fill_8 FILLER_126_976 ();
 sg13g2_fill_8 FILLER_126_984 ();
 sg13g2_fill_8 FILLER_126_992 ();
 sg13g2_fill_8 FILLER_126_1000 ();
 sg13g2_fill_8 FILLER_126_1008 ();
 sg13g2_fill_8 FILLER_126_1016 ();
 sg13g2_fill_8 FILLER_126_1024 ();
 sg13g2_fill_8 FILLER_126_1032 ();
 sg13g2_fill_8 FILLER_126_1040 ();
 sg13g2_fill_8 FILLER_126_1048 ();
 sg13g2_fill_8 FILLER_126_1056 ();
 sg13g2_fill_8 FILLER_126_1064 ();
 sg13g2_fill_8 FILLER_126_1072 ();
 sg13g2_fill_8 FILLER_126_1080 ();
 sg13g2_fill_8 FILLER_126_1088 ();
 sg13g2_fill_8 FILLER_126_1096 ();
 sg13g2_fill_8 FILLER_126_1104 ();
 sg13g2_fill_8 FILLER_126_1112 ();
 sg13g2_fill_8 FILLER_126_1120 ();
 sg13g2_fill_8 FILLER_126_1128 ();
 sg13g2_fill_8 FILLER_126_1136 ();
 sg13g2_fill_8 FILLER_126_1144 ();
 sg13g2_fill_8 FILLER_126_1152 ();
 sg13g2_fill_4 FILLER_126_1160 ();
 sg13g2_fill_2 FILLER_126_1164 ();
 sg13g2_fill_8 FILLER_127_0 ();
 sg13g2_fill_8 FILLER_127_8 ();
 sg13g2_fill_8 FILLER_127_16 ();
 sg13g2_fill_8 FILLER_127_24 ();
 sg13g2_fill_8 FILLER_127_32 ();
 sg13g2_fill_8 FILLER_127_40 ();
 sg13g2_fill_8 FILLER_127_48 ();
 sg13g2_fill_8 FILLER_127_56 ();
 sg13g2_fill_8 FILLER_127_64 ();
 sg13g2_fill_8 FILLER_127_72 ();
 sg13g2_fill_8 FILLER_127_80 ();
 sg13g2_fill_8 FILLER_127_88 ();
 sg13g2_fill_8 FILLER_127_96 ();
 sg13g2_fill_8 FILLER_127_104 ();
 sg13g2_fill_8 FILLER_127_112 ();
 sg13g2_fill_8 FILLER_127_120 ();
 sg13g2_fill_8 FILLER_127_128 ();
 sg13g2_fill_8 FILLER_127_136 ();
 sg13g2_fill_8 FILLER_127_144 ();
 sg13g2_fill_8 FILLER_127_152 ();
 sg13g2_fill_8 FILLER_127_160 ();
 sg13g2_fill_8 FILLER_127_168 ();
 sg13g2_fill_8 FILLER_127_176 ();
 sg13g2_fill_8 FILLER_127_184 ();
 sg13g2_fill_8 FILLER_127_192 ();
 sg13g2_fill_8 FILLER_127_200 ();
 sg13g2_fill_8 FILLER_127_208 ();
 sg13g2_fill_8 FILLER_127_216 ();
 sg13g2_fill_8 FILLER_127_224 ();
 sg13g2_fill_8 FILLER_127_232 ();
 sg13g2_fill_8 FILLER_127_240 ();
 sg13g2_fill_8 FILLER_127_248 ();
 sg13g2_fill_8 FILLER_127_256 ();
 sg13g2_fill_8 FILLER_127_264 ();
 sg13g2_fill_8 FILLER_127_272 ();
 sg13g2_fill_8 FILLER_127_280 ();
 sg13g2_fill_8 FILLER_127_288 ();
 sg13g2_fill_8 FILLER_127_296 ();
 sg13g2_fill_8 FILLER_127_304 ();
 sg13g2_fill_8 FILLER_127_312 ();
 sg13g2_fill_8 FILLER_127_320 ();
 sg13g2_fill_8 FILLER_127_328 ();
 sg13g2_fill_8 FILLER_127_336 ();
 sg13g2_fill_8 FILLER_127_344 ();
 sg13g2_fill_8 FILLER_127_352 ();
 sg13g2_fill_8 FILLER_127_360 ();
 sg13g2_fill_8 FILLER_127_368 ();
 sg13g2_fill_8 FILLER_127_376 ();
 sg13g2_fill_8 FILLER_127_384 ();
 sg13g2_fill_8 FILLER_127_392 ();
 sg13g2_fill_8 FILLER_127_400 ();
 sg13g2_fill_8 FILLER_127_408 ();
 sg13g2_fill_8 FILLER_127_416 ();
 sg13g2_fill_8 FILLER_127_424 ();
 sg13g2_fill_8 FILLER_127_432 ();
 sg13g2_fill_8 FILLER_127_440 ();
 sg13g2_fill_8 FILLER_127_448 ();
 sg13g2_fill_8 FILLER_127_456 ();
 sg13g2_fill_8 FILLER_127_464 ();
 sg13g2_fill_8 FILLER_127_472 ();
 sg13g2_fill_8 FILLER_127_480 ();
 sg13g2_fill_8 FILLER_127_488 ();
 sg13g2_fill_8 FILLER_127_496 ();
 sg13g2_fill_8 FILLER_127_504 ();
 sg13g2_fill_8 FILLER_127_512 ();
 sg13g2_fill_8 FILLER_127_520 ();
 sg13g2_fill_8 FILLER_127_528 ();
 sg13g2_fill_8 FILLER_127_536 ();
 sg13g2_fill_8 FILLER_127_544 ();
 sg13g2_fill_8 FILLER_127_552 ();
 sg13g2_fill_8 FILLER_127_560 ();
 sg13g2_fill_8 FILLER_127_568 ();
 sg13g2_fill_8 FILLER_127_576 ();
 sg13g2_fill_8 FILLER_127_584 ();
 sg13g2_fill_8 FILLER_127_592 ();
 sg13g2_fill_8 FILLER_127_600 ();
 sg13g2_fill_8 FILLER_127_608 ();
 sg13g2_fill_8 FILLER_127_616 ();
 sg13g2_fill_8 FILLER_127_624 ();
 sg13g2_fill_8 FILLER_127_632 ();
 sg13g2_fill_8 FILLER_127_640 ();
 sg13g2_fill_8 FILLER_127_648 ();
 sg13g2_fill_8 FILLER_127_656 ();
 sg13g2_fill_8 FILLER_127_664 ();
 sg13g2_fill_8 FILLER_127_672 ();
 sg13g2_fill_8 FILLER_127_680 ();
 sg13g2_fill_8 FILLER_127_688 ();
 sg13g2_fill_8 FILLER_127_696 ();
 sg13g2_fill_8 FILLER_127_704 ();
 sg13g2_fill_8 FILLER_127_712 ();
 sg13g2_fill_8 FILLER_127_720 ();
 sg13g2_fill_8 FILLER_127_728 ();
 sg13g2_fill_8 FILLER_127_736 ();
 sg13g2_fill_8 FILLER_127_744 ();
 sg13g2_fill_8 FILLER_127_752 ();
 sg13g2_fill_8 FILLER_127_760 ();
 sg13g2_fill_8 FILLER_127_768 ();
 sg13g2_fill_8 FILLER_127_776 ();
 sg13g2_fill_8 FILLER_127_784 ();
 sg13g2_fill_8 FILLER_127_792 ();
 sg13g2_fill_8 FILLER_127_800 ();
 sg13g2_fill_8 FILLER_127_808 ();
 sg13g2_fill_8 FILLER_127_816 ();
 sg13g2_fill_8 FILLER_127_824 ();
 sg13g2_fill_8 FILLER_127_832 ();
 sg13g2_fill_8 FILLER_127_840 ();
 sg13g2_fill_8 FILLER_127_848 ();
 sg13g2_fill_8 FILLER_127_856 ();
 sg13g2_fill_8 FILLER_127_864 ();
 sg13g2_fill_8 FILLER_127_872 ();
 sg13g2_fill_8 FILLER_127_880 ();
 sg13g2_fill_8 FILLER_127_888 ();
 sg13g2_fill_8 FILLER_127_896 ();
 sg13g2_fill_8 FILLER_127_904 ();
 sg13g2_fill_8 FILLER_127_912 ();
 sg13g2_fill_8 FILLER_127_920 ();
 sg13g2_fill_8 FILLER_127_928 ();
 sg13g2_fill_8 FILLER_127_936 ();
 sg13g2_fill_8 FILLER_127_944 ();
 sg13g2_fill_8 FILLER_127_952 ();
 sg13g2_fill_8 FILLER_127_960 ();
 sg13g2_fill_8 FILLER_127_968 ();
 sg13g2_fill_8 FILLER_127_976 ();
 sg13g2_fill_8 FILLER_127_984 ();
 sg13g2_fill_8 FILLER_127_992 ();
 sg13g2_fill_8 FILLER_127_1000 ();
 sg13g2_fill_8 FILLER_127_1008 ();
 sg13g2_fill_8 FILLER_127_1016 ();
 sg13g2_fill_8 FILLER_127_1024 ();
 sg13g2_fill_8 FILLER_127_1032 ();
 sg13g2_fill_8 FILLER_127_1040 ();
 sg13g2_fill_8 FILLER_127_1048 ();
 sg13g2_fill_8 FILLER_127_1056 ();
 sg13g2_fill_8 FILLER_127_1064 ();
 sg13g2_fill_8 FILLER_127_1072 ();
 sg13g2_fill_8 FILLER_127_1080 ();
 sg13g2_fill_8 FILLER_127_1088 ();
 sg13g2_fill_8 FILLER_127_1096 ();
 sg13g2_fill_8 FILLER_127_1104 ();
 sg13g2_fill_8 FILLER_127_1112 ();
 sg13g2_fill_8 FILLER_127_1120 ();
 sg13g2_fill_8 FILLER_127_1128 ();
 sg13g2_fill_8 FILLER_127_1136 ();
 sg13g2_fill_8 FILLER_127_1144 ();
 sg13g2_fill_8 FILLER_127_1152 ();
 sg13g2_fill_4 FILLER_127_1160 ();
 sg13g2_fill_2 FILLER_127_1164 ();
 sg13g2_fill_8 FILLER_128_0 ();
 sg13g2_fill_8 FILLER_128_8 ();
 sg13g2_fill_8 FILLER_128_16 ();
 sg13g2_fill_8 FILLER_128_24 ();
 sg13g2_fill_8 FILLER_128_32 ();
 sg13g2_fill_8 FILLER_128_40 ();
 sg13g2_fill_8 FILLER_128_48 ();
 sg13g2_fill_8 FILLER_128_56 ();
 sg13g2_fill_8 FILLER_128_64 ();
 sg13g2_fill_8 FILLER_128_72 ();
 sg13g2_fill_8 FILLER_128_80 ();
 sg13g2_fill_8 FILLER_128_88 ();
 sg13g2_fill_8 FILLER_128_96 ();
 sg13g2_fill_8 FILLER_128_104 ();
 sg13g2_fill_8 FILLER_128_112 ();
 sg13g2_fill_8 FILLER_128_120 ();
 sg13g2_fill_8 FILLER_128_128 ();
 sg13g2_fill_8 FILLER_128_136 ();
 sg13g2_fill_8 FILLER_128_144 ();
 sg13g2_fill_8 FILLER_128_152 ();
 sg13g2_fill_8 FILLER_128_160 ();
 sg13g2_fill_8 FILLER_128_168 ();
 sg13g2_fill_8 FILLER_128_176 ();
 sg13g2_fill_8 FILLER_128_184 ();
 sg13g2_fill_8 FILLER_128_192 ();
 sg13g2_fill_8 FILLER_128_200 ();
 sg13g2_fill_8 FILLER_128_208 ();
 sg13g2_fill_8 FILLER_128_216 ();
 sg13g2_fill_8 FILLER_128_224 ();
 sg13g2_fill_8 FILLER_128_232 ();
 sg13g2_fill_8 FILLER_128_240 ();
 sg13g2_fill_8 FILLER_128_248 ();
 sg13g2_fill_8 FILLER_128_256 ();
 sg13g2_fill_8 FILLER_128_264 ();
 sg13g2_fill_8 FILLER_128_272 ();
 sg13g2_fill_8 FILLER_128_280 ();
 sg13g2_fill_8 FILLER_128_288 ();
 sg13g2_fill_8 FILLER_128_296 ();
 sg13g2_fill_8 FILLER_128_304 ();
 sg13g2_fill_8 FILLER_128_312 ();
 sg13g2_fill_8 FILLER_128_320 ();
 sg13g2_fill_8 FILLER_128_328 ();
 sg13g2_fill_8 FILLER_128_336 ();
 sg13g2_fill_8 FILLER_128_344 ();
 sg13g2_fill_8 FILLER_128_352 ();
 sg13g2_fill_8 FILLER_128_360 ();
 sg13g2_fill_8 FILLER_128_368 ();
 sg13g2_fill_8 FILLER_128_376 ();
 sg13g2_fill_8 FILLER_128_384 ();
 sg13g2_fill_8 FILLER_128_392 ();
 sg13g2_fill_8 FILLER_128_400 ();
 sg13g2_fill_8 FILLER_128_408 ();
 sg13g2_fill_8 FILLER_128_416 ();
 sg13g2_fill_8 FILLER_128_424 ();
 sg13g2_fill_8 FILLER_128_432 ();
 sg13g2_fill_8 FILLER_128_440 ();
 sg13g2_fill_8 FILLER_128_448 ();
 sg13g2_fill_8 FILLER_128_456 ();
 sg13g2_fill_8 FILLER_128_464 ();
 sg13g2_fill_8 FILLER_128_472 ();
 sg13g2_fill_8 FILLER_128_480 ();
 sg13g2_fill_8 FILLER_128_488 ();
 sg13g2_fill_8 FILLER_128_496 ();
 sg13g2_fill_8 FILLER_128_504 ();
 sg13g2_fill_8 FILLER_128_512 ();
 sg13g2_fill_8 FILLER_128_520 ();
 sg13g2_fill_8 FILLER_128_528 ();
 sg13g2_fill_8 FILLER_128_536 ();
 sg13g2_fill_8 FILLER_128_544 ();
 sg13g2_fill_8 FILLER_128_552 ();
 sg13g2_fill_8 FILLER_128_560 ();
 sg13g2_fill_8 FILLER_128_568 ();
 sg13g2_fill_8 FILLER_128_576 ();
 sg13g2_fill_8 FILLER_128_584 ();
 sg13g2_fill_8 FILLER_128_592 ();
 sg13g2_fill_8 FILLER_128_600 ();
 sg13g2_fill_8 FILLER_128_608 ();
 sg13g2_fill_8 FILLER_128_616 ();
 sg13g2_fill_8 FILLER_128_624 ();
 sg13g2_fill_8 FILLER_128_632 ();
 sg13g2_fill_8 FILLER_128_640 ();
 sg13g2_fill_8 FILLER_128_648 ();
 sg13g2_fill_8 FILLER_128_656 ();
 sg13g2_fill_8 FILLER_128_664 ();
 sg13g2_fill_8 FILLER_128_672 ();
 sg13g2_fill_8 FILLER_128_680 ();
 sg13g2_fill_8 FILLER_128_688 ();
 sg13g2_fill_8 FILLER_128_696 ();
 sg13g2_fill_8 FILLER_128_704 ();
 sg13g2_fill_8 FILLER_128_712 ();
 sg13g2_fill_8 FILLER_128_720 ();
 sg13g2_fill_8 FILLER_128_728 ();
 sg13g2_fill_8 FILLER_128_736 ();
 sg13g2_fill_8 FILLER_128_744 ();
 sg13g2_fill_8 FILLER_128_752 ();
 sg13g2_fill_8 FILLER_128_760 ();
 sg13g2_fill_8 FILLER_128_768 ();
 sg13g2_fill_8 FILLER_128_776 ();
 sg13g2_fill_8 FILLER_128_784 ();
 sg13g2_fill_8 FILLER_128_792 ();
 sg13g2_fill_8 FILLER_128_800 ();
 sg13g2_fill_8 FILLER_128_808 ();
 sg13g2_fill_8 FILLER_128_816 ();
 sg13g2_fill_8 FILLER_128_824 ();
 sg13g2_fill_8 FILLER_128_832 ();
 sg13g2_fill_8 FILLER_128_840 ();
 sg13g2_fill_8 FILLER_128_848 ();
 sg13g2_fill_8 FILLER_128_856 ();
 sg13g2_fill_8 FILLER_128_864 ();
 sg13g2_fill_8 FILLER_128_872 ();
 sg13g2_fill_8 FILLER_128_880 ();
 sg13g2_fill_8 FILLER_128_888 ();
 sg13g2_fill_8 FILLER_128_896 ();
 sg13g2_fill_8 FILLER_128_904 ();
 sg13g2_fill_8 FILLER_128_912 ();
 sg13g2_fill_8 FILLER_128_920 ();
 sg13g2_fill_8 FILLER_128_928 ();
 sg13g2_fill_8 FILLER_128_936 ();
 sg13g2_fill_8 FILLER_128_944 ();
 sg13g2_fill_8 FILLER_128_952 ();
 sg13g2_fill_8 FILLER_128_960 ();
 sg13g2_fill_8 FILLER_128_968 ();
 sg13g2_fill_8 FILLER_128_976 ();
 sg13g2_fill_8 FILLER_128_984 ();
 sg13g2_fill_8 FILLER_128_992 ();
 sg13g2_fill_8 FILLER_128_1000 ();
 sg13g2_fill_8 FILLER_128_1008 ();
 sg13g2_fill_8 FILLER_128_1016 ();
 sg13g2_fill_8 FILLER_128_1024 ();
 sg13g2_fill_8 FILLER_128_1032 ();
 sg13g2_fill_8 FILLER_128_1040 ();
 sg13g2_fill_8 FILLER_128_1048 ();
 sg13g2_fill_8 FILLER_128_1056 ();
 sg13g2_fill_8 FILLER_128_1064 ();
 sg13g2_fill_8 FILLER_128_1072 ();
 sg13g2_fill_8 FILLER_128_1080 ();
 sg13g2_fill_8 FILLER_128_1088 ();
 sg13g2_fill_8 FILLER_128_1096 ();
 sg13g2_fill_8 FILLER_128_1104 ();
 sg13g2_fill_8 FILLER_128_1112 ();
 sg13g2_fill_8 FILLER_128_1120 ();
 sg13g2_fill_8 FILLER_128_1128 ();
 sg13g2_fill_8 FILLER_128_1136 ();
 sg13g2_fill_8 FILLER_128_1144 ();
 sg13g2_fill_8 FILLER_128_1152 ();
 sg13g2_fill_4 FILLER_128_1160 ();
 sg13g2_fill_2 FILLER_128_1164 ();
 sg13g2_fill_8 FILLER_129_0 ();
 sg13g2_fill_8 FILLER_129_8 ();
 sg13g2_fill_8 FILLER_129_16 ();
 sg13g2_fill_8 FILLER_129_24 ();
 sg13g2_fill_8 FILLER_129_32 ();
 sg13g2_fill_8 FILLER_129_40 ();
 sg13g2_fill_8 FILLER_129_48 ();
 sg13g2_fill_8 FILLER_129_56 ();
 sg13g2_fill_8 FILLER_129_64 ();
 sg13g2_fill_8 FILLER_129_72 ();
 sg13g2_fill_8 FILLER_129_80 ();
 sg13g2_fill_8 FILLER_129_88 ();
 sg13g2_fill_8 FILLER_129_96 ();
 sg13g2_fill_8 FILLER_129_104 ();
 sg13g2_fill_8 FILLER_129_112 ();
 sg13g2_fill_8 FILLER_129_120 ();
 sg13g2_fill_8 FILLER_129_128 ();
 sg13g2_fill_8 FILLER_129_136 ();
 sg13g2_fill_8 FILLER_129_144 ();
 sg13g2_fill_8 FILLER_129_152 ();
 sg13g2_fill_8 FILLER_129_160 ();
 sg13g2_fill_8 FILLER_129_168 ();
 sg13g2_fill_8 FILLER_129_176 ();
 sg13g2_fill_8 FILLER_129_184 ();
 sg13g2_fill_8 FILLER_129_192 ();
 sg13g2_fill_8 FILLER_129_200 ();
 sg13g2_fill_8 FILLER_129_208 ();
 sg13g2_fill_8 FILLER_129_216 ();
 sg13g2_fill_8 FILLER_129_224 ();
 sg13g2_fill_8 FILLER_129_232 ();
 sg13g2_fill_8 FILLER_129_240 ();
 sg13g2_fill_8 FILLER_129_248 ();
 sg13g2_fill_8 FILLER_129_256 ();
 sg13g2_fill_8 FILLER_129_264 ();
 sg13g2_fill_8 FILLER_129_272 ();
 sg13g2_fill_8 FILLER_129_280 ();
 sg13g2_fill_8 FILLER_129_288 ();
 sg13g2_fill_8 FILLER_129_296 ();
 sg13g2_fill_8 FILLER_129_304 ();
 sg13g2_fill_8 FILLER_129_312 ();
 sg13g2_fill_8 FILLER_129_320 ();
 sg13g2_fill_8 FILLER_129_328 ();
 sg13g2_fill_8 FILLER_129_336 ();
 sg13g2_fill_8 FILLER_129_344 ();
 sg13g2_fill_8 FILLER_129_352 ();
 sg13g2_fill_8 FILLER_129_360 ();
 sg13g2_fill_8 FILLER_129_368 ();
 sg13g2_fill_8 FILLER_129_376 ();
 sg13g2_fill_8 FILLER_129_384 ();
 sg13g2_fill_8 FILLER_129_392 ();
 sg13g2_fill_8 FILLER_129_400 ();
 sg13g2_fill_8 FILLER_129_408 ();
 sg13g2_fill_8 FILLER_129_416 ();
 sg13g2_fill_8 FILLER_129_424 ();
 sg13g2_fill_8 FILLER_129_432 ();
 sg13g2_fill_8 FILLER_129_440 ();
 sg13g2_fill_8 FILLER_129_448 ();
 sg13g2_fill_8 FILLER_129_456 ();
 sg13g2_fill_8 FILLER_129_464 ();
 sg13g2_fill_8 FILLER_129_472 ();
 sg13g2_fill_8 FILLER_129_480 ();
 sg13g2_fill_8 FILLER_129_488 ();
 sg13g2_fill_8 FILLER_129_496 ();
 sg13g2_fill_8 FILLER_129_504 ();
 sg13g2_fill_8 FILLER_129_512 ();
 sg13g2_fill_8 FILLER_129_520 ();
 sg13g2_fill_8 FILLER_129_528 ();
 sg13g2_fill_8 FILLER_129_536 ();
 sg13g2_fill_8 FILLER_129_544 ();
 sg13g2_fill_8 FILLER_129_552 ();
 sg13g2_fill_8 FILLER_129_560 ();
 sg13g2_fill_8 FILLER_129_568 ();
 sg13g2_fill_8 FILLER_129_576 ();
 sg13g2_fill_8 FILLER_129_584 ();
 sg13g2_fill_8 FILLER_129_592 ();
 sg13g2_fill_8 FILLER_129_600 ();
 sg13g2_fill_8 FILLER_129_608 ();
 sg13g2_fill_8 FILLER_129_616 ();
 sg13g2_fill_8 FILLER_129_624 ();
 sg13g2_fill_8 FILLER_129_632 ();
 sg13g2_fill_8 FILLER_129_640 ();
 sg13g2_fill_8 FILLER_129_648 ();
 sg13g2_fill_8 FILLER_129_656 ();
 sg13g2_fill_8 FILLER_129_664 ();
 sg13g2_fill_8 FILLER_129_672 ();
 sg13g2_fill_8 FILLER_129_680 ();
 sg13g2_fill_8 FILLER_129_688 ();
 sg13g2_fill_8 FILLER_129_696 ();
 sg13g2_fill_8 FILLER_129_704 ();
 sg13g2_fill_8 FILLER_129_712 ();
 sg13g2_fill_8 FILLER_129_720 ();
 sg13g2_fill_8 FILLER_129_728 ();
 sg13g2_fill_8 FILLER_129_736 ();
 sg13g2_fill_8 FILLER_129_744 ();
 sg13g2_fill_8 FILLER_129_752 ();
 sg13g2_fill_8 FILLER_129_760 ();
 sg13g2_fill_8 FILLER_129_768 ();
 sg13g2_fill_8 FILLER_129_776 ();
 sg13g2_fill_8 FILLER_129_784 ();
 sg13g2_fill_8 FILLER_129_792 ();
 sg13g2_fill_8 FILLER_129_800 ();
 sg13g2_fill_8 FILLER_129_808 ();
 sg13g2_fill_8 FILLER_129_816 ();
 sg13g2_fill_8 FILLER_129_824 ();
 sg13g2_fill_8 FILLER_129_832 ();
 sg13g2_fill_8 FILLER_129_840 ();
 sg13g2_fill_8 FILLER_129_848 ();
 sg13g2_fill_8 FILLER_129_856 ();
 sg13g2_fill_8 FILLER_129_864 ();
 sg13g2_fill_8 FILLER_129_872 ();
 sg13g2_fill_8 FILLER_129_880 ();
 sg13g2_fill_8 FILLER_129_888 ();
 sg13g2_fill_8 FILLER_129_896 ();
 sg13g2_fill_8 FILLER_129_904 ();
 sg13g2_fill_8 FILLER_129_912 ();
 sg13g2_fill_8 FILLER_129_920 ();
 sg13g2_fill_8 FILLER_129_928 ();
 sg13g2_fill_8 FILLER_129_936 ();
 sg13g2_fill_8 FILLER_129_944 ();
 sg13g2_fill_8 FILLER_129_952 ();
 sg13g2_fill_8 FILLER_129_960 ();
 sg13g2_fill_8 FILLER_129_968 ();
 sg13g2_fill_8 FILLER_129_976 ();
 sg13g2_fill_8 FILLER_129_984 ();
 sg13g2_fill_8 FILLER_129_992 ();
 sg13g2_fill_8 FILLER_129_1000 ();
 sg13g2_fill_8 FILLER_129_1008 ();
 sg13g2_fill_8 FILLER_129_1016 ();
 sg13g2_fill_8 FILLER_129_1024 ();
 sg13g2_fill_8 FILLER_129_1032 ();
 sg13g2_fill_8 FILLER_129_1040 ();
 sg13g2_fill_8 FILLER_129_1048 ();
 sg13g2_fill_8 FILLER_129_1056 ();
 sg13g2_fill_8 FILLER_129_1064 ();
 sg13g2_fill_8 FILLER_129_1072 ();
 sg13g2_fill_8 FILLER_129_1080 ();
 sg13g2_fill_8 FILLER_129_1088 ();
 sg13g2_fill_8 FILLER_129_1096 ();
 sg13g2_fill_8 FILLER_129_1104 ();
 sg13g2_fill_8 FILLER_129_1112 ();
 sg13g2_fill_8 FILLER_129_1120 ();
 sg13g2_fill_8 FILLER_129_1128 ();
 sg13g2_fill_8 FILLER_129_1136 ();
 sg13g2_fill_8 FILLER_129_1144 ();
 sg13g2_fill_8 FILLER_129_1152 ();
 sg13g2_fill_4 FILLER_129_1160 ();
 sg13g2_fill_2 FILLER_129_1164 ();
 sg13g2_fill_8 FILLER_130_0 ();
 sg13g2_fill_8 FILLER_130_8 ();
 sg13g2_fill_8 FILLER_130_16 ();
 sg13g2_fill_8 FILLER_130_24 ();
 sg13g2_fill_8 FILLER_130_32 ();
 sg13g2_fill_8 FILLER_130_40 ();
 sg13g2_fill_8 FILLER_130_48 ();
 sg13g2_fill_8 FILLER_130_56 ();
 sg13g2_fill_8 FILLER_130_64 ();
 sg13g2_fill_8 FILLER_130_72 ();
 sg13g2_fill_8 FILLER_130_80 ();
 sg13g2_fill_8 FILLER_130_88 ();
 sg13g2_fill_8 FILLER_130_96 ();
 sg13g2_fill_8 FILLER_130_104 ();
 sg13g2_fill_8 FILLER_130_112 ();
 sg13g2_fill_8 FILLER_130_120 ();
 sg13g2_fill_8 FILLER_130_128 ();
 sg13g2_fill_8 FILLER_130_136 ();
 sg13g2_fill_8 FILLER_130_144 ();
 sg13g2_fill_8 FILLER_130_152 ();
 sg13g2_fill_8 FILLER_130_160 ();
 sg13g2_fill_8 FILLER_130_168 ();
 sg13g2_fill_8 FILLER_130_176 ();
 sg13g2_fill_8 FILLER_130_184 ();
 sg13g2_fill_8 FILLER_130_192 ();
 sg13g2_fill_8 FILLER_130_200 ();
 sg13g2_fill_8 FILLER_130_208 ();
 sg13g2_fill_8 FILLER_130_216 ();
 sg13g2_fill_8 FILLER_130_224 ();
 sg13g2_fill_8 FILLER_130_232 ();
 sg13g2_fill_8 FILLER_130_240 ();
 sg13g2_fill_8 FILLER_130_248 ();
 sg13g2_fill_8 FILLER_130_256 ();
 sg13g2_fill_8 FILLER_130_264 ();
 sg13g2_fill_8 FILLER_130_272 ();
 sg13g2_fill_8 FILLER_130_280 ();
 sg13g2_fill_8 FILLER_130_288 ();
 sg13g2_fill_8 FILLER_130_296 ();
 sg13g2_fill_8 FILLER_130_304 ();
 sg13g2_fill_8 FILLER_130_312 ();
 sg13g2_fill_8 FILLER_130_320 ();
 sg13g2_fill_8 FILLER_130_328 ();
 sg13g2_fill_8 FILLER_130_336 ();
 sg13g2_fill_8 FILLER_130_344 ();
 sg13g2_fill_8 FILLER_130_352 ();
 sg13g2_fill_8 FILLER_130_360 ();
 sg13g2_fill_8 FILLER_130_368 ();
 sg13g2_fill_8 FILLER_130_376 ();
 sg13g2_fill_8 FILLER_130_384 ();
 sg13g2_fill_8 FILLER_130_392 ();
 sg13g2_fill_8 FILLER_130_400 ();
 sg13g2_fill_8 FILLER_130_408 ();
 sg13g2_fill_8 FILLER_130_416 ();
 sg13g2_fill_8 FILLER_130_424 ();
 sg13g2_fill_8 FILLER_130_432 ();
 sg13g2_fill_8 FILLER_130_440 ();
 sg13g2_fill_8 FILLER_130_448 ();
 sg13g2_fill_8 FILLER_130_456 ();
 sg13g2_fill_8 FILLER_130_464 ();
 sg13g2_fill_8 FILLER_130_472 ();
 sg13g2_fill_8 FILLER_130_480 ();
 sg13g2_fill_8 FILLER_130_488 ();
 sg13g2_fill_8 FILLER_130_496 ();
 sg13g2_fill_8 FILLER_130_504 ();
 sg13g2_fill_8 FILLER_130_512 ();
 sg13g2_fill_8 FILLER_130_520 ();
 sg13g2_fill_8 FILLER_130_528 ();
 sg13g2_fill_8 FILLER_130_536 ();
 sg13g2_fill_8 FILLER_130_544 ();
 sg13g2_fill_8 FILLER_130_552 ();
 sg13g2_fill_8 FILLER_130_560 ();
 sg13g2_fill_8 FILLER_130_568 ();
 sg13g2_fill_8 FILLER_130_576 ();
 sg13g2_fill_8 FILLER_130_584 ();
 sg13g2_fill_8 FILLER_130_592 ();
 sg13g2_fill_8 FILLER_130_600 ();
 sg13g2_fill_8 FILLER_130_608 ();
 sg13g2_fill_8 FILLER_130_616 ();
 sg13g2_fill_8 FILLER_130_624 ();
 sg13g2_fill_8 FILLER_130_632 ();
 sg13g2_fill_8 FILLER_130_640 ();
 sg13g2_fill_8 FILLER_130_648 ();
 sg13g2_fill_8 FILLER_130_656 ();
 sg13g2_fill_8 FILLER_130_664 ();
 sg13g2_fill_8 FILLER_130_672 ();
 sg13g2_fill_8 FILLER_130_680 ();
 sg13g2_fill_8 FILLER_130_688 ();
 sg13g2_fill_8 FILLER_130_696 ();
 sg13g2_fill_8 FILLER_130_704 ();
 sg13g2_fill_8 FILLER_130_712 ();
 sg13g2_fill_8 FILLER_130_720 ();
 sg13g2_fill_8 FILLER_130_728 ();
 sg13g2_fill_8 FILLER_130_736 ();
 sg13g2_fill_8 FILLER_130_744 ();
 sg13g2_fill_8 FILLER_130_752 ();
 sg13g2_fill_8 FILLER_130_760 ();
 sg13g2_fill_8 FILLER_130_768 ();
 sg13g2_fill_8 FILLER_130_776 ();
 sg13g2_fill_8 FILLER_130_784 ();
 sg13g2_fill_8 FILLER_130_792 ();
 sg13g2_fill_8 FILLER_130_800 ();
 sg13g2_fill_8 FILLER_130_808 ();
 sg13g2_fill_8 FILLER_130_816 ();
 sg13g2_fill_8 FILLER_130_824 ();
 sg13g2_fill_8 FILLER_130_832 ();
 sg13g2_fill_8 FILLER_130_840 ();
 sg13g2_fill_8 FILLER_130_848 ();
 sg13g2_fill_8 FILLER_130_856 ();
 sg13g2_fill_8 FILLER_130_864 ();
 sg13g2_fill_8 FILLER_130_872 ();
 sg13g2_fill_8 FILLER_130_880 ();
 sg13g2_fill_8 FILLER_130_888 ();
 sg13g2_fill_8 FILLER_130_896 ();
 sg13g2_fill_8 FILLER_130_904 ();
 sg13g2_fill_8 FILLER_130_912 ();
 sg13g2_fill_8 FILLER_130_920 ();
 sg13g2_fill_8 FILLER_130_928 ();
 sg13g2_fill_8 FILLER_130_936 ();
 sg13g2_fill_8 FILLER_130_944 ();
 sg13g2_fill_8 FILLER_130_952 ();
 sg13g2_fill_8 FILLER_130_960 ();
 sg13g2_fill_8 FILLER_130_968 ();
 sg13g2_fill_8 FILLER_130_976 ();
 sg13g2_fill_8 FILLER_130_984 ();
 sg13g2_fill_8 FILLER_130_992 ();
 sg13g2_fill_8 FILLER_130_1000 ();
 sg13g2_fill_8 FILLER_130_1008 ();
 sg13g2_fill_8 FILLER_130_1016 ();
 sg13g2_fill_8 FILLER_130_1024 ();
 sg13g2_fill_8 FILLER_130_1032 ();
 sg13g2_fill_8 FILLER_130_1040 ();
 sg13g2_fill_8 FILLER_130_1048 ();
 sg13g2_fill_8 FILLER_130_1056 ();
 sg13g2_fill_8 FILLER_130_1064 ();
 sg13g2_fill_8 FILLER_130_1072 ();
 sg13g2_fill_8 FILLER_130_1080 ();
 sg13g2_fill_8 FILLER_130_1088 ();
 sg13g2_fill_8 FILLER_130_1096 ();
 sg13g2_fill_8 FILLER_130_1104 ();
 sg13g2_fill_8 FILLER_130_1112 ();
 sg13g2_fill_8 FILLER_130_1120 ();
 sg13g2_fill_8 FILLER_130_1128 ();
 sg13g2_fill_8 FILLER_130_1136 ();
 sg13g2_fill_8 FILLER_130_1144 ();
 sg13g2_fill_8 FILLER_130_1152 ();
 sg13g2_fill_4 FILLER_130_1160 ();
 sg13g2_fill_2 FILLER_130_1164 ();
 sg13g2_fill_8 FILLER_131_0 ();
 sg13g2_fill_8 FILLER_131_8 ();
 sg13g2_fill_8 FILLER_131_16 ();
 sg13g2_fill_8 FILLER_131_24 ();
 sg13g2_fill_8 FILLER_131_32 ();
 sg13g2_fill_8 FILLER_131_40 ();
 sg13g2_fill_8 FILLER_131_48 ();
 sg13g2_fill_8 FILLER_131_56 ();
 sg13g2_fill_8 FILLER_131_64 ();
 sg13g2_fill_8 FILLER_131_72 ();
 sg13g2_fill_8 FILLER_131_80 ();
 sg13g2_fill_8 FILLER_131_88 ();
 sg13g2_fill_8 FILLER_131_96 ();
 sg13g2_fill_8 FILLER_131_104 ();
 sg13g2_fill_8 FILLER_131_112 ();
 sg13g2_fill_8 FILLER_131_120 ();
 sg13g2_fill_8 FILLER_131_128 ();
 sg13g2_fill_8 FILLER_131_136 ();
 sg13g2_fill_8 FILLER_131_144 ();
 sg13g2_fill_8 FILLER_131_152 ();
 sg13g2_fill_8 FILLER_131_160 ();
 sg13g2_fill_8 FILLER_131_168 ();
 sg13g2_fill_8 FILLER_131_176 ();
 sg13g2_fill_8 FILLER_131_184 ();
 sg13g2_fill_8 FILLER_131_192 ();
 sg13g2_fill_8 FILLER_131_200 ();
 sg13g2_fill_8 FILLER_131_208 ();
 sg13g2_fill_8 FILLER_131_216 ();
 sg13g2_fill_8 FILLER_131_224 ();
 sg13g2_fill_8 FILLER_131_232 ();
 sg13g2_fill_8 FILLER_131_240 ();
 sg13g2_fill_8 FILLER_131_248 ();
 sg13g2_fill_8 FILLER_131_256 ();
 sg13g2_fill_8 FILLER_131_264 ();
 sg13g2_fill_8 FILLER_131_272 ();
 sg13g2_fill_8 FILLER_131_280 ();
 sg13g2_fill_8 FILLER_131_288 ();
 sg13g2_fill_8 FILLER_131_296 ();
 sg13g2_fill_8 FILLER_131_304 ();
 sg13g2_fill_8 FILLER_131_312 ();
 sg13g2_fill_8 FILLER_131_320 ();
 sg13g2_fill_8 FILLER_131_328 ();
 sg13g2_fill_8 FILLER_131_336 ();
 sg13g2_fill_8 FILLER_131_344 ();
 sg13g2_fill_8 FILLER_131_352 ();
 sg13g2_fill_8 FILLER_131_360 ();
 sg13g2_fill_8 FILLER_131_368 ();
 sg13g2_fill_8 FILLER_131_376 ();
 sg13g2_fill_8 FILLER_131_384 ();
 sg13g2_fill_8 FILLER_131_392 ();
 sg13g2_fill_8 FILLER_131_400 ();
 sg13g2_fill_8 FILLER_131_408 ();
 sg13g2_fill_8 FILLER_131_416 ();
 sg13g2_fill_8 FILLER_131_424 ();
 sg13g2_fill_8 FILLER_131_432 ();
 sg13g2_fill_8 FILLER_131_440 ();
 sg13g2_fill_8 FILLER_131_448 ();
 sg13g2_fill_8 FILLER_131_456 ();
 sg13g2_fill_8 FILLER_131_464 ();
 sg13g2_fill_8 FILLER_131_472 ();
 sg13g2_fill_8 FILLER_131_480 ();
 sg13g2_fill_8 FILLER_131_488 ();
 sg13g2_fill_8 FILLER_131_496 ();
 sg13g2_fill_8 FILLER_131_504 ();
 sg13g2_fill_8 FILLER_131_512 ();
 sg13g2_fill_8 FILLER_131_520 ();
 sg13g2_fill_8 FILLER_131_528 ();
 sg13g2_fill_8 FILLER_131_536 ();
 sg13g2_fill_8 FILLER_131_544 ();
 sg13g2_fill_8 FILLER_131_552 ();
 sg13g2_fill_8 FILLER_131_560 ();
 sg13g2_fill_8 FILLER_131_568 ();
 sg13g2_fill_8 FILLER_131_576 ();
 sg13g2_fill_8 FILLER_131_584 ();
 sg13g2_fill_8 FILLER_131_592 ();
 sg13g2_fill_8 FILLER_131_600 ();
 sg13g2_fill_8 FILLER_131_608 ();
 sg13g2_fill_8 FILLER_131_616 ();
 sg13g2_fill_8 FILLER_131_624 ();
 sg13g2_fill_8 FILLER_131_632 ();
 sg13g2_fill_8 FILLER_131_640 ();
 sg13g2_fill_8 FILLER_131_648 ();
 sg13g2_fill_8 FILLER_131_656 ();
 sg13g2_fill_8 FILLER_131_664 ();
 sg13g2_fill_8 FILLER_131_672 ();
 sg13g2_fill_8 FILLER_131_680 ();
 sg13g2_fill_8 FILLER_131_688 ();
 sg13g2_fill_8 FILLER_131_696 ();
 sg13g2_fill_8 FILLER_131_704 ();
 sg13g2_fill_8 FILLER_131_712 ();
 sg13g2_fill_8 FILLER_131_720 ();
 sg13g2_fill_8 FILLER_131_728 ();
 sg13g2_fill_8 FILLER_131_736 ();
 sg13g2_fill_8 FILLER_131_744 ();
 sg13g2_fill_8 FILLER_131_752 ();
 sg13g2_fill_8 FILLER_131_760 ();
 sg13g2_fill_8 FILLER_131_768 ();
 sg13g2_fill_8 FILLER_131_776 ();
 sg13g2_fill_8 FILLER_131_784 ();
 sg13g2_fill_8 FILLER_131_792 ();
 sg13g2_fill_8 FILLER_131_800 ();
 sg13g2_fill_8 FILLER_131_808 ();
 sg13g2_fill_8 FILLER_131_816 ();
 sg13g2_fill_8 FILLER_131_824 ();
 sg13g2_fill_8 FILLER_131_832 ();
 sg13g2_fill_8 FILLER_131_840 ();
 sg13g2_fill_8 FILLER_131_848 ();
 sg13g2_fill_8 FILLER_131_856 ();
 sg13g2_fill_8 FILLER_131_864 ();
 sg13g2_fill_8 FILLER_131_872 ();
 sg13g2_fill_8 FILLER_131_880 ();
 sg13g2_fill_8 FILLER_131_888 ();
 sg13g2_fill_8 FILLER_131_896 ();
 sg13g2_fill_8 FILLER_131_904 ();
 sg13g2_fill_8 FILLER_131_912 ();
 sg13g2_fill_8 FILLER_131_920 ();
 sg13g2_fill_8 FILLER_131_928 ();
 sg13g2_fill_8 FILLER_131_936 ();
 sg13g2_fill_8 FILLER_131_944 ();
 sg13g2_fill_8 FILLER_131_952 ();
 sg13g2_fill_8 FILLER_131_960 ();
 sg13g2_fill_8 FILLER_131_968 ();
 sg13g2_fill_8 FILLER_131_976 ();
 sg13g2_fill_8 FILLER_131_984 ();
 sg13g2_fill_8 FILLER_131_992 ();
 sg13g2_fill_8 FILLER_131_1000 ();
 sg13g2_fill_8 FILLER_131_1008 ();
 sg13g2_fill_8 FILLER_131_1016 ();
 sg13g2_fill_8 FILLER_131_1024 ();
 sg13g2_fill_8 FILLER_131_1032 ();
 sg13g2_fill_8 FILLER_131_1040 ();
 sg13g2_fill_8 FILLER_131_1048 ();
 sg13g2_fill_8 FILLER_131_1056 ();
 sg13g2_fill_8 FILLER_131_1064 ();
 sg13g2_fill_8 FILLER_131_1072 ();
 sg13g2_fill_8 FILLER_131_1080 ();
 sg13g2_fill_8 FILLER_131_1088 ();
 sg13g2_fill_8 FILLER_131_1096 ();
 sg13g2_fill_8 FILLER_131_1104 ();
 sg13g2_fill_8 FILLER_131_1112 ();
 sg13g2_fill_8 FILLER_131_1120 ();
 sg13g2_fill_8 FILLER_131_1128 ();
 sg13g2_fill_8 FILLER_131_1136 ();
 sg13g2_fill_8 FILLER_131_1144 ();
 sg13g2_fill_8 FILLER_131_1152 ();
 sg13g2_fill_4 FILLER_131_1160 ();
 sg13g2_fill_2 FILLER_131_1164 ();
 sg13g2_fill_8 FILLER_132_0 ();
 sg13g2_fill_8 FILLER_132_8 ();
 sg13g2_fill_8 FILLER_132_16 ();
 sg13g2_fill_8 FILLER_132_24 ();
 sg13g2_fill_8 FILLER_132_32 ();
 sg13g2_fill_8 FILLER_132_40 ();
 sg13g2_fill_8 FILLER_132_48 ();
 sg13g2_fill_8 FILLER_132_56 ();
 sg13g2_fill_8 FILLER_132_64 ();
 sg13g2_fill_8 FILLER_132_72 ();
 sg13g2_fill_8 FILLER_132_80 ();
 sg13g2_fill_8 FILLER_132_88 ();
 sg13g2_fill_8 FILLER_132_96 ();
 sg13g2_fill_8 FILLER_132_104 ();
 sg13g2_fill_8 FILLER_132_112 ();
 sg13g2_fill_8 FILLER_132_120 ();
 sg13g2_fill_8 FILLER_132_128 ();
 sg13g2_fill_8 FILLER_132_136 ();
 sg13g2_fill_8 FILLER_132_144 ();
 sg13g2_fill_8 FILLER_132_152 ();
 sg13g2_fill_8 FILLER_132_160 ();
 sg13g2_fill_8 FILLER_132_168 ();
 sg13g2_fill_8 FILLER_132_176 ();
 sg13g2_fill_8 FILLER_132_184 ();
 sg13g2_fill_8 FILLER_132_192 ();
 sg13g2_fill_8 FILLER_132_200 ();
 sg13g2_fill_8 FILLER_132_208 ();
 sg13g2_fill_8 FILLER_132_216 ();
 sg13g2_fill_8 FILLER_132_224 ();
 sg13g2_fill_8 FILLER_132_232 ();
 sg13g2_fill_8 FILLER_132_240 ();
 sg13g2_fill_8 FILLER_132_248 ();
 sg13g2_fill_8 FILLER_132_256 ();
 sg13g2_fill_8 FILLER_132_264 ();
 sg13g2_fill_8 FILLER_132_272 ();
 sg13g2_fill_8 FILLER_132_280 ();
 sg13g2_fill_8 FILLER_132_288 ();
 sg13g2_fill_8 FILLER_132_296 ();
 sg13g2_fill_8 FILLER_132_304 ();
 sg13g2_fill_8 FILLER_132_312 ();
 sg13g2_fill_8 FILLER_132_320 ();
 sg13g2_fill_8 FILLER_132_328 ();
 sg13g2_fill_8 FILLER_132_336 ();
 sg13g2_fill_8 FILLER_132_344 ();
 sg13g2_fill_8 FILLER_132_352 ();
 sg13g2_fill_8 FILLER_132_360 ();
 sg13g2_fill_8 FILLER_132_368 ();
 sg13g2_fill_8 FILLER_132_376 ();
 sg13g2_fill_8 FILLER_132_384 ();
 sg13g2_fill_8 FILLER_132_392 ();
 sg13g2_fill_8 FILLER_132_400 ();
 sg13g2_fill_8 FILLER_132_408 ();
 sg13g2_fill_8 FILLER_132_416 ();
 sg13g2_fill_8 FILLER_132_424 ();
 sg13g2_fill_8 FILLER_132_432 ();
 sg13g2_fill_8 FILLER_132_440 ();
 sg13g2_fill_8 FILLER_132_448 ();
 sg13g2_fill_8 FILLER_132_456 ();
 sg13g2_fill_8 FILLER_132_464 ();
 sg13g2_fill_8 FILLER_132_472 ();
 sg13g2_fill_8 FILLER_132_480 ();
 sg13g2_fill_8 FILLER_132_488 ();
 sg13g2_fill_8 FILLER_132_496 ();
 sg13g2_fill_8 FILLER_132_504 ();
 sg13g2_fill_8 FILLER_132_512 ();
 sg13g2_fill_8 FILLER_132_520 ();
 sg13g2_fill_8 FILLER_132_528 ();
 sg13g2_fill_8 FILLER_132_536 ();
 sg13g2_fill_8 FILLER_132_544 ();
 sg13g2_fill_8 FILLER_132_552 ();
 sg13g2_fill_8 FILLER_132_560 ();
 sg13g2_fill_8 FILLER_132_568 ();
 sg13g2_fill_8 FILLER_132_576 ();
 sg13g2_fill_8 FILLER_132_584 ();
 sg13g2_fill_8 FILLER_132_592 ();
 sg13g2_fill_8 FILLER_132_600 ();
 sg13g2_fill_8 FILLER_132_608 ();
 sg13g2_fill_8 FILLER_132_616 ();
 sg13g2_fill_8 FILLER_132_624 ();
 sg13g2_fill_8 FILLER_132_632 ();
 sg13g2_fill_8 FILLER_132_640 ();
 sg13g2_fill_8 FILLER_132_648 ();
 sg13g2_fill_8 FILLER_132_656 ();
 sg13g2_fill_8 FILLER_132_664 ();
 sg13g2_fill_8 FILLER_132_672 ();
 sg13g2_fill_8 FILLER_132_680 ();
 sg13g2_fill_8 FILLER_132_688 ();
 sg13g2_fill_8 FILLER_132_696 ();
 sg13g2_fill_8 FILLER_132_704 ();
 sg13g2_fill_8 FILLER_132_712 ();
 sg13g2_fill_8 FILLER_132_720 ();
 sg13g2_fill_8 FILLER_132_728 ();
 sg13g2_fill_8 FILLER_132_736 ();
 sg13g2_fill_8 FILLER_132_744 ();
 sg13g2_fill_8 FILLER_132_752 ();
 sg13g2_fill_8 FILLER_132_760 ();
 sg13g2_fill_8 FILLER_132_768 ();
 sg13g2_fill_8 FILLER_132_776 ();
 sg13g2_fill_8 FILLER_132_784 ();
 sg13g2_fill_8 FILLER_132_792 ();
 sg13g2_fill_8 FILLER_132_800 ();
 sg13g2_fill_8 FILLER_132_808 ();
 sg13g2_fill_8 FILLER_132_816 ();
 sg13g2_fill_8 FILLER_132_824 ();
 sg13g2_fill_8 FILLER_132_832 ();
 sg13g2_fill_8 FILLER_132_840 ();
 sg13g2_fill_8 FILLER_132_848 ();
 sg13g2_fill_8 FILLER_132_856 ();
 sg13g2_fill_8 FILLER_132_864 ();
 sg13g2_fill_8 FILLER_132_872 ();
 sg13g2_fill_8 FILLER_132_880 ();
 sg13g2_fill_8 FILLER_132_888 ();
 sg13g2_fill_8 FILLER_132_896 ();
 sg13g2_fill_8 FILLER_132_904 ();
 sg13g2_fill_8 FILLER_132_912 ();
 sg13g2_fill_8 FILLER_132_920 ();
 sg13g2_fill_8 FILLER_132_928 ();
 sg13g2_fill_8 FILLER_132_936 ();
 sg13g2_fill_8 FILLER_132_944 ();
 sg13g2_fill_8 FILLER_132_952 ();
 sg13g2_fill_8 FILLER_132_960 ();
 sg13g2_fill_8 FILLER_132_968 ();
 sg13g2_fill_8 FILLER_132_976 ();
 sg13g2_fill_8 FILLER_132_984 ();
 sg13g2_fill_8 FILLER_132_992 ();
 sg13g2_fill_8 FILLER_132_1000 ();
 sg13g2_fill_8 FILLER_132_1008 ();
 sg13g2_fill_8 FILLER_132_1016 ();
 sg13g2_fill_8 FILLER_132_1024 ();
 sg13g2_fill_8 FILLER_132_1032 ();
 sg13g2_fill_8 FILLER_132_1040 ();
 sg13g2_fill_8 FILLER_132_1048 ();
 sg13g2_fill_8 FILLER_132_1056 ();
 sg13g2_fill_8 FILLER_132_1064 ();
 sg13g2_fill_8 FILLER_132_1072 ();
 sg13g2_fill_8 FILLER_132_1080 ();
 sg13g2_fill_8 FILLER_132_1088 ();
 sg13g2_fill_8 FILLER_132_1096 ();
 sg13g2_fill_8 FILLER_132_1104 ();
 sg13g2_fill_8 FILLER_132_1112 ();
 sg13g2_fill_8 FILLER_132_1120 ();
 sg13g2_fill_8 FILLER_132_1128 ();
 sg13g2_fill_8 FILLER_132_1136 ();
 sg13g2_fill_8 FILLER_132_1144 ();
 sg13g2_fill_8 FILLER_132_1152 ();
 sg13g2_fill_4 FILLER_132_1160 ();
 sg13g2_fill_2 FILLER_132_1164 ();
 sg13g2_fill_8 FILLER_133_0 ();
 sg13g2_fill_8 FILLER_133_8 ();
 sg13g2_fill_8 FILLER_133_16 ();
 sg13g2_fill_8 FILLER_133_24 ();
 sg13g2_fill_8 FILLER_133_32 ();
 sg13g2_fill_8 FILLER_133_40 ();
 sg13g2_fill_8 FILLER_133_48 ();
 sg13g2_fill_8 FILLER_133_56 ();
 sg13g2_fill_8 FILLER_133_64 ();
 sg13g2_fill_8 FILLER_133_72 ();
 sg13g2_fill_8 FILLER_133_80 ();
 sg13g2_fill_8 FILLER_133_88 ();
 sg13g2_fill_8 FILLER_133_96 ();
 sg13g2_fill_8 FILLER_133_104 ();
 sg13g2_fill_8 FILLER_133_112 ();
 sg13g2_fill_8 FILLER_133_120 ();
 sg13g2_fill_8 FILLER_133_128 ();
 sg13g2_fill_8 FILLER_133_136 ();
 sg13g2_fill_8 FILLER_133_144 ();
 sg13g2_fill_8 FILLER_133_152 ();
 sg13g2_fill_8 FILLER_133_160 ();
 sg13g2_fill_8 FILLER_133_168 ();
 sg13g2_fill_8 FILLER_133_176 ();
 sg13g2_fill_8 FILLER_133_184 ();
 sg13g2_fill_8 FILLER_133_192 ();
 sg13g2_fill_8 FILLER_133_200 ();
 sg13g2_fill_8 FILLER_133_208 ();
 sg13g2_fill_8 FILLER_133_216 ();
 sg13g2_fill_8 FILLER_133_224 ();
 sg13g2_fill_8 FILLER_133_232 ();
 sg13g2_fill_8 FILLER_133_240 ();
 sg13g2_fill_8 FILLER_133_248 ();
 sg13g2_fill_8 FILLER_133_256 ();
 sg13g2_fill_8 FILLER_133_264 ();
 sg13g2_fill_8 FILLER_133_272 ();
 sg13g2_fill_8 FILLER_133_280 ();
 sg13g2_fill_8 FILLER_133_288 ();
 sg13g2_fill_8 FILLER_133_296 ();
 sg13g2_fill_8 FILLER_133_304 ();
 sg13g2_fill_8 FILLER_133_312 ();
 sg13g2_fill_8 FILLER_133_320 ();
 sg13g2_fill_8 FILLER_133_328 ();
 sg13g2_fill_8 FILLER_133_336 ();
 sg13g2_fill_8 FILLER_133_344 ();
 sg13g2_fill_8 FILLER_133_352 ();
 sg13g2_fill_8 FILLER_133_360 ();
 sg13g2_fill_8 FILLER_133_368 ();
 sg13g2_fill_8 FILLER_133_376 ();
 sg13g2_fill_8 FILLER_133_384 ();
 sg13g2_fill_8 FILLER_133_392 ();
 sg13g2_fill_8 FILLER_133_400 ();
 sg13g2_fill_8 FILLER_133_408 ();
 sg13g2_fill_8 FILLER_133_416 ();
 sg13g2_fill_8 FILLER_133_424 ();
 sg13g2_fill_8 FILLER_133_432 ();
 sg13g2_fill_8 FILLER_133_440 ();
 sg13g2_fill_8 FILLER_133_448 ();
 sg13g2_fill_8 FILLER_133_456 ();
 sg13g2_fill_8 FILLER_133_464 ();
 sg13g2_fill_8 FILLER_133_472 ();
 sg13g2_fill_8 FILLER_133_480 ();
 sg13g2_fill_8 FILLER_133_488 ();
 sg13g2_fill_8 FILLER_133_496 ();
 sg13g2_fill_8 FILLER_133_504 ();
 sg13g2_fill_8 FILLER_133_512 ();
 sg13g2_fill_8 FILLER_133_520 ();
 sg13g2_fill_8 FILLER_133_528 ();
 sg13g2_fill_8 FILLER_133_536 ();
 sg13g2_fill_8 FILLER_133_544 ();
 sg13g2_fill_8 FILLER_133_552 ();
 sg13g2_fill_8 FILLER_133_560 ();
 sg13g2_fill_8 FILLER_133_568 ();
 sg13g2_fill_8 FILLER_133_576 ();
 sg13g2_fill_8 FILLER_133_584 ();
 sg13g2_fill_8 FILLER_133_592 ();
 sg13g2_fill_8 FILLER_133_600 ();
 sg13g2_fill_8 FILLER_133_608 ();
 sg13g2_fill_8 FILLER_133_616 ();
 sg13g2_fill_8 FILLER_133_624 ();
 sg13g2_fill_8 FILLER_133_632 ();
 sg13g2_fill_8 FILLER_133_640 ();
 sg13g2_fill_8 FILLER_133_648 ();
 sg13g2_fill_8 FILLER_133_656 ();
 sg13g2_fill_8 FILLER_133_664 ();
 sg13g2_fill_8 FILLER_133_672 ();
 sg13g2_fill_8 FILLER_133_680 ();
 sg13g2_fill_8 FILLER_133_688 ();
 sg13g2_fill_8 FILLER_133_696 ();
 sg13g2_fill_8 FILLER_133_704 ();
 sg13g2_fill_8 FILLER_133_712 ();
 sg13g2_fill_8 FILLER_133_720 ();
 sg13g2_fill_8 FILLER_133_728 ();
 sg13g2_fill_8 FILLER_133_736 ();
 sg13g2_fill_8 FILLER_133_744 ();
 sg13g2_fill_8 FILLER_133_752 ();
 sg13g2_fill_8 FILLER_133_760 ();
 sg13g2_fill_8 FILLER_133_768 ();
 sg13g2_fill_8 FILLER_133_776 ();
 sg13g2_fill_8 FILLER_133_784 ();
 sg13g2_fill_8 FILLER_133_792 ();
 sg13g2_fill_8 FILLER_133_800 ();
 sg13g2_fill_8 FILLER_133_808 ();
 sg13g2_fill_8 FILLER_133_816 ();
 sg13g2_fill_8 FILLER_133_824 ();
 sg13g2_fill_8 FILLER_133_832 ();
 sg13g2_fill_8 FILLER_133_840 ();
 sg13g2_fill_8 FILLER_133_848 ();
 sg13g2_fill_8 FILLER_133_856 ();
 sg13g2_fill_8 FILLER_133_864 ();
 sg13g2_fill_8 FILLER_133_872 ();
 sg13g2_fill_8 FILLER_133_880 ();
 sg13g2_fill_8 FILLER_133_888 ();
 sg13g2_fill_8 FILLER_133_896 ();
 sg13g2_fill_8 FILLER_133_904 ();
 sg13g2_fill_8 FILLER_133_912 ();
 sg13g2_fill_8 FILLER_133_920 ();
 sg13g2_fill_8 FILLER_133_928 ();
 sg13g2_fill_8 FILLER_133_936 ();
 sg13g2_fill_8 FILLER_133_944 ();
 sg13g2_fill_8 FILLER_133_952 ();
 sg13g2_fill_8 FILLER_133_960 ();
 sg13g2_fill_8 FILLER_133_968 ();
 sg13g2_fill_8 FILLER_133_976 ();
 sg13g2_fill_8 FILLER_133_984 ();
 sg13g2_fill_8 FILLER_133_992 ();
 sg13g2_fill_8 FILLER_133_1000 ();
 sg13g2_fill_8 FILLER_133_1008 ();
 sg13g2_fill_8 FILLER_133_1016 ();
 sg13g2_fill_8 FILLER_133_1024 ();
 sg13g2_fill_8 FILLER_133_1032 ();
 sg13g2_fill_8 FILLER_133_1040 ();
 sg13g2_fill_8 FILLER_133_1048 ();
 sg13g2_fill_8 FILLER_133_1056 ();
 sg13g2_fill_8 FILLER_133_1064 ();
 sg13g2_fill_8 FILLER_133_1072 ();
 sg13g2_fill_8 FILLER_133_1080 ();
 sg13g2_fill_8 FILLER_133_1088 ();
 sg13g2_fill_8 FILLER_133_1096 ();
 sg13g2_fill_8 FILLER_133_1104 ();
 sg13g2_fill_8 FILLER_133_1112 ();
 sg13g2_fill_8 FILLER_133_1120 ();
 sg13g2_fill_8 FILLER_133_1128 ();
 sg13g2_fill_8 FILLER_133_1136 ();
 sg13g2_fill_8 FILLER_133_1144 ();
 sg13g2_fill_8 FILLER_133_1152 ();
 sg13g2_fill_4 FILLER_133_1160 ();
 sg13g2_fill_2 FILLER_133_1164 ();
 sg13g2_fill_8 FILLER_134_0 ();
 sg13g2_fill_8 FILLER_134_8 ();
 sg13g2_fill_8 FILLER_134_16 ();
 sg13g2_fill_8 FILLER_134_24 ();
 sg13g2_fill_8 FILLER_134_32 ();
 sg13g2_fill_8 FILLER_134_40 ();
 sg13g2_fill_8 FILLER_134_48 ();
 sg13g2_fill_8 FILLER_134_56 ();
 sg13g2_fill_8 FILLER_134_64 ();
 sg13g2_fill_8 FILLER_134_72 ();
 sg13g2_fill_8 FILLER_134_80 ();
 sg13g2_fill_8 FILLER_134_88 ();
 sg13g2_fill_8 FILLER_134_96 ();
 sg13g2_fill_8 FILLER_134_104 ();
 sg13g2_fill_8 FILLER_134_112 ();
 sg13g2_fill_8 FILLER_134_120 ();
 sg13g2_fill_8 FILLER_134_128 ();
 sg13g2_fill_8 FILLER_134_136 ();
 sg13g2_fill_8 FILLER_134_144 ();
 sg13g2_fill_8 FILLER_134_152 ();
 sg13g2_fill_8 FILLER_134_160 ();
 sg13g2_fill_8 FILLER_134_168 ();
 sg13g2_fill_8 FILLER_134_176 ();
 sg13g2_fill_8 FILLER_134_184 ();
 sg13g2_fill_8 FILLER_134_192 ();
 sg13g2_fill_8 FILLER_134_200 ();
 sg13g2_fill_8 FILLER_134_208 ();
 sg13g2_fill_8 FILLER_134_216 ();
 sg13g2_fill_8 FILLER_134_224 ();
 sg13g2_fill_8 FILLER_134_232 ();
 sg13g2_fill_8 FILLER_134_240 ();
 sg13g2_fill_8 FILLER_134_248 ();
 sg13g2_fill_8 FILLER_134_256 ();
 sg13g2_fill_8 FILLER_134_264 ();
 sg13g2_fill_8 FILLER_134_272 ();
 sg13g2_fill_8 FILLER_134_280 ();
 sg13g2_fill_8 FILLER_134_288 ();
 sg13g2_fill_8 FILLER_134_296 ();
 sg13g2_fill_8 FILLER_134_304 ();
 sg13g2_fill_8 FILLER_134_312 ();
 sg13g2_fill_8 FILLER_134_320 ();
 sg13g2_fill_8 FILLER_134_328 ();
 sg13g2_fill_8 FILLER_134_336 ();
 sg13g2_fill_8 FILLER_134_344 ();
 sg13g2_fill_8 FILLER_134_352 ();
 sg13g2_fill_8 FILLER_134_360 ();
 sg13g2_fill_8 FILLER_134_368 ();
 sg13g2_fill_8 FILLER_134_376 ();
 sg13g2_fill_8 FILLER_134_384 ();
 sg13g2_fill_8 FILLER_134_392 ();
 sg13g2_fill_8 FILLER_134_400 ();
 sg13g2_fill_8 FILLER_134_408 ();
 sg13g2_fill_8 FILLER_134_416 ();
 sg13g2_fill_8 FILLER_134_424 ();
 sg13g2_fill_8 FILLER_134_432 ();
 sg13g2_fill_8 FILLER_134_440 ();
 sg13g2_fill_8 FILLER_134_448 ();
 sg13g2_fill_8 FILLER_134_456 ();
 sg13g2_fill_8 FILLER_134_464 ();
 sg13g2_fill_8 FILLER_134_472 ();
 sg13g2_fill_8 FILLER_134_480 ();
 sg13g2_fill_8 FILLER_134_488 ();
 sg13g2_fill_8 FILLER_134_496 ();
 sg13g2_fill_8 FILLER_134_504 ();
 sg13g2_fill_8 FILLER_134_512 ();
 sg13g2_fill_8 FILLER_134_520 ();
 sg13g2_fill_8 FILLER_134_528 ();
 sg13g2_fill_8 FILLER_134_536 ();
 sg13g2_fill_8 FILLER_134_544 ();
 sg13g2_fill_8 FILLER_134_552 ();
 sg13g2_fill_8 FILLER_134_560 ();
 sg13g2_fill_8 FILLER_134_568 ();
 sg13g2_fill_8 FILLER_134_576 ();
 sg13g2_fill_8 FILLER_134_584 ();
 sg13g2_fill_8 FILLER_134_592 ();
 sg13g2_fill_8 FILLER_134_600 ();
 sg13g2_fill_8 FILLER_134_608 ();
 sg13g2_fill_8 FILLER_134_616 ();
 sg13g2_fill_8 FILLER_134_624 ();
 sg13g2_fill_8 FILLER_134_632 ();
 sg13g2_fill_8 FILLER_134_640 ();
 sg13g2_fill_8 FILLER_134_648 ();
 sg13g2_fill_8 FILLER_134_656 ();
 sg13g2_fill_8 FILLER_134_664 ();
 sg13g2_fill_8 FILLER_134_672 ();
 sg13g2_fill_8 FILLER_134_680 ();
 sg13g2_fill_8 FILLER_134_688 ();
 sg13g2_fill_8 FILLER_134_696 ();
 sg13g2_fill_8 FILLER_134_704 ();
 sg13g2_fill_8 FILLER_134_712 ();
 sg13g2_fill_8 FILLER_134_720 ();
 sg13g2_fill_8 FILLER_134_728 ();
 sg13g2_fill_8 FILLER_134_736 ();
 sg13g2_fill_8 FILLER_134_744 ();
 sg13g2_fill_8 FILLER_134_752 ();
 sg13g2_fill_8 FILLER_134_760 ();
 sg13g2_fill_8 FILLER_134_768 ();
 sg13g2_fill_8 FILLER_134_776 ();
 sg13g2_fill_8 FILLER_134_784 ();
 sg13g2_fill_8 FILLER_134_792 ();
 sg13g2_fill_8 FILLER_134_800 ();
 sg13g2_fill_8 FILLER_134_808 ();
 sg13g2_fill_8 FILLER_134_816 ();
 sg13g2_fill_8 FILLER_134_824 ();
 sg13g2_fill_8 FILLER_134_832 ();
 sg13g2_fill_8 FILLER_134_840 ();
 sg13g2_fill_8 FILLER_134_848 ();
 sg13g2_fill_8 FILLER_134_856 ();
 sg13g2_fill_8 FILLER_134_864 ();
 sg13g2_fill_8 FILLER_134_872 ();
 sg13g2_fill_8 FILLER_134_880 ();
 sg13g2_fill_8 FILLER_134_888 ();
 sg13g2_fill_8 FILLER_134_896 ();
 sg13g2_fill_8 FILLER_134_904 ();
 sg13g2_fill_8 FILLER_134_912 ();
 sg13g2_fill_8 FILLER_134_920 ();
 sg13g2_fill_8 FILLER_134_928 ();
 sg13g2_fill_8 FILLER_134_936 ();
 sg13g2_fill_8 FILLER_134_944 ();
 sg13g2_fill_8 FILLER_134_952 ();
 sg13g2_fill_8 FILLER_134_960 ();
 sg13g2_fill_8 FILLER_134_968 ();
 sg13g2_fill_8 FILLER_134_976 ();
 sg13g2_fill_8 FILLER_134_984 ();
 sg13g2_fill_8 FILLER_134_992 ();
 sg13g2_fill_8 FILLER_134_1000 ();
 sg13g2_fill_8 FILLER_134_1008 ();
 sg13g2_fill_8 FILLER_134_1016 ();
 sg13g2_fill_8 FILLER_134_1024 ();
 sg13g2_fill_8 FILLER_134_1032 ();
 sg13g2_fill_8 FILLER_134_1040 ();
 sg13g2_fill_8 FILLER_134_1048 ();
 sg13g2_fill_8 FILLER_134_1056 ();
 sg13g2_fill_8 FILLER_134_1064 ();
 sg13g2_fill_8 FILLER_134_1072 ();
 sg13g2_fill_8 FILLER_134_1080 ();
 sg13g2_fill_8 FILLER_134_1088 ();
 sg13g2_fill_8 FILLER_134_1096 ();
 sg13g2_fill_8 FILLER_134_1104 ();
 sg13g2_fill_8 FILLER_134_1112 ();
 sg13g2_fill_8 FILLER_134_1120 ();
 sg13g2_fill_8 FILLER_134_1128 ();
 sg13g2_fill_8 FILLER_134_1136 ();
 sg13g2_fill_8 FILLER_134_1144 ();
 sg13g2_fill_8 FILLER_134_1152 ();
 sg13g2_fill_4 FILLER_134_1160 ();
 sg13g2_fill_2 FILLER_134_1164 ();
 sg13g2_fill_8 FILLER_135_0 ();
 sg13g2_fill_8 FILLER_135_8 ();
 sg13g2_fill_8 FILLER_135_16 ();
 sg13g2_fill_8 FILLER_135_24 ();
 sg13g2_fill_8 FILLER_135_32 ();
 sg13g2_fill_8 FILLER_135_40 ();
 sg13g2_fill_8 FILLER_135_48 ();
 sg13g2_fill_8 FILLER_135_56 ();
 sg13g2_fill_8 FILLER_135_64 ();
 sg13g2_fill_8 FILLER_135_72 ();
 sg13g2_fill_8 FILLER_135_80 ();
 sg13g2_fill_8 FILLER_135_88 ();
 sg13g2_fill_8 FILLER_135_96 ();
 sg13g2_fill_8 FILLER_135_104 ();
 sg13g2_fill_8 FILLER_135_112 ();
 sg13g2_fill_8 FILLER_135_120 ();
 sg13g2_fill_8 FILLER_135_128 ();
 sg13g2_fill_8 FILLER_135_136 ();
 sg13g2_fill_8 FILLER_135_144 ();
 sg13g2_fill_8 FILLER_135_152 ();
 sg13g2_fill_8 FILLER_135_160 ();
 sg13g2_fill_8 FILLER_135_168 ();
 sg13g2_fill_8 FILLER_135_176 ();
 sg13g2_fill_8 FILLER_135_184 ();
 sg13g2_fill_8 FILLER_135_192 ();
 sg13g2_fill_8 FILLER_135_200 ();
 sg13g2_fill_8 FILLER_135_208 ();
 sg13g2_fill_8 FILLER_135_216 ();
 sg13g2_fill_8 FILLER_135_224 ();
 sg13g2_fill_8 FILLER_135_232 ();
 sg13g2_fill_8 FILLER_135_240 ();
 sg13g2_fill_8 FILLER_135_248 ();
 sg13g2_fill_8 FILLER_135_256 ();
 sg13g2_fill_8 FILLER_135_264 ();
 sg13g2_fill_8 FILLER_135_272 ();
 sg13g2_fill_8 FILLER_135_280 ();
 sg13g2_fill_8 FILLER_135_288 ();
 sg13g2_fill_8 FILLER_135_296 ();
 sg13g2_fill_8 FILLER_135_304 ();
 sg13g2_fill_8 FILLER_135_312 ();
 sg13g2_fill_8 FILLER_135_320 ();
 sg13g2_fill_8 FILLER_135_328 ();
 sg13g2_fill_8 FILLER_135_336 ();
 sg13g2_fill_8 FILLER_135_344 ();
 sg13g2_fill_8 FILLER_135_352 ();
 sg13g2_fill_8 FILLER_135_360 ();
 sg13g2_fill_8 FILLER_135_368 ();
 sg13g2_fill_8 FILLER_135_376 ();
 sg13g2_fill_8 FILLER_135_384 ();
 sg13g2_fill_8 FILLER_135_392 ();
 sg13g2_fill_8 FILLER_135_400 ();
 sg13g2_fill_8 FILLER_135_408 ();
 sg13g2_fill_8 FILLER_135_416 ();
 sg13g2_fill_8 FILLER_135_424 ();
 sg13g2_fill_8 FILLER_135_432 ();
 sg13g2_fill_8 FILLER_135_440 ();
 sg13g2_fill_8 FILLER_135_448 ();
 sg13g2_fill_8 FILLER_135_456 ();
 sg13g2_fill_8 FILLER_135_464 ();
 sg13g2_fill_8 FILLER_135_472 ();
 sg13g2_fill_8 FILLER_135_480 ();
 sg13g2_fill_8 FILLER_135_488 ();
 sg13g2_fill_8 FILLER_135_496 ();
 sg13g2_fill_8 FILLER_135_504 ();
 sg13g2_fill_8 FILLER_135_512 ();
 sg13g2_fill_8 FILLER_135_520 ();
 sg13g2_fill_8 FILLER_135_528 ();
 sg13g2_fill_8 FILLER_135_536 ();
 sg13g2_fill_8 FILLER_135_544 ();
 sg13g2_fill_8 FILLER_135_552 ();
 sg13g2_fill_8 FILLER_135_560 ();
 sg13g2_fill_8 FILLER_135_568 ();
 sg13g2_fill_8 FILLER_135_576 ();
 sg13g2_fill_8 FILLER_135_584 ();
 sg13g2_fill_8 FILLER_135_592 ();
 sg13g2_fill_8 FILLER_135_600 ();
 sg13g2_fill_8 FILLER_135_608 ();
 sg13g2_fill_8 FILLER_135_616 ();
 sg13g2_fill_8 FILLER_135_624 ();
 sg13g2_fill_8 FILLER_135_632 ();
 sg13g2_fill_8 FILLER_135_640 ();
 sg13g2_fill_8 FILLER_135_648 ();
 sg13g2_fill_8 FILLER_135_656 ();
 sg13g2_fill_8 FILLER_135_664 ();
 sg13g2_fill_8 FILLER_135_672 ();
 sg13g2_fill_8 FILLER_135_680 ();
 sg13g2_fill_8 FILLER_135_688 ();
 sg13g2_fill_8 FILLER_135_696 ();
 sg13g2_fill_8 FILLER_135_704 ();
 sg13g2_fill_8 FILLER_135_712 ();
 sg13g2_fill_8 FILLER_135_720 ();
 sg13g2_fill_8 FILLER_135_728 ();
 sg13g2_fill_8 FILLER_135_736 ();
 sg13g2_fill_8 FILLER_135_744 ();
 sg13g2_fill_8 FILLER_135_752 ();
 sg13g2_fill_8 FILLER_135_760 ();
 sg13g2_fill_8 FILLER_135_768 ();
 sg13g2_fill_8 FILLER_135_776 ();
 sg13g2_fill_8 FILLER_135_784 ();
 sg13g2_fill_8 FILLER_135_792 ();
 sg13g2_fill_8 FILLER_135_800 ();
 sg13g2_fill_8 FILLER_135_808 ();
 sg13g2_fill_8 FILLER_135_816 ();
 sg13g2_fill_8 FILLER_135_824 ();
 sg13g2_fill_8 FILLER_135_832 ();
 sg13g2_fill_8 FILLER_135_840 ();
 sg13g2_fill_8 FILLER_135_848 ();
 sg13g2_fill_8 FILLER_135_856 ();
 sg13g2_fill_8 FILLER_135_864 ();
 sg13g2_fill_8 FILLER_135_872 ();
 sg13g2_fill_8 FILLER_135_880 ();
 sg13g2_fill_8 FILLER_135_888 ();
 sg13g2_fill_8 FILLER_135_896 ();
 sg13g2_fill_8 FILLER_135_904 ();
 sg13g2_fill_8 FILLER_135_912 ();
 sg13g2_fill_8 FILLER_135_920 ();
 sg13g2_fill_8 FILLER_135_928 ();
 sg13g2_fill_8 FILLER_135_936 ();
 sg13g2_fill_8 FILLER_135_944 ();
 sg13g2_fill_8 FILLER_135_952 ();
 sg13g2_fill_8 FILLER_135_960 ();
 sg13g2_fill_8 FILLER_135_968 ();
 sg13g2_fill_8 FILLER_135_976 ();
 sg13g2_fill_8 FILLER_135_984 ();
 sg13g2_fill_8 FILLER_135_992 ();
 sg13g2_fill_8 FILLER_135_1000 ();
 sg13g2_fill_8 FILLER_135_1008 ();
 sg13g2_fill_8 FILLER_135_1016 ();
 sg13g2_fill_8 FILLER_135_1024 ();
 sg13g2_fill_8 FILLER_135_1032 ();
 sg13g2_fill_8 FILLER_135_1040 ();
 sg13g2_fill_8 FILLER_135_1048 ();
 sg13g2_fill_8 FILLER_135_1056 ();
 sg13g2_fill_8 FILLER_135_1064 ();
 sg13g2_fill_8 FILLER_135_1072 ();
 sg13g2_fill_8 FILLER_135_1080 ();
 sg13g2_fill_8 FILLER_135_1088 ();
 sg13g2_fill_8 FILLER_135_1096 ();
 sg13g2_fill_8 FILLER_135_1104 ();
 sg13g2_fill_8 FILLER_135_1112 ();
 sg13g2_fill_8 FILLER_135_1120 ();
 sg13g2_fill_8 FILLER_135_1128 ();
 sg13g2_fill_8 FILLER_135_1136 ();
 sg13g2_fill_8 FILLER_135_1144 ();
 sg13g2_fill_8 FILLER_135_1152 ();
 sg13g2_fill_4 FILLER_135_1160 ();
 sg13g2_fill_2 FILLER_135_1164 ();
 sg13g2_fill_8 FILLER_136_0 ();
 sg13g2_fill_8 FILLER_136_8 ();
 sg13g2_fill_8 FILLER_136_16 ();
 sg13g2_fill_8 FILLER_136_24 ();
 sg13g2_fill_8 FILLER_136_32 ();
 sg13g2_fill_8 FILLER_136_40 ();
 sg13g2_fill_8 FILLER_136_48 ();
 sg13g2_fill_8 FILLER_136_56 ();
 sg13g2_fill_8 FILLER_136_64 ();
 sg13g2_fill_8 FILLER_136_72 ();
 sg13g2_fill_8 FILLER_136_80 ();
 sg13g2_fill_8 FILLER_136_88 ();
 sg13g2_fill_8 FILLER_136_96 ();
 sg13g2_fill_8 FILLER_136_104 ();
 sg13g2_fill_8 FILLER_136_112 ();
 sg13g2_fill_8 FILLER_136_120 ();
 sg13g2_fill_8 FILLER_136_128 ();
 sg13g2_fill_8 FILLER_136_136 ();
 sg13g2_fill_8 FILLER_136_144 ();
 sg13g2_fill_8 FILLER_136_152 ();
 sg13g2_fill_8 FILLER_136_160 ();
 sg13g2_fill_8 FILLER_136_168 ();
 sg13g2_fill_8 FILLER_136_176 ();
 sg13g2_fill_8 FILLER_136_184 ();
 sg13g2_fill_8 FILLER_136_192 ();
 sg13g2_fill_8 FILLER_136_200 ();
 sg13g2_fill_8 FILLER_136_208 ();
 sg13g2_fill_8 FILLER_136_216 ();
 sg13g2_fill_8 FILLER_136_224 ();
 sg13g2_fill_8 FILLER_136_232 ();
 sg13g2_fill_8 FILLER_136_240 ();
 sg13g2_fill_8 FILLER_136_248 ();
 sg13g2_fill_8 FILLER_136_256 ();
 sg13g2_fill_8 FILLER_136_264 ();
 sg13g2_fill_8 FILLER_136_272 ();
 sg13g2_fill_8 FILLER_136_280 ();
 sg13g2_fill_8 FILLER_136_288 ();
 sg13g2_fill_8 FILLER_136_296 ();
 sg13g2_fill_8 FILLER_136_304 ();
 sg13g2_fill_8 FILLER_136_312 ();
 sg13g2_fill_8 FILLER_136_320 ();
 sg13g2_fill_8 FILLER_136_328 ();
 sg13g2_fill_8 FILLER_136_336 ();
 sg13g2_fill_8 FILLER_136_344 ();
 sg13g2_fill_8 FILLER_136_352 ();
 sg13g2_fill_8 FILLER_136_360 ();
 sg13g2_fill_8 FILLER_136_368 ();
 sg13g2_fill_8 FILLER_136_376 ();
 sg13g2_fill_8 FILLER_136_384 ();
 sg13g2_fill_8 FILLER_136_392 ();
 sg13g2_fill_8 FILLER_136_400 ();
 sg13g2_fill_8 FILLER_136_408 ();
 sg13g2_fill_8 FILLER_136_416 ();
 sg13g2_fill_8 FILLER_136_424 ();
 sg13g2_fill_8 FILLER_136_432 ();
 sg13g2_fill_8 FILLER_136_440 ();
 sg13g2_fill_8 FILLER_136_448 ();
 sg13g2_fill_8 FILLER_136_456 ();
 sg13g2_fill_8 FILLER_136_464 ();
 sg13g2_fill_8 FILLER_136_472 ();
 sg13g2_fill_8 FILLER_136_480 ();
 sg13g2_fill_8 FILLER_136_488 ();
 sg13g2_fill_8 FILLER_136_496 ();
 sg13g2_fill_8 FILLER_136_504 ();
 sg13g2_fill_8 FILLER_136_512 ();
 sg13g2_fill_8 FILLER_136_520 ();
 sg13g2_fill_8 FILLER_136_528 ();
 sg13g2_fill_8 FILLER_136_536 ();
 sg13g2_fill_8 FILLER_136_544 ();
 sg13g2_fill_8 FILLER_136_552 ();
 sg13g2_fill_8 FILLER_136_560 ();
 sg13g2_fill_8 FILLER_136_568 ();
 sg13g2_fill_8 FILLER_136_576 ();
 sg13g2_fill_8 FILLER_136_584 ();
 sg13g2_fill_8 FILLER_136_592 ();
 sg13g2_fill_8 FILLER_136_600 ();
 sg13g2_fill_8 FILLER_136_608 ();
 sg13g2_fill_8 FILLER_136_616 ();
 sg13g2_fill_8 FILLER_136_624 ();
 sg13g2_fill_8 FILLER_136_632 ();
 sg13g2_fill_8 FILLER_136_640 ();
 sg13g2_fill_8 FILLER_136_648 ();
 sg13g2_fill_8 FILLER_136_656 ();
 sg13g2_fill_8 FILLER_136_664 ();
 sg13g2_fill_8 FILLER_136_672 ();
 sg13g2_fill_8 FILLER_136_680 ();
 sg13g2_fill_8 FILLER_136_688 ();
 sg13g2_fill_8 FILLER_136_696 ();
 sg13g2_fill_8 FILLER_136_704 ();
 sg13g2_fill_8 FILLER_136_712 ();
 sg13g2_fill_8 FILLER_136_720 ();
 sg13g2_fill_8 FILLER_136_728 ();
 sg13g2_fill_8 FILLER_136_736 ();
 sg13g2_fill_8 FILLER_136_744 ();
 sg13g2_fill_8 FILLER_136_752 ();
 sg13g2_fill_8 FILLER_136_760 ();
 sg13g2_fill_8 FILLER_136_768 ();
 sg13g2_fill_8 FILLER_136_776 ();
 sg13g2_fill_8 FILLER_136_784 ();
 sg13g2_fill_8 FILLER_136_792 ();
 sg13g2_fill_8 FILLER_136_800 ();
 sg13g2_fill_8 FILLER_136_808 ();
 sg13g2_fill_8 FILLER_136_816 ();
 sg13g2_fill_8 FILLER_136_824 ();
 sg13g2_fill_8 FILLER_136_832 ();
 sg13g2_fill_8 FILLER_136_840 ();
 sg13g2_fill_8 FILLER_136_848 ();
 sg13g2_fill_8 FILLER_136_856 ();
 sg13g2_fill_8 FILLER_136_864 ();
 sg13g2_fill_8 FILLER_136_872 ();
 sg13g2_fill_8 FILLER_136_880 ();
 sg13g2_fill_8 FILLER_136_888 ();
 sg13g2_fill_8 FILLER_136_896 ();
 sg13g2_fill_8 FILLER_136_904 ();
 sg13g2_fill_8 FILLER_136_912 ();
 sg13g2_fill_8 FILLER_136_920 ();
 sg13g2_fill_8 FILLER_136_928 ();
 sg13g2_fill_8 FILLER_136_936 ();
 sg13g2_fill_8 FILLER_136_944 ();
 sg13g2_fill_8 FILLER_136_952 ();
 sg13g2_fill_8 FILLER_136_960 ();
 sg13g2_fill_8 FILLER_136_968 ();
 sg13g2_fill_8 FILLER_136_976 ();
 sg13g2_fill_8 FILLER_136_984 ();
 sg13g2_fill_8 FILLER_136_992 ();
 sg13g2_fill_8 FILLER_136_1000 ();
 sg13g2_fill_8 FILLER_136_1008 ();
 sg13g2_fill_8 FILLER_136_1016 ();
 sg13g2_fill_8 FILLER_136_1024 ();
 sg13g2_fill_8 FILLER_136_1032 ();
 sg13g2_fill_8 FILLER_136_1040 ();
 sg13g2_fill_8 FILLER_136_1048 ();
 sg13g2_fill_8 FILLER_136_1056 ();
 sg13g2_fill_8 FILLER_136_1064 ();
 sg13g2_fill_8 FILLER_136_1072 ();
 sg13g2_fill_8 FILLER_136_1080 ();
 sg13g2_fill_8 FILLER_136_1088 ();
 sg13g2_fill_8 FILLER_136_1096 ();
 sg13g2_fill_8 FILLER_136_1104 ();
 sg13g2_fill_8 FILLER_136_1112 ();
 sg13g2_fill_8 FILLER_136_1120 ();
 sg13g2_fill_8 FILLER_136_1128 ();
 sg13g2_fill_8 FILLER_136_1136 ();
 sg13g2_fill_8 FILLER_136_1144 ();
 sg13g2_fill_8 FILLER_136_1152 ();
 sg13g2_fill_4 FILLER_136_1160 ();
 sg13g2_fill_2 FILLER_136_1164 ();
 sg13g2_fill_8 FILLER_137_0 ();
 sg13g2_fill_8 FILLER_137_8 ();
 sg13g2_fill_8 FILLER_137_16 ();
 sg13g2_fill_8 FILLER_137_24 ();
 sg13g2_fill_8 FILLER_137_32 ();
 sg13g2_fill_8 FILLER_137_40 ();
 sg13g2_fill_8 FILLER_137_48 ();
 sg13g2_fill_8 FILLER_137_56 ();
 sg13g2_fill_8 FILLER_137_64 ();
 sg13g2_fill_8 FILLER_137_72 ();
 sg13g2_fill_8 FILLER_137_80 ();
 sg13g2_fill_8 FILLER_137_88 ();
 sg13g2_fill_8 FILLER_137_96 ();
 sg13g2_fill_8 FILLER_137_104 ();
 sg13g2_fill_8 FILLER_137_112 ();
 sg13g2_fill_8 FILLER_137_120 ();
 sg13g2_fill_8 FILLER_137_128 ();
 sg13g2_fill_8 FILLER_137_136 ();
 sg13g2_fill_8 FILLER_137_144 ();
 sg13g2_fill_8 FILLER_137_152 ();
 sg13g2_fill_8 FILLER_137_160 ();
 sg13g2_fill_8 FILLER_137_168 ();
 sg13g2_fill_8 FILLER_137_176 ();
 sg13g2_fill_8 FILLER_137_184 ();
 sg13g2_fill_8 FILLER_137_192 ();
 sg13g2_fill_8 FILLER_137_200 ();
 sg13g2_fill_8 FILLER_137_208 ();
 sg13g2_fill_8 FILLER_137_216 ();
 sg13g2_fill_8 FILLER_137_224 ();
 sg13g2_fill_8 FILLER_137_232 ();
 sg13g2_fill_8 FILLER_137_240 ();
 sg13g2_fill_8 FILLER_137_248 ();
 sg13g2_fill_8 FILLER_137_256 ();
 sg13g2_fill_8 FILLER_137_264 ();
 sg13g2_fill_8 FILLER_137_272 ();
 sg13g2_fill_8 FILLER_137_280 ();
 sg13g2_fill_8 FILLER_137_288 ();
 sg13g2_fill_8 FILLER_137_296 ();
 sg13g2_fill_8 FILLER_137_304 ();
 sg13g2_fill_8 FILLER_137_312 ();
 sg13g2_fill_8 FILLER_137_320 ();
 sg13g2_fill_8 FILLER_137_328 ();
 sg13g2_fill_8 FILLER_137_336 ();
 sg13g2_fill_8 FILLER_137_344 ();
 sg13g2_fill_8 FILLER_137_352 ();
 sg13g2_fill_8 FILLER_137_360 ();
 sg13g2_fill_8 FILLER_137_368 ();
 sg13g2_fill_8 FILLER_137_376 ();
 sg13g2_fill_8 FILLER_137_384 ();
 sg13g2_fill_8 FILLER_137_392 ();
 sg13g2_fill_8 FILLER_137_400 ();
 sg13g2_fill_8 FILLER_137_408 ();
 sg13g2_fill_8 FILLER_137_416 ();
 sg13g2_fill_8 FILLER_137_424 ();
 sg13g2_fill_8 FILLER_137_432 ();
 sg13g2_fill_8 FILLER_137_440 ();
 sg13g2_fill_8 FILLER_137_448 ();
 sg13g2_fill_8 FILLER_137_456 ();
 sg13g2_fill_8 FILLER_137_464 ();
 sg13g2_fill_8 FILLER_137_472 ();
 sg13g2_fill_8 FILLER_137_480 ();
 sg13g2_fill_8 FILLER_137_488 ();
 sg13g2_fill_8 FILLER_137_496 ();
 sg13g2_fill_8 FILLER_137_504 ();
 sg13g2_fill_8 FILLER_137_512 ();
 sg13g2_fill_8 FILLER_137_520 ();
 sg13g2_fill_8 FILLER_137_528 ();
 sg13g2_fill_8 FILLER_137_536 ();
 sg13g2_fill_8 FILLER_137_544 ();
 sg13g2_fill_8 FILLER_137_552 ();
 sg13g2_fill_8 FILLER_137_560 ();
 sg13g2_fill_8 FILLER_137_568 ();
 sg13g2_fill_8 FILLER_137_576 ();
 sg13g2_fill_8 FILLER_137_584 ();
 sg13g2_fill_8 FILLER_137_592 ();
 sg13g2_fill_8 FILLER_137_600 ();
 sg13g2_fill_8 FILLER_137_608 ();
 sg13g2_fill_8 FILLER_137_616 ();
 sg13g2_fill_8 FILLER_137_624 ();
 sg13g2_fill_8 FILLER_137_632 ();
 sg13g2_fill_8 FILLER_137_640 ();
 sg13g2_fill_8 FILLER_137_648 ();
 sg13g2_fill_8 FILLER_137_656 ();
 sg13g2_fill_8 FILLER_137_664 ();
 sg13g2_fill_8 FILLER_137_672 ();
 sg13g2_fill_8 FILLER_137_680 ();
 sg13g2_fill_8 FILLER_137_688 ();
 sg13g2_fill_8 FILLER_137_696 ();
 sg13g2_fill_8 FILLER_137_704 ();
 sg13g2_fill_8 FILLER_137_712 ();
 sg13g2_fill_8 FILLER_137_720 ();
 sg13g2_fill_8 FILLER_137_728 ();
 sg13g2_fill_8 FILLER_137_736 ();
 sg13g2_fill_8 FILLER_137_744 ();
 sg13g2_fill_8 FILLER_137_752 ();
 sg13g2_fill_8 FILLER_137_760 ();
 sg13g2_fill_8 FILLER_137_768 ();
 sg13g2_fill_8 FILLER_137_776 ();
 sg13g2_fill_8 FILLER_137_784 ();
 sg13g2_fill_8 FILLER_137_792 ();
 sg13g2_fill_8 FILLER_137_800 ();
 sg13g2_fill_8 FILLER_137_808 ();
 sg13g2_fill_8 FILLER_137_816 ();
 sg13g2_fill_8 FILLER_137_824 ();
 sg13g2_fill_8 FILLER_137_832 ();
 sg13g2_fill_8 FILLER_137_840 ();
 sg13g2_fill_8 FILLER_137_848 ();
 sg13g2_fill_8 FILLER_137_856 ();
 sg13g2_fill_8 FILLER_137_864 ();
 sg13g2_fill_8 FILLER_137_872 ();
 sg13g2_fill_8 FILLER_137_880 ();
 sg13g2_fill_8 FILLER_137_888 ();
 sg13g2_fill_8 FILLER_137_896 ();
 sg13g2_fill_8 FILLER_137_904 ();
 sg13g2_fill_8 FILLER_137_912 ();
 sg13g2_fill_8 FILLER_137_920 ();
 sg13g2_fill_8 FILLER_137_928 ();
 sg13g2_fill_8 FILLER_137_936 ();
 sg13g2_fill_8 FILLER_137_944 ();
 sg13g2_fill_8 FILLER_137_952 ();
 sg13g2_fill_8 FILLER_137_960 ();
 sg13g2_fill_8 FILLER_137_968 ();
 sg13g2_fill_8 FILLER_137_976 ();
 sg13g2_fill_8 FILLER_137_984 ();
 sg13g2_fill_8 FILLER_137_992 ();
 sg13g2_fill_8 FILLER_137_1000 ();
 sg13g2_fill_8 FILLER_137_1008 ();
 sg13g2_fill_8 FILLER_137_1016 ();
 sg13g2_fill_8 FILLER_137_1024 ();
 sg13g2_fill_8 FILLER_137_1032 ();
 sg13g2_fill_8 FILLER_137_1040 ();
 sg13g2_fill_8 FILLER_137_1048 ();
 sg13g2_fill_8 FILLER_137_1056 ();
 sg13g2_fill_8 FILLER_137_1064 ();
 sg13g2_fill_8 FILLER_137_1072 ();
 sg13g2_fill_8 FILLER_137_1080 ();
 sg13g2_fill_8 FILLER_137_1088 ();
 sg13g2_fill_8 FILLER_137_1096 ();
 sg13g2_fill_8 FILLER_137_1104 ();
 sg13g2_fill_8 FILLER_137_1112 ();
 sg13g2_fill_8 FILLER_137_1120 ();
 sg13g2_fill_8 FILLER_137_1128 ();
 sg13g2_fill_8 FILLER_137_1136 ();
 sg13g2_fill_8 FILLER_137_1144 ();
 sg13g2_fill_8 FILLER_137_1152 ();
 sg13g2_fill_4 FILLER_137_1160 ();
 sg13g2_fill_2 FILLER_137_1164 ();
 sg13g2_fill_8 FILLER_138_0 ();
 sg13g2_fill_8 FILLER_138_8 ();
 sg13g2_fill_8 FILLER_138_16 ();
 sg13g2_fill_8 FILLER_138_24 ();
 sg13g2_fill_8 FILLER_138_32 ();
 sg13g2_fill_8 FILLER_138_40 ();
 sg13g2_fill_8 FILLER_138_48 ();
 sg13g2_fill_8 FILLER_138_56 ();
 sg13g2_fill_8 FILLER_138_64 ();
 sg13g2_fill_8 FILLER_138_72 ();
 sg13g2_fill_8 FILLER_138_80 ();
 sg13g2_fill_8 FILLER_138_88 ();
 sg13g2_fill_8 FILLER_138_96 ();
 sg13g2_fill_8 FILLER_138_104 ();
 sg13g2_fill_8 FILLER_138_112 ();
 sg13g2_fill_8 FILLER_138_120 ();
 sg13g2_fill_8 FILLER_138_128 ();
 sg13g2_fill_8 FILLER_138_136 ();
 sg13g2_fill_8 FILLER_138_144 ();
 sg13g2_fill_8 FILLER_138_152 ();
 sg13g2_fill_8 FILLER_138_160 ();
 sg13g2_fill_8 FILLER_138_168 ();
 sg13g2_fill_8 FILLER_138_176 ();
 sg13g2_fill_8 FILLER_138_184 ();
 sg13g2_fill_8 FILLER_138_192 ();
 sg13g2_fill_8 FILLER_138_200 ();
 sg13g2_fill_8 FILLER_138_208 ();
 sg13g2_fill_8 FILLER_138_216 ();
 sg13g2_fill_8 FILLER_138_224 ();
 sg13g2_fill_8 FILLER_138_232 ();
 sg13g2_fill_8 FILLER_138_240 ();
 sg13g2_fill_8 FILLER_138_248 ();
 sg13g2_fill_8 FILLER_138_256 ();
 sg13g2_fill_8 FILLER_138_264 ();
 sg13g2_fill_8 FILLER_138_272 ();
 sg13g2_fill_8 FILLER_138_280 ();
 sg13g2_fill_8 FILLER_138_288 ();
 sg13g2_fill_8 FILLER_138_296 ();
 sg13g2_fill_8 FILLER_138_304 ();
 sg13g2_fill_8 FILLER_138_312 ();
 sg13g2_fill_8 FILLER_138_320 ();
 sg13g2_fill_8 FILLER_138_328 ();
 sg13g2_fill_8 FILLER_138_336 ();
 sg13g2_fill_8 FILLER_138_344 ();
 sg13g2_fill_8 FILLER_138_352 ();
 sg13g2_fill_8 FILLER_138_360 ();
 sg13g2_fill_8 FILLER_138_368 ();
 sg13g2_fill_8 FILLER_138_376 ();
 sg13g2_fill_8 FILLER_138_384 ();
 sg13g2_fill_8 FILLER_138_392 ();
 sg13g2_fill_8 FILLER_138_400 ();
 sg13g2_fill_8 FILLER_138_408 ();
 sg13g2_fill_8 FILLER_138_416 ();
 sg13g2_fill_8 FILLER_138_424 ();
 sg13g2_fill_8 FILLER_138_432 ();
 sg13g2_fill_8 FILLER_138_440 ();
 sg13g2_fill_8 FILLER_138_448 ();
 sg13g2_fill_8 FILLER_138_456 ();
 sg13g2_fill_8 FILLER_138_464 ();
 sg13g2_fill_8 FILLER_138_472 ();
 sg13g2_fill_8 FILLER_138_480 ();
 sg13g2_fill_8 FILLER_138_488 ();
 sg13g2_fill_8 FILLER_138_496 ();
 sg13g2_fill_8 FILLER_138_504 ();
 sg13g2_fill_8 FILLER_138_512 ();
 sg13g2_fill_8 FILLER_138_520 ();
 sg13g2_fill_8 FILLER_138_528 ();
 sg13g2_fill_8 FILLER_138_536 ();
 sg13g2_fill_8 FILLER_138_544 ();
 sg13g2_fill_8 FILLER_138_552 ();
 sg13g2_fill_8 FILLER_138_560 ();
 sg13g2_fill_8 FILLER_138_568 ();
 sg13g2_fill_8 FILLER_138_576 ();
 sg13g2_fill_8 FILLER_138_584 ();
 sg13g2_fill_8 FILLER_138_592 ();
 sg13g2_fill_8 FILLER_138_600 ();
 sg13g2_fill_8 FILLER_138_608 ();
 sg13g2_fill_8 FILLER_138_616 ();
 sg13g2_fill_8 FILLER_138_624 ();
 sg13g2_fill_8 FILLER_138_632 ();
 sg13g2_fill_8 FILLER_138_640 ();
 sg13g2_fill_8 FILLER_138_648 ();
 sg13g2_fill_8 FILLER_138_656 ();
 sg13g2_fill_8 FILLER_138_664 ();
 sg13g2_fill_8 FILLER_138_672 ();
 sg13g2_fill_8 FILLER_138_680 ();
 sg13g2_fill_8 FILLER_138_688 ();
 sg13g2_fill_8 FILLER_138_696 ();
 sg13g2_fill_8 FILLER_138_704 ();
 sg13g2_fill_8 FILLER_138_712 ();
 sg13g2_fill_8 FILLER_138_720 ();
 sg13g2_fill_8 FILLER_138_728 ();
 sg13g2_fill_8 FILLER_138_736 ();
 sg13g2_fill_8 FILLER_138_744 ();
 sg13g2_fill_8 FILLER_138_752 ();
 sg13g2_fill_8 FILLER_138_760 ();
 sg13g2_fill_8 FILLER_138_768 ();
 sg13g2_fill_8 FILLER_138_776 ();
 sg13g2_fill_8 FILLER_138_784 ();
 sg13g2_fill_8 FILLER_138_792 ();
 sg13g2_fill_8 FILLER_138_800 ();
 sg13g2_fill_8 FILLER_138_808 ();
 sg13g2_fill_8 FILLER_138_816 ();
 sg13g2_fill_8 FILLER_138_824 ();
 sg13g2_fill_8 FILLER_138_832 ();
 sg13g2_fill_8 FILLER_138_840 ();
 sg13g2_fill_8 FILLER_138_848 ();
 sg13g2_fill_8 FILLER_138_856 ();
 sg13g2_fill_8 FILLER_138_864 ();
 sg13g2_fill_8 FILLER_138_872 ();
 sg13g2_fill_8 FILLER_138_880 ();
 sg13g2_fill_8 FILLER_138_888 ();
 sg13g2_fill_8 FILLER_138_896 ();
 sg13g2_fill_8 FILLER_138_904 ();
 sg13g2_fill_8 FILLER_138_912 ();
 sg13g2_fill_8 FILLER_138_920 ();
 sg13g2_fill_8 FILLER_138_928 ();
 sg13g2_fill_8 FILLER_138_936 ();
 sg13g2_fill_8 FILLER_138_944 ();
 sg13g2_fill_8 FILLER_138_952 ();
 sg13g2_fill_8 FILLER_138_960 ();
 sg13g2_fill_8 FILLER_138_968 ();
 sg13g2_fill_8 FILLER_138_976 ();
 sg13g2_fill_8 FILLER_138_984 ();
 sg13g2_fill_8 FILLER_138_992 ();
 sg13g2_fill_8 FILLER_138_1000 ();
 sg13g2_fill_8 FILLER_138_1008 ();
 sg13g2_fill_8 FILLER_138_1016 ();
 sg13g2_fill_8 FILLER_138_1024 ();
 sg13g2_fill_8 FILLER_138_1032 ();
 sg13g2_fill_8 FILLER_138_1040 ();
 sg13g2_fill_8 FILLER_138_1048 ();
 sg13g2_fill_8 FILLER_138_1056 ();
 sg13g2_fill_8 FILLER_138_1064 ();
 sg13g2_fill_8 FILLER_138_1072 ();
 sg13g2_fill_8 FILLER_138_1080 ();
 sg13g2_fill_8 FILLER_138_1088 ();
 sg13g2_fill_8 FILLER_138_1096 ();
 sg13g2_fill_8 FILLER_138_1104 ();
 sg13g2_fill_8 FILLER_138_1112 ();
 sg13g2_fill_8 FILLER_138_1120 ();
 sg13g2_fill_8 FILLER_138_1128 ();
 sg13g2_fill_8 FILLER_138_1136 ();
 sg13g2_fill_8 FILLER_138_1144 ();
 sg13g2_fill_8 FILLER_138_1152 ();
 sg13g2_fill_4 FILLER_138_1160 ();
 sg13g2_fill_2 FILLER_138_1164 ();
 sg13g2_fill_8 FILLER_139_0 ();
 sg13g2_fill_8 FILLER_139_8 ();
 sg13g2_fill_8 FILLER_139_16 ();
 sg13g2_fill_8 FILLER_139_24 ();
 sg13g2_fill_8 FILLER_139_32 ();
 sg13g2_fill_8 FILLER_139_40 ();
 sg13g2_fill_8 FILLER_139_48 ();
 sg13g2_fill_8 FILLER_139_56 ();
 sg13g2_fill_8 FILLER_139_64 ();
 sg13g2_fill_8 FILLER_139_72 ();
 sg13g2_fill_8 FILLER_139_80 ();
 sg13g2_fill_8 FILLER_139_88 ();
 sg13g2_fill_8 FILLER_139_96 ();
 sg13g2_fill_8 FILLER_139_104 ();
 sg13g2_fill_8 FILLER_139_112 ();
 sg13g2_fill_8 FILLER_139_120 ();
 sg13g2_fill_8 FILLER_139_128 ();
 sg13g2_fill_8 FILLER_139_136 ();
 sg13g2_fill_8 FILLER_139_144 ();
 sg13g2_fill_8 FILLER_139_152 ();
 sg13g2_fill_8 FILLER_139_160 ();
 sg13g2_fill_8 FILLER_139_168 ();
 sg13g2_fill_8 FILLER_139_176 ();
 sg13g2_fill_8 FILLER_139_184 ();
 sg13g2_fill_8 FILLER_139_192 ();
 sg13g2_fill_8 FILLER_139_200 ();
 sg13g2_fill_8 FILLER_139_208 ();
 sg13g2_fill_8 FILLER_139_216 ();
 sg13g2_fill_8 FILLER_139_224 ();
 sg13g2_fill_8 FILLER_139_232 ();
 sg13g2_fill_8 FILLER_139_240 ();
 sg13g2_fill_8 FILLER_139_248 ();
 sg13g2_fill_8 FILLER_139_256 ();
 sg13g2_fill_8 FILLER_139_264 ();
 sg13g2_fill_8 FILLER_139_272 ();
 sg13g2_fill_8 FILLER_139_280 ();
 sg13g2_fill_8 FILLER_139_288 ();
 sg13g2_fill_8 FILLER_139_296 ();
 sg13g2_fill_8 FILLER_139_304 ();
 sg13g2_fill_8 FILLER_139_312 ();
 sg13g2_fill_8 FILLER_139_320 ();
 sg13g2_fill_8 FILLER_139_328 ();
 sg13g2_fill_8 FILLER_139_336 ();
 sg13g2_fill_8 FILLER_139_344 ();
 sg13g2_fill_8 FILLER_139_352 ();
 sg13g2_fill_8 FILLER_139_360 ();
 sg13g2_fill_8 FILLER_139_368 ();
 sg13g2_fill_8 FILLER_139_376 ();
 sg13g2_fill_8 FILLER_139_384 ();
 sg13g2_fill_8 FILLER_139_392 ();
 sg13g2_fill_8 FILLER_139_400 ();
 sg13g2_fill_8 FILLER_139_408 ();
 sg13g2_fill_8 FILLER_139_416 ();
 sg13g2_fill_8 FILLER_139_424 ();
 sg13g2_fill_8 FILLER_139_432 ();
 sg13g2_fill_8 FILLER_139_440 ();
 sg13g2_fill_8 FILLER_139_448 ();
 sg13g2_fill_8 FILLER_139_456 ();
 sg13g2_fill_8 FILLER_139_464 ();
 sg13g2_fill_8 FILLER_139_472 ();
 sg13g2_fill_8 FILLER_139_480 ();
 sg13g2_fill_8 FILLER_139_488 ();
 sg13g2_fill_8 FILLER_139_496 ();
 sg13g2_fill_8 FILLER_139_504 ();
 sg13g2_fill_8 FILLER_139_512 ();
 sg13g2_fill_8 FILLER_139_520 ();
 sg13g2_fill_8 FILLER_139_528 ();
 sg13g2_fill_8 FILLER_139_536 ();
 sg13g2_fill_8 FILLER_139_544 ();
 sg13g2_fill_8 FILLER_139_552 ();
 sg13g2_fill_8 FILLER_139_560 ();
 sg13g2_fill_8 FILLER_139_568 ();
 sg13g2_fill_8 FILLER_139_576 ();
 sg13g2_fill_8 FILLER_139_584 ();
 sg13g2_fill_8 FILLER_139_592 ();
 sg13g2_fill_8 FILLER_139_600 ();
 sg13g2_fill_8 FILLER_139_608 ();
 sg13g2_fill_8 FILLER_139_616 ();
 sg13g2_fill_8 FILLER_139_624 ();
 sg13g2_fill_8 FILLER_139_632 ();
 sg13g2_fill_8 FILLER_139_640 ();
 sg13g2_fill_8 FILLER_139_648 ();
 sg13g2_fill_8 FILLER_139_656 ();
 sg13g2_fill_8 FILLER_139_664 ();
 sg13g2_fill_8 FILLER_139_672 ();
 sg13g2_fill_8 FILLER_139_680 ();
 sg13g2_fill_8 FILLER_139_688 ();
 sg13g2_fill_8 FILLER_139_696 ();
 sg13g2_fill_8 FILLER_139_704 ();
 sg13g2_fill_8 FILLER_139_712 ();
 sg13g2_fill_8 FILLER_139_720 ();
 sg13g2_fill_8 FILLER_139_728 ();
 sg13g2_fill_8 FILLER_139_736 ();
 sg13g2_fill_8 FILLER_139_744 ();
 sg13g2_fill_8 FILLER_139_752 ();
 sg13g2_fill_8 FILLER_139_760 ();
 sg13g2_fill_8 FILLER_139_768 ();
 sg13g2_fill_8 FILLER_139_776 ();
 sg13g2_fill_8 FILLER_139_784 ();
 sg13g2_fill_8 FILLER_139_792 ();
 sg13g2_fill_8 FILLER_139_800 ();
 sg13g2_fill_8 FILLER_139_808 ();
 sg13g2_fill_8 FILLER_139_816 ();
 sg13g2_fill_8 FILLER_139_824 ();
 sg13g2_fill_8 FILLER_139_832 ();
 sg13g2_fill_8 FILLER_139_840 ();
 sg13g2_fill_8 FILLER_139_848 ();
 sg13g2_fill_8 FILLER_139_856 ();
 sg13g2_fill_8 FILLER_139_864 ();
 sg13g2_fill_8 FILLER_139_872 ();
 sg13g2_fill_8 FILLER_139_880 ();
 sg13g2_fill_8 FILLER_139_888 ();
 sg13g2_fill_8 FILLER_139_896 ();
 sg13g2_fill_8 FILLER_139_904 ();
 sg13g2_fill_8 FILLER_139_912 ();
 sg13g2_fill_8 FILLER_139_920 ();
 sg13g2_fill_8 FILLER_139_928 ();
 sg13g2_fill_8 FILLER_139_936 ();
 sg13g2_fill_8 FILLER_139_944 ();
 sg13g2_fill_8 FILLER_139_952 ();
 sg13g2_fill_8 FILLER_139_960 ();
 sg13g2_fill_8 FILLER_139_968 ();
 sg13g2_fill_8 FILLER_139_976 ();
 sg13g2_fill_8 FILLER_139_984 ();
 sg13g2_fill_8 FILLER_139_992 ();
 sg13g2_fill_8 FILLER_139_1000 ();
 sg13g2_fill_8 FILLER_139_1008 ();
 sg13g2_fill_8 FILLER_139_1016 ();
 sg13g2_fill_8 FILLER_139_1024 ();
 sg13g2_fill_8 FILLER_139_1032 ();
 sg13g2_fill_8 FILLER_139_1040 ();
 sg13g2_fill_8 FILLER_139_1048 ();
 sg13g2_fill_8 FILLER_139_1056 ();
 sg13g2_fill_8 FILLER_139_1064 ();
 sg13g2_fill_8 FILLER_139_1072 ();
 sg13g2_fill_8 FILLER_139_1080 ();
 sg13g2_fill_8 FILLER_139_1088 ();
 sg13g2_fill_8 FILLER_139_1096 ();
 sg13g2_fill_8 FILLER_139_1104 ();
 sg13g2_fill_8 FILLER_139_1112 ();
 sg13g2_fill_8 FILLER_139_1120 ();
 sg13g2_fill_8 FILLER_139_1128 ();
 sg13g2_fill_8 FILLER_139_1136 ();
 sg13g2_fill_8 FILLER_139_1144 ();
 sg13g2_fill_8 FILLER_139_1152 ();
 sg13g2_fill_4 FILLER_139_1160 ();
 sg13g2_fill_2 FILLER_139_1164 ();
 sg13g2_fill_8 FILLER_140_0 ();
 sg13g2_fill_8 FILLER_140_8 ();
 sg13g2_fill_8 FILLER_140_16 ();
 sg13g2_fill_8 FILLER_140_24 ();
 sg13g2_fill_8 FILLER_140_32 ();
 sg13g2_fill_8 FILLER_140_40 ();
 sg13g2_fill_8 FILLER_140_48 ();
 sg13g2_fill_8 FILLER_140_56 ();
 sg13g2_fill_8 FILLER_140_64 ();
 sg13g2_fill_8 FILLER_140_72 ();
 sg13g2_fill_8 FILLER_140_80 ();
 sg13g2_fill_8 FILLER_140_88 ();
 sg13g2_fill_8 FILLER_140_96 ();
 sg13g2_fill_8 FILLER_140_104 ();
 sg13g2_fill_8 FILLER_140_112 ();
 sg13g2_fill_8 FILLER_140_120 ();
 sg13g2_fill_8 FILLER_140_128 ();
 sg13g2_fill_8 FILLER_140_136 ();
 sg13g2_fill_8 FILLER_140_144 ();
 sg13g2_fill_8 FILLER_140_152 ();
 sg13g2_fill_8 FILLER_140_160 ();
 sg13g2_fill_8 FILLER_140_168 ();
 sg13g2_fill_8 FILLER_140_176 ();
 sg13g2_fill_8 FILLER_140_184 ();
 sg13g2_fill_8 FILLER_140_192 ();
 sg13g2_fill_8 FILLER_140_200 ();
 sg13g2_fill_8 FILLER_140_208 ();
 sg13g2_fill_8 FILLER_140_216 ();
 sg13g2_fill_8 FILLER_140_224 ();
 sg13g2_fill_8 FILLER_140_232 ();
 sg13g2_fill_8 FILLER_140_240 ();
 sg13g2_fill_8 FILLER_140_248 ();
 sg13g2_fill_8 FILLER_140_256 ();
 sg13g2_fill_8 FILLER_140_264 ();
 sg13g2_fill_8 FILLER_140_272 ();
 sg13g2_fill_8 FILLER_140_280 ();
 sg13g2_fill_8 FILLER_140_288 ();
 sg13g2_fill_8 FILLER_140_296 ();
 sg13g2_fill_8 FILLER_140_304 ();
 sg13g2_fill_8 FILLER_140_312 ();
 sg13g2_fill_8 FILLER_140_320 ();
 sg13g2_fill_8 FILLER_140_328 ();
 sg13g2_fill_8 FILLER_140_336 ();
 sg13g2_fill_8 FILLER_140_344 ();
 sg13g2_fill_8 FILLER_140_352 ();
 sg13g2_fill_8 FILLER_140_360 ();
 sg13g2_fill_8 FILLER_140_368 ();
 sg13g2_fill_8 FILLER_140_376 ();
 sg13g2_fill_8 FILLER_140_384 ();
 sg13g2_fill_8 FILLER_140_392 ();
 sg13g2_fill_8 FILLER_140_400 ();
 sg13g2_fill_8 FILLER_140_408 ();
 sg13g2_fill_8 FILLER_140_416 ();
 sg13g2_fill_8 FILLER_140_424 ();
 sg13g2_fill_8 FILLER_140_432 ();
 sg13g2_fill_8 FILLER_140_440 ();
 sg13g2_fill_8 FILLER_140_448 ();
 sg13g2_fill_8 FILLER_140_456 ();
 sg13g2_fill_8 FILLER_140_464 ();
 sg13g2_fill_8 FILLER_140_472 ();
 sg13g2_fill_8 FILLER_140_480 ();
 sg13g2_fill_8 FILLER_140_488 ();
 sg13g2_fill_8 FILLER_140_496 ();
 sg13g2_fill_8 FILLER_140_504 ();
 sg13g2_fill_8 FILLER_140_512 ();
 sg13g2_fill_8 FILLER_140_520 ();
 sg13g2_fill_8 FILLER_140_528 ();
 sg13g2_fill_8 FILLER_140_536 ();
 sg13g2_fill_8 FILLER_140_544 ();
 sg13g2_fill_8 FILLER_140_552 ();
 sg13g2_fill_8 FILLER_140_560 ();
 sg13g2_fill_8 FILLER_140_568 ();
 sg13g2_fill_8 FILLER_140_576 ();
 sg13g2_fill_8 FILLER_140_584 ();
 sg13g2_fill_8 FILLER_140_592 ();
 sg13g2_fill_8 FILLER_140_600 ();
 sg13g2_fill_8 FILLER_140_608 ();
 sg13g2_fill_8 FILLER_140_616 ();
 sg13g2_fill_8 FILLER_140_624 ();
 sg13g2_fill_8 FILLER_140_632 ();
 sg13g2_fill_8 FILLER_140_640 ();
 sg13g2_fill_8 FILLER_140_648 ();
 sg13g2_fill_8 FILLER_140_656 ();
 sg13g2_fill_8 FILLER_140_664 ();
 sg13g2_fill_8 FILLER_140_672 ();
 sg13g2_fill_8 FILLER_140_680 ();
 sg13g2_fill_8 FILLER_140_688 ();
 sg13g2_fill_8 FILLER_140_696 ();
 sg13g2_fill_8 FILLER_140_704 ();
 sg13g2_fill_8 FILLER_140_712 ();
 sg13g2_fill_8 FILLER_140_720 ();
 sg13g2_fill_8 FILLER_140_728 ();
 sg13g2_fill_8 FILLER_140_736 ();
 sg13g2_fill_8 FILLER_140_744 ();
 sg13g2_fill_8 FILLER_140_752 ();
 sg13g2_fill_8 FILLER_140_760 ();
 sg13g2_fill_8 FILLER_140_768 ();
 sg13g2_fill_8 FILLER_140_776 ();
 sg13g2_fill_8 FILLER_140_784 ();
 sg13g2_fill_8 FILLER_140_792 ();
 sg13g2_fill_8 FILLER_140_800 ();
 sg13g2_fill_8 FILLER_140_808 ();
 sg13g2_fill_8 FILLER_140_816 ();
 sg13g2_fill_8 FILLER_140_824 ();
 sg13g2_fill_8 FILLER_140_832 ();
 sg13g2_fill_8 FILLER_140_840 ();
 sg13g2_fill_8 FILLER_140_848 ();
 sg13g2_fill_8 FILLER_140_856 ();
 sg13g2_fill_8 FILLER_140_864 ();
 sg13g2_fill_8 FILLER_140_872 ();
 sg13g2_fill_8 FILLER_140_880 ();
 sg13g2_fill_8 FILLER_140_888 ();
 sg13g2_fill_8 FILLER_140_896 ();
 sg13g2_fill_8 FILLER_140_904 ();
 sg13g2_fill_8 FILLER_140_912 ();
 sg13g2_fill_8 FILLER_140_920 ();
 sg13g2_fill_8 FILLER_140_928 ();
 sg13g2_fill_8 FILLER_140_936 ();
 sg13g2_fill_8 FILLER_140_944 ();
 sg13g2_fill_8 FILLER_140_952 ();
 sg13g2_fill_8 FILLER_140_960 ();
 sg13g2_fill_8 FILLER_140_968 ();
 sg13g2_fill_8 FILLER_140_976 ();
 sg13g2_fill_8 FILLER_140_984 ();
 sg13g2_fill_8 FILLER_140_992 ();
 sg13g2_fill_8 FILLER_140_1000 ();
 sg13g2_fill_8 FILLER_140_1008 ();
 sg13g2_fill_8 FILLER_140_1016 ();
 sg13g2_fill_8 FILLER_140_1024 ();
 sg13g2_fill_8 FILLER_140_1032 ();
 sg13g2_fill_8 FILLER_140_1040 ();
 sg13g2_fill_8 FILLER_140_1048 ();
 sg13g2_fill_8 FILLER_140_1056 ();
 sg13g2_fill_8 FILLER_140_1064 ();
 sg13g2_fill_8 FILLER_140_1072 ();
 sg13g2_fill_8 FILLER_140_1080 ();
 sg13g2_fill_8 FILLER_140_1088 ();
 sg13g2_fill_8 FILLER_140_1096 ();
 sg13g2_fill_8 FILLER_140_1104 ();
 sg13g2_fill_8 FILLER_140_1112 ();
 sg13g2_fill_8 FILLER_140_1120 ();
 sg13g2_fill_8 FILLER_140_1128 ();
 sg13g2_fill_8 FILLER_140_1136 ();
 sg13g2_fill_8 FILLER_140_1144 ();
 sg13g2_fill_8 FILLER_140_1152 ();
 sg13g2_fill_4 FILLER_140_1160 ();
 sg13g2_fill_2 FILLER_140_1164 ();
 sg13g2_fill_8 FILLER_141_0 ();
 sg13g2_fill_8 FILLER_141_8 ();
 sg13g2_fill_8 FILLER_141_16 ();
 sg13g2_fill_8 FILLER_141_24 ();
 sg13g2_fill_8 FILLER_141_32 ();
 sg13g2_fill_8 FILLER_141_40 ();
 sg13g2_fill_8 FILLER_141_48 ();
 sg13g2_fill_8 FILLER_141_56 ();
 sg13g2_fill_8 FILLER_141_64 ();
 sg13g2_fill_8 FILLER_141_72 ();
 sg13g2_fill_8 FILLER_141_80 ();
 sg13g2_fill_8 FILLER_141_88 ();
 sg13g2_fill_8 FILLER_141_96 ();
 sg13g2_fill_8 FILLER_141_104 ();
 sg13g2_fill_8 FILLER_141_112 ();
 sg13g2_fill_8 FILLER_141_120 ();
 sg13g2_fill_8 FILLER_141_128 ();
 sg13g2_fill_8 FILLER_141_136 ();
 sg13g2_fill_8 FILLER_141_144 ();
 sg13g2_fill_8 FILLER_141_152 ();
 sg13g2_fill_8 FILLER_141_160 ();
 sg13g2_fill_8 FILLER_141_168 ();
 sg13g2_fill_8 FILLER_141_176 ();
 sg13g2_fill_8 FILLER_141_184 ();
 sg13g2_fill_8 FILLER_141_192 ();
 sg13g2_fill_8 FILLER_141_200 ();
 sg13g2_fill_8 FILLER_141_208 ();
 sg13g2_fill_8 FILLER_141_216 ();
 sg13g2_fill_8 FILLER_141_224 ();
 sg13g2_fill_8 FILLER_141_232 ();
 sg13g2_fill_8 FILLER_141_240 ();
 sg13g2_fill_8 FILLER_141_248 ();
 sg13g2_fill_8 FILLER_141_256 ();
 sg13g2_fill_8 FILLER_141_264 ();
 sg13g2_fill_8 FILLER_141_272 ();
 sg13g2_fill_8 FILLER_141_280 ();
 sg13g2_fill_8 FILLER_141_288 ();
 sg13g2_fill_8 FILLER_141_296 ();
 sg13g2_fill_8 FILLER_141_304 ();
 sg13g2_fill_8 FILLER_141_312 ();
 sg13g2_fill_8 FILLER_141_320 ();
 sg13g2_fill_8 FILLER_141_328 ();
 sg13g2_fill_8 FILLER_141_336 ();
 sg13g2_fill_8 FILLER_141_344 ();
 sg13g2_fill_8 FILLER_141_352 ();
 sg13g2_fill_8 FILLER_141_360 ();
 sg13g2_fill_8 FILLER_141_368 ();
 sg13g2_fill_8 FILLER_141_376 ();
 sg13g2_fill_8 FILLER_141_384 ();
 sg13g2_fill_8 FILLER_141_392 ();
 sg13g2_fill_8 FILLER_141_400 ();
 sg13g2_fill_8 FILLER_141_408 ();
 sg13g2_fill_8 FILLER_141_416 ();
 sg13g2_fill_8 FILLER_141_424 ();
 sg13g2_fill_8 FILLER_141_432 ();
 sg13g2_fill_8 FILLER_141_440 ();
 sg13g2_fill_8 FILLER_141_448 ();
 sg13g2_fill_8 FILLER_141_456 ();
 sg13g2_fill_8 FILLER_141_464 ();
 sg13g2_fill_8 FILLER_141_472 ();
 sg13g2_fill_8 FILLER_141_480 ();
 sg13g2_fill_8 FILLER_141_488 ();
 sg13g2_fill_8 FILLER_141_496 ();
 sg13g2_fill_8 FILLER_141_504 ();
 sg13g2_fill_8 FILLER_141_512 ();
 sg13g2_fill_8 FILLER_141_520 ();
 sg13g2_fill_8 FILLER_141_528 ();
 sg13g2_fill_8 FILLER_141_536 ();
 sg13g2_fill_8 FILLER_141_544 ();
 sg13g2_fill_8 FILLER_141_552 ();
 sg13g2_fill_8 FILLER_141_560 ();
 sg13g2_fill_8 FILLER_141_568 ();
 sg13g2_fill_8 FILLER_141_576 ();
 sg13g2_fill_8 FILLER_141_584 ();
 sg13g2_fill_8 FILLER_141_592 ();
 sg13g2_fill_8 FILLER_141_600 ();
 sg13g2_fill_8 FILLER_141_608 ();
 sg13g2_fill_8 FILLER_141_616 ();
 sg13g2_fill_8 FILLER_141_624 ();
 sg13g2_fill_8 FILLER_141_632 ();
 sg13g2_fill_8 FILLER_141_640 ();
 sg13g2_fill_8 FILLER_141_648 ();
 sg13g2_fill_8 FILLER_141_656 ();
 sg13g2_fill_8 FILLER_141_664 ();
 sg13g2_fill_8 FILLER_141_672 ();
 sg13g2_fill_8 FILLER_141_680 ();
 sg13g2_fill_8 FILLER_141_688 ();
 sg13g2_fill_8 FILLER_141_696 ();
 sg13g2_fill_8 FILLER_141_704 ();
 sg13g2_fill_8 FILLER_141_712 ();
 sg13g2_fill_8 FILLER_141_720 ();
 sg13g2_fill_8 FILLER_141_728 ();
 sg13g2_fill_8 FILLER_141_736 ();
 sg13g2_fill_8 FILLER_141_744 ();
 sg13g2_fill_8 FILLER_141_752 ();
 sg13g2_fill_8 FILLER_141_760 ();
 sg13g2_fill_8 FILLER_141_768 ();
 sg13g2_fill_8 FILLER_141_776 ();
 sg13g2_fill_8 FILLER_141_784 ();
 sg13g2_fill_8 FILLER_141_792 ();
 sg13g2_fill_8 FILLER_141_800 ();
 sg13g2_fill_8 FILLER_141_808 ();
 sg13g2_fill_8 FILLER_141_816 ();
 sg13g2_fill_8 FILLER_141_824 ();
 sg13g2_fill_8 FILLER_141_832 ();
 sg13g2_fill_8 FILLER_141_840 ();
 sg13g2_fill_8 FILLER_141_848 ();
 sg13g2_fill_8 FILLER_141_856 ();
 sg13g2_fill_8 FILLER_141_864 ();
 sg13g2_fill_8 FILLER_141_872 ();
 sg13g2_fill_8 FILLER_141_880 ();
 sg13g2_fill_8 FILLER_141_888 ();
 sg13g2_fill_8 FILLER_141_896 ();
 sg13g2_fill_8 FILLER_141_904 ();
 sg13g2_fill_8 FILLER_141_912 ();
 sg13g2_fill_8 FILLER_141_920 ();
 sg13g2_fill_8 FILLER_141_928 ();
 sg13g2_fill_8 FILLER_141_936 ();
 sg13g2_fill_8 FILLER_141_944 ();
 sg13g2_fill_8 FILLER_141_952 ();
 sg13g2_fill_8 FILLER_141_960 ();
 sg13g2_fill_8 FILLER_141_968 ();
 sg13g2_fill_8 FILLER_141_976 ();
 sg13g2_fill_8 FILLER_141_984 ();
 sg13g2_fill_8 FILLER_141_992 ();
 sg13g2_fill_8 FILLER_141_1000 ();
 sg13g2_fill_8 FILLER_141_1008 ();
 sg13g2_fill_8 FILLER_141_1016 ();
 sg13g2_fill_8 FILLER_141_1024 ();
 sg13g2_fill_8 FILLER_141_1032 ();
 sg13g2_fill_8 FILLER_141_1040 ();
 sg13g2_fill_8 FILLER_141_1048 ();
 sg13g2_fill_8 FILLER_141_1056 ();
 sg13g2_fill_8 FILLER_141_1064 ();
 sg13g2_fill_8 FILLER_141_1072 ();
 sg13g2_fill_8 FILLER_141_1080 ();
 sg13g2_fill_8 FILLER_141_1088 ();
 sg13g2_fill_8 FILLER_141_1096 ();
 sg13g2_fill_8 FILLER_141_1104 ();
 sg13g2_fill_8 FILLER_141_1112 ();
 sg13g2_fill_8 FILLER_141_1120 ();
 sg13g2_fill_8 FILLER_141_1128 ();
 sg13g2_fill_8 FILLER_141_1136 ();
 sg13g2_fill_8 FILLER_141_1144 ();
 sg13g2_fill_8 FILLER_141_1152 ();
 sg13g2_fill_4 FILLER_141_1160 ();
 sg13g2_fill_2 FILLER_141_1164 ();
 sg13g2_fill_8 FILLER_142_0 ();
 sg13g2_fill_8 FILLER_142_8 ();
 sg13g2_fill_8 FILLER_142_16 ();
 sg13g2_fill_8 FILLER_142_24 ();
 sg13g2_fill_8 FILLER_142_32 ();
 sg13g2_fill_8 FILLER_142_40 ();
 sg13g2_fill_8 FILLER_142_48 ();
 sg13g2_fill_8 FILLER_142_56 ();
 sg13g2_fill_8 FILLER_142_64 ();
 sg13g2_fill_8 FILLER_142_72 ();
 sg13g2_fill_8 FILLER_142_80 ();
 sg13g2_fill_8 FILLER_142_88 ();
 sg13g2_fill_8 FILLER_142_96 ();
 sg13g2_fill_8 FILLER_142_104 ();
 sg13g2_fill_8 FILLER_142_112 ();
 sg13g2_fill_8 FILLER_142_120 ();
 sg13g2_fill_8 FILLER_142_128 ();
 sg13g2_fill_8 FILLER_142_136 ();
 sg13g2_fill_8 FILLER_142_144 ();
 sg13g2_fill_8 FILLER_142_152 ();
 sg13g2_fill_8 FILLER_142_160 ();
 sg13g2_fill_8 FILLER_142_168 ();
 sg13g2_fill_8 FILLER_142_176 ();
 sg13g2_fill_8 FILLER_142_184 ();
 sg13g2_fill_8 FILLER_142_192 ();
 sg13g2_fill_8 FILLER_142_200 ();
 sg13g2_fill_8 FILLER_142_208 ();
 sg13g2_fill_8 FILLER_142_216 ();
 sg13g2_fill_8 FILLER_142_224 ();
 sg13g2_fill_8 FILLER_142_232 ();
 sg13g2_fill_8 FILLER_142_240 ();
 sg13g2_fill_8 FILLER_142_248 ();
 sg13g2_fill_8 FILLER_142_256 ();
 sg13g2_fill_8 FILLER_142_264 ();
 sg13g2_fill_8 FILLER_142_272 ();
 sg13g2_fill_8 FILLER_142_280 ();
 sg13g2_fill_8 FILLER_142_288 ();
 sg13g2_fill_8 FILLER_142_296 ();
 sg13g2_fill_8 FILLER_142_304 ();
 sg13g2_fill_8 FILLER_142_312 ();
 sg13g2_fill_8 FILLER_142_320 ();
 sg13g2_fill_8 FILLER_142_328 ();
 sg13g2_fill_8 FILLER_142_336 ();
 sg13g2_fill_8 FILLER_142_344 ();
 sg13g2_fill_8 FILLER_142_352 ();
 sg13g2_fill_8 FILLER_142_360 ();
 sg13g2_fill_8 FILLER_142_368 ();
 sg13g2_fill_8 FILLER_142_376 ();
 sg13g2_fill_8 FILLER_142_384 ();
 sg13g2_fill_8 FILLER_142_392 ();
 sg13g2_fill_8 FILLER_142_400 ();
 sg13g2_fill_8 FILLER_142_408 ();
 sg13g2_fill_8 FILLER_142_416 ();
 sg13g2_fill_8 FILLER_142_424 ();
 sg13g2_fill_8 FILLER_142_432 ();
 sg13g2_fill_8 FILLER_142_440 ();
 sg13g2_fill_8 FILLER_142_448 ();
 sg13g2_fill_8 FILLER_142_456 ();
 sg13g2_fill_8 FILLER_142_464 ();
 sg13g2_fill_8 FILLER_142_472 ();
 sg13g2_fill_8 FILLER_142_480 ();
 sg13g2_fill_8 FILLER_142_488 ();
 sg13g2_fill_8 FILLER_142_496 ();
 sg13g2_fill_8 FILLER_142_504 ();
 sg13g2_fill_8 FILLER_142_512 ();
 sg13g2_fill_8 FILLER_142_520 ();
 sg13g2_fill_8 FILLER_142_528 ();
 sg13g2_fill_8 FILLER_142_536 ();
 sg13g2_fill_8 FILLER_142_544 ();
 sg13g2_fill_8 FILLER_142_552 ();
 sg13g2_fill_8 FILLER_142_560 ();
 sg13g2_fill_8 FILLER_142_568 ();
 sg13g2_fill_8 FILLER_142_576 ();
 sg13g2_fill_8 FILLER_142_584 ();
 sg13g2_fill_8 FILLER_142_592 ();
 sg13g2_fill_8 FILLER_142_600 ();
 sg13g2_fill_8 FILLER_142_608 ();
 sg13g2_fill_8 FILLER_142_616 ();
 sg13g2_fill_8 FILLER_142_624 ();
 sg13g2_fill_8 FILLER_142_632 ();
 sg13g2_fill_8 FILLER_142_640 ();
 sg13g2_fill_8 FILLER_142_648 ();
 sg13g2_fill_8 FILLER_142_656 ();
 sg13g2_fill_8 FILLER_142_664 ();
 sg13g2_fill_8 FILLER_142_672 ();
 sg13g2_fill_8 FILLER_142_680 ();
 sg13g2_fill_8 FILLER_142_688 ();
 sg13g2_fill_8 FILLER_142_696 ();
 sg13g2_fill_8 FILLER_142_704 ();
 sg13g2_fill_8 FILLER_142_712 ();
 sg13g2_fill_8 FILLER_142_720 ();
 sg13g2_fill_8 FILLER_142_728 ();
 sg13g2_fill_8 FILLER_142_736 ();
 sg13g2_fill_8 FILLER_142_744 ();
 sg13g2_fill_8 FILLER_142_752 ();
 sg13g2_fill_8 FILLER_142_760 ();
 sg13g2_fill_8 FILLER_142_768 ();
 sg13g2_fill_8 FILLER_142_776 ();
 sg13g2_fill_8 FILLER_142_784 ();
 sg13g2_fill_8 FILLER_142_792 ();
 sg13g2_fill_8 FILLER_142_800 ();
 sg13g2_fill_8 FILLER_142_808 ();
 sg13g2_fill_8 FILLER_142_816 ();
 sg13g2_fill_8 FILLER_142_824 ();
 sg13g2_fill_8 FILLER_142_832 ();
 sg13g2_fill_8 FILLER_142_840 ();
 sg13g2_fill_8 FILLER_142_848 ();
 sg13g2_fill_8 FILLER_142_856 ();
 sg13g2_fill_8 FILLER_142_864 ();
 sg13g2_fill_8 FILLER_142_872 ();
 sg13g2_fill_8 FILLER_142_880 ();
 sg13g2_fill_8 FILLER_142_888 ();
 sg13g2_fill_8 FILLER_142_896 ();
 sg13g2_fill_8 FILLER_142_904 ();
 sg13g2_fill_8 FILLER_142_912 ();
 sg13g2_fill_8 FILLER_142_920 ();
 sg13g2_fill_8 FILLER_142_928 ();
 sg13g2_fill_8 FILLER_142_936 ();
 sg13g2_fill_8 FILLER_142_944 ();
 sg13g2_fill_8 FILLER_142_952 ();
 sg13g2_fill_8 FILLER_142_960 ();
 sg13g2_fill_8 FILLER_142_968 ();
 sg13g2_fill_8 FILLER_142_976 ();
 sg13g2_fill_8 FILLER_142_984 ();
 sg13g2_fill_8 FILLER_142_992 ();
 sg13g2_fill_8 FILLER_142_1000 ();
 sg13g2_fill_8 FILLER_142_1008 ();
 sg13g2_fill_8 FILLER_142_1016 ();
 sg13g2_fill_8 FILLER_142_1024 ();
 sg13g2_fill_8 FILLER_142_1032 ();
 sg13g2_fill_8 FILLER_142_1040 ();
 sg13g2_fill_8 FILLER_142_1048 ();
 sg13g2_fill_8 FILLER_142_1056 ();
 sg13g2_fill_8 FILLER_142_1064 ();
 sg13g2_fill_8 FILLER_142_1072 ();
 sg13g2_fill_8 FILLER_142_1080 ();
 sg13g2_fill_8 FILLER_142_1088 ();
 sg13g2_fill_8 FILLER_142_1096 ();
 sg13g2_fill_8 FILLER_142_1104 ();
 sg13g2_fill_8 FILLER_142_1112 ();
 sg13g2_fill_8 FILLER_142_1120 ();
 sg13g2_fill_8 FILLER_142_1128 ();
 sg13g2_fill_8 FILLER_142_1136 ();
 sg13g2_fill_8 FILLER_142_1144 ();
 sg13g2_fill_8 FILLER_142_1152 ();
 sg13g2_fill_4 FILLER_142_1160 ();
 sg13g2_fill_2 FILLER_142_1164 ();
 sg13g2_fill_8 FILLER_143_0 ();
 sg13g2_fill_8 FILLER_143_8 ();
 sg13g2_fill_8 FILLER_143_16 ();
 sg13g2_fill_8 FILLER_143_24 ();
 sg13g2_fill_8 FILLER_143_32 ();
 sg13g2_fill_8 FILLER_143_40 ();
 sg13g2_fill_8 FILLER_143_48 ();
 sg13g2_fill_8 FILLER_143_56 ();
 sg13g2_fill_8 FILLER_143_64 ();
 sg13g2_fill_8 FILLER_143_72 ();
 sg13g2_fill_8 FILLER_143_80 ();
 sg13g2_fill_8 FILLER_143_88 ();
 sg13g2_fill_8 FILLER_143_96 ();
 sg13g2_fill_8 FILLER_143_104 ();
 sg13g2_fill_8 FILLER_143_112 ();
 sg13g2_fill_8 FILLER_143_120 ();
 sg13g2_fill_8 FILLER_143_128 ();
 sg13g2_fill_8 FILLER_143_136 ();
 sg13g2_fill_8 FILLER_143_144 ();
 sg13g2_fill_8 FILLER_143_152 ();
 sg13g2_fill_8 FILLER_143_160 ();
 sg13g2_fill_8 FILLER_143_168 ();
 sg13g2_fill_8 FILLER_143_176 ();
 sg13g2_fill_8 FILLER_143_184 ();
 sg13g2_fill_8 FILLER_143_192 ();
 sg13g2_fill_8 FILLER_143_200 ();
 sg13g2_fill_8 FILLER_143_208 ();
 sg13g2_fill_8 FILLER_143_216 ();
 sg13g2_fill_8 FILLER_143_224 ();
 sg13g2_fill_8 FILLER_143_232 ();
 sg13g2_fill_8 FILLER_143_240 ();
 sg13g2_fill_8 FILLER_143_248 ();
 sg13g2_fill_8 FILLER_143_256 ();
 sg13g2_fill_8 FILLER_143_264 ();
 sg13g2_fill_8 FILLER_143_272 ();
 sg13g2_fill_8 FILLER_143_280 ();
 sg13g2_fill_8 FILLER_143_288 ();
 sg13g2_fill_8 FILLER_143_296 ();
 sg13g2_fill_8 FILLER_143_304 ();
 sg13g2_fill_8 FILLER_143_312 ();
 sg13g2_fill_8 FILLER_143_320 ();
 sg13g2_fill_8 FILLER_143_328 ();
 sg13g2_fill_8 FILLER_143_336 ();
 sg13g2_fill_8 FILLER_143_344 ();
 sg13g2_fill_8 FILLER_143_352 ();
 sg13g2_fill_8 FILLER_143_360 ();
 sg13g2_fill_8 FILLER_143_368 ();
 sg13g2_fill_8 FILLER_143_376 ();
 sg13g2_fill_8 FILLER_143_384 ();
 sg13g2_fill_8 FILLER_143_392 ();
 sg13g2_fill_8 FILLER_143_400 ();
 sg13g2_fill_8 FILLER_143_408 ();
 sg13g2_fill_8 FILLER_143_416 ();
 sg13g2_fill_8 FILLER_143_424 ();
 sg13g2_fill_8 FILLER_143_432 ();
 sg13g2_fill_8 FILLER_143_440 ();
 sg13g2_fill_8 FILLER_143_448 ();
 sg13g2_fill_8 FILLER_143_456 ();
 sg13g2_fill_8 FILLER_143_464 ();
 sg13g2_fill_8 FILLER_143_472 ();
 sg13g2_fill_8 FILLER_143_480 ();
 sg13g2_fill_8 FILLER_143_488 ();
 sg13g2_fill_8 FILLER_143_496 ();
 sg13g2_fill_8 FILLER_143_504 ();
 sg13g2_fill_8 FILLER_143_512 ();
 sg13g2_fill_8 FILLER_143_520 ();
 sg13g2_fill_8 FILLER_143_528 ();
 sg13g2_fill_8 FILLER_143_536 ();
 sg13g2_fill_8 FILLER_143_544 ();
 sg13g2_fill_8 FILLER_143_552 ();
 sg13g2_fill_8 FILLER_143_560 ();
 sg13g2_fill_8 FILLER_143_568 ();
 sg13g2_fill_8 FILLER_143_576 ();
 sg13g2_fill_8 FILLER_143_584 ();
 sg13g2_fill_8 FILLER_143_592 ();
 sg13g2_fill_8 FILLER_143_600 ();
 sg13g2_fill_8 FILLER_143_608 ();
 sg13g2_fill_8 FILLER_143_616 ();
 sg13g2_fill_8 FILLER_143_624 ();
 sg13g2_fill_8 FILLER_143_632 ();
 sg13g2_fill_8 FILLER_143_640 ();
 sg13g2_fill_8 FILLER_143_648 ();
 sg13g2_fill_8 FILLER_143_656 ();
 sg13g2_fill_8 FILLER_143_664 ();
 sg13g2_fill_8 FILLER_143_672 ();
 sg13g2_fill_8 FILLER_143_680 ();
 sg13g2_fill_8 FILLER_143_688 ();
 sg13g2_fill_8 FILLER_143_696 ();
 sg13g2_fill_8 FILLER_143_704 ();
 sg13g2_fill_8 FILLER_143_712 ();
 sg13g2_fill_8 FILLER_143_720 ();
 sg13g2_fill_8 FILLER_143_728 ();
 sg13g2_fill_8 FILLER_143_736 ();
 sg13g2_fill_8 FILLER_143_744 ();
 sg13g2_fill_8 FILLER_143_752 ();
 sg13g2_fill_8 FILLER_143_760 ();
 sg13g2_fill_8 FILLER_143_768 ();
 sg13g2_fill_8 FILLER_143_776 ();
 sg13g2_fill_8 FILLER_143_784 ();
 sg13g2_fill_8 FILLER_143_792 ();
 sg13g2_fill_8 FILLER_143_800 ();
 sg13g2_fill_8 FILLER_143_808 ();
 sg13g2_fill_8 FILLER_143_816 ();
 sg13g2_fill_8 FILLER_143_824 ();
 sg13g2_fill_8 FILLER_143_832 ();
 sg13g2_fill_8 FILLER_143_840 ();
 sg13g2_fill_8 FILLER_143_848 ();
 sg13g2_fill_8 FILLER_143_856 ();
 sg13g2_fill_8 FILLER_143_864 ();
 sg13g2_fill_8 FILLER_143_872 ();
 sg13g2_fill_8 FILLER_143_880 ();
 sg13g2_fill_8 FILLER_143_888 ();
 sg13g2_fill_8 FILLER_143_896 ();
 sg13g2_fill_8 FILLER_143_904 ();
 sg13g2_fill_8 FILLER_143_912 ();
 sg13g2_fill_8 FILLER_143_920 ();
 sg13g2_fill_8 FILLER_143_928 ();
 sg13g2_fill_8 FILLER_143_936 ();
 sg13g2_fill_8 FILLER_143_944 ();
 sg13g2_fill_8 FILLER_143_952 ();
 sg13g2_fill_8 FILLER_143_960 ();
 sg13g2_fill_8 FILLER_143_968 ();
 sg13g2_fill_8 FILLER_143_976 ();
 sg13g2_fill_8 FILLER_143_984 ();
 sg13g2_fill_8 FILLER_143_992 ();
 sg13g2_fill_8 FILLER_143_1000 ();
 sg13g2_fill_8 FILLER_143_1008 ();
 sg13g2_fill_8 FILLER_143_1016 ();
 sg13g2_fill_8 FILLER_143_1024 ();
 sg13g2_fill_8 FILLER_143_1032 ();
 sg13g2_fill_8 FILLER_143_1040 ();
 sg13g2_fill_8 FILLER_143_1048 ();
 sg13g2_fill_8 FILLER_143_1056 ();
 sg13g2_fill_8 FILLER_143_1064 ();
 sg13g2_fill_8 FILLER_143_1072 ();
 sg13g2_fill_8 FILLER_143_1080 ();
 sg13g2_fill_8 FILLER_143_1088 ();
 sg13g2_fill_8 FILLER_143_1096 ();
 sg13g2_fill_8 FILLER_143_1104 ();
 sg13g2_fill_8 FILLER_143_1112 ();
 sg13g2_fill_8 FILLER_143_1120 ();
 sg13g2_fill_8 FILLER_143_1128 ();
 sg13g2_fill_8 FILLER_143_1136 ();
 sg13g2_fill_8 FILLER_143_1144 ();
 sg13g2_fill_8 FILLER_143_1152 ();
 sg13g2_fill_4 FILLER_143_1160 ();
 sg13g2_fill_2 FILLER_143_1164 ();
 sg13g2_fill_8 FILLER_144_0 ();
 sg13g2_fill_8 FILLER_144_8 ();
 sg13g2_fill_8 FILLER_144_16 ();
 sg13g2_fill_8 FILLER_144_24 ();
 sg13g2_fill_8 FILLER_144_32 ();
 sg13g2_fill_8 FILLER_144_40 ();
 sg13g2_fill_8 FILLER_144_48 ();
 sg13g2_fill_8 FILLER_144_56 ();
 sg13g2_fill_8 FILLER_144_64 ();
 sg13g2_fill_8 FILLER_144_72 ();
 sg13g2_fill_8 FILLER_144_80 ();
 sg13g2_fill_8 FILLER_144_88 ();
 sg13g2_fill_8 FILLER_144_96 ();
 sg13g2_fill_8 FILLER_144_104 ();
 sg13g2_fill_8 FILLER_144_112 ();
 sg13g2_fill_8 FILLER_144_120 ();
 sg13g2_fill_8 FILLER_144_128 ();
 sg13g2_fill_8 FILLER_144_136 ();
 sg13g2_fill_8 FILLER_144_144 ();
 sg13g2_fill_8 FILLER_144_152 ();
 sg13g2_fill_8 FILLER_144_160 ();
 sg13g2_fill_8 FILLER_144_168 ();
 sg13g2_fill_8 FILLER_144_176 ();
 sg13g2_fill_8 FILLER_144_184 ();
 sg13g2_fill_8 FILLER_144_192 ();
 sg13g2_fill_8 FILLER_144_200 ();
 sg13g2_fill_8 FILLER_144_208 ();
 sg13g2_fill_8 FILLER_144_216 ();
 sg13g2_fill_8 FILLER_144_224 ();
 sg13g2_fill_8 FILLER_144_232 ();
 sg13g2_fill_8 FILLER_144_240 ();
 sg13g2_fill_8 FILLER_144_248 ();
 sg13g2_fill_8 FILLER_144_256 ();
 sg13g2_fill_8 FILLER_144_264 ();
 sg13g2_fill_8 FILLER_144_272 ();
 sg13g2_fill_8 FILLER_144_280 ();
 sg13g2_fill_8 FILLER_144_288 ();
 sg13g2_fill_8 FILLER_144_296 ();
 sg13g2_fill_8 FILLER_144_304 ();
 sg13g2_fill_8 FILLER_144_312 ();
 sg13g2_fill_8 FILLER_144_320 ();
 sg13g2_fill_8 FILLER_144_328 ();
 sg13g2_fill_8 FILLER_144_336 ();
 sg13g2_fill_8 FILLER_144_344 ();
 sg13g2_fill_8 FILLER_144_352 ();
 sg13g2_fill_8 FILLER_144_360 ();
 sg13g2_fill_8 FILLER_144_368 ();
 sg13g2_fill_8 FILLER_144_376 ();
 sg13g2_fill_8 FILLER_144_384 ();
 sg13g2_fill_8 FILLER_144_392 ();
 sg13g2_fill_8 FILLER_144_400 ();
 sg13g2_fill_8 FILLER_144_408 ();
 sg13g2_fill_8 FILLER_144_416 ();
 sg13g2_fill_8 FILLER_144_424 ();
 sg13g2_fill_8 FILLER_144_432 ();
 sg13g2_fill_8 FILLER_144_440 ();
 sg13g2_fill_8 FILLER_144_448 ();
 sg13g2_fill_8 FILLER_144_456 ();
 sg13g2_fill_8 FILLER_144_464 ();
 sg13g2_fill_8 FILLER_144_472 ();
 sg13g2_fill_8 FILLER_144_480 ();
 sg13g2_fill_8 FILLER_144_488 ();
 sg13g2_fill_8 FILLER_144_496 ();
 sg13g2_fill_8 FILLER_144_504 ();
 sg13g2_fill_8 FILLER_144_512 ();
 sg13g2_fill_8 FILLER_144_520 ();
 sg13g2_fill_8 FILLER_144_528 ();
 sg13g2_fill_8 FILLER_144_536 ();
 sg13g2_fill_8 FILLER_144_544 ();
 sg13g2_fill_8 FILLER_144_552 ();
 sg13g2_fill_8 FILLER_144_560 ();
 sg13g2_fill_8 FILLER_144_568 ();
 sg13g2_fill_8 FILLER_144_576 ();
 sg13g2_fill_8 FILLER_144_584 ();
 sg13g2_fill_8 FILLER_144_592 ();
 sg13g2_fill_8 FILLER_144_600 ();
 sg13g2_fill_8 FILLER_144_608 ();
 sg13g2_fill_8 FILLER_144_616 ();
 sg13g2_fill_8 FILLER_144_624 ();
 sg13g2_fill_8 FILLER_144_632 ();
 sg13g2_fill_8 FILLER_144_640 ();
 sg13g2_fill_8 FILLER_144_648 ();
 sg13g2_fill_8 FILLER_144_656 ();
 sg13g2_fill_8 FILLER_144_664 ();
 sg13g2_fill_8 FILLER_144_672 ();
 sg13g2_fill_8 FILLER_144_680 ();
 sg13g2_fill_8 FILLER_144_688 ();
 sg13g2_fill_8 FILLER_144_696 ();
 sg13g2_fill_8 FILLER_144_704 ();
 sg13g2_fill_8 FILLER_144_712 ();
 sg13g2_fill_8 FILLER_144_720 ();
 sg13g2_fill_8 FILLER_144_728 ();
 sg13g2_fill_8 FILLER_144_736 ();
 sg13g2_fill_8 FILLER_144_744 ();
 sg13g2_fill_8 FILLER_144_752 ();
 sg13g2_fill_8 FILLER_144_760 ();
 sg13g2_fill_8 FILLER_144_768 ();
 sg13g2_fill_8 FILLER_144_776 ();
 sg13g2_fill_8 FILLER_144_784 ();
 sg13g2_fill_8 FILLER_144_792 ();
 sg13g2_fill_8 FILLER_144_800 ();
 sg13g2_fill_8 FILLER_144_808 ();
 sg13g2_fill_8 FILLER_144_816 ();
 sg13g2_fill_8 FILLER_144_824 ();
 sg13g2_fill_8 FILLER_144_832 ();
 sg13g2_fill_8 FILLER_144_840 ();
 sg13g2_fill_8 FILLER_144_848 ();
 sg13g2_fill_8 FILLER_144_856 ();
 sg13g2_fill_8 FILLER_144_864 ();
 sg13g2_fill_8 FILLER_144_872 ();
 sg13g2_fill_8 FILLER_144_880 ();
 sg13g2_fill_8 FILLER_144_888 ();
 sg13g2_fill_8 FILLER_144_896 ();
 sg13g2_fill_8 FILLER_144_904 ();
 sg13g2_fill_8 FILLER_144_912 ();
 sg13g2_fill_8 FILLER_144_920 ();
 sg13g2_fill_8 FILLER_144_928 ();
 sg13g2_fill_8 FILLER_144_936 ();
 sg13g2_fill_8 FILLER_144_944 ();
 sg13g2_fill_8 FILLER_144_952 ();
 sg13g2_fill_8 FILLER_144_960 ();
 sg13g2_fill_8 FILLER_144_968 ();
 sg13g2_fill_8 FILLER_144_976 ();
 sg13g2_fill_8 FILLER_144_984 ();
 sg13g2_fill_8 FILLER_144_992 ();
 sg13g2_fill_8 FILLER_144_1000 ();
 sg13g2_fill_8 FILLER_144_1008 ();
 sg13g2_fill_8 FILLER_144_1016 ();
 sg13g2_fill_8 FILLER_144_1024 ();
 sg13g2_fill_8 FILLER_144_1032 ();
 sg13g2_fill_8 FILLER_144_1040 ();
 sg13g2_fill_8 FILLER_144_1048 ();
 sg13g2_fill_8 FILLER_144_1056 ();
 sg13g2_fill_8 FILLER_144_1064 ();
 sg13g2_fill_8 FILLER_144_1072 ();
 sg13g2_fill_8 FILLER_144_1080 ();
 sg13g2_fill_8 FILLER_144_1088 ();
 sg13g2_fill_8 FILLER_144_1096 ();
 sg13g2_fill_8 FILLER_144_1104 ();
 sg13g2_fill_8 FILLER_144_1112 ();
 sg13g2_fill_8 FILLER_144_1120 ();
 sg13g2_fill_8 FILLER_144_1128 ();
 sg13g2_fill_8 FILLER_144_1136 ();
 sg13g2_fill_8 FILLER_144_1144 ();
 sg13g2_fill_8 FILLER_144_1152 ();
 sg13g2_fill_4 FILLER_144_1160 ();
 sg13g2_fill_2 FILLER_144_1164 ();
 sg13g2_fill_8 FILLER_145_0 ();
 sg13g2_fill_8 FILLER_145_8 ();
 sg13g2_fill_8 FILLER_145_16 ();
 sg13g2_fill_8 FILLER_145_24 ();
 sg13g2_fill_8 FILLER_145_32 ();
 sg13g2_fill_8 FILLER_145_40 ();
 sg13g2_fill_8 FILLER_145_48 ();
 sg13g2_fill_8 FILLER_145_56 ();
 sg13g2_fill_8 FILLER_145_64 ();
 sg13g2_fill_8 FILLER_145_72 ();
 sg13g2_fill_8 FILLER_145_80 ();
 sg13g2_fill_8 FILLER_145_88 ();
 sg13g2_fill_8 FILLER_145_96 ();
 sg13g2_fill_8 FILLER_145_104 ();
 sg13g2_fill_8 FILLER_145_112 ();
 sg13g2_fill_8 FILLER_145_120 ();
 sg13g2_fill_8 FILLER_145_128 ();
 sg13g2_fill_8 FILLER_145_136 ();
 sg13g2_fill_8 FILLER_145_144 ();
 sg13g2_fill_8 FILLER_145_152 ();
 sg13g2_fill_8 FILLER_145_160 ();
 sg13g2_fill_8 FILLER_145_168 ();
 sg13g2_fill_8 FILLER_145_176 ();
 sg13g2_fill_8 FILLER_145_184 ();
 sg13g2_fill_8 FILLER_145_192 ();
 sg13g2_fill_8 FILLER_145_200 ();
 sg13g2_fill_8 FILLER_145_208 ();
 sg13g2_fill_8 FILLER_145_216 ();
 sg13g2_fill_8 FILLER_145_224 ();
 sg13g2_fill_8 FILLER_145_232 ();
 sg13g2_fill_8 FILLER_145_240 ();
 sg13g2_fill_8 FILLER_145_248 ();
 sg13g2_fill_8 FILLER_145_256 ();
 sg13g2_fill_8 FILLER_145_264 ();
 sg13g2_fill_8 FILLER_145_272 ();
 sg13g2_fill_8 FILLER_145_280 ();
 sg13g2_fill_8 FILLER_145_288 ();
 sg13g2_fill_8 FILLER_145_296 ();
 sg13g2_fill_8 FILLER_145_304 ();
 sg13g2_fill_8 FILLER_145_312 ();
 sg13g2_fill_8 FILLER_145_320 ();
 sg13g2_fill_8 FILLER_145_328 ();
 sg13g2_fill_8 FILLER_145_336 ();
 sg13g2_fill_8 FILLER_145_344 ();
 sg13g2_fill_8 FILLER_145_352 ();
 sg13g2_fill_8 FILLER_145_360 ();
 sg13g2_fill_8 FILLER_145_368 ();
 sg13g2_fill_8 FILLER_145_376 ();
 sg13g2_fill_8 FILLER_145_384 ();
 sg13g2_fill_8 FILLER_145_392 ();
 sg13g2_fill_8 FILLER_145_400 ();
 sg13g2_fill_8 FILLER_145_408 ();
 sg13g2_fill_8 FILLER_145_416 ();
 sg13g2_fill_8 FILLER_145_424 ();
 sg13g2_fill_8 FILLER_145_432 ();
 sg13g2_fill_8 FILLER_145_440 ();
 sg13g2_fill_8 FILLER_145_448 ();
 sg13g2_fill_8 FILLER_145_456 ();
 sg13g2_fill_8 FILLER_145_464 ();
 sg13g2_fill_8 FILLER_145_472 ();
 sg13g2_fill_8 FILLER_145_480 ();
 sg13g2_fill_8 FILLER_145_488 ();
 sg13g2_fill_8 FILLER_145_496 ();
 sg13g2_fill_8 FILLER_145_504 ();
 sg13g2_fill_8 FILLER_145_512 ();
 sg13g2_fill_8 FILLER_145_520 ();
 sg13g2_fill_8 FILLER_145_528 ();
 sg13g2_fill_8 FILLER_145_536 ();
 sg13g2_fill_8 FILLER_145_544 ();
 sg13g2_fill_8 FILLER_145_552 ();
 sg13g2_fill_8 FILLER_145_560 ();
 sg13g2_fill_8 FILLER_145_568 ();
 sg13g2_fill_8 FILLER_145_576 ();
 sg13g2_fill_8 FILLER_145_584 ();
 sg13g2_fill_8 FILLER_145_592 ();
 sg13g2_fill_8 FILLER_145_600 ();
 sg13g2_fill_8 FILLER_145_608 ();
 sg13g2_fill_8 FILLER_145_616 ();
 sg13g2_fill_8 FILLER_145_624 ();
 sg13g2_fill_8 FILLER_145_632 ();
 sg13g2_fill_8 FILLER_145_640 ();
 sg13g2_fill_8 FILLER_145_648 ();
 sg13g2_fill_8 FILLER_145_656 ();
 sg13g2_fill_8 FILLER_145_664 ();
 sg13g2_fill_8 FILLER_145_672 ();
 sg13g2_fill_8 FILLER_145_680 ();
 sg13g2_fill_8 FILLER_145_688 ();
 sg13g2_fill_8 FILLER_145_696 ();
 sg13g2_fill_8 FILLER_145_704 ();
 sg13g2_fill_8 FILLER_145_712 ();
 sg13g2_fill_8 FILLER_145_720 ();
 sg13g2_fill_8 FILLER_145_728 ();
 sg13g2_fill_8 FILLER_145_736 ();
 sg13g2_fill_8 FILLER_145_744 ();
 sg13g2_fill_8 FILLER_145_752 ();
 sg13g2_fill_8 FILLER_145_760 ();
 sg13g2_fill_8 FILLER_145_768 ();
 sg13g2_fill_8 FILLER_145_776 ();
 sg13g2_fill_8 FILLER_145_784 ();
 sg13g2_fill_8 FILLER_145_792 ();
 sg13g2_fill_8 FILLER_145_800 ();
 sg13g2_fill_8 FILLER_145_808 ();
 sg13g2_fill_8 FILLER_145_816 ();
 sg13g2_fill_8 FILLER_145_824 ();
 sg13g2_fill_8 FILLER_145_832 ();
 sg13g2_fill_8 FILLER_145_840 ();
 sg13g2_fill_8 FILLER_145_848 ();
 sg13g2_fill_8 FILLER_145_856 ();
 sg13g2_fill_8 FILLER_145_864 ();
 sg13g2_fill_8 FILLER_145_872 ();
 sg13g2_fill_8 FILLER_145_880 ();
 sg13g2_fill_8 FILLER_145_888 ();
 sg13g2_fill_8 FILLER_145_896 ();
 sg13g2_fill_8 FILLER_145_904 ();
 sg13g2_fill_8 FILLER_145_912 ();
 sg13g2_fill_8 FILLER_145_920 ();
 sg13g2_fill_8 FILLER_145_928 ();
 sg13g2_fill_8 FILLER_145_936 ();
 sg13g2_fill_8 FILLER_145_944 ();
 sg13g2_fill_8 FILLER_145_952 ();
 sg13g2_fill_8 FILLER_145_960 ();
 sg13g2_fill_8 FILLER_145_968 ();
 sg13g2_fill_8 FILLER_145_976 ();
 sg13g2_fill_8 FILLER_145_984 ();
 sg13g2_fill_8 FILLER_145_992 ();
 sg13g2_fill_8 FILLER_145_1000 ();
 sg13g2_fill_8 FILLER_145_1008 ();
 sg13g2_fill_8 FILLER_145_1016 ();
 sg13g2_fill_8 FILLER_145_1024 ();
 sg13g2_fill_8 FILLER_145_1032 ();
 sg13g2_fill_8 FILLER_145_1040 ();
 sg13g2_fill_8 FILLER_145_1048 ();
 sg13g2_fill_8 FILLER_145_1056 ();
 sg13g2_fill_8 FILLER_145_1064 ();
 sg13g2_fill_8 FILLER_145_1072 ();
 sg13g2_fill_8 FILLER_145_1080 ();
 sg13g2_fill_8 FILLER_145_1088 ();
 sg13g2_fill_8 FILLER_145_1096 ();
 sg13g2_fill_8 FILLER_145_1104 ();
 sg13g2_fill_8 FILLER_145_1112 ();
 sg13g2_fill_8 FILLER_145_1120 ();
 sg13g2_fill_8 FILLER_145_1128 ();
 sg13g2_fill_8 FILLER_145_1136 ();
 sg13g2_fill_8 FILLER_145_1144 ();
 sg13g2_fill_8 FILLER_145_1152 ();
 sg13g2_fill_4 FILLER_145_1160 ();
 sg13g2_fill_2 FILLER_145_1164 ();
 sg13g2_fill_8 FILLER_146_0 ();
 sg13g2_fill_8 FILLER_146_8 ();
 sg13g2_fill_8 FILLER_146_16 ();
 sg13g2_fill_8 FILLER_146_24 ();
 sg13g2_fill_8 FILLER_146_32 ();
 sg13g2_fill_8 FILLER_146_40 ();
 sg13g2_fill_8 FILLER_146_48 ();
 sg13g2_fill_8 FILLER_146_56 ();
 sg13g2_fill_8 FILLER_146_64 ();
 sg13g2_fill_8 FILLER_146_72 ();
 sg13g2_fill_8 FILLER_146_80 ();
 sg13g2_fill_8 FILLER_146_88 ();
 sg13g2_fill_8 FILLER_146_96 ();
 sg13g2_fill_8 FILLER_146_104 ();
 sg13g2_fill_8 FILLER_146_112 ();
 sg13g2_fill_8 FILLER_146_120 ();
 sg13g2_fill_8 FILLER_146_128 ();
 sg13g2_fill_8 FILLER_146_136 ();
 sg13g2_fill_8 FILLER_146_144 ();
 sg13g2_fill_8 FILLER_146_152 ();
 sg13g2_fill_8 FILLER_146_160 ();
 sg13g2_fill_8 FILLER_146_168 ();
 sg13g2_fill_8 FILLER_146_176 ();
 sg13g2_fill_8 FILLER_146_184 ();
 sg13g2_fill_8 FILLER_146_192 ();
 sg13g2_fill_8 FILLER_146_200 ();
 sg13g2_fill_8 FILLER_146_208 ();
 sg13g2_fill_8 FILLER_146_216 ();
 sg13g2_fill_8 FILLER_146_224 ();
 sg13g2_fill_8 FILLER_146_232 ();
 sg13g2_fill_8 FILLER_146_240 ();
 sg13g2_fill_8 FILLER_146_248 ();
 sg13g2_fill_8 FILLER_146_256 ();
 sg13g2_fill_8 FILLER_146_264 ();
 sg13g2_fill_8 FILLER_146_272 ();
 sg13g2_fill_8 FILLER_146_280 ();
 sg13g2_fill_8 FILLER_146_288 ();
 sg13g2_fill_8 FILLER_146_296 ();
 sg13g2_fill_8 FILLER_146_304 ();
 sg13g2_fill_8 FILLER_146_312 ();
 sg13g2_fill_8 FILLER_146_320 ();
 sg13g2_fill_8 FILLER_146_328 ();
 sg13g2_fill_8 FILLER_146_336 ();
 sg13g2_fill_8 FILLER_146_344 ();
 sg13g2_fill_8 FILLER_146_352 ();
 sg13g2_fill_8 FILLER_146_360 ();
 sg13g2_fill_8 FILLER_146_368 ();
 sg13g2_fill_8 FILLER_146_376 ();
 sg13g2_fill_8 FILLER_146_384 ();
 sg13g2_fill_8 FILLER_146_392 ();
 sg13g2_fill_8 FILLER_146_400 ();
 sg13g2_fill_8 FILLER_146_408 ();
 sg13g2_fill_8 FILLER_146_416 ();
 sg13g2_fill_8 FILLER_146_424 ();
 sg13g2_fill_8 FILLER_146_432 ();
 sg13g2_fill_8 FILLER_146_440 ();
 sg13g2_fill_8 FILLER_146_448 ();
 sg13g2_fill_8 FILLER_146_456 ();
 sg13g2_fill_8 FILLER_146_464 ();
 sg13g2_fill_8 FILLER_146_472 ();
 sg13g2_fill_8 FILLER_146_480 ();
 sg13g2_fill_8 FILLER_146_488 ();
 sg13g2_fill_8 FILLER_146_496 ();
 sg13g2_fill_8 FILLER_146_504 ();
 sg13g2_fill_8 FILLER_146_512 ();
 sg13g2_fill_8 FILLER_146_520 ();
 sg13g2_fill_8 FILLER_146_528 ();
 sg13g2_fill_8 FILLER_146_536 ();
 sg13g2_fill_8 FILLER_146_544 ();
 sg13g2_fill_8 FILLER_146_552 ();
 sg13g2_fill_8 FILLER_146_560 ();
 sg13g2_fill_8 FILLER_146_568 ();
 sg13g2_fill_8 FILLER_146_576 ();
 sg13g2_fill_8 FILLER_146_584 ();
 sg13g2_fill_8 FILLER_146_592 ();
 sg13g2_fill_8 FILLER_146_600 ();
 sg13g2_fill_8 FILLER_146_608 ();
 sg13g2_fill_8 FILLER_146_616 ();
 sg13g2_fill_8 FILLER_146_624 ();
 sg13g2_fill_8 FILLER_146_632 ();
 sg13g2_fill_8 FILLER_146_640 ();
 sg13g2_fill_8 FILLER_146_648 ();
 sg13g2_fill_8 FILLER_146_656 ();
 sg13g2_fill_8 FILLER_146_664 ();
 sg13g2_fill_8 FILLER_146_672 ();
 sg13g2_fill_8 FILLER_146_680 ();
 sg13g2_fill_8 FILLER_146_688 ();
 sg13g2_fill_8 FILLER_146_696 ();
 sg13g2_fill_8 FILLER_146_704 ();
 sg13g2_fill_8 FILLER_146_712 ();
 sg13g2_fill_8 FILLER_146_720 ();
 sg13g2_fill_8 FILLER_146_728 ();
 sg13g2_fill_8 FILLER_146_736 ();
 sg13g2_fill_8 FILLER_146_744 ();
 sg13g2_fill_8 FILLER_146_752 ();
 sg13g2_fill_8 FILLER_146_760 ();
 sg13g2_fill_8 FILLER_146_768 ();
 sg13g2_fill_8 FILLER_146_776 ();
 sg13g2_fill_8 FILLER_146_784 ();
 sg13g2_fill_8 FILLER_146_792 ();
 sg13g2_fill_8 FILLER_146_800 ();
 sg13g2_fill_8 FILLER_146_808 ();
 sg13g2_fill_8 FILLER_146_816 ();
 sg13g2_fill_8 FILLER_146_824 ();
 sg13g2_fill_8 FILLER_146_832 ();
 sg13g2_fill_8 FILLER_146_840 ();
 sg13g2_fill_8 FILLER_146_848 ();
 sg13g2_fill_8 FILLER_146_856 ();
 sg13g2_fill_8 FILLER_146_864 ();
 sg13g2_fill_8 FILLER_146_872 ();
 sg13g2_fill_8 FILLER_146_880 ();
 sg13g2_fill_8 FILLER_146_888 ();
 sg13g2_fill_8 FILLER_146_896 ();
 sg13g2_fill_8 FILLER_146_904 ();
 sg13g2_fill_8 FILLER_146_912 ();
 sg13g2_fill_8 FILLER_146_920 ();
 sg13g2_fill_8 FILLER_146_928 ();
 sg13g2_fill_8 FILLER_146_936 ();
 sg13g2_fill_8 FILLER_146_944 ();
 sg13g2_fill_8 FILLER_146_952 ();
 sg13g2_fill_8 FILLER_146_960 ();
 sg13g2_fill_8 FILLER_146_968 ();
 sg13g2_fill_8 FILLER_146_976 ();
 sg13g2_fill_8 FILLER_146_984 ();
 sg13g2_fill_8 FILLER_146_992 ();
 sg13g2_fill_8 FILLER_146_1000 ();
 sg13g2_fill_8 FILLER_146_1008 ();
 sg13g2_fill_8 FILLER_146_1016 ();
 sg13g2_fill_8 FILLER_146_1024 ();
 sg13g2_fill_8 FILLER_146_1032 ();
 sg13g2_fill_8 FILLER_146_1040 ();
 sg13g2_fill_8 FILLER_146_1048 ();
 sg13g2_fill_8 FILLER_146_1056 ();
 sg13g2_fill_8 FILLER_146_1064 ();
 sg13g2_fill_8 FILLER_146_1072 ();
 sg13g2_fill_8 FILLER_146_1080 ();
 sg13g2_fill_8 FILLER_146_1088 ();
 sg13g2_fill_8 FILLER_146_1096 ();
 sg13g2_fill_8 FILLER_146_1104 ();
 sg13g2_fill_8 FILLER_146_1112 ();
 sg13g2_fill_8 FILLER_146_1120 ();
 sg13g2_fill_8 FILLER_146_1128 ();
 sg13g2_fill_8 FILLER_146_1136 ();
 sg13g2_fill_8 FILLER_146_1144 ();
 sg13g2_fill_8 FILLER_146_1152 ();
 sg13g2_fill_4 FILLER_146_1160 ();
 sg13g2_fill_2 FILLER_146_1164 ();
endmodule
