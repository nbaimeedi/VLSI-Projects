//Latest Update Date: 10th Aug, 2025
//Owner: B Nithin Reddy


//Interface
interface spi_master_if;
  
  logic clk, newd, rst;
  logic [11:0] din;
  logic mosi,cs,sclk;
  
endinterface
