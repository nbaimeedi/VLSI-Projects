module dmi_jtag (clk_i,
    dmi_req_o_0_,
    dmi_req_o_10_,
    dmi_req_o_11_,
    dmi_req_o_12_,
    dmi_req_o_13_,
    dmi_req_o_14_,
    dmi_req_o_15_,
    dmi_req_o_16_,
    dmi_req_o_17_,
    dmi_req_o_18_,
    dmi_req_o_19_,
    dmi_req_o_1_,
    dmi_req_o_20_,
    dmi_req_o_21_,
    dmi_req_o_22_,
    dmi_req_o_23_,
    dmi_req_o_24_,
    dmi_req_o_25_,
    dmi_req_o_26_,
    dmi_req_o_27_,
    dmi_req_o_28_,
    dmi_req_o_29_,
    dmi_req_o_2_,
    dmi_req_o_30_,
    dmi_req_o_31_,
    dmi_req_o_32_,
    dmi_req_o_33_,
    dmi_req_o_34_,
    dmi_req_o_35_,
    dmi_req_o_36_,
    dmi_req_o_37_,
    dmi_req_o_38_,
    dmi_req_o_39_,
    dmi_req_o_3_,
    dmi_req_o_40_,
    dmi_req_o_4_,
    dmi_req_o_5_,
    dmi_req_o_6_,
    dmi_req_o_7_,
    dmi_req_o_8_,
    dmi_req_o_9_,
    dmi_req_ready_i,
    dmi_req_valid_o,
    dmi_resp_i_0_,
    dmi_resp_i_10_,
    dmi_resp_i_11_,
    dmi_resp_i_12_,
    dmi_resp_i_13_,
    dmi_resp_i_14_,
    dmi_resp_i_15_,
    dmi_resp_i_16_,
    dmi_resp_i_17_,
    dmi_resp_i_18_,
    dmi_resp_i_19_,
    dmi_resp_i_1_,
    dmi_resp_i_20_,
    dmi_resp_i_21_,
    dmi_resp_i_22_,
    dmi_resp_i_23_,
    dmi_resp_i_24_,
    dmi_resp_i_25_,
    dmi_resp_i_26_,
    dmi_resp_i_27_,
    dmi_resp_i_28_,
    dmi_resp_i_29_,
    dmi_resp_i_2_,
    dmi_resp_i_30_,
    dmi_resp_i_31_,
    dmi_resp_i_32_,
    dmi_resp_i_33_,
    dmi_resp_i_3_,
    dmi_resp_i_4_,
    dmi_resp_i_5_,
    dmi_resp_i_6_,
    dmi_resp_i_7_,
    dmi_resp_i_8_,
    dmi_resp_i_9_,
    dmi_resp_ready_o,
    dmi_resp_valid_i,
    dmi_rst_no,
    rst_ni,
    tck_i,
    td_i,
    td_o,
    tdo_oe_o,
    testmode_i,
    tms_i,
    trst_ni);
 input clk_i;
 output dmi_req_o_0_;
 output dmi_req_o_10_;
 output dmi_req_o_11_;
 output dmi_req_o_12_;
 output dmi_req_o_13_;
 output dmi_req_o_14_;
 output dmi_req_o_15_;
 output dmi_req_o_16_;
 output dmi_req_o_17_;
 output dmi_req_o_18_;
 output dmi_req_o_19_;
 output dmi_req_o_1_;
 output dmi_req_o_20_;
 output dmi_req_o_21_;
 output dmi_req_o_22_;
 output dmi_req_o_23_;
 output dmi_req_o_24_;
 output dmi_req_o_25_;
 output dmi_req_o_26_;
 output dmi_req_o_27_;
 output dmi_req_o_28_;
 output dmi_req_o_29_;
 output dmi_req_o_2_;
 output dmi_req_o_30_;
 output dmi_req_o_31_;
 output dmi_req_o_32_;
 output dmi_req_o_33_;
 output dmi_req_o_34_;
 output dmi_req_o_35_;
 output dmi_req_o_36_;
 output dmi_req_o_37_;
 output dmi_req_o_38_;
 output dmi_req_o_39_;
 output dmi_req_o_3_;
 output dmi_req_o_40_;
 output dmi_req_o_4_;
 output dmi_req_o_5_;
 output dmi_req_o_6_;
 output dmi_req_o_7_;
 output dmi_req_o_8_;
 output dmi_req_o_9_;
 input dmi_req_ready_i;
 output dmi_req_valid_o;
 input dmi_resp_i_0_;
 input dmi_resp_i_10_;
 input dmi_resp_i_11_;
 input dmi_resp_i_12_;
 input dmi_resp_i_13_;
 input dmi_resp_i_14_;
 input dmi_resp_i_15_;
 input dmi_resp_i_16_;
 input dmi_resp_i_17_;
 input dmi_resp_i_18_;
 input dmi_resp_i_19_;
 input dmi_resp_i_1_;
 input dmi_resp_i_20_;
 input dmi_resp_i_21_;
 input dmi_resp_i_22_;
 input dmi_resp_i_23_;
 input dmi_resp_i_24_;
 input dmi_resp_i_25_;
 input dmi_resp_i_26_;
 input dmi_resp_i_27_;
 input dmi_resp_i_28_;
 input dmi_resp_i_29_;
 input dmi_resp_i_2_;
 input dmi_resp_i_30_;
 input dmi_resp_i_31_;
 input dmi_resp_i_32_;
 input dmi_resp_i_33_;
 input dmi_resp_i_3_;
 input dmi_resp_i_4_;
 input dmi_resp_i_5_;
 input dmi_resp_i_6_;
 input dmi_resp_i_7_;
 input dmi_resp_i_8_;
 input dmi_resp_i_9_;
 output dmi_resp_ready_o;
 input dmi_resp_valid_i;
 output dmi_rst_no;
 input rst_ni;
 input tck_i;
 input td_i;
 output td_o;
 output tdo_oe_o;
 input testmode_i;
 input tms_i;
 input trst_ni;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire net219;
 wire _0099_;
 wire net218;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire net217;
 wire _0114_;
 wire _0115_;
 wire net216;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire net215;
 wire _0126_;
 wire _0127_;
 wire net214;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire net213;
 wire net212;
 wire _0157_;
 wire _0158_;
 wire net211;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire net210;
 wire _0167_;
 wire _0168_;
 wire net209;
 wire _0170_;
 wire _0171_;
 wire net208;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire net207;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire net206;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire net282;
 wire _0238_;
 wire net281;
 wire net280;
 wire net279;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire net278;
 wire _0246_;
 wire net277;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire net276;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire net275;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire net274;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire net273;
 wire net272;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire net271;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire net270;
 wire net268;
 wire net267;
 wire net266;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire net265;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire net264;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire net263;
 wire _0346_;
 wire _0347_;
 wire net262;
 wire net261;
 wire net260;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire net259;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire net258;
 wire net257;
 wire _0360_;
 wire net256;
 wire net255;
 wire _0363_;
 wire net254;
 wire net253;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire net252;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire net251;
 wire _0393_;
 wire _0394_;
 wire net250;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire net249;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire net248;
 wire _0409_;
 wire net247;
 wire net246;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire net245;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire net244;
 wire net243;
 wire net242;
 wire _0529_;
 wire net241;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire net240;
 wire _0547_;
 wire _0548_;
 wire net239;
 wire net238;
 wire _0551_;
 wire _0552_;
 wire net237;
 wire net236;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire net235;
 wire _0575_;
 wire _0576_;
 wire net234;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire net233;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire net232;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire net231;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire net230;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire net229;
 wire _0634_;
 wire _0635_;
 wire net228;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire net227;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire net226;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire net225;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire net224;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire net223;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire net222;
 wire _0697_;
 wire net221;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire net220;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire net4;
 wire net3;
 wire address_q_0_;
 wire address_q_1_;
 wire address_q_2_;
 wire address_q_3_;
 wire address_q_4_;
 wire address_q_5_;
 wire address_q_6_;
 wire data_q_0_;
 wire data_q_10_;
 wire data_q_11_;
 wire data_q_12_;
 wire data_q_13_;
 wire data_q_14_;
 wire data_q_15_;
 wire data_q_16_;
 wire data_q_17_;
 wire data_q_18_;
 wire data_q_19_;
 wire data_q_1_;
 wire data_q_20_;
 wire data_q_21_;
 wire data_q_22_;
 wire data_q_23_;
 wire data_q_24_;
 wire data_q_25_;
 wire data_q_26_;
 wire data_q_27_;
 wire data_q_28_;
 wire data_q_29_;
 wire data_q_2_;
 wire data_q_30_;
 wire data_q_31_;
 wire data_q_3_;
 wire data_q_4_;
 wire data_q_5_;
 wire data_q_6_;
 wire data_q_7_;
 wire data_q_8_;
 wire data_q_9_;
 wire dmi_0_;
 wire dmi_10_;
 wire dmi_11_;
 wire dmi_12_;
 wire dmi_13_;
 wire dmi_14_;
 wire dmi_15_;
 wire dmi_16_;
 wire dmi_17_;
 wire dmi_18_;
 wire dmi_19_;
 wire dmi_1_;
 wire dmi_20_;
 wire dmi_21_;
 wire dmi_22_;
 wire dmi_23_;
 wire dmi_24_;
 wire dmi_25_;
 wire dmi_26_;
 wire dmi_27_;
 wire dmi_28_;
 wire dmi_29_;
 wire dmi_2_;
 wire dmi_30_;
 wire dmi_31_;
 wire dmi_32_;
 wire dmi_33_;
 wire dmi_34_;
 wire dmi_35_;
 wire dmi_36_;
 wire dmi_37_;
 wire dmi_38_;
 wire dmi_39_;
 wire dmi_3_;
 wire dmi_40_;
 wire dmi_4_;
 wire dmi_5_;
 wire dmi_6_;
 wire dmi_7_;
 wire dmi_8_;
 wire dmi_9_;
 wire net269;
 wire dmi_req_32_;
 wire dmi_req_33_;
 wire dmi_req_ready;
 wire dmi_req_valid;
 wire dmi_resp_0_;
 wire dmi_resp_10_;
 wire dmi_resp_11_;
 wire dmi_resp_12_;
 wire dmi_resp_13_;
 wire dmi_resp_14_;
 wire dmi_resp_15_;
 wire dmi_resp_16_;
 wire dmi_resp_17_;
 wire dmi_resp_18_;
 wire dmi_resp_19_;
 wire dmi_resp_1_;
 wire dmi_resp_20_;
 wire dmi_resp_21_;
 wire dmi_resp_22_;
 wire dmi_resp_23_;
 wire dmi_resp_24_;
 wire dmi_resp_25_;
 wire dmi_resp_26_;
 wire dmi_resp_27_;
 wire dmi_resp_28_;
 wire dmi_resp_29_;
 wire dmi_resp_2_;
 wire dmi_resp_30_;
 wire dmi_resp_31_;
 wire dmi_resp_32_;
 wire dmi_resp_33_;
 wire dmi_resp_3_;
 wire dmi_resp_4_;
 wire dmi_resp_5_;
 wire dmi_resp_6_;
 wire dmi_resp_7_;
 wire dmi_resp_8_;
 wire dmi_resp_9_;
 wire dmi_resp_valid;
 wire dr_d_0_;
 wire dr_d_10_;
 wire dr_d_11_;
 wire dr_d_12_;
 wire dr_d_13_;
 wire dr_d_14_;
 wire dr_d_15_;
 wire dr_d_16_;
 wire dr_d_17_;
 wire dr_d_18_;
 wire dr_d_19_;
 wire dr_d_1_;
 wire dr_d_20_;
 wire dr_d_21_;
 wire dr_d_22_;
 wire dr_d_23_;
 wire dr_d_24_;
 wire dr_d_25_;
 wire dr_d_26_;
 wire dr_d_27_;
 wire dr_d_28_;
 wire dr_d_29_;
 wire dr_d_2_;
 wire dr_d_30_;
 wire dr_d_31_;
 wire dr_d_32_;
 wire dr_d_33_;
 wire dr_d_34_;
 wire dr_d_35_;
 wire dr_d_36_;
 wire dr_d_37_;
 wire dr_d_38_;
 wire dr_d_39_;
 wire dr_d_3_;
 wire dr_d_40_;
 wire dr_d_4_;
 wire dr_d_5_;
 wire dr_d_6_;
 wire dr_d_7_;
 wire dr_d_8_;
 wire dr_d_9_;
 wire dtmcs_d_0_;
 wire dtmcs_d_10_;
 wire dtmcs_d_11_;
 wire dtmcs_d_12_;
 wire dtmcs_d_13_;
 wire dtmcs_d_14_;
 wire dtmcs_d_15_;
 wire dtmcs_d_16_;
 wire dtmcs_d_17_;
 wire dtmcs_d_18_;
 wire dtmcs_d_19_;
 wire dtmcs_d_1_;
 wire dtmcs_d_20_;
 wire dtmcs_d_21_;
 wire dtmcs_d_22_;
 wire dtmcs_d_23_;
 wire dtmcs_d_24_;
 wire dtmcs_d_25_;
 wire dtmcs_d_26_;
 wire dtmcs_d_27_;
 wire dtmcs_d_28_;
 wire dtmcs_d_29_;
 wire dtmcs_d_2_;
 wire dtmcs_d_30_;
 wire dtmcs_d_31_;
 wire dtmcs_d_3_;
 wire dtmcs_d_4_;
 wire dtmcs_d_5_;
 wire dtmcs_d_6_;
 wire dtmcs_d_7_;
 wire dtmcs_d_8_;
 wire dtmcs_d_9_;
 wire dtmcs_q_0_;
 wire dtmcs_q_10_;
 wire dtmcs_q_11_;
 wire dtmcs_q_12_;
 wire dtmcs_q_13_;
 wire dtmcs_q_14_;
 wire dtmcs_q_15_;
 wire dtmcs_q_16_;
 wire dtmcs_q_17_;
 wire dtmcs_q_18_;
 wire dtmcs_q_19_;
 wire dtmcs_q_1_;
 wire dtmcs_q_20_;
 wire dtmcs_q_21_;
 wire dtmcs_q_22_;
 wire dtmcs_q_23_;
 wire dtmcs_q_24_;
 wire dtmcs_q_25_;
 wire dtmcs_q_26_;
 wire dtmcs_q_27_;
 wire dtmcs_q_28_;
 wire dtmcs_q_29_;
 wire dtmcs_q_2_;
 wire dtmcs_q_30_;
 wire dtmcs_q_31_;
 wire dtmcs_q_3_;
 wire dtmcs_q_4_;
 wire dtmcs_q_5_;
 wire dtmcs_q_6_;
 wire dtmcs_q_7_;
 wire dtmcs_q_8_;
 wire dtmcs_q_9_;
 wire error_q_0_;
 wire \error_q_0__$_NOT__A_Y ;
 wire error_q_1_;
 wire \error_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.clear_pending_rise_edge_detect_$_AND__Y_A ;
 wire \i_dmi_cdc.core_clear_pending ;
 wire \i_dmi_cdc.core_clear_pending_q ;
 wire \i_dmi_jtag_tap.bypass_d ;
 wire \i_dmi_jtag_tap.bypass_q ;
 wire \i_dmi_jtag_tap.idcode_d_12_ ;
 wire \i_dmi_jtag_tap.idcode_d_13_ ;
 wire \i_dmi_jtag_tap.idcode_d_14_ ;
 wire \i_dmi_jtag_tap.idcode_d_15_ ;
 wire \i_dmi_jtag_tap.idcode_d_16_ ;
 wire \i_dmi_jtag_tap.idcode_d_17_ ;
 wire \i_dmi_jtag_tap.idcode_d_18_ ;
 wire \i_dmi_jtag_tap.idcode_d_19_ ;
 wire \i_dmi_jtag_tap.idcode_d_20_ ;
 wire \i_dmi_jtag_tap.idcode_d_21_ ;
 wire \i_dmi_jtag_tap.idcode_d_22_ ;
 wire \i_dmi_jtag_tap.idcode_d_23_ ;
 wire \i_dmi_jtag_tap.idcode_d_24_ ;
 wire \i_dmi_jtag_tap.idcode_d_25_ ;
 wire \i_dmi_jtag_tap.idcode_d_26_ ;
 wire \i_dmi_jtag_tap.idcode_d_27_ ;
 wire \i_dmi_jtag_tap.idcode_d_28_ ;
 wire \i_dmi_jtag_tap.idcode_d_29_ ;
 wire \i_dmi_jtag_tap.idcode_d_2_ ;
 wire \i_dmi_jtag_tap.idcode_d_30_ ;
 wire \i_dmi_jtag_tap.idcode_d_31_ ;
 wire \i_dmi_jtag_tap.idcode_d_3_ ;
 wire \i_dmi_jtag_tap.idcode_d_6_ ;
 wire \i_dmi_jtag_tap.idcode_d_9_ ;
 wire \i_dmi_jtag_tap.idcode_q_0_ ;
 wire \i_dmi_jtag_tap.idcode_q_10_ ;
 wire \i_dmi_jtag_tap.idcode_q_11_ ;
 wire \i_dmi_jtag_tap.idcode_q_12_ ;
 wire \i_dmi_jtag_tap.idcode_q_13_ ;
 wire \i_dmi_jtag_tap.idcode_q_14_ ;
 wire \i_dmi_jtag_tap.idcode_q_15_ ;
 wire \i_dmi_jtag_tap.idcode_q_16_ ;
 wire \i_dmi_jtag_tap.idcode_q_17_ ;
 wire \i_dmi_jtag_tap.idcode_q_18_ ;
 wire \i_dmi_jtag_tap.idcode_q_19_ ;
 wire \i_dmi_jtag_tap.idcode_q_1_ ;
 wire \i_dmi_jtag_tap.idcode_q_20_ ;
 wire \i_dmi_jtag_tap.idcode_q_21_ ;
 wire \i_dmi_jtag_tap.idcode_q_22_ ;
 wire \i_dmi_jtag_tap.idcode_q_23_ ;
 wire \i_dmi_jtag_tap.idcode_q_24_ ;
 wire \i_dmi_jtag_tap.idcode_q_25_ ;
 wire \i_dmi_jtag_tap.idcode_q_26_ ;
 wire \i_dmi_jtag_tap.idcode_q_27_ ;
 wire \i_dmi_jtag_tap.idcode_q_28_ ;
 wire \i_dmi_jtag_tap.idcode_q_29_ ;
 wire \i_dmi_jtag_tap.idcode_q_2_ ;
 wire \i_dmi_jtag_tap.idcode_q_30_ ;
 wire \i_dmi_jtag_tap.idcode_q_31_ ;
 wire \i_dmi_jtag_tap.idcode_q_3_ ;
 wire \i_dmi_jtag_tap.idcode_q_4_ ;
 wire \i_dmi_jtag_tap.idcode_q_5_ ;
 wire \i_dmi_jtag_tap.idcode_q_6_ ;
 wire \i_dmi_jtag_tap.idcode_q_7_ ;
 wire \i_dmi_jtag_tap.idcode_q_8_ ;
 wire \i_dmi_jtag_tap.idcode_q_9_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_0_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_1_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_2_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_3_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_4_ ;
 wire \i_dmi_jtag_tap.jtag_ir_q_4__$_NOT__A_Y ;
 wire \i_dmi_jtag_tap.jtag_ir_shift_q_0_ ;
 wire \i_dmi_jtag_tap.jtag_ir_shift_q_1_ ;
 wire \i_dmi_jtag_tap.jtag_ir_shift_q_2_ ;
 wire \i_dmi_jtag_tap.jtag_ir_shift_q_3_ ;
 wire \i_dmi_jtag_tap.jtag_ir_shift_q_4_ ;
 wire \i_dmi_jtag_tap.tap_state_d_1_ ;
 wire \i_dmi_jtag_tap.tap_state_d_2_ ;
 wire \i_dmi_jtag_tap.tap_state_d_3_ ;
 wire \i_dmi_jtag_tap.tap_state_q_0_ ;
 wire \i_dmi_jtag_tap.tap_state_q_1_ ;
 wire \i_dmi_jtag_tap.tap_state_q_1__$_NOT__A_Y ;
 wire \i_dmi_jtag_tap.tap_state_q_2_ ;
 wire \i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ;
 wire \i_dmi_jtag_tap.tap_state_q_3_ ;
 wire \i_dmi_jtag_tap.tap_state_q_3__$_NOT__A_Y ;
 wire \i_dmi_jtag_tap.tck_n ;
 wire \i_dmi_jtag_tap.tck_ni ;
 wire \i_dmi_jtag_tap.tdo_mux ;
 wire \state_d_1__$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_OR__Y_A ;
 wire state_q_0_;
 wire \state_q_0__$_NOT__A_Y ;
 wire \state_q_0__$_OR__A_Y_$_OR__A_1_B ;
 wire \state_q_0__reg_E_$_AND__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B ;
 wire state_q_1_;
 wire \state_q_1__$_NOT__A_Y ;
 wire state_q_2_;
 wire tdo_oe_o_reg_D;
 wire \i_dmi_cdc.i_cdc_req/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/_2_ ;
 wire \i_dmi_cdc.i_cdc_req/_3_ ;
 wire \i_dmi_cdc.i_cdc_req/async_ack ;
 wire \i_dmi_cdc.i_cdc_req/async_data_0_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_10_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_11_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_12_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_13_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_14_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_15_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_16_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_17_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_18_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_19_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_1_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_20_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_21_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_22_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_23_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_24_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_25_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_26_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_27_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_28_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_29_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_2_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_30_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_31_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_32_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_33_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_34_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_35_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_36_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_37_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_38_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_39_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_3_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_40_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_4_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_5_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_6_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_7_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_8_ ;
 wire \i_dmi_cdc.i_cdc_req/async_data_9_ ;
 wire \i_dmi_cdc.i_cdc_req/async_req ;
 wire \i_dmi_cdc.i_cdc_req/i_dst_ready_i ;
 wire \i_dmi_cdc.i_cdc_req/i_src_valid_i ;
 wire \i_dmi_cdc.i_cdc_req/s_dst_clear_ack_q ;
 wire \i_dmi_cdc.i_cdc_req/s_dst_clear_req ;
 wire \i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ;
 wire \i_dmi_cdc.i_cdc_req/s_dst_valid ;
 wire \i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ;
 wire \i_dmi_cdc.i_cdc_req/s_src_clear_req ;
 wire \i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ;
 wire \i_dmi_cdc.i_cdc_req/s_src_ready ;
 wire \i_dmi_cdc.i_cdc_req/src_clear_pending_o ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_012_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_013_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_015_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ;
 wire net205;
 wire net204;
 wire net203;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ;
 wire net202;
 wire net201;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ;
 wire net200;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_072_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_073_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_074_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_075_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_076_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_077_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_078_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_079_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_01_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_20_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ;
 wire net199;
 wire net198;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ;
 wire net197;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ;
 wire net196;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_01_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_20_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_000_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_001_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_002_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_003_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_004_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_005_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_006_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_007_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_008_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_009_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_010_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_011_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_012_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_013_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_014_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_015_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_016_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_017_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_018_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_019_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_020_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_021_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_022_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_023_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_024_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_025_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_026_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_027_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_028_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_029_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_030_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_031_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_032_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_033_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_034_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_035_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_036_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_037_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_038_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_039_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_040_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_041_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_042_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_043_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_044_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_045_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_046_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_047_ ;
 wire net195;
 wire net194;
 wire net193;
 wire net192;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire net187;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_057_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_058_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_059_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_060_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_061_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_062_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_063_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_064_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_065_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_066_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_067_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_068_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_069_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_070_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_071_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_072_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_073_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_074_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_075_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_076_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_077_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_078_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_079_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_080_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_081_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_082_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_083_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_084_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_085_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_086_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_087_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_088_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_089_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_090_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_091_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_092_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_093_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_094_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_095_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_096_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_097_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/_098_ ;
 wire net45;
 wire \i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d_$_MUX__Y_A ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_13_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_14_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_15_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_16_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_17_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_18_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_19_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_20_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_21_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_22_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_23_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_24_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_25_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_26_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_27_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_28_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_29_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_30_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_31_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_32_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_33_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_34_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_35_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_36_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_37_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_38_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_39_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_3_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_40_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_4_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_5_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_6_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_7_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_8_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_9_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/i_sync/_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_000_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_001_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_002_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_003_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_004_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_005_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_006_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_007_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_008_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_009_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_010_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_011_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_012_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_013_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_014_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_015_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_016_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_017_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_018_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_019_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_020_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_021_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_022_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_023_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_024_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_025_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_026_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_027_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_028_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_029_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_030_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_031_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_032_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_033_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_034_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_035_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_036_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_037_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_038_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_039_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_040_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_041_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_042_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_043_ ;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire net182;
 wire net181;
 wire \i_dmi_cdc.i_cdc_req/i_src/_050_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_051_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_052_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_053_ ;
 wire net180;
 wire net179;
 wire net178;
 wire \i_dmi_cdc.i_cdc_req/i_src/_057_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_058_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_059_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_060_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_061_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_062_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_063_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_064_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_065_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_066_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_067_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_068_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_069_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_070_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_071_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_072_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_073_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_074_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_075_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_076_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_077_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_078_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_079_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_080_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_081_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_082_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_083_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_084_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_085_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_086_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_087_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_088_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_089_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_090_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_091_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_092_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_093_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_094_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_095_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_096_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/_097_ ;
 wire net86;
 wire \i_dmi_cdc.i_cdc_req/i_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_10_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_11_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_12_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_13_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_14_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_15_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_16_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_17_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_18_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_19_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_20_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_21_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_22_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_23_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_24_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_25_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_26_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_27_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_28_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_29_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_30_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_31_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_32_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_33_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_34_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_35_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_36_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_37_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_38_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_39_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_3_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_40_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_4_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_5_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_6_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_7_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_8_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/data_src_d_9_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_req/i_src/req_src_d_$_MUX__Y_A ;
 wire \i_dmi_cdc.i_cdc_req/i_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/i_sync/_2_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_ack ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_13_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_14_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_15_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_16_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_17_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_18_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_19_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_20_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_21_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_22_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_23_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_24_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_25_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_26_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_27_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_28_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_29_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_30_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_31_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_32_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_33_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_4_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_5_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_6_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_7_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_8_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_data_9_ ;
 wire \i_dmi_cdc.i_cdc_resp/async_req ;
 wire \i_dmi_cdc.i_cdc_resp/dst_clear_pending_o ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst_ready_i ;
 wire \i_dmi_cdc.i_cdc_resp/i_src_valid_i ;
 wire \i_dmi_cdc.i_cdc_resp/s_dst_clear_ack_q ;
 wire \i_dmi_cdc.i_cdc_resp/s_dst_clear_req ;
 wire \i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ;
 wire \i_dmi_cdc.i_cdc_resp/s_dst_valid ;
 wire \i_dmi_cdc.i_cdc_resp/s_src_clear_ack_q ;
 wire \i_dmi_cdc.i_cdc_resp/s_src_clear_req ;
 wire \i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ;
 wire \i_dmi_cdc.i_cdc_resp/s_src_ready ;
 wire \i_dmi_cdc.i_cdc_resp/src_clear_pending_o ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ;
 wire net177;
 wire net176;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ;
 wire net175;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_022_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_023_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ;
 wire net174;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_026_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_027_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_032_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_01_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_20_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ;
 wire net173;
 wire net172;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ;
 wire net171;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ;
 wire net170;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_01_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_20_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_000_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_001_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_002_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_003_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_004_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_005_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_006_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_007_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_008_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_009_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_010_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_011_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_012_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_013_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_014_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_015_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_016_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_017_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_018_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_019_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_020_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_021_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_022_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_023_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_024_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_025_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_026_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_027_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_028_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_029_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_030_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_031_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_032_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_033_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_034_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_035_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_036_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_037_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_038_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_039_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_040_ ;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire net162;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_049_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_050_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_051_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_052_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_053_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_054_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_055_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_056_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_057_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_058_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_059_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_060_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_061_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_062_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_063_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_064_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_065_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_066_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_067_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_068_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_069_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_070_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_071_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_072_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_073_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_074_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_075_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_076_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_077_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_078_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_079_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_080_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_081_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_082_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/_083_ ;
 wire net120;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d_$_MUX__Y_A ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_13_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_14_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_15_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_16_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_17_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_18_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_19_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_20_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_21_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_22_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_23_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_24_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_25_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_26_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_27_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_28_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_29_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_30_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_31_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_32_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_33_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_4_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_5_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_6_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_7_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_8_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_9_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/req_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_000_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_001_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_002_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_003_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_004_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_005_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_006_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_007_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_008_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_009_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_010_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_011_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_012_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_013_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_014_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_015_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_016_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_017_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_018_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_019_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_020_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_021_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_022_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_023_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_024_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_025_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_026_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_027_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_028_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_029_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_030_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_031_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_032_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_033_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_034_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_035_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_036_ ;
 wire net161;
 wire net160;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_043_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_044_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_045_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_046_ ;
 wire net155;
 wire net154;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_049_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_050_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_051_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_052_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_053_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_054_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_055_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_056_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_057_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_058_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_059_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_060_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_061_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_062_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_063_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_064_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_065_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_066_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_067_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_068_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_069_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_070_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_071_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_072_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_073_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_074_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_075_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_076_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_077_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_078_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_079_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_080_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_081_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/_082_ ;
 wire net283;
 wire \i_dmi_cdc.i_cdc_resp/i_src/ack_synced ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_10_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_11_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_12_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_13_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_14_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_15_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_16_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_17_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_18_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_19_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_20_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_21_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_22_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_23_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_24_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_25_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_26_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_27_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_28_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_29_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_30_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_31_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_32_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_33_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_3_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_4_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_5_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_6_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_7_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_8_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/data_src_d_9_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/req_src_d ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/req_src_d_$_MUX__Y_A ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/i_sync/_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/i_sync/_1_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/i_sync/_2_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_0_ ;
 wire \i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_1_ ;
 wire net1;
 wire net2;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire clknet_0_clk_i;
 wire clknet_4_0_0_clk_i;
 wire clknet_4_1_0_clk_i;
 wire clknet_4_2_0_clk_i;
 wire clknet_4_3_0_clk_i;
 wire clknet_4_4_0_clk_i;
 wire clknet_4_5_0_clk_i;
 wire clknet_4_6_0_clk_i;
 wire clknet_4_7_0_clk_i;
 wire clknet_4_8_0_clk_i;
 wire clknet_4_9_0_clk_i;
 wire clknet_4_10_0_clk_i;
 wire clknet_4_11_0_clk_i;
 wire clknet_4_12_0_clk_i;
 wire clknet_4_13_0_clk_i;
 wire clknet_4_14_0_clk_i;
 wire clknet_4_15_0_clk_i;
 wire clknet_5_0__leaf_clk_i;
 wire clknet_5_1__leaf_clk_i;
 wire clknet_5_2__leaf_clk_i;
 wire clknet_5_3__leaf_clk_i;
 wire clknet_5_4__leaf_clk_i;
 wire clknet_5_5__leaf_clk_i;
 wire clknet_5_6__leaf_clk_i;
 wire clknet_5_7__leaf_clk_i;
 wire clknet_5_8__leaf_clk_i;
 wire clknet_5_9__leaf_clk_i;
 wire clknet_5_10__leaf_clk_i;
 wire clknet_5_11__leaf_clk_i;
 wire clknet_5_12__leaf_clk_i;
 wire clknet_5_13__leaf_clk_i;
 wire clknet_5_14__leaf_clk_i;
 wire clknet_5_15__leaf_clk_i;
 wire clknet_5_16__leaf_clk_i;
 wire clknet_5_17__leaf_clk_i;
 wire clknet_5_18__leaf_clk_i;
 wire clknet_5_19__leaf_clk_i;
 wire clknet_5_20__leaf_clk_i;
 wire clknet_5_21__leaf_clk_i;
 wire clknet_5_22__leaf_clk_i;
 wire clknet_5_23__leaf_clk_i;
 wire clknet_5_24__leaf_clk_i;
 wire clknet_5_25__leaf_clk_i;
 wire clknet_5_26__leaf_clk_i;
 wire clknet_5_27__leaf_clk_i;
 wire clknet_5_28__leaf_clk_i;
 wire clknet_5_29__leaf_clk_i;
 wire clknet_5_30__leaf_clk_i;
 wire clknet_5_31__leaf_clk_i;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;

 sg13g2_buf_4 fanout282 (.X(net282),
    .A(net283));
 sg13g2_or2_2 _0896_ (.X(_0238_),
    .B(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .A(\i_dmi_jtag_tap.tap_state_q_1_ ));
 sg13g2_buf_2 fanout281 (.A(net282),
    .X(net281));
 sg13g2_buf_4 fanout280 (.X(net280),
    .A(net282));
 sg13g2_buf_4 fanout279 (.X(net279),
    .A(net283));
 sg13g2_or2_1 _0900_ (.X(_0242_),
    .B(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .A(net319));
 sg13g2_nand2_1 _0901_ (.Y(_0243_),
    .A(\i_dmi_jtag_tap.tap_state_q_2_ ),
    .B(_0242_));
 sg13g2_nand2b_1 _0902_ (.Y(_0244_),
    .B(_0243_),
    .A_N(net317));
 sg13g2_buf_4 fanout278 (.X(net278),
    .A(net279));
 sg13g2_a21oi_1 _0904_ (.A1(_0238_),
    .A2(_0244_),
    .Y(_0246_),
    .B1(net314));
 sg13g2_buf_2 fanout277 (.A(_0342_),
    .X(net277));
 sg13g2_or2_2 _0906_ (.X(_0248_),
    .B(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .A(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ));
 sg13g2_nor2_1 _0907_ (.A(net317),
    .B(_0248_),
    .Y(_0249_));
 sg13g2_or2_2 _0908_ (.X(_0250_),
    .B(net316),
    .A(net317));
 sg13g2_buf_2 fanout276 (.A(net277),
    .X(net276));
 sg13g2_a21oi_1 _0910_ (.A1(_0238_),
    .A2(_0250_),
    .Y(_0252_),
    .B1(\i_dmi_jtag_tap.tap_state_q_3_ ));
 sg13g2_nand2b_1 _0911_ (.Y(_0253_),
    .B(net319),
    .A_N(\i_dmi_jtag_tap.tap_state_q_1_ ));
 sg13g2_nor3_1 _0912_ (.A(\i_dmi_jtag_tap.tap_state_q_2_ ),
    .B(net314),
    .C(_0253_),
    .Y(_0254_));
 sg13g2_nor3_1 _0913_ (.A(_0249_),
    .B(_0252_),
    .C(_0254_),
    .Y(_0255_));
 sg13g2_inv_1 _0914_ (.Y(_0256_),
    .A(_0255_));
 sg13g2_nand2b_2 _0915_ (.Y(_0257_),
    .B(net319),
    .A_N(\i_dmi_jtag_tap.tap_state_q_1__$_NOT__A_Y ));
 sg13g2_nor3_1 _0916_ (.A(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .B(net315),
    .C(_0257_),
    .Y(_0258_));
 sg13g2_mux2_1 _0917_ (.A0(net314),
    .A1(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .S(net319),
    .X(_0259_));
 sg13g2_nor3_1 _0918_ (.A(\i_dmi_jtag_tap.tap_state_q_1_ ),
    .B(net316),
    .C(_0259_),
    .Y(_0260_));
 sg13g2_nor2_1 _0919_ (.A(_0258_),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_o21ai_1 _0920_ (.B1(_0261_),
    .Y(_0262_),
    .A1(_0246_),
    .A2(_0256_));
 sg13g2_nor2b_1 _0921_ (.A(tms_i),
    .B_N(_0262_),
    .Y(_0263_));
 sg13g2_nor2_1 _0922_ (.A(net314),
    .B(_0238_),
    .Y(_0264_));
 sg13g2_buf_2 fanout275 (.A(net276),
    .X(net275));
 sg13g2_nand2_1 _0924_ (.Y(_0266_),
    .A(tms_i),
    .B(net320));
 sg13g2_nand2_1 _0925_ (.Y(_0267_),
    .A(_0264_),
    .B(_0266_));
 sg13g2_mux2_1 _0926_ (.A0(_0238_),
    .A1(_0250_),
    .S(net318),
    .X(_0268_));
 sg13g2_nor2_2 _0927_ (.A(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nor3_1 _0928_ (.A(net320),
    .B(net317),
    .C(_0248_),
    .Y(_0270_));
 sg13g2_o21ai_1 _0929_ (.B1(tms_i),
    .Y(_0271_),
    .A1(_0269_),
    .A2(_0270_));
 sg13g2_o21ai_1 _0930_ (.B1(_0242_),
    .Y(_0272_),
    .A1(net174),
    .A2(net316));
 sg13g2_nor2_1 _0931_ (.A(net317),
    .B(net315),
    .Y(_0273_));
 sg13g2_and2_1 _0932_ (.A(_0272_),
    .B(_0273_),
    .X(_0274_));
 sg13g2_nor3_1 _0933_ (.A(net318),
    .B(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .C(_0250_),
    .Y(_0275_));
 sg13g2_nor2_1 _0934_ (.A(_0274_),
    .B(_0275_),
    .Y(_0276_));
 sg13g2_nand3_1 _0935_ (.B(_0271_),
    .C(_0276_),
    .A(_0267_),
    .Y(_0277_));
 sg13g2_nand2_1 _0936_ (.Y(_0278_),
    .A(_0261_),
    .B(_0255_));
 sg13g2_nor2_1 _0937_ (.A(_0246_),
    .B(_0278_),
    .Y(_0279_));
 sg13g2_nand2_1 _0938_ (.Y(_0280_),
    .A(net174),
    .B(_0279_));
 sg13g2_o21ai_1 _0939_ (.B1(_0280_),
    .Y(_0011_),
    .A1(_0263_),
    .A2(_0277_));
 sg13g2_nand2b_1 _0940_ (.Y(_0281_),
    .B(\i_dmi_jtag_tap.jtag_ir_q_0_ ),
    .A_N(\i_dmi_jtag_tap.jtag_ir_q_4_ ));
 sg13g2_nor3_1 _0941_ (.A(\i_dmi_jtag_tap.jtag_ir_q_1_ ),
    .B(\i_dmi_jtag_tap.jtag_ir_q_2_ ),
    .C(\i_dmi_jtag_tap.jtag_ir_q_3_ ),
    .Y(_0282_));
 sg13g2_nor2b_1 _0942_ (.A(_0281_),
    .B_N(_0282_),
    .Y(_0283_));
 sg13g2_nand2_1 _0943_ (.Y(_0284_),
    .A(_0269_),
    .B(_0283_));
 sg13g2_buf_2 fanout274 (.A(net276),
    .X(net274));
 sg13g2_nand2b_1 _0945_ (.Y(_0286_),
    .B(net252),
    .A_N(\i_dmi_jtag_tap.idcode_q_8_ ));
 sg13g2_nor3_2 _0946_ (.A(net319),
    .B(\i_dmi_jtag_tap.tap_state_q_1_ ),
    .C(_0248_),
    .Y(_0287_));
 sg13g2_and2_1 _0947_ (.A(_0283_),
    .B(net154),
    .X(_0288_));
 sg13g2_buf_2 fanout273 (.A(net277),
    .X(net273));
 sg13g2_buf_2 fanout272 (.A(net277),
    .X(net272));
 sg13g2_nand2b_1 _0950_ (.Y(_0291_),
    .B(net263),
    .A_N(\i_dmi_jtag_tap.idcode_q_9_ ));
 sg13g2_a21o_1 _0951_ (.A2(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .A1(net316),
    .B1(net317),
    .X(_0292_));
 sg13g2_a21oi_1 _0952_ (.A1(_0238_),
    .A2(_0292_),
    .Y(_0293_),
    .B1(net315));
 sg13g2_nor3_1 _0953_ (.A(_0260_),
    .B(_0256_),
    .C(_0293_),
    .Y(_0294_));
 sg13g2_buf_4 fanout271 (.X(net271),
    .A(net277));
 sg13g2_a21oi_1 _0955_ (.A1(_0286_),
    .A2(_0291_),
    .Y(_0020_),
    .B1(net238));
 sg13g2_nand2b_1 _0956_ (.Y(_0296_),
    .B(net252),
    .A_N(\i_dmi_jtag_tap.idcode_q_7_ ));
 sg13g2_nand2b_1 _0957_ (.Y(_0297_),
    .B(net264),
    .A_N(\i_dmi_jtag_tap.idcode_q_8_ ));
 sg13g2_a21oi_1 _0958_ (.A1(_0296_),
    .A2(_0297_),
    .Y(_0019_),
    .B1(net238));
 sg13g2_nand2b_1 _0959_ (.Y(_0298_),
    .B(net252),
    .A_N(\i_dmi_jtag_tap.idcode_q_5_ ));
 sg13g2_nand2b_1 _0960_ (.Y(_0299_),
    .B(net264),
    .A_N(\i_dmi_jtag_tap.idcode_q_6_ ));
 sg13g2_a21oi_1 _0961_ (.A1(_0298_),
    .A2(_0299_),
    .Y(_0018_),
    .B1(net242));
 sg13g2_nand2b_1 _0962_ (.Y(_0300_),
    .B(net252),
    .A_N(\i_dmi_jtag_tap.idcode_q_4_ ));
 sg13g2_nand2b_1 _0963_ (.Y(_0301_),
    .B(net264),
    .A_N(\i_dmi_jtag_tap.idcode_q_5_ ));
 sg13g2_a21oi_1 _0964_ (.A1(_0300_),
    .A2(_0301_),
    .Y(_0017_),
    .B1(net242));
 sg13g2_nand2b_1 _0965_ (.Y(_0302_),
    .B(net252),
    .A_N(\i_dmi_jtag_tap.idcode_q_1_ ));
 sg13g2_nand2b_1 _0966_ (.Y(_0303_),
    .B(net264),
    .A_N(\i_dmi_jtag_tap.idcode_q_2_ ));
 sg13g2_a21oi_1 _0967_ (.A1(_0302_),
    .A2(_0303_),
    .Y(_0016_),
    .B1(net242));
 sg13g2_nand2b_1 _0968_ (.Y(_0304_),
    .B(net249),
    .A_N(\i_dmi_jtag_tap.idcode_q_11_ ));
 sg13g2_nand2b_1 _0969_ (.Y(_0305_),
    .B(net261),
    .A_N(\i_dmi_jtag_tap.idcode_q_12_ ));
 sg13g2_a21oi_1 _0970_ (.A1(_0304_),
    .A2(_0305_),
    .Y(_0015_),
    .B1(net237));
 sg13g2_nand2b_1 _0971_ (.Y(_0306_),
    .B(net249),
    .A_N(\i_dmi_jtag_tap.idcode_q_10_ ));
 sg13g2_nand2b_1 _0972_ (.Y(_0307_),
    .B(net261),
    .A_N(\i_dmi_jtag_tap.idcode_q_11_ ));
 sg13g2_a21oi_1 _0973_ (.A1(_0306_),
    .A2(_0307_),
    .Y(_0014_),
    .B1(net237));
 sg13g2_nand2b_1 _0974_ (.Y(_0308_),
    .B(net253),
    .A_N(\i_dmi_jtag_tap.idcode_q_0_ ));
 sg13g2_nand2b_1 _0975_ (.Y(_0309_),
    .B(net265),
    .A_N(\i_dmi_jtag_tap.idcode_q_1_ ));
 sg13g2_a21oi_1 _0976_ (.A1(_0308_),
    .A2(_0309_),
    .Y(_0013_),
    .B1(net242));
 sg13g2_and2_1 _0977_ (.A(net448),
    .B(\i_dmi_cdc.core_clear_pending ),
    .X(_0012_));
 sg13g2_or4_1 _0978_ (.A(net319),
    .B(\i_dmi_jtag_tap.tap_state_q_1_ ),
    .C(net316),
    .D(net315),
    .X(_0310_));
 sg13g2_nor4_2 _0979_ (.A(\i_dmi_jtag_tap.jtag_ir_q_4__$_NOT__A_Y ),
    .B(\i_dmi_jtag_tap.jtag_ir_q_1_ ),
    .C(\i_dmi_jtag_tap.jtag_ir_q_2_ ),
    .Y(_0311_),
    .D(\i_dmi_jtag_tap.jtag_ir_q_3_ ));
 sg13g2_nand2b_1 _0980_ (.Y(_0312_),
    .B(_0311_),
    .A_N(\i_dmi_jtag_tap.jtag_ir_q_0_ ));
 sg13g2_nor2_1 _0981_ (.A(_0310_),
    .B(_0312_),
    .Y(_0313_));
 sg13g2_a21o_2 _0982_ (.A2(_0313_),
    .A1(dtmcs_q_17_),
    .B1(net241),
    .X(_0314_));
 sg13g2_buf_2 fanout270 (.A(_0353_),
    .X(net270));
 sg13g2_buf_2 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_1 fanout268 (.A(net270),
    .X(net268));
 sg13g2_buf_2 fanout267 (.A(net270),
    .X(net267));
 sg13g2_buf_2 fanout266 (.A(_0412_),
    .X(net266));
 sg13g2_and2_1 _0988_ (.A(\i_dmi_jtag_tap.jtag_ir_q_0_ ),
    .B(_0311_),
    .X(_0319_));
 sg13g2_nor2_2 _0989_ (.A(error_q_0_),
    .B(error_q_1_),
    .Y(_0320_));
 sg13g2_nand3b_1 _0990_ (.B(net173),
    .C(_0320_),
    .Y(_0321_),
    .A_N(_0310_));
 sg13g2_nor4_2 _0991_ (.A(state_q_2_),
    .B(state_q_0_),
    .C(state_q_1_),
    .Y(_0322_),
    .D(_0321_));
 sg13g2_buf_2 fanout265 (.A(_0288_),
    .X(net265));
 sg13g2_nor2b_1 _0993_ (.A(net259),
    .B_N(address_q_0_),
    .Y(_0324_));
 sg13g2_a21oi_1 _0994_ (.A1(dmi_34_),
    .A2(net259),
    .Y(_0325_),
    .B1(_0324_));
 sg13g2_nor2_1 _0995_ (.A(net233),
    .B(_0325_),
    .Y(_0027_));
 sg13g2_nor2b_1 _0996_ (.A(net259),
    .B_N(address_q_1_),
    .Y(_0326_));
 sg13g2_a21oi_1 _0997_ (.A1(dmi_35_),
    .A2(net259),
    .Y(_0327_),
    .B1(_0326_));
 sg13g2_nor2_1 _0998_ (.A(net233),
    .B(_0327_),
    .Y(_0028_));
 sg13g2_buf_2 fanout264 (.A(net265),
    .X(net264));
 sg13g2_nor2b_1 _1000_ (.A(net260),
    .B_N(address_q_2_),
    .Y(_0329_));
 sg13g2_a21oi_1 _1001_ (.A1(dmi_36_),
    .A2(net260),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_nor2_1 _1002_ (.A(net236),
    .B(_0330_),
    .Y(_0029_));
 sg13g2_nor2b_1 _1003_ (.A(net259),
    .B_N(address_q_3_),
    .Y(_0331_));
 sg13g2_a21oi_1 _1004_ (.A1(dmi_37_),
    .A2(net259),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_nor2_1 _1005_ (.A(net234),
    .B(_0332_),
    .Y(_0030_));
 sg13g2_nor2b_1 _1006_ (.A(net259),
    .B_N(address_q_4_),
    .Y(_0333_));
 sg13g2_a21oi_1 _1007_ (.A1(dmi_38_),
    .A2(net259),
    .Y(_0334_),
    .B1(_0333_));
 sg13g2_nor2_1 _1008_ (.A(net234),
    .B(_0334_),
    .Y(_0031_));
 sg13g2_nor2b_1 _1009_ (.A(net260),
    .B_N(address_q_5_),
    .Y(_0335_));
 sg13g2_a21oi_1 _1010_ (.A1(dmi_39_),
    .A2(net260),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_nor2_1 _1011_ (.A(net236),
    .B(_0336_),
    .Y(_0032_));
 sg13g2_nor2b_1 _1012_ (.A(net260),
    .B_N(address_q_6_),
    .Y(_0337_));
 sg13g2_a21oi_1 _1013_ (.A1(dmi_40_),
    .A2(net260),
    .Y(_0338_),
    .B1(_0337_));
 sg13g2_nor2_1 _1014_ (.A(net235),
    .B(_0338_),
    .Y(_0033_));
 sg13g2_nor3_2 _1015_ (.A(state_q_2_),
    .B(state_q_0_),
    .C(state_q_1_),
    .Y(_0339_));
 sg13g2_nand2_2 _1016_ (.Y(_0340_),
    .A(_0339_),
    .B(_0321_));
 sg13g2_nor2_1 _1017_ (.A(state_q_2_),
    .B(\state_q_1__$_NOT__A_Y ),
    .Y(_0341_));
 sg13g2_nand2b_1 _1018_ (.Y(_0342_),
    .B(_0341_),
    .A_N(state_q_0_));
 sg13g2_mux2_1 _1019_ (.A0(dmi_resp_valid),
    .A1(_0339_),
    .S(net273),
    .X(_0343_));
 sg13g2_nand2_1 _1020_ (.Y(_0344_),
    .A(_0340_),
    .B(_0343_));
 sg13g2_buf_2 fanout263 (.A(net265),
    .X(net263));
 sg13g2_nand2_1 _1022_ (.Y(_0346_),
    .A(data_q_0_),
    .B(net217));
 sg13g2_inv_1 _1023_ (.Y(_0347_),
    .A(dmi_resp_0_));
 sg13g2_buf_2 fanout262 (.A(net263),
    .X(net262));
 sg13g2_buf_2 fanout261 (.A(net263),
    .X(net261));
 sg13g2_buf_1 fanout260 (.A(_0322_),
    .X(net260));
 sg13g2_a21oi_1 _1027_ (.A1(net312),
    .A2(dmi_resp_2_),
    .Y(_0351_),
    .B1(net321));
 sg13g2_or2_1 _1028_ (.X(_0352_),
    .B(\state_q_1__$_NOT__A_Y ),
    .A(state_q_2_));
 sg13g2_nor2_1 _1029_ (.A(state_q_0_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_buf_2 fanout259 (.A(_0322_),
    .X(net259));
 sg13g2_nor2_1 _1031_ (.A(dmi_2_),
    .B(net267),
    .Y(_0355_));
 sg13g2_a21oi_1 _1032_ (.A1(_0351_),
    .A2(net267),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_and2_1 _1033_ (.A(_0340_),
    .B(_0343_),
    .X(_0357_));
 sg13g2_buf_2 fanout258 (.A(_0097_),
    .X(net258));
 sg13g2_buf_2 fanout257 (.A(net258),
    .X(net257));
 sg13g2_nand2_1 _1036_ (.Y(_0360_),
    .A(_0356_),
    .B(net211));
 sg13g2_a21oi_1 _1037_ (.A1(_0346_),
    .A2(_0360_),
    .Y(_0034_),
    .B1(net223));
 sg13g2_buf_2 fanout256 (.A(net258),
    .X(net256));
 sg13g2_buf_2 fanout255 (.A(net256),
    .X(net255));
 sg13g2_nor2_1 _1040_ (.A(data_q_10_),
    .B(net210),
    .Y(_0363_));
 sg13g2_buf_2 fanout254 (.A(net256),
    .X(net254));
 sg13g2_buf_1 fanout253 (.A(_0284_),
    .X(net253));
 sg13g2_o21ai_1 _1043_ (.B1(net313),
    .Y(_0366_),
    .A1(dmi_resp_12_),
    .A2(net322));
 sg13g2_nor2_1 _1044_ (.A(net273),
    .B(_0366_),
    .Y(_0367_));
 sg13g2_a21oi_1 _1045_ (.A1(dmi_12_),
    .A2(net272),
    .Y(_0368_),
    .B1(_0367_));
 sg13g2_and2_1 _1046_ (.A(net210),
    .B(_0368_),
    .X(_0369_));
 sg13g2_nor3_1 _1047_ (.A(net222),
    .B(_0363_),
    .C(_0369_),
    .Y(_0035_));
 sg13g2_nor2_1 _1048_ (.A(data_q_11_),
    .B(net210),
    .Y(_0370_));
 sg13g2_o21ai_1 _1049_ (.B1(net312),
    .Y(_0371_),
    .A1(dmi_resp_13_),
    .A2(net321));
 sg13g2_nor2_1 _1050_ (.A(net272),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_a21oi_1 _1051_ (.A1(dmi_13_),
    .A2(net272),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_and2_1 _1052_ (.A(net210),
    .B(_0373_),
    .X(_0374_));
 sg13g2_nor3_1 _1053_ (.A(net221),
    .B(_0370_),
    .C(_0374_),
    .Y(_0036_));
 sg13g2_nand2_1 _1054_ (.Y(_0375_),
    .A(data_q_12_),
    .B(net216));
 sg13g2_a21oi_1 _1055_ (.A1(net313),
    .A2(dmi_resp_14_),
    .Y(_0376_),
    .B1(net322));
 sg13g2_nor2_1 _1056_ (.A(dmi_14_),
    .B(net268),
    .Y(_0377_));
 sg13g2_a21oi_1 _1057_ (.A1(net268),
    .A2(_0376_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_nand2_1 _1058_ (.Y(_0379_),
    .A(net212),
    .B(_0378_));
 sg13g2_a21oi_1 _1059_ (.A1(_0375_),
    .A2(_0379_),
    .Y(_0037_),
    .B1(net221));
 sg13g2_nand2_1 _1060_ (.Y(_0380_),
    .A(data_q_13_),
    .B(net216));
 sg13g2_a21oi_1 _1061_ (.A1(net313),
    .A2(dmi_resp_15_),
    .Y(_0381_),
    .B1(net322));
 sg13g2_buf_2 fanout252 (.A(net253),
    .X(net252));
 sg13g2_nor2_1 _1063_ (.A(dmi_15_),
    .B(net268),
    .Y(_0383_));
 sg13g2_a21oi_1 _1064_ (.A1(net267),
    .A2(_0381_),
    .Y(_0384_),
    .B1(_0383_));
 sg13g2_nand2_1 _1065_ (.Y(_0385_),
    .A(net212),
    .B(_0384_));
 sg13g2_a21oi_1 _1066_ (.A1(_0380_),
    .A2(_0385_),
    .Y(_0038_),
    .B1(net224));
 sg13g2_nor2_1 _1067_ (.A(data_q_14_),
    .B(net213),
    .Y(_0386_));
 sg13g2_nor2_2 _1068_ (.A(dmi_resp_0_),
    .B(dmi_resp_16_),
    .Y(_0387_));
 sg13g2_nor3_2 _1069_ (.A(net323),
    .B(net271),
    .C(_0387_),
    .Y(_0388_));
 sg13g2_a21oi_1 _1070_ (.A1(dmi_16_),
    .A2(net273),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_and2_1 _1071_ (.A(net212),
    .B(_0389_),
    .X(_0390_));
 sg13g2_nor3_1 _1072_ (.A(net225),
    .B(_0386_),
    .C(_0390_),
    .Y(_0039_));
 sg13g2_nand2_1 _1073_ (.Y(_0391_),
    .A(data_q_15_),
    .B(net216));
 sg13g2_buf_2 fanout251 (.A(_0284_),
    .X(net251));
 sg13g2_nor2_1 _1075_ (.A(dmi_17_),
    .B(net270),
    .Y(_0393_));
 sg13g2_or2_1 _1076_ (.X(_0394_),
    .B(net323),
    .A(dmi_resp_0_));
 sg13g2_buf_2 fanout250 (.A(net251),
    .X(net250));
 sg13g2_nor3_2 _1078_ (.A(dmi_resp_17_),
    .B(net271),
    .C(net311),
    .Y(_0396_));
 sg13g2_or3_1 _1079_ (.A(net216),
    .B(_0393_),
    .C(_0396_),
    .X(_0397_));
 sg13g2_a21oi_1 _1080_ (.A1(_0391_),
    .A2(_0397_),
    .Y(_0040_),
    .B1(net224));
 sg13g2_nand2_1 _1081_ (.Y(_0398_),
    .A(data_q_16_),
    .B(net218));
 sg13g2_nor2_1 _1082_ (.A(dmi_18_),
    .B(net270),
    .Y(_0399_));
 sg13g2_nor3_2 _1083_ (.A(dmi_resp_18_),
    .B(net271),
    .C(net310),
    .Y(_0400_));
 sg13g2_or3_1 _1084_ (.A(net218),
    .B(_0399_),
    .C(_0400_),
    .X(_0401_));
 sg13g2_a21oi_1 _1085_ (.A1(_0398_),
    .A2(_0401_),
    .Y(_0041_),
    .B1(net228));
 sg13g2_nor2_1 _1086_ (.A(data_q_17_),
    .B(net214),
    .Y(_0402_));
 sg13g2_buf_2 fanout249 (.A(net251),
    .X(net249));
 sg13g2_nand2_1 _1088_ (.Y(_0404_),
    .A(dmi_19_),
    .B(net275));
 sg13g2_nor2_2 _1089_ (.A(dmi_resp_0_),
    .B(net321),
    .Y(_0405_));
 sg13g2_nand3_1 _1090_ (.B(net267),
    .C(_0405_),
    .A(dmi_resp_19_),
    .Y(_0406_));
 sg13g2_and3_1 _1091_ (.X(_0407_),
    .A(net212),
    .B(_0404_),
    .C(_0406_));
 sg13g2_nor3_1 _1092_ (.A(net230),
    .B(_0402_),
    .C(_0407_),
    .Y(_0042_));
 sg13g2_buf_1 fanout248 (.A(_0099_),
    .X(net248));
 sg13g2_nor2_1 _1094_ (.A(data_q_18_),
    .B(net212),
    .Y(_0409_));
 sg13g2_buf_2 fanout247 (.A(net248),
    .X(net247));
 sg13g2_buf_2 fanout246 (.A(net248),
    .X(net246));
 sg13g2_nand2_1 _1097_ (.Y(_0412_),
    .A(dmi_resp_0_),
    .B(net323));
 sg13g2_o21ai_1 _1098_ (.B1(net266),
    .Y(_0413_),
    .A1(dmi_resp_20_),
    .A2(net311));
 sg13g2_nand2_1 _1099_ (.Y(_0414_),
    .A(dmi_20_),
    .B(net273));
 sg13g2_o21ai_1 _1100_ (.B1(_0414_),
    .Y(_0415_),
    .A1(net273),
    .A2(_0413_));
 sg13g2_nor2_1 _1101_ (.A(net217),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nor3_1 _1102_ (.A(net225),
    .B(_0409_),
    .C(_0416_),
    .Y(_0043_));
 sg13g2_nor2_1 _1103_ (.A(data_q_19_),
    .B(net211),
    .Y(_0417_));
 sg13g2_o21ai_1 _1104_ (.B1(net266),
    .Y(_0418_),
    .A1(dmi_resp_21_),
    .A2(net310));
 sg13g2_nand2_1 _1105_ (.Y(_0419_),
    .A(dmi_21_),
    .B(net274));
 sg13g2_o21ai_1 _1106_ (.B1(_0419_),
    .Y(_0420_),
    .A1(net274),
    .A2(_0418_));
 sg13g2_nor2_1 _1107_ (.A(net217),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_nor3_1 _1108_ (.A(net228),
    .B(_0417_),
    .C(_0421_),
    .Y(_0044_));
 sg13g2_nor2_1 _1109_ (.A(data_q_1_),
    .B(net214),
    .Y(_0422_));
 sg13g2_o21ai_1 _1110_ (.B1(net266),
    .Y(_0423_),
    .A1(dmi_resp_3_),
    .A2(net310));
 sg13g2_nand2_1 _1111_ (.Y(_0424_),
    .A(dmi_3_),
    .B(net274));
 sg13g2_o21ai_1 _1112_ (.B1(_0424_),
    .Y(_0425_),
    .A1(net276),
    .A2(_0423_));
 sg13g2_nor2_1 _1113_ (.A(net219),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_nor3_1 _1114_ (.A(net233),
    .B(_0422_),
    .C(_0426_),
    .Y(_0045_));
 sg13g2_nand2_1 _1115_ (.Y(_0427_),
    .A(data_q_20_),
    .B(net217));
 sg13g2_and2_1 _1116_ (.A(dmi_resp_0_),
    .B(net321),
    .X(_0428_));
 sg13g2_a21oi_1 _1117_ (.A1(dmi_resp_22_),
    .A2(_0405_),
    .Y(_0429_),
    .B1(_0428_));
 sg13g2_nor2_1 _1118_ (.A(dmi_22_),
    .B(net269),
    .Y(_0430_));
 sg13g2_a21oi_1 _1119_ (.A1(net269),
    .A2(_0429_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_nand2_1 _1120_ (.Y(_0432_),
    .A(net211),
    .B(_0431_));
 sg13g2_a21oi_1 _1121_ (.A1(_0427_),
    .A2(_0432_),
    .Y(_0046_),
    .B1(net223));
 sg13g2_nor2_1 _1122_ (.A(data_q_21_),
    .B(net212),
    .Y(_0433_));
 sg13g2_o21ai_1 _1123_ (.B1(net266),
    .Y(_0434_),
    .A1(dmi_resp_23_),
    .A2(net311));
 sg13g2_nand2_1 _1124_ (.Y(_0435_),
    .A(dmi_23_),
    .B(net273));
 sg13g2_o21ai_1 _1125_ (.B1(_0435_),
    .Y(_0436_),
    .A1(net273),
    .A2(_0434_));
 sg13g2_nor2_1 _1126_ (.A(net216),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_nor3_1 _1127_ (.A(net225),
    .B(_0433_),
    .C(_0437_),
    .Y(_0047_));
 sg13g2_nand2_1 _1128_ (.Y(_0438_),
    .A(data_q_22_),
    .B(net218));
 sg13g2_a21oi_1 _1129_ (.A1(dmi_resp_24_),
    .A2(_0405_),
    .Y(_0439_),
    .B1(_0428_));
 sg13g2_nor2_1 _1130_ (.A(dmi_24_),
    .B(net269),
    .Y(_0440_));
 sg13g2_a21oi_1 _1131_ (.A1(net269),
    .A2(_0439_),
    .Y(_0441_),
    .B1(_0440_));
 sg13g2_nand2_1 _1132_ (.Y(_0442_),
    .A(net212),
    .B(_0441_));
 sg13g2_a21oi_1 _1133_ (.A1(_0438_),
    .A2(_0442_),
    .Y(_0048_),
    .B1(net230));
 sg13g2_nor2_1 _1134_ (.A(data_q_23_),
    .B(net214),
    .Y(_0443_));
 sg13g2_o21ai_1 _1135_ (.B1(net266),
    .Y(_0444_),
    .A1(dmi_resp_25_),
    .A2(net310));
 sg13g2_nand2_1 _1136_ (.Y(_0445_),
    .A(dmi_25_),
    .B(net274));
 sg13g2_o21ai_1 _1137_ (.B1(_0445_),
    .Y(_0446_),
    .A1(net276),
    .A2(_0444_));
 sg13g2_nor2_1 _1138_ (.A(net219),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_nor3_1 _1139_ (.A(net229),
    .B(_0443_),
    .C(_0447_),
    .Y(_0049_));
 sg13g2_nor2_1 _1140_ (.A(data_q_24_),
    .B(net214),
    .Y(_0448_));
 sg13g2_nand2_1 _1141_ (.Y(_0449_),
    .A(dmi_26_),
    .B(net274));
 sg13g2_nand3_1 _1142_ (.B(net267),
    .C(_0405_),
    .A(dmi_resp_26_),
    .Y(_0450_));
 sg13g2_and3_1 _1143_ (.X(_0451_),
    .A(net214),
    .B(_0449_),
    .C(_0450_));
 sg13g2_nor3_1 _1144_ (.A(net229),
    .B(_0448_),
    .C(_0451_),
    .Y(_0050_));
 sg13g2_buf_2 fanout245 (.A(net246),
    .X(net245));
 sg13g2_nor2_1 _1146_ (.A(data_q_25_),
    .B(net215),
    .Y(_0453_));
 sg13g2_o21ai_1 _1147_ (.B1(net266),
    .Y(_0454_),
    .A1(dmi_resp_27_),
    .A2(net311));
 sg13g2_nand2_1 _1148_ (.Y(_0455_),
    .A(dmi_27_),
    .B(net275));
 sg13g2_o21ai_1 _1149_ (.B1(_0455_),
    .Y(_0456_),
    .A1(net276),
    .A2(_0454_));
 sg13g2_nor2_1 _1150_ (.A(net219),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor3_1 _1151_ (.A(net235),
    .B(_0453_),
    .C(_0457_),
    .Y(_0051_));
 sg13g2_nor2_1 _1152_ (.A(data_q_26_),
    .B(net215),
    .Y(_0458_));
 sg13g2_o21ai_1 _1153_ (.B1(net313),
    .Y(_0459_),
    .A1(net322),
    .A2(dmi_resp_28_));
 sg13g2_nor2_1 _1154_ (.A(net275),
    .B(_0459_),
    .Y(_0460_));
 sg13g2_a21oi_1 _1155_ (.A1(dmi_28_),
    .A2(net275),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_and2_1 _1156_ (.A(net214),
    .B(_0461_),
    .X(_0462_));
 sg13g2_nor3_1 _1157_ (.A(net231),
    .B(_0458_),
    .C(_0462_),
    .Y(_0052_));
 sg13g2_nor2_1 _1158_ (.A(data_q_27_),
    .B(net215),
    .Y(_0463_));
 sg13g2_o21ai_1 _1159_ (.B1(_0412_),
    .Y(_0464_),
    .A1(dmi_resp_29_),
    .A2(net311));
 sg13g2_nand2_1 _1160_ (.Y(_0465_),
    .A(dmi_29_),
    .B(net275));
 sg13g2_o21ai_1 _1161_ (.B1(_0465_),
    .Y(_0466_),
    .A1(net275),
    .A2(_0464_));
 sg13g2_nor2_1 _1162_ (.A(net220),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_nor3_1 _1163_ (.A(net235),
    .B(_0463_),
    .C(_0467_),
    .Y(_0053_));
 sg13g2_nand2_1 _1164_ (.Y(_0468_),
    .A(data_q_28_),
    .B(net218));
 sg13g2_nor2_1 _1165_ (.A(dmi_30_),
    .B(net269),
    .Y(_0469_));
 sg13g2_nor3_2 _1166_ (.A(dmi_resp_30_),
    .B(net271),
    .C(net310),
    .Y(_0470_));
 sg13g2_or3_1 _1167_ (.A(net218),
    .B(_0469_),
    .C(_0470_),
    .X(_0471_));
 sg13g2_a21oi_1 _1168_ (.A1(_0468_),
    .A2(_0471_),
    .Y(_0054_),
    .B1(net230));
 sg13g2_nand2_1 _1169_ (.Y(_0472_),
    .A(data_q_29_),
    .B(net218));
 sg13g2_nand2b_2 _1170_ (.Y(_0473_),
    .B(dmi_resp_31_),
    .A_N(net324));
 sg13g2_nand3_1 _1171_ (.B(net267),
    .C(_0473_),
    .A(net312),
    .Y(_0474_));
 sg13g2_o21ai_1 _1172_ (.B1(_0474_),
    .Y(_0475_),
    .A1(dmi_31_),
    .A2(net269));
 sg13g2_or2_1 _1173_ (.X(_0476_),
    .B(_0475_),
    .A(net218));
 sg13g2_a21oi_1 _1174_ (.A1(_0472_),
    .A2(_0476_),
    .Y(_0055_),
    .B1(net230));
 sg13g2_nor2_1 _1175_ (.A(data_q_2_),
    .B(net215),
    .Y(_0477_));
 sg13g2_o21ai_1 _1176_ (.B1(_0412_),
    .Y(_0478_),
    .A1(dmi_resp_4_),
    .A2(net311));
 sg13g2_nand2_1 _1177_ (.Y(_0479_),
    .A(dmi_4_),
    .B(net275));
 sg13g2_o21ai_1 _1178_ (.B1(_0479_),
    .Y(_0480_),
    .A1(net275),
    .A2(_0478_));
 sg13g2_nor2_1 _1179_ (.A(net220),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_nor3_1 _1180_ (.A(net233),
    .B(_0477_),
    .C(_0481_),
    .Y(_0056_));
 sg13g2_nor2_1 _1181_ (.A(data_q_30_),
    .B(net214),
    .Y(_0482_));
 sg13g2_o21ai_1 _1182_ (.B1(net312),
    .Y(_0483_),
    .A1(net321),
    .A2(dmi_resp_32_));
 sg13g2_nor2_1 _1183_ (.A(net277),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_a21oi_1 _1184_ (.A1(dmi_32_),
    .A2(net274),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_and2_1 _1185_ (.A(net214),
    .B(_0485_),
    .X(_0486_));
 sg13g2_nor3_1 _1186_ (.A(net228),
    .B(_0482_),
    .C(_0486_),
    .Y(_0057_));
 sg13g2_nand2_1 _1187_ (.Y(_0487_),
    .A(data_q_31_),
    .B(net219));
 sg13g2_nor2_1 _1188_ (.A(dmi_33_),
    .B(net269),
    .Y(_0488_));
 sg13g2_nor3_2 _1189_ (.A(dmi_resp_33_),
    .B(net271),
    .C(net310),
    .Y(_0489_));
 sg13g2_or3_1 _1190_ (.A(net219),
    .B(_0488_),
    .C(_0489_),
    .X(_0490_));
 sg13g2_a21oi_1 _1191_ (.A1(_0487_),
    .A2(_0490_),
    .Y(_0058_),
    .B1(net229));
 sg13g2_nor2_1 _1192_ (.A(data_q_3_),
    .B(net215),
    .Y(_0491_));
 sg13g2_o21ai_1 _1193_ (.B1(net266),
    .Y(_0492_),
    .A1(dmi_resp_5_),
    .A2(net310));
 sg13g2_nand2_1 _1194_ (.Y(_0493_),
    .A(dmi_5_),
    .B(net274));
 sg13g2_o21ai_1 _1195_ (.B1(_0493_),
    .Y(_0494_),
    .A1(net274),
    .A2(_0492_));
 sg13g2_nor2_1 _1196_ (.A(net218),
    .B(_0494_),
    .Y(_0495_));
 sg13g2_nor3_1 _1197_ (.A(net235),
    .B(_0491_),
    .C(_0495_),
    .Y(_0059_));
 sg13g2_nand2_1 _1198_ (.Y(_0496_),
    .A(data_q_4_),
    .B(net219));
 sg13g2_nand2b_2 _1199_ (.Y(_0497_),
    .B(dmi_resp_6_),
    .A_N(net324));
 sg13g2_nand3_1 _1200_ (.B(net267),
    .C(_0497_),
    .A(net312),
    .Y(_0498_));
 sg13g2_o21ai_1 _1201_ (.B1(_0498_),
    .Y(_0499_),
    .A1(dmi_6_),
    .A2(net269));
 sg13g2_or2_1 _1202_ (.X(_0500_),
    .B(_0499_),
    .A(net219));
 sg13g2_a21oi_1 _1203_ (.A1(_0496_),
    .A2(_0500_),
    .Y(_0060_),
    .B1(net228));
 sg13g2_nor2_1 _1204_ (.A(data_q_5_),
    .B(net211),
    .Y(_0501_));
 sg13g2_o21ai_1 _1205_ (.B1(net312),
    .Y(_0502_),
    .A1(net321),
    .A2(dmi_resp_7_));
 sg13g2_nor2_1 _1206_ (.A(net271),
    .B(_0502_),
    .Y(_0503_));
 sg13g2_a21oi_1 _1207_ (.A1(dmi_7_),
    .A2(net272),
    .Y(_0504_),
    .B1(_0503_));
 sg13g2_and2_1 _1208_ (.A(net210),
    .B(_0504_),
    .X(_0505_));
 sg13g2_nor3_1 _1209_ (.A(net223),
    .B(_0501_),
    .C(_0505_),
    .Y(_0061_));
 sg13g2_nand2_1 _1210_ (.Y(_0506_),
    .A(data_q_6_),
    .B(net216));
 sg13g2_nor2_1 _1211_ (.A(dmi_8_),
    .B(net268),
    .Y(_0507_));
 sg13g2_nor3_2 _1212_ (.A(dmi_resp_8_),
    .B(net271),
    .C(net311),
    .Y(_0508_));
 sg13g2_or3_1 _1213_ (.A(net216),
    .B(_0507_),
    .C(_0508_),
    .X(_0509_));
 sg13g2_a21oi_1 _1214_ (.A1(_0506_),
    .A2(_0509_),
    .Y(_0062_),
    .B1(net224));
 sg13g2_nor2_1 _1215_ (.A(data_q_7_),
    .B(net212),
    .Y(_0510_));
 sg13g2_o21ai_1 _1216_ (.B1(net266),
    .Y(_0511_),
    .A1(dmi_resp_9_),
    .A2(net310));
 sg13g2_nand2_1 _1217_ (.Y(_0512_),
    .A(dmi_9_),
    .B(net272));
 sg13g2_o21ai_1 _1218_ (.B1(_0512_),
    .Y(_0513_),
    .A1(net272),
    .A2(_0511_));
 sg13g2_nor2_1 _1219_ (.A(net216),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_nor3_1 _1220_ (.A(net224),
    .B(_0510_),
    .C(_0514_),
    .Y(_0063_));
 sg13g2_nor2_1 _1221_ (.A(data_q_8_),
    .B(net210),
    .Y(_0515_));
 sg13g2_nand2_1 _1222_ (.Y(_0516_),
    .A(dmi_10_),
    .B(net272));
 sg13g2_nand3_1 _1223_ (.B(net267),
    .C(_0405_),
    .A(dmi_resp_10_),
    .Y(_0517_));
 sg13g2_and3_1 _1224_ (.X(_0518_),
    .A(net210),
    .B(_0516_),
    .C(_0517_));
 sg13g2_nor3_1 _1225_ (.A(net222),
    .B(_0515_),
    .C(_0518_),
    .Y(_0064_));
 sg13g2_nor2_1 _1226_ (.A(data_q_9_),
    .B(net211),
    .Y(_0519_));
 sg13g2_o21ai_1 _1227_ (.B1(net312),
    .Y(_0520_),
    .A1(dmi_resp_11_),
    .A2(net321));
 sg13g2_nor2_1 _1228_ (.A(net271),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_a21oi_1 _1229_ (.A1(dmi_11_),
    .A2(net272),
    .Y(_0522_),
    .B1(_0521_));
 sg13g2_and2_1 _1230_ (.A(net210),
    .B(_0522_),
    .X(_0523_));
 sg13g2_nor3_1 _1231_ (.A(net222),
    .B(_0519_),
    .C(_0523_),
    .Y(_0065_));
 sg13g2_nor2_2 _1232_ (.A(\state_q_0__$_NOT__A_Y ),
    .B(_0352_),
    .Y(dmi_req_33_));
 sg13g2_inv_1 _1233_ (.Y(dmi_req_32_),
    .A(dmi_req_33_));
 sg13g2_and2_1 _1234_ (.A(\state_q_1__$_NOT__A_Y ),
    .B(state_q_1_),
    .X(_0524_));
 sg13g2_or3_1 _1235_ (.A(state_q_2_),
    .B(\state_q_0__$_NOT__A_Y ),
    .C(_0524_),
    .X(_0525_));
 sg13g2_nor2_1 _1236_ (.A(net224),
    .B(_0525_),
    .Y(dmi_req_valid));
 sg13g2_buf_2 fanout244 (.A(net246),
    .X(net244));
 sg13g2_buf_1 fanout243 (.A(_0294_),
    .X(net243));
 sg13g2_buf_2 fanout242 (.A(net243),
    .X(net242));
 sg13g2_nand3_1 _1240_ (.B(net154),
    .C(net168),
    .A(dmi_1_),
    .Y(_0529_));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_nor3_2 _1242_ (.A(net316),
    .B(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .C(_0257_),
    .Y(_0531_));
 sg13g2_or2_1 _1243_ (.X(_0532_),
    .B(state_q_0_),
    .A(\state_q_1__$_NOT__A_Y ));
 sg13g2_or2_1 _1244_ (.X(_0533_),
    .B(state_q_1_),
    .A(\state_q_0__$_NOT__A_Y ));
 sg13g2_a21oi_1 _1245_ (.A1(_0532_),
    .A2(_0533_),
    .Y(_0534_),
    .B1(state_q_2_));
 sg13g2_or2_1 _1246_ (.X(_0535_),
    .B(\state_q_0__$_OR__A_Y_$_OR__A_1_B ),
    .A(state_q_1_));
 sg13g2_nand2b_1 _1247_ (.Y(_0536_),
    .B(dmi_resp_valid),
    .A_N(state_q_0_));
 sg13g2_a21oi_1 _1248_ (.A1(_0352_),
    .A2(_0535_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_nor2_1 _1249_ (.A(_0310_),
    .B(_0339_),
    .Y(_0538_));
 sg13g2_a221oi_1 _1250_ (.B2(_0428_),
    .C1(_0538_),
    .B1(_0537_),
    .A1(_0531_),
    .Y(_0539_),
    .A2(_0534_));
 sg13g2_or2_1 _1251_ (.X(_0540_),
    .B(\error_q_1__$_NOT__A_Y ),
    .A(\error_q_0__$_NOT__A_Y ));
 sg13g2_nand2_1 _1252_ (.Y(_0541_),
    .A(net172),
    .B(_0531_));
 sg13g2_a21oi_1 _1253_ (.A1(_0539_),
    .A2(_0540_),
    .Y(_0542_),
    .B1(_0541_));
 sg13g2_nand4_1 _1254_ (.B(_0320_),
    .C(_0531_),
    .A(net173),
    .Y(_0543_),
    .D(_0539_));
 sg13g2_o21ai_1 _1255_ (.B1(_0543_),
    .Y(_0544_),
    .A1(dmi_0_),
    .A2(_0542_));
 sg13g2_a21o_1 _1256_ (.A2(net173),
    .A1(net161),
    .B1(_0544_),
    .X(_0545_));
 sg13g2_a21oi_1 _1257_ (.A1(_0529_),
    .A2(_0545_),
    .Y(dr_d_0_),
    .B1(net221));
 sg13g2_buf_2 fanout240 (.A(net243),
    .X(net240));
 sg13g2_nor2b_1 _1259_ (.A(_0320_),
    .B_N(_0540_),
    .Y(_0547_));
 sg13g2_a21oi_1 _1260_ (.A1(_0539_),
    .A2(_0547_),
    .Y(_0548_),
    .B1(_0541_));
 sg13g2_buf_2 fanout239 (.A(net240),
    .X(net239));
 sg13g2_buf_2 fanout238 (.A(net243),
    .X(net238));
 sg13g2_mux2_1 _1263_ (.A0(dmi_10_),
    .A1(data_q_8_),
    .S(net192),
    .X(_0551_));
 sg13g2_nand2_1 _1264_ (.Y(_0552_),
    .A(\i_dmi_jtag_tap.jtag_ir_q_0_ ),
    .B(_0311_));
 sg13g2_buf_2 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_2 fanout236 (.A(_0314_),
    .X(net236));
 sg13g2_nand2_1 _1267_ (.Y(_0555_),
    .A(dmi_10_),
    .B(net303));
 sg13g2_nand2_1 _1268_ (.Y(_0556_),
    .A(dmi_11_),
    .B(net168));
 sg13g2_nand3_1 _1269_ (.B(_0555_),
    .C(_0556_),
    .A(net160),
    .Y(_0557_));
 sg13g2_o21ai_1 _1270_ (.B1(_0557_),
    .Y(_0558_),
    .A1(net156),
    .A2(_0551_));
 sg13g2_nor2_1 _1271_ (.A(net222),
    .B(_0558_),
    .Y(dr_d_10_));
 sg13g2_mux2_1 _1272_ (.A0(dmi_11_),
    .A1(data_q_9_),
    .S(net192),
    .X(_0559_));
 sg13g2_nand2_1 _1273_ (.Y(_0560_),
    .A(dmi_12_),
    .B(net168));
 sg13g2_nand2_1 _1274_ (.Y(_0561_),
    .A(dmi_11_),
    .B(net303));
 sg13g2_nand3_1 _1275_ (.B(_0560_),
    .C(_0561_),
    .A(net160),
    .Y(_0562_));
 sg13g2_o21ai_1 _1276_ (.B1(_0562_),
    .Y(_0563_),
    .A1(net156),
    .A2(_0559_));
 sg13g2_nor2_1 _1277_ (.A(net222),
    .B(_0563_),
    .Y(dr_d_11_));
 sg13g2_mux2_1 _1278_ (.A0(dmi_12_),
    .A1(data_q_10_),
    .S(net192),
    .X(_0564_));
 sg13g2_nand2_1 _1279_ (.Y(_0565_),
    .A(dmi_12_),
    .B(net303));
 sg13g2_nand2_1 _1280_ (.Y(_0566_),
    .A(dmi_13_),
    .B(net167));
 sg13g2_nand3_1 _1281_ (.B(_0565_),
    .C(_0566_),
    .A(net160),
    .Y(_0567_));
 sg13g2_o21ai_1 _1282_ (.B1(_0567_),
    .Y(_0568_),
    .A1(net155),
    .A2(_0564_));
 sg13g2_nor2_1 _1283_ (.A(net222),
    .B(_0568_),
    .Y(dr_d_12_));
 sg13g2_mux2_1 _1284_ (.A0(dmi_13_),
    .A1(data_q_11_),
    .S(net192),
    .X(_0569_));
 sg13g2_nand2_1 _1285_ (.Y(_0570_),
    .A(dmi_13_),
    .B(net303));
 sg13g2_nand2_1 _1286_ (.Y(_0571_),
    .A(dmi_14_),
    .B(net167));
 sg13g2_nand3_1 _1287_ (.B(_0570_),
    .C(_0571_),
    .A(net160),
    .Y(_0572_));
 sg13g2_o21ai_1 _1288_ (.B1(_0572_),
    .Y(_0573_),
    .A1(net155),
    .A2(_0569_));
 sg13g2_nor2_1 _1289_ (.A(net222),
    .B(_0573_),
    .Y(dr_d_13_));
 sg13g2_buf_2 fanout235 (.A(net236),
    .X(net235));
 sg13g2_mux2_1 _1291_ (.A0(dmi_14_),
    .A1(data_q_12_),
    .S(net193),
    .X(_0575_));
 sg13g2_nand2_1 _1292_ (.Y(_0576_),
    .A(dmi_14_),
    .B(net306));
 sg13g2_buf_2 fanout234 (.A(net236),
    .X(net234));
 sg13g2_nand2_1 _1294_ (.Y(_0578_),
    .A(dmi_15_),
    .B(net169));
 sg13g2_nand3_1 _1295_ (.B(_0576_),
    .C(_0578_),
    .A(net160),
    .Y(_0579_));
 sg13g2_o21ai_1 _1296_ (.B1(_0579_),
    .Y(_0580_),
    .A1(net155),
    .A2(_0575_));
 sg13g2_nor2_1 _1297_ (.A(net224),
    .B(_0580_),
    .Y(dr_d_14_));
 sg13g2_mux2_1 _1298_ (.A0(dmi_15_),
    .A1(data_q_13_),
    .S(net193),
    .X(_0581_));
 sg13g2_buf_2 fanout233 (.A(net236),
    .X(net233));
 sg13g2_nand2_1 _1300_ (.Y(_0583_),
    .A(dmi_15_),
    .B(net306));
 sg13g2_nand2_1 _1301_ (.Y(_0584_),
    .A(dmi_16_),
    .B(net169));
 sg13g2_nand3_1 _1302_ (.B(_0583_),
    .C(_0584_),
    .A(net162),
    .Y(_0585_));
 sg13g2_o21ai_1 _1303_ (.B1(_0585_),
    .Y(_0586_),
    .A1(net155),
    .A2(_0581_));
 sg13g2_nor2_1 _1304_ (.A(net224),
    .B(_0586_),
    .Y(dr_d_15_));
 sg13g2_mux2_1 _1305_ (.A0(dmi_16_),
    .A1(data_q_14_),
    .S(net193),
    .X(_0587_));
 sg13g2_nand2_1 _1306_ (.Y(_0588_),
    .A(dmi_16_),
    .B(net303));
 sg13g2_nand2_1 _1307_ (.Y(_0589_),
    .A(dmi_17_),
    .B(net169));
 sg13g2_nand3_1 _1308_ (.B(_0588_),
    .C(_0589_),
    .A(net162),
    .Y(_0590_));
 sg13g2_o21ai_1 _1309_ (.B1(_0590_),
    .Y(_0591_),
    .A1(net155),
    .A2(_0587_));
 sg13g2_nor2_1 _1310_ (.A(net224),
    .B(_0591_),
    .Y(dr_d_16_));
 sg13g2_buf_1 fanout232 (.A(_0314_),
    .X(net232));
 sg13g2_mux2_1 _1312_ (.A0(dmi_17_),
    .A1(data_q_15_),
    .S(net193),
    .X(_0593_));
 sg13g2_nand2_1 _1313_ (.Y(_0594_),
    .A(dmi_17_),
    .B(net305));
 sg13g2_nand2_1 _1314_ (.Y(_0595_),
    .A(dmi_18_),
    .B(net169));
 sg13g2_nand3_1 _1315_ (.B(_0594_),
    .C(_0595_),
    .A(net162),
    .Y(_0596_));
 sg13g2_o21ai_1 _1316_ (.B1(_0596_),
    .Y(_0597_),
    .A1(net157),
    .A2(_0593_));
 sg13g2_nor2_1 _1317_ (.A(net230),
    .B(_0597_),
    .Y(dr_d_17_));
 sg13g2_mux2_1 _1318_ (.A0(dmi_18_),
    .A1(data_q_16_),
    .S(net193),
    .X(_0598_));
 sg13g2_nand2_1 _1319_ (.Y(_0599_),
    .A(dmi_18_),
    .B(net304));
 sg13g2_nand2_1 _1320_ (.Y(_0600_),
    .A(dmi_19_),
    .B(net169));
 sg13g2_nand3_1 _1321_ (.B(_0599_),
    .C(_0600_),
    .A(net162),
    .Y(_0601_));
 sg13g2_o21ai_1 _1322_ (.B1(_0601_),
    .Y(_0602_),
    .A1(net157),
    .A2(_0598_));
 sg13g2_nor2_1 _1323_ (.A(net230),
    .B(_0602_),
    .Y(dr_d_18_));
 sg13g2_mux2_1 _1324_ (.A0(dmi_19_),
    .A1(data_q_17_),
    .S(net193),
    .X(_0603_));
 sg13g2_nand2_1 _1325_ (.Y(_0604_),
    .A(dmi_19_),
    .B(net304));
 sg13g2_nand2_1 _1326_ (.Y(_0605_),
    .A(dmi_20_),
    .B(net168));
 sg13g2_nand3_1 _1327_ (.B(_0604_),
    .C(_0605_),
    .A(net162),
    .Y(_0606_));
 sg13g2_o21ai_1 _1328_ (.B1(_0606_),
    .Y(_0607_),
    .A1(net157),
    .A2(_0603_));
 sg13g2_nor2_1 _1329_ (.A(net230),
    .B(_0607_),
    .Y(dr_d_19_));
 sg13g2_nand3_1 _1330_ (.B(net154),
    .C(net167),
    .A(dmi_2_),
    .Y(_0608_));
 sg13g2_o21ai_1 _1331_ (.B1(_0543_),
    .Y(_0609_),
    .A1(dmi_1_),
    .A2(_0542_));
 sg13g2_a21o_1 _1332_ (.A2(net173),
    .A1(net161),
    .B1(_0609_),
    .X(_0610_));
 sg13g2_a21oi_1 _1333_ (.A1(_0608_),
    .A2(_0610_),
    .Y(dr_d_1_),
    .B1(net221));
 sg13g2_buf_1 fanout231 (.A(net232),
    .X(net231));
 sg13g2_mux2_1 _1335_ (.A0(dmi_20_),
    .A1(data_q_18_),
    .S(net194),
    .X(_0612_));
 sg13g2_nand2_1 _1336_ (.Y(_0613_),
    .A(dmi_20_),
    .B(net304));
 sg13g2_nand2_1 _1337_ (.Y(_0614_),
    .A(dmi_21_),
    .B(net168));
 sg13g2_nand3_1 _1338_ (.B(_0613_),
    .C(_0614_),
    .A(net161),
    .Y(_0615_));
 sg13g2_o21ai_1 _1339_ (.B1(_0615_),
    .Y(_0616_),
    .A1(net157),
    .A2(_0612_));
 sg13g2_nor2_1 _1340_ (.A(net225),
    .B(_0616_),
    .Y(dr_d_20_));
 sg13g2_mux2_1 _1341_ (.A0(dmi_21_),
    .A1(data_q_19_),
    .S(net192),
    .X(_0617_));
 sg13g2_buf_2 fanout230 (.A(net232),
    .X(net230));
 sg13g2_nand2_1 _1343_ (.Y(_0619_),
    .A(dmi_21_),
    .B(net304));
 sg13g2_nand2_1 _1344_ (.Y(_0620_),
    .A(dmi_22_),
    .B(net168));
 sg13g2_nand3_1 _1345_ (.B(_0619_),
    .C(_0620_),
    .A(net161),
    .Y(_0621_));
 sg13g2_o21ai_1 _1346_ (.B1(_0621_),
    .Y(_0622_),
    .A1(net156),
    .A2(_0617_));
 sg13g2_nor2_1 _1347_ (.A(net223),
    .B(_0622_),
    .Y(dr_d_21_));
 sg13g2_mux2_1 _1348_ (.A0(dmi_22_),
    .A1(data_q_20_),
    .S(net192),
    .X(_0623_));
 sg13g2_nand2_1 _1349_ (.Y(_0624_),
    .A(dmi_22_),
    .B(net304));
 sg13g2_nand2_1 _1350_ (.Y(_0625_),
    .A(dmi_23_),
    .B(net168));
 sg13g2_nand3_1 _1351_ (.B(_0624_),
    .C(_0625_),
    .A(net161),
    .Y(_0626_));
 sg13g2_o21ai_1 _1352_ (.B1(_0626_),
    .Y(_0627_),
    .A1(net156),
    .A2(_0623_));
 sg13g2_nor2_1 _1353_ (.A(net223),
    .B(_0627_),
    .Y(dr_d_22_));
 sg13g2_mux2_1 _1354_ (.A0(dmi_23_),
    .A1(data_q_21_),
    .S(net194),
    .X(_0628_));
 sg13g2_nand2_1 _1355_ (.Y(_0629_),
    .A(dmi_23_),
    .B(net305));
 sg13g2_nand2_1 _1356_ (.Y(_0630_),
    .A(dmi_24_),
    .B(net168));
 sg13g2_nand3_1 _1357_ (.B(_0629_),
    .C(_0630_),
    .A(net161),
    .Y(_0631_));
 sg13g2_o21ai_1 _1358_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net156),
    .A2(_0628_));
 sg13g2_nor2_1 _1359_ (.A(net223),
    .B(_0632_),
    .Y(dr_d_23_));
 sg13g2_buf_2 fanout229 (.A(net232),
    .X(net229));
 sg13g2_mux2_1 _1361_ (.A0(dmi_24_),
    .A1(data_q_22_),
    .S(net193),
    .X(_0634_));
 sg13g2_nand2_1 _1362_ (.Y(_0635_),
    .A(dmi_24_),
    .B(net305));
 sg13g2_buf_2 fanout228 (.A(net232),
    .X(net228));
 sg13g2_nand2_1 _1364_ (.Y(_0637_),
    .A(dmi_25_),
    .B(net170));
 sg13g2_nand3_1 _1365_ (.B(_0635_),
    .C(_0637_),
    .A(net161),
    .Y(_0638_));
 sg13g2_o21ai_1 _1366_ (.B1(_0638_),
    .Y(_0639_),
    .A1(net156),
    .A2(_0634_));
 sg13g2_nor2_1 _1367_ (.A(net228),
    .B(_0639_),
    .Y(dr_d_24_));
 sg13g2_mux2_1 _1368_ (.A0(dmi_25_),
    .A1(data_q_23_),
    .S(net195),
    .X(_0640_));
 sg13g2_buf_2 fanout227 (.A(_0314_),
    .X(net227));
 sg13g2_nand2_1 _1370_ (.Y(_0642_),
    .A(dmi_25_),
    .B(net308));
 sg13g2_nand2_1 _1371_ (.Y(_0643_),
    .A(dmi_26_),
    .B(net170));
 sg13g2_nand3_1 _1372_ (.B(_0642_),
    .C(_0643_),
    .A(net163),
    .Y(_0644_));
 sg13g2_o21ai_1 _1373_ (.B1(_0644_),
    .Y(_0645_),
    .A1(net156),
    .A2(_0640_));
 sg13g2_nor2_1 _1374_ (.A(net229),
    .B(_0645_),
    .Y(dr_d_25_));
 sg13g2_mux2_1 _1375_ (.A0(dmi_26_),
    .A1(data_q_24_),
    .S(net195),
    .X(_0646_));
 sg13g2_nand2_1 _1376_ (.Y(_0647_),
    .A(dmi_26_),
    .B(net308));
 sg13g2_nand2_1 _1377_ (.Y(_0648_),
    .A(dmi_27_),
    .B(net170));
 sg13g2_nand3_1 _1378_ (.B(_0647_),
    .C(_0648_),
    .A(net163),
    .Y(_0649_));
 sg13g2_o21ai_1 _1379_ (.B1(_0649_),
    .Y(_0650_),
    .A1(net156),
    .A2(_0646_));
 sg13g2_nor2_1 _1380_ (.A(net229),
    .B(_0650_),
    .Y(dr_d_26_));
 sg13g2_buf_1 fanout226 (.A(net227),
    .X(net226));
 sg13g2_mux2_1 _1382_ (.A0(dmi_27_),
    .A1(data_q_25_),
    .S(net197),
    .X(_0652_));
 sg13g2_nand2_1 _1383_ (.Y(_0653_),
    .A(dmi_27_),
    .B(net308));
 sg13g2_nand2_1 _1384_ (.Y(_0654_),
    .A(dmi_28_),
    .B(net170));
 sg13g2_nand3_1 _1385_ (.B(_0653_),
    .C(_0654_),
    .A(net163),
    .Y(_0655_));
 sg13g2_o21ai_1 _1386_ (.B1(_0655_),
    .Y(_0656_),
    .A1(net158),
    .A2(_0652_));
 sg13g2_nor2_1 _1387_ (.A(net231),
    .B(_0656_),
    .Y(dr_d_27_));
 sg13g2_mux2_1 _1388_ (.A0(dmi_28_),
    .A1(data_q_26_),
    .S(net197),
    .X(_0657_));
 sg13g2_nand2_1 _1389_ (.Y(_0658_),
    .A(dmi_28_),
    .B(net308));
 sg13g2_nand2_1 _1390_ (.Y(_0659_),
    .A(dmi_29_),
    .B(net170));
 sg13g2_nand3_1 _1391_ (.B(_0658_),
    .C(_0659_),
    .A(net163),
    .Y(_0660_));
 sg13g2_o21ai_1 _1392_ (.B1(_0660_),
    .Y(_0661_),
    .A1(net158),
    .A2(_0657_));
 sg13g2_nor2_1 _1393_ (.A(net231),
    .B(_0661_),
    .Y(dr_d_28_));
 sg13g2_mux2_1 _1394_ (.A0(dmi_29_),
    .A1(data_q_27_),
    .S(net197),
    .X(_0662_));
 sg13g2_nand2_1 _1395_ (.Y(_0663_),
    .A(dmi_29_),
    .B(net308));
 sg13g2_nand2_1 _1396_ (.Y(_0664_),
    .A(dmi_30_),
    .B(net170));
 sg13g2_nand3_1 _1397_ (.B(_0663_),
    .C(_0664_),
    .A(net163),
    .Y(_0665_));
 sg13g2_o21ai_1 _1398_ (.B1(_0665_),
    .Y(_0666_),
    .A1(net158),
    .A2(_0662_));
 sg13g2_nor2_1 _1399_ (.A(net235),
    .B(_0666_),
    .Y(dr_d_29_));
 sg13g2_buf_1 fanout225 (.A(net226),
    .X(net225));
 sg13g2_mux2_1 _1401_ (.A0(dmi_2_),
    .A1(data_q_0_),
    .S(net195),
    .X(_0668_));
 sg13g2_nand2_1 _1402_ (.Y(_0669_),
    .A(dmi_2_),
    .B(net308));
 sg13g2_nand2_1 _1403_ (.Y(_0670_),
    .A(dmi_3_),
    .B(net170));
 sg13g2_nand3_1 _1404_ (.B(_0669_),
    .C(_0670_),
    .A(net163),
    .Y(_0671_));
 sg13g2_o21ai_1 _1405_ (.B1(_0671_),
    .Y(_0672_),
    .A1(net158),
    .A2(_0668_));
 sg13g2_nor2_1 _1406_ (.A(net229),
    .B(_0672_),
    .Y(dr_d_2_));
 sg13g2_mux2_1 _1407_ (.A0(dmi_30_),
    .A1(data_q_28_),
    .S(net198),
    .X(_0673_));
 sg13g2_buf_2 fanout224 (.A(net226),
    .X(net224));
 sg13g2_nand2_1 _1409_ (.Y(_0675_),
    .A(dmi_30_),
    .B(net308));
 sg13g2_nand2_1 _1410_ (.Y(_0676_),
    .A(dmi_31_),
    .B(net169));
 sg13g2_nand3_1 _1411_ (.B(_0675_),
    .C(_0676_),
    .A(net163),
    .Y(_0677_));
 sg13g2_o21ai_1 _1412_ (.B1(_0677_),
    .Y(_0678_),
    .A1(net158),
    .A2(_0673_));
 sg13g2_nor2_1 _1413_ (.A(net231),
    .B(_0678_),
    .Y(dr_d_30_));
 sg13g2_mux2_1 _1414_ (.A0(dmi_31_),
    .A1(data_q_29_),
    .S(net198),
    .X(_0679_));
 sg13g2_nand2_1 _1415_ (.Y(_0680_),
    .A(dmi_31_),
    .B(net305));
 sg13g2_nand2_1 _1416_ (.Y(_0681_),
    .A(dmi_32_),
    .B(net169));
 sg13g2_nand3_1 _1417_ (.B(_0680_),
    .C(_0681_),
    .A(net162),
    .Y(_0682_));
 sg13g2_o21ai_1 _1418_ (.B1(_0682_),
    .Y(_0683_),
    .A1(net158),
    .A2(_0679_));
 sg13g2_nor2_1 _1419_ (.A(net230),
    .B(_0683_),
    .Y(dr_d_31_));
 sg13g2_mux2_1 _1420_ (.A0(dmi_32_),
    .A1(data_q_30_),
    .S(net194),
    .X(_0684_));
 sg13g2_nand2_1 _1421_ (.Y(_0685_),
    .A(dmi_32_),
    .B(net304));
 sg13g2_nand2_1 _1422_ (.Y(_0686_),
    .A(dmi_33_),
    .B(net169));
 sg13g2_nand3_1 _1423_ (.B(_0685_),
    .C(_0686_),
    .A(net162),
    .Y(_0687_));
 sg13g2_o21ai_1 _1424_ (.B1(_0687_),
    .Y(_0688_),
    .A1(net157),
    .A2(_0684_));
 sg13g2_nor2_1 _1425_ (.A(net228),
    .B(_0688_),
    .Y(dr_d_32_));
 sg13g2_buf_2 fanout223 (.A(net226),
    .X(net223));
 sg13g2_mux2_1 _1427_ (.A0(dmi_33_),
    .A1(data_q_31_),
    .S(net195),
    .X(_0690_));
 sg13g2_nand2_1 _1428_ (.Y(_0691_),
    .A(dmi_34_),
    .B(net167));
 sg13g2_nand2_1 _1429_ (.Y(_0692_),
    .A(dmi_33_),
    .B(net304));
 sg13g2_nand3_1 _1430_ (.B(_0691_),
    .C(_0692_),
    .A(net162),
    .Y(_0693_));
 sg13g2_o21ai_1 _1431_ (.B1(_0693_),
    .Y(_0694_),
    .A1(net157),
    .A2(_0690_));
 sg13g2_nor2_1 _1432_ (.A(net228),
    .B(_0694_),
    .Y(dr_d_33_));
 sg13g2_mux2_1 _1433_ (.A0(dmi_34_),
    .A1(address_q_0_),
    .S(net196),
    .X(_0695_));
 sg13g2_buf_2 fanout222 (.A(net226),
    .X(net222));
 sg13g2_nand2_1 _1435_ (.Y(_0697_),
    .A(dmi_34_),
    .B(net307));
 sg13g2_buf_2 fanout221 (.A(net227),
    .X(net221));
 sg13g2_nand2_1 _1437_ (.Y(_0699_),
    .A(dmi_35_),
    .B(net172));
 sg13g2_nand3_1 _1438_ (.B(_0697_),
    .C(_0699_),
    .A(net166),
    .Y(_0700_));
 sg13g2_o21ai_1 _1439_ (.B1(_0700_),
    .Y(_0701_),
    .A1(net157),
    .A2(_0695_));
 sg13g2_nor2_1 _1440_ (.A(net233),
    .B(_0701_),
    .Y(dr_d_34_));
 sg13g2_mux2_1 _1441_ (.A0(dmi_35_),
    .A1(address_q_1_),
    .S(net196),
    .X(_0702_));
 sg13g2_nand2_1 _1442_ (.Y(_0703_),
    .A(dmi_35_),
    .B(net307));
 sg13g2_nand2_1 _1443_ (.Y(_0704_),
    .A(dmi_36_),
    .B(net171));
 sg13g2_nand3_1 _1444_ (.B(_0703_),
    .C(_0704_),
    .A(net164),
    .Y(_0705_));
 sg13g2_o21ai_1 _1445_ (.B1(_0705_),
    .Y(_0706_),
    .A1(net157),
    .A2(_0702_));
 sg13g2_nor2_1 _1446_ (.A(net234),
    .B(_0706_),
    .Y(dr_d_35_));
 sg13g2_buf_2 fanout220 (.A(_0344_),
    .X(net220));
 sg13g2_mux2_1 _1448_ (.A0(dmi_36_),
    .A1(address_q_2_),
    .S(net197),
    .X(_0708_));
 sg13g2_nand2_1 _1449_ (.Y(_0709_),
    .A(dmi_36_),
    .B(net309));
 sg13g2_nand2_1 _1450_ (.Y(_0710_),
    .A(dmi_37_),
    .B(net171));
 sg13g2_nand3_1 _1451_ (.B(_0709_),
    .C(_0710_),
    .A(net164),
    .Y(_0711_));
 sg13g2_o21ai_1 _1452_ (.B1(_0711_),
    .Y(_0712_),
    .A1(net159),
    .A2(_0708_));
 sg13g2_nor2_1 _1453_ (.A(net236),
    .B(_0712_),
    .Y(dr_d_36_));
 sg13g2_mux2_1 _1454_ (.A0(dmi_37_),
    .A1(address_q_3_),
    .S(net196),
    .X(_0713_));
 sg13g2_nand2_1 _1455_ (.Y(_0714_),
    .A(dmi_37_),
    .B(net307));
 sg13g2_nand2_1 _1456_ (.Y(_0715_),
    .A(dmi_38_),
    .B(net171));
 sg13g2_nand3_1 _1457_ (.B(_0714_),
    .C(_0715_),
    .A(net164),
    .Y(_0716_));
 sg13g2_o21ai_1 _1458_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net159),
    .A2(_0713_));
 sg13g2_nor2_1 _1459_ (.A(net234),
    .B(_0717_),
    .Y(dr_d_37_));
 sg13g2_mux2_1 _1460_ (.A0(dmi_38_),
    .A1(address_q_4_),
    .S(net196),
    .X(_0718_));
 sg13g2_nand2_1 _1461_ (.Y(_0719_),
    .A(dmi_38_),
    .B(net307));
 sg13g2_nand2_1 _1462_ (.Y(_0720_),
    .A(dmi_39_),
    .B(net171));
 sg13g2_nand3_1 _1463_ (.B(_0719_),
    .C(_0720_),
    .A(net164),
    .Y(_0721_));
 sg13g2_o21ai_1 _1464_ (.B1(_0721_),
    .Y(_0722_),
    .A1(net159),
    .A2(_0718_));
 sg13g2_nor2_1 _1465_ (.A(net234),
    .B(_0722_),
    .Y(dr_d_38_));
 sg13g2_mux2_1 _1466_ (.A0(dmi_39_),
    .A1(address_q_5_),
    .S(net197),
    .X(_0723_));
 sg13g2_nand2_1 _1467_ (.Y(_0724_),
    .A(dmi_39_),
    .B(net307));
 sg13g2_nand2_1 _1468_ (.Y(_0725_),
    .A(dmi_40_),
    .B(net171));
 sg13g2_nand3_1 _1469_ (.B(_0724_),
    .C(_0725_),
    .A(net164),
    .Y(_0726_));
 sg13g2_o21ai_1 _1470_ (.B1(_0726_),
    .Y(_0727_),
    .A1(net159),
    .A2(_0723_));
 sg13g2_nor2_1 _1471_ (.A(net234),
    .B(_0727_),
    .Y(dr_d_39_));
 sg13g2_mux2_1 _1472_ (.A0(dmi_3_),
    .A1(data_q_1_),
    .S(net195),
    .X(_0728_));
 sg13g2_nand2_1 _1473_ (.Y(_0729_),
    .A(dmi_3_),
    .B(net307));
 sg13g2_nand2_1 _1474_ (.Y(_0730_),
    .A(dmi_4_),
    .B(net171));
 sg13g2_nand3_1 _1475_ (.B(_0729_),
    .C(_0730_),
    .A(net164),
    .Y(_0731_));
 sg13g2_o21ai_1 _1476_ (.B1(_0731_),
    .Y(_0732_),
    .A1(net159),
    .A2(_0728_));
 sg13g2_nor2_1 _1477_ (.A(net233),
    .B(_0732_),
    .Y(dr_d_3_));
 sg13g2_mux2_1 _1478_ (.A0(dmi_40_),
    .A1(address_q_6_),
    .S(net197),
    .X(_0733_));
 sg13g2_nand2_1 _1479_ (.Y(_0734_),
    .A(dmi_40_),
    .B(net307));
 sg13g2_nand2_1 _1480_ (.Y(_0735_),
    .A(td_i),
    .B(net171));
 sg13g2_nand3_1 _1481_ (.B(_0734_),
    .C(_0735_),
    .A(net164),
    .Y(_0736_));
 sg13g2_o21ai_1 _1482_ (.B1(_0736_),
    .Y(_0737_),
    .A1(net159),
    .A2(_0733_));
 sg13g2_nor2_1 _1483_ (.A(net235),
    .B(_0737_),
    .Y(dr_d_40_));
 sg13g2_mux2_1 _1484_ (.A0(dmi_4_),
    .A1(data_q_2_),
    .S(net195),
    .X(_0738_));
 sg13g2_nand2_1 _1485_ (.Y(_0739_),
    .A(dmi_4_),
    .B(net307));
 sg13g2_nand2_1 _1486_ (.Y(_0740_),
    .A(dmi_5_),
    .B(net171));
 sg13g2_nand3_1 _1487_ (.B(_0739_),
    .C(_0740_),
    .A(net164),
    .Y(_0741_));
 sg13g2_o21ai_1 _1488_ (.B1(_0741_),
    .Y(_0742_),
    .A1(net159),
    .A2(_0738_));
 sg13g2_nor2_1 _1489_ (.A(net233),
    .B(_0742_),
    .Y(dr_d_4_));
 sg13g2_mux2_1 _1490_ (.A0(dmi_5_),
    .A1(data_q_3_),
    .S(net195),
    .X(_0743_));
 sg13g2_nand2_1 _1491_ (.Y(_0744_),
    .A(dmi_5_),
    .B(net308));
 sg13g2_nand2_1 _1492_ (.Y(_0745_),
    .A(dmi_6_),
    .B(net170));
 sg13g2_nand3_1 _1493_ (.B(_0744_),
    .C(_0745_),
    .A(net163),
    .Y(_0746_));
 sg13g2_o21ai_1 _1494_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net159),
    .A2(_0743_));
 sg13g2_nor2_1 _1495_ (.A(net233),
    .B(_0747_),
    .Y(dr_d_5_));
 sg13g2_mux2_1 _1496_ (.A0(dmi_6_),
    .A1(data_q_4_),
    .S(net195),
    .X(_0075_));
 sg13g2_nand2_1 _1497_ (.Y(_0076_),
    .A(dmi_6_),
    .B(net304));
 sg13g2_nand2_1 _1498_ (.Y(_0077_),
    .A(dmi_7_),
    .B(net167));
 sg13g2_nand3_1 _1499_ (.B(_0076_),
    .C(_0077_),
    .A(net161),
    .Y(_0078_));
 sg13g2_o21ai_1 _1500_ (.B1(_0078_),
    .Y(_0079_),
    .A1(net158),
    .A2(_0075_));
 sg13g2_nor2_1 _1501_ (.A(net228),
    .B(_0079_),
    .Y(dr_d_6_));
 sg13g2_mux2_1 _1502_ (.A0(dmi_7_),
    .A1(data_q_5_),
    .S(net192),
    .X(_0080_));
 sg13g2_nand2_1 _1503_ (.Y(_0081_),
    .A(dmi_7_),
    .B(net303));
 sg13g2_nand2_1 _1504_ (.Y(_0082_),
    .A(dmi_8_),
    .B(net167));
 sg13g2_nand3_1 _1505_ (.B(_0081_),
    .C(_0082_),
    .A(net160),
    .Y(_0083_));
 sg13g2_o21ai_1 _1506_ (.B1(_0083_),
    .Y(_0084_),
    .A1(net158),
    .A2(_0080_));
 sg13g2_nor2_1 _1507_ (.A(net223),
    .B(_0084_),
    .Y(dr_d_7_));
 sg13g2_mux2_1 _1508_ (.A0(dmi_8_),
    .A1(data_q_6_),
    .S(net193),
    .X(_0085_));
 sg13g2_nand2_1 _1509_ (.Y(_0086_),
    .A(dmi_8_),
    .B(net303));
 sg13g2_nand2_1 _1510_ (.Y(_0087_),
    .A(dmi_9_),
    .B(net167));
 sg13g2_nand3_1 _1511_ (.B(_0086_),
    .C(_0087_),
    .A(net160),
    .Y(_0088_));
 sg13g2_o21ai_1 _1512_ (.B1(_0088_),
    .Y(_0089_),
    .A1(net154),
    .A2(_0085_));
 sg13g2_nor2_1 _1513_ (.A(net222),
    .B(_0089_),
    .Y(dr_d_8_));
 sg13g2_mux2_1 _1514_ (.A0(dmi_9_),
    .A1(data_q_7_),
    .S(net192),
    .X(_0090_));
 sg13g2_nand2_1 _1515_ (.Y(_0091_),
    .A(dmi_9_),
    .B(net303));
 sg13g2_nand2_1 _1516_ (.Y(_0092_),
    .A(dmi_10_),
    .B(net167));
 sg13g2_nand3_1 _1517_ (.B(_0091_),
    .C(_0092_),
    .A(net160),
    .Y(_0093_));
 sg13g2_o21ai_1 _1518_ (.B1(_0093_),
    .Y(_0094_),
    .A1(net154),
    .A2(_0090_));
 sg13g2_nor2_1 _1519_ (.A(net221),
    .B(_0094_),
    .Y(dr_d_9_));
 sg13g2_inv_1 _1520_ (.Y(_0095_),
    .A(dtmcs_q_1_));
 sg13g2_nor2b_1 _1521_ (.A(\i_dmi_jtag_tap.jtag_ir_q_0_ ),
    .B_N(_0311_),
    .Y(_0096_));
 sg13g2_and2_1 _1522_ (.A(net154),
    .B(_0096_),
    .X(_0097_));
 sg13g2_buf_2 fanout219 (.A(net220),
    .X(net219));
 sg13g2_nand2_1 _1524_ (.Y(_0099_),
    .A(_0269_),
    .B(_0096_));
 sg13g2_buf_2 fanout218 (.A(net219),
    .X(net218));
 sg13g2_inv_1 _1526_ (.Y(_0101_),
    .A(dtmcs_q_0_));
 sg13g2_a22oi_1 _1527_ (.Y(dtmcs_d_0_),
    .B1(net247),
    .B2(_0101_),
    .A2(net258),
    .A1(_0095_));
 sg13g2_or3_1 _1528_ (.A(net316),
    .B(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .C(_0257_),
    .X(_0102_));
 sg13g2_nor2_1 _1529_ (.A(_0312_),
    .B(_0102_),
    .Y(_0103_));
 sg13g2_a22oi_1 _1530_ (.Y(_0104_),
    .B1(_0103_),
    .B2(error_q_0_),
    .A2(_0102_),
    .A1(dtmcs_q_10_));
 sg13g2_a22oi_1 _1531_ (.Y(_0105_),
    .B1(net258),
    .B2(dtmcs_q_11_),
    .A2(_0312_),
    .A1(dtmcs_q_10_));
 sg13g2_o21ai_1 _1532_ (.B1(_0105_),
    .Y(dtmcs_d_10_),
    .A1(net155),
    .A2(_0104_));
 sg13g2_a22oi_1 _1533_ (.Y(_0106_),
    .B1(_0103_),
    .B2(error_q_1_),
    .A2(_0102_),
    .A1(dtmcs_q_11_));
 sg13g2_a22oi_1 _1534_ (.Y(_0107_),
    .B1(net257),
    .B2(dtmcs_q_12_),
    .A2(_0312_),
    .A1(dtmcs_q_11_));
 sg13g2_o21ai_1 _1535_ (.B1(_0107_),
    .Y(dtmcs_d_11_),
    .A1(net155),
    .A2(_0106_));
 sg13g2_inv_1 _1536_ (.Y(_0108_),
    .A(dtmcs_q_13_));
 sg13g2_inv_1 _1537_ (.Y(_0109_),
    .A(dtmcs_q_12_));
 sg13g2_a22oi_1 _1538_ (.Y(dtmcs_d_12_),
    .B1(net247),
    .B2(_0109_),
    .A2(net257),
    .A1(_0108_));
 sg13g2_a22oi_1 _1539_ (.Y(_0110_),
    .B1(net247),
    .B2(dtmcs_q_13_),
    .A2(net257),
    .A1(dtmcs_q_14_));
 sg13g2_inv_1 _1540_ (.Y(dtmcs_d_13_),
    .A(_0110_));
 sg13g2_a22oi_1 _1541_ (.Y(_0111_),
    .B1(net247),
    .B2(dtmcs_q_14_),
    .A2(net257),
    .A1(dtmcs_q_15_));
 sg13g2_inv_1 _1542_ (.Y(dtmcs_d_14_),
    .A(_0111_));
 sg13g2_a22oi_1 _1543_ (.Y(_0112_),
    .B1(net247),
    .B2(dtmcs_q_15_),
    .A2(net257),
    .A1(dtmcs_q_16_));
 sg13g2_inv_1 _1544_ (.Y(dtmcs_d_15_),
    .A(_0112_));
 sg13g2_buf_2 fanout217 (.A(net220),
    .X(net217));
 sg13g2_a22oi_1 _1546_ (.Y(_0114_),
    .B1(net247),
    .B2(dtmcs_q_16_),
    .A2(net257),
    .A1(dtmcs_q_17_));
 sg13g2_inv_1 _1547_ (.Y(dtmcs_d_16_),
    .A(_0114_));
 sg13g2_a22oi_1 _1548_ (.Y(_0115_),
    .B1(net247),
    .B2(dtmcs_q_17_),
    .A2(net257),
    .A1(dtmcs_q_18_));
 sg13g2_inv_1 _1549_ (.Y(dtmcs_d_17_),
    .A(_0115_));
 sg13g2_buf_2 fanout216 (.A(net217),
    .X(net216));
 sg13g2_a22oi_1 _1551_ (.Y(_0117_),
    .B1(net244),
    .B2(dtmcs_q_18_),
    .A2(net256),
    .A1(dtmcs_q_19_));
 sg13g2_inv_1 _1552_ (.Y(dtmcs_d_18_),
    .A(_0117_));
 sg13g2_a22oi_1 _1553_ (.Y(_0118_),
    .B1(net244),
    .B2(dtmcs_q_19_),
    .A2(net254),
    .A1(dtmcs_q_20_));
 sg13g2_inv_1 _1554_ (.Y(dtmcs_d_19_),
    .A(_0118_));
 sg13g2_a22oi_1 _1555_ (.Y(_0119_),
    .B1(net248),
    .B2(dtmcs_q_1_),
    .A2(net258),
    .A1(dtmcs_q_2_));
 sg13g2_inv_1 _1556_ (.Y(dtmcs_d_1_),
    .A(_0119_));
 sg13g2_a22oi_1 _1557_ (.Y(_0120_),
    .B1(net244),
    .B2(dtmcs_q_20_),
    .A2(net254),
    .A1(dtmcs_q_21_));
 sg13g2_inv_1 _1558_ (.Y(dtmcs_d_20_),
    .A(_0120_));
 sg13g2_a22oi_1 _1559_ (.Y(_0121_),
    .B1(net245),
    .B2(dtmcs_q_21_),
    .A2(net255),
    .A1(dtmcs_q_22_));
 sg13g2_inv_1 _1560_ (.Y(dtmcs_d_21_),
    .A(_0121_));
 sg13g2_a22oi_1 _1561_ (.Y(_0122_),
    .B1(net245),
    .B2(dtmcs_q_22_),
    .A2(net255),
    .A1(dtmcs_q_23_));
 sg13g2_inv_1 _1562_ (.Y(dtmcs_d_22_),
    .A(_0122_));
 sg13g2_a22oi_1 _1563_ (.Y(_0123_),
    .B1(net244),
    .B2(dtmcs_q_23_),
    .A2(net254),
    .A1(dtmcs_q_24_));
 sg13g2_inv_1 _1564_ (.Y(dtmcs_d_23_),
    .A(_0123_));
 sg13g2_a22oi_1 _1565_ (.Y(_0124_),
    .B1(net244),
    .B2(dtmcs_q_24_),
    .A2(net254),
    .A1(dtmcs_q_25_));
 sg13g2_inv_1 _1566_ (.Y(dtmcs_d_24_),
    .A(_0124_));
 sg13g2_buf_1 fanout215 (.A(_0357_),
    .X(net215));
 sg13g2_a22oi_1 _1568_ (.Y(_0126_),
    .B1(net244),
    .B2(dtmcs_q_25_),
    .A2(net254),
    .A1(dtmcs_q_26_));
 sg13g2_inv_1 _1569_ (.Y(dtmcs_d_25_),
    .A(_0126_));
 sg13g2_a22oi_1 _1570_ (.Y(_0127_),
    .B1(net244),
    .B2(dtmcs_q_26_),
    .A2(net254),
    .A1(dtmcs_q_27_));
 sg13g2_inv_1 _1571_ (.Y(dtmcs_d_26_),
    .A(_0127_));
 sg13g2_buf_2 fanout214 (.A(_0357_),
    .X(net214));
 sg13g2_a22oi_1 _1573_ (.Y(_0129_),
    .B1(net244),
    .B2(dtmcs_q_27_),
    .A2(net254),
    .A1(dtmcs_q_28_));
 sg13g2_inv_1 _1574_ (.Y(dtmcs_d_27_),
    .A(_0129_));
 sg13g2_a22oi_1 _1575_ (.Y(_0130_),
    .B1(net246),
    .B2(dtmcs_q_28_),
    .A2(net254),
    .A1(dtmcs_q_29_));
 sg13g2_inv_1 _1576_ (.Y(dtmcs_d_28_),
    .A(_0130_));
 sg13g2_a22oi_1 _1577_ (.Y(_0131_),
    .B1(net246),
    .B2(dtmcs_q_29_),
    .A2(net256),
    .A1(dtmcs_q_30_));
 sg13g2_inv_1 _1578_ (.Y(dtmcs_d_29_),
    .A(_0131_));
 sg13g2_a22oi_1 _1579_ (.Y(_0132_),
    .B1(net248),
    .B2(dtmcs_q_2_),
    .A2(net256),
    .A1(dtmcs_q_3_));
 sg13g2_inv_1 _1580_ (.Y(dtmcs_d_2_),
    .A(_0132_));
 sg13g2_a22oi_1 _1581_ (.Y(_0133_),
    .B1(net246),
    .B2(dtmcs_q_30_),
    .A2(net256),
    .A1(dtmcs_q_31_));
 sg13g2_inv_1 _1582_ (.Y(dtmcs_d_30_),
    .A(_0133_));
 sg13g2_a22oi_1 _1583_ (.Y(_0134_),
    .B1(net247),
    .B2(dtmcs_q_31_),
    .A2(net257),
    .A1(td_i));
 sg13g2_inv_1 _1584_ (.Y(dtmcs_d_31_),
    .A(_0134_));
 sg13g2_a22oi_1 _1585_ (.Y(_0135_),
    .B1(net246),
    .B2(dtmcs_q_3_),
    .A2(net256),
    .A1(dtmcs_q_4_));
 sg13g2_inv_1 _1586_ (.Y(dtmcs_d_3_),
    .A(_0135_));
 sg13g2_inv_1 _1587_ (.Y(_0136_),
    .A(dtmcs_q_5_));
 sg13g2_inv_1 _1588_ (.Y(_0137_),
    .A(dtmcs_q_4_));
 sg13g2_a22oi_1 _1589_ (.Y(dtmcs_d_4_),
    .B1(net245),
    .B2(_0137_),
    .A2(net255),
    .A1(_0136_));
 sg13g2_inv_1 _1590_ (.Y(_0138_),
    .A(dtmcs_q_6_));
 sg13g2_a22oi_1 _1591_ (.Y(dtmcs_d_5_),
    .B1(net245),
    .B2(_0136_),
    .A2(net255),
    .A1(_0138_));
 sg13g2_inv_1 _1592_ (.Y(_0139_),
    .A(dtmcs_q_7_));
 sg13g2_a22oi_1 _1593_ (.Y(dtmcs_d_6_),
    .B1(net245),
    .B2(_0138_),
    .A2(net255),
    .A1(_0139_));
 sg13g2_a22oi_1 _1594_ (.Y(_0140_),
    .B1(net245),
    .B2(dtmcs_q_7_),
    .A2(net255),
    .A1(dtmcs_q_8_));
 sg13g2_inv_1 _1595_ (.Y(dtmcs_d_7_),
    .A(_0140_));
 sg13g2_a22oi_1 _1596_ (.Y(_0141_),
    .B1(net245),
    .B2(dtmcs_q_8_),
    .A2(net255),
    .A1(dtmcs_q_9_));
 sg13g2_inv_1 _1597_ (.Y(dtmcs_d_8_),
    .A(_0141_));
 sg13g2_a22oi_1 _1598_ (.Y(_0142_),
    .B1(net245),
    .B2(dtmcs_q_9_),
    .A2(net255),
    .A1(dtmcs_q_10_));
 sg13g2_inv_1 _1599_ (.Y(dtmcs_d_9_),
    .A(_0142_));
 sg13g2_nand2_1 _1600_ (.Y(_0143_),
    .A(dtmcs_q_16_),
    .B(_0313_));
 sg13g2_nand4_1 _1601_ (.B(net321),
    .C(_0320_),
    .A(net312),
    .Y(_0144_),
    .D(_0537_));
 sg13g2_nand2_1 _1602_ (.Y(_0145_),
    .A(_0143_),
    .B(_0144_));
 sg13g2_nor2_1 _1603_ (.A(error_q_1_),
    .B(_0539_),
    .Y(_0146_));
 sg13g2_nor2_1 _1604_ (.A(error_q_0_),
    .B(_0146_),
    .Y(_0147_));
 sg13g2_nor3_1 _1605_ (.A(net221),
    .B(_0145_),
    .C(_0147_),
    .Y(_0066_));
 sg13g2_nor2_1 _1606_ (.A(error_q_0_),
    .B(_0539_),
    .Y(_0148_));
 sg13g2_nor2_1 _1607_ (.A(error_q_1_),
    .B(_0148_),
    .Y(_0149_));
 sg13g2_a221oi_1 _1608_ (.B2(_0149_),
    .C1(net221),
    .B1(_0144_),
    .A1(dtmcs_q_16_),
    .Y(_0067_),
    .A2(_0313_));
 sg13g2_nand2_1 _1609_ (.Y(_0150_),
    .A(\i_dmi_jtag_tap.jtag_ir_q_4__$_NOT__A_Y ),
    .B(_0281_));
 sg13g2_nand2_1 _1610_ (.Y(_0151_),
    .A(_0282_),
    .B(_0150_));
 sg13g2_o21ai_1 _1611_ (.B1(_0151_),
    .Y(_0152_),
    .A1(net154),
    .A2(_0531_));
 sg13g2_nand2_1 _1612_ (.Y(_0153_),
    .A(\i_dmi_jtag_tap.bypass_q ),
    .B(_0152_));
 sg13g2_nand3_1 _1613_ (.B(net154),
    .C(_0151_),
    .A(td_i),
    .Y(_0154_));
 sg13g2_a21oi_1 _1614_ (.A1(_0153_),
    .A2(_0154_),
    .Y(\i_dmi_jtag_tap.bypass_d ),
    .B1(net241));
 sg13g2_buf_2 fanout213 (.A(_0357_),
    .X(net213));
 sg13g2_buf_2 fanout212 (.A(net213),
    .X(net212));
 sg13g2_a22oi_1 _1617_ (.Y(_0157_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_13_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_12_ ));
 sg13g2_nor2_1 _1618_ (.A(net237),
    .B(_0157_),
    .Y(\i_dmi_jtag_tap.idcode_d_12_ ));
 sg13g2_a22oi_1 _1619_ (.Y(_0158_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_14_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_13_ ));
 sg13g2_nor2_1 _1620_ (.A(net237),
    .B(_0158_),
    .Y(\i_dmi_jtag_tap.idcode_d_13_ ));
 sg13g2_buf_1 fanout211 (.A(net213),
    .X(net211));
 sg13g2_a22oi_1 _1622_ (.Y(_0160_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_15_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_14_ ));
 sg13g2_nor2_1 _1623_ (.A(net237),
    .B(_0160_),
    .Y(\i_dmi_jtag_tap.idcode_d_14_ ));
 sg13g2_a22oi_1 _1624_ (.Y(_0161_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_16_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_15_ ));
 sg13g2_nor2_1 _1625_ (.A(net237),
    .B(_0161_),
    .Y(\i_dmi_jtag_tap.idcode_d_15_ ));
 sg13g2_a22oi_1 _1626_ (.Y(_0162_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_17_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_16_ ));
 sg13g2_nor2_1 _1627_ (.A(net237),
    .B(_0162_),
    .Y(\i_dmi_jtag_tap.idcode_d_16_ ));
 sg13g2_a22oi_1 _1628_ (.Y(_0163_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_18_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_17_ ));
 sg13g2_nor2_1 _1629_ (.A(net237),
    .B(_0163_),
    .Y(\i_dmi_jtag_tap.idcode_d_17_ ));
 sg13g2_a22oi_1 _1630_ (.Y(_0164_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_19_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_18_ ));
 sg13g2_nor2_1 _1631_ (.A(net239),
    .B(_0164_),
    .Y(\i_dmi_jtag_tap.idcode_d_18_ ));
 sg13g2_a22oi_1 _1632_ (.Y(_0165_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_20_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_19_ ));
 sg13g2_nor2_1 _1633_ (.A(net239),
    .B(_0165_),
    .Y(\i_dmi_jtag_tap.idcode_d_19_ ));
 sg13g2_buf_2 fanout210 (.A(net213),
    .X(net210));
 sg13g2_a22oi_1 _1635_ (.Y(_0167_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_21_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_20_ ));
 sg13g2_nor2_1 _1636_ (.A(net239),
    .B(_0167_),
    .Y(\i_dmi_jtag_tap.idcode_d_20_ ));
 sg13g2_a22oi_1 _1637_ (.Y(_0168_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_22_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_21_ ));
 sg13g2_nor2_1 _1638_ (.A(net240),
    .B(_0168_),
    .Y(\i_dmi_jtag_tap.idcode_d_21_ ));
 sg13g2_buf_2 fanout209 (.A(\i_dmi_cdc.i_cdc_resp/i_src/_036_ ),
    .X(net209));
 sg13g2_a22oi_1 _1640_ (.Y(_0170_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_23_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_22_ ));
 sg13g2_nor2_1 _1641_ (.A(net239),
    .B(_0170_),
    .Y(\i_dmi_jtag_tap.idcode_d_22_ ));
 sg13g2_a22oi_1 _1642_ (.Y(_0171_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_24_ ),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_23_ ));
 sg13g2_nor2_1 _1643_ (.A(net239),
    .B(_0171_),
    .Y(\i_dmi_jtag_tap.idcode_d_23_ ));
 sg13g2_buf_4 fanout208 (.X(net208),
    .A(net209));
 sg13g2_a22oi_1 _1645_ (.Y(_0173_),
    .B1(net263),
    .B2(\i_dmi_jtag_tap.idcode_q_25_ ),
    .A2(net251),
    .A1(\i_dmi_jtag_tap.idcode_q_24_ ));
 sg13g2_nor2_1 _1646_ (.A(net239),
    .B(_0173_),
    .Y(\i_dmi_jtag_tap.idcode_d_24_ ));
 sg13g2_a22oi_1 _1647_ (.Y(_0174_),
    .B1(net263),
    .B2(\i_dmi_jtag_tap.idcode_q_26_ ),
    .A2(net251),
    .A1(\i_dmi_jtag_tap.idcode_q_25_ ));
 sg13g2_nor2_1 _1648_ (.A(net239),
    .B(_0174_),
    .Y(\i_dmi_jtag_tap.idcode_d_25_ ));
 sg13g2_a22oi_1 _1649_ (.Y(_0175_),
    .B1(net262),
    .B2(\i_dmi_jtag_tap.idcode_q_27_ ),
    .A2(net251),
    .A1(\i_dmi_jtag_tap.idcode_q_26_ ));
 sg13g2_nor2_1 _1650_ (.A(net239),
    .B(_0175_),
    .Y(\i_dmi_jtag_tap.idcode_d_26_ ));
 sg13g2_a22oi_1 _1651_ (.Y(_0176_),
    .B1(net263),
    .B2(\i_dmi_jtag_tap.idcode_q_28_ ),
    .A2(net251),
    .A1(\i_dmi_jtag_tap.idcode_q_27_ ));
 sg13g2_nor2_1 _1652_ (.A(net238),
    .B(_0176_),
    .Y(\i_dmi_jtag_tap.idcode_d_27_ ));
 sg13g2_a22oi_1 _1653_ (.Y(_0177_),
    .B1(net263),
    .B2(\i_dmi_jtag_tap.idcode_q_29_ ),
    .A2(net251),
    .A1(\i_dmi_jtag_tap.idcode_q_28_ ));
 sg13g2_nor2_1 _1654_ (.A(net238),
    .B(_0177_),
    .Y(\i_dmi_jtag_tap.idcode_d_28_ ));
 sg13g2_a22oi_1 _1655_ (.Y(_0178_),
    .B1(net264),
    .B2(\i_dmi_jtag_tap.idcode_q_30_ ),
    .A2(net252),
    .A1(\i_dmi_jtag_tap.idcode_q_29_ ));
 sg13g2_nor2_1 _1656_ (.A(net238),
    .B(_0178_),
    .Y(\i_dmi_jtag_tap.idcode_d_29_ ));
 sg13g2_buf_4 fanout207 (.X(net207),
    .A(net209));
 sg13g2_a22oi_1 _1658_ (.Y(_0180_),
    .B1(net264),
    .B2(\i_dmi_jtag_tap.idcode_q_3_ ),
    .A2(net253),
    .A1(\i_dmi_jtag_tap.idcode_q_2_ ));
 sg13g2_nor2_1 _1659_ (.A(net242),
    .B(_0180_),
    .Y(\i_dmi_jtag_tap.idcode_d_2_ ));
 sg13g2_a22oi_1 _1660_ (.Y(_0181_),
    .B1(net265),
    .B2(\i_dmi_jtag_tap.idcode_q_31_ ),
    .A2(net253),
    .A1(\i_dmi_jtag_tap.idcode_q_30_ ));
 sg13g2_nor2_1 _1661_ (.A(net238),
    .B(_0181_),
    .Y(\i_dmi_jtag_tap.idcode_d_30_ ));
 sg13g2_a22oi_1 _1662_ (.Y(_0182_),
    .B1(net265),
    .B2(td_i),
    .A2(net250),
    .A1(\i_dmi_jtag_tap.idcode_q_31_ ));
 sg13g2_nor2_1 _1663_ (.A(net240),
    .B(_0182_),
    .Y(\i_dmi_jtag_tap.idcode_d_31_ ));
 sg13g2_a22oi_1 _1664_ (.Y(_0183_),
    .B1(net264),
    .B2(\i_dmi_jtag_tap.idcode_q_4_ ),
    .A2(net252),
    .A1(\i_dmi_jtag_tap.idcode_q_3_ ));
 sg13g2_nor2_1 _1665_ (.A(net242),
    .B(_0183_),
    .Y(\i_dmi_jtag_tap.idcode_d_3_ ));
 sg13g2_a22oi_1 _1666_ (.Y(_0184_),
    .B1(net264),
    .B2(\i_dmi_jtag_tap.idcode_q_7_ ),
    .A2(net252),
    .A1(\i_dmi_jtag_tap.idcode_q_6_ ));
 sg13g2_nor2_1 _1667_ (.A(net242),
    .B(_0184_),
    .Y(\i_dmi_jtag_tap.idcode_d_6_ ));
 sg13g2_a22oi_1 _1668_ (.Y(_0185_),
    .B1(net261),
    .B2(\i_dmi_jtag_tap.idcode_q_10_ ),
    .A2(net249),
    .A1(\i_dmi_jtag_tap.idcode_q_9_ ));
 sg13g2_nor2_1 _1669_ (.A(net238),
    .B(_0185_),
    .Y(\i_dmi_jtag_tap.idcode_d_9_ ));
 sg13g2_or3_2 _1670_ (.A(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .B(net315),
    .C(_0257_),
    .X(_0186_));
 sg13g2_buf_2 fanout206 (.A(net209),
    .X(net206));
 sg13g2_nand3b_1 _1672_ (.B(_0010_),
    .C(_0186_),
    .Y(_0188_),
    .A_N(net243));
 sg13g2_o21ai_1 _1673_ (.B1(_0188_),
    .Y(_0068_),
    .A1(\i_dmi_jtag_tap.jtag_ir_shift_q_0_ ),
    .A2(_0186_));
 sg13g2_nor2b_1 _1674_ (.A(net241),
    .B_N(\i_dmi_jtag_tap.jtag_ir_q_1_ ),
    .Y(_0189_));
 sg13g2_mux2_1 _1675_ (.A0(\i_dmi_jtag_tap.jtag_ir_shift_q_1_ ),
    .A1(_0189_),
    .S(_0186_),
    .X(_0069_));
 sg13g2_nor2b_1 _1676_ (.A(net241),
    .B_N(\i_dmi_jtag_tap.jtag_ir_q_2_ ),
    .Y(_0190_));
 sg13g2_mux2_1 _1677_ (.A0(\i_dmi_jtag_tap.jtag_ir_shift_q_2_ ),
    .A1(_0190_),
    .S(_0186_),
    .X(_0070_));
 sg13g2_nor2b_1 _1678_ (.A(net241),
    .B_N(\i_dmi_jtag_tap.jtag_ir_q_3_ ),
    .Y(_0191_));
 sg13g2_mux2_1 _1679_ (.A0(\i_dmi_jtag_tap.jtag_ir_shift_q_3_ ),
    .A1(_0191_),
    .S(_0186_),
    .X(_0071_));
 sg13g2_nor2b_1 _1680_ (.A(net241),
    .B_N(\i_dmi_jtag_tap.jtag_ir_q_4_ ),
    .Y(_0192_));
 sg13g2_mux2_1 _1681_ (.A0(\i_dmi_jtag_tap.jtag_ir_shift_q_4_ ),
    .A1(_0192_),
    .S(_0186_),
    .X(_0072_));
 sg13g2_nor2_2 _1682_ (.A(net314),
    .B(_0250_),
    .Y(_0193_));
 sg13g2_nand3b_1 _1683_ (.B(net319),
    .C(_0193_),
    .Y(_0194_),
    .A_N(\i_dmi_jtag_tap.jtag_ir_shift_q_1_ ));
 sg13g2_o21ai_1 _1684_ (.B1(_0194_),
    .Y(_0195_),
    .A1(\i_dmi_jtag_tap.jtag_ir_shift_q_0_ ),
    .A2(_0193_));
 sg13g2_nor2_1 _1685_ (.A(net241),
    .B(_0195_),
    .Y(_0073_));
 sg13g2_o21ai_1 _1686_ (.B1(\i_dmi_jtag_tap.jtag_ir_shift_q_1_ ),
    .Y(_0196_),
    .A1(net314),
    .A2(_0250_));
 sg13g2_nand3_1 _1687_ (.B(net318),
    .C(_0193_),
    .A(\i_dmi_jtag_tap.jtag_ir_shift_q_2_ ),
    .Y(_0197_));
 sg13g2_a21oi_1 _1688_ (.A1(_0196_),
    .A2(_0197_),
    .Y(_0074_),
    .B1(net241));
 sg13g2_nand3b_1 _1689_ (.B(net318),
    .C(_0193_),
    .Y(_0198_),
    .A_N(\i_dmi_jtag_tap.jtag_ir_shift_q_3_ ));
 sg13g2_o21ai_1 _1690_ (.B1(_0198_),
    .Y(_0199_),
    .A1(\i_dmi_jtag_tap.jtag_ir_shift_q_2_ ),
    .A2(_0193_));
 sg13g2_nor2_1 _1691_ (.A(net240),
    .B(_0199_),
    .Y(_0021_));
 sg13g2_o21ai_1 _1692_ (.B1(\i_dmi_jtag_tap.jtag_ir_shift_q_3_ ),
    .Y(_0200_),
    .A1(net314),
    .A2(_0250_));
 sg13g2_nand3_1 _1693_ (.B(net318),
    .C(_0193_),
    .A(\i_dmi_jtag_tap.jtag_ir_shift_q_4_ ),
    .Y(_0201_));
 sg13g2_a21oi_1 _1694_ (.A1(_0200_),
    .A2(_0201_),
    .Y(_0022_),
    .B1(net240));
 sg13g2_o21ai_1 _1695_ (.B1(\i_dmi_jtag_tap.jtag_ir_shift_q_4_ ),
    .Y(_0202_),
    .A1(net314),
    .A2(_0250_));
 sg13g2_nand3_1 _1696_ (.B(net318),
    .C(_0193_),
    .A(td_i),
    .Y(_0203_));
 sg13g2_a21oi_1 _1697_ (.A1(_0202_),
    .A2(_0203_),
    .Y(_0023_),
    .B1(net240));
 sg13g2_nor3_1 _1698_ (.A(_0264_),
    .B(_0258_),
    .C(_0260_),
    .Y(_0204_));
 sg13g2_mux2_1 _1699_ (.A0(_0250_),
    .A1(_0238_),
    .S(net318),
    .X(_0205_));
 sg13g2_nor2_1 _1700_ (.A(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_nor3_1 _1701_ (.A(net174),
    .B(_0254_),
    .C(_0206_),
    .Y(_0207_));
 sg13g2_a21oi_1 _1702_ (.A1(net174),
    .A2(_0204_),
    .Y(_0208_),
    .B1(_0207_));
 sg13g2_nor3_1 _1703_ (.A(_0274_),
    .B(_0270_),
    .C(_0208_),
    .Y(_0209_));
 sg13g2_nor2_1 _1704_ (.A(_0279_),
    .B(_0209_),
    .Y(\i_dmi_jtag_tap.tap_state_d_1_ ));
 sg13g2_a221oi_1 _1705_ (.B2(_0253_),
    .C1(_0248_),
    .B1(net317),
    .A1(net174),
    .Y(_0210_),
    .A2(net320));
 sg13g2_and3_1 _1706_ (.X(_0211_),
    .A(net174),
    .B(_0273_),
    .C(_0243_));
 sg13g2_nor4_1 _1707_ (.A(_0264_),
    .B(_0269_),
    .C(_0210_),
    .D(_0211_),
    .Y(_0212_));
 sg13g2_nor2_1 _1708_ (.A(_0279_),
    .B(_0212_),
    .Y(\i_dmi_jtag_tap.tap_state_d_2_ ));
 sg13g2_o21ai_1 _1709_ (.B1(net174),
    .Y(_0213_),
    .A1(net317),
    .A2(_0248_));
 sg13g2_a21o_1 _1710_ (.A2(_0213_),
    .A1(net318),
    .B1(_0206_),
    .X(_0214_));
 sg13g2_o21ai_1 _1711_ (.B1(_0214_),
    .Y(_0215_),
    .A1(net174),
    .A2(_0254_));
 sg13g2_nor2b_1 _1712_ (.A(_0215_),
    .B_N(_0278_),
    .Y(_0216_));
 sg13g2_or2_1 _1713_ (.X(\i_dmi_jtag_tap.tap_state_d_3_ ),
    .B(_0216_),
    .A(_0246_));
 sg13g2_nor3_1 _1714_ (.A(net316),
    .B(net315),
    .C(_0257_),
    .Y(_0217_));
 sg13g2_a221oi_1 _1715_ (.B2(\i_dmi_jtag_tap.bypass_q ),
    .C1(_0217_),
    .B1(_0151_),
    .A1(\i_dmi_jtag_tap.idcode_q_0_ ),
    .Y(_0218_),
    .A2(_0283_));
 sg13g2_a22oi_1 _1716_ (.Y(_0219_),
    .B1(net172),
    .B2(dmi_0_),
    .A2(_0096_),
    .A1(dtmcs_q_0_));
 sg13g2_nand2_1 _1717_ (.Y(_0220_),
    .A(net319),
    .B(_0193_));
 sg13g2_nor2_1 _1718_ (.A(\i_dmi_jtag_tap.jtag_ir_shift_q_0_ ),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_a21oi_1 _1719_ (.A1(_0218_),
    .A2(_0219_),
    .Y(\i_dmi_jtag_tap.tdo_mux ),
    .B1(_0221_));
 sg13g2_nor2_1 _1720_ (.A(dmi_resp_valid),
    .B(_0339_),
    .Y(_0222_));
 sg13g2_nor2_1 _1721_ (.A(dmi_1_),
    .B(\state_d_1__$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_OR__Y_A ),
    .Y(_0223_));
 sg13g2_nor2_1 _1722_ (.A(dmi_0_),
    .B(\state_q_0__reg_E_$_AND__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B ),
    .Y(_0224_));
 sg13g2_nor2_1 _1723_ (.A(_0223_),
    .B(_0224_),
    .Y(_0225_));
 sg13g2_nor2_1 _1724_ (.A(dmi_req_ready),
    .B(_0525_),
    .Y(_0226_));
 sg13g2_a221oi_1 _1725_ (.B2(_0322_),
    .C1(_0226_),
    .B1(_0225_),
    .A1(_0525_),
    .Y(_0227_),
    .A2(_0222_));
 sg13g2_nand2b_1 _1726_ (.Y(_0228_),
    .B(state_q_0_),
    .A_N(_0227_));
 sg13g2_nand3_1 _1727_ (.B(_0340_),
    .C(_0227_),
    .A(_0339_),
    .Y(_0229_));
 sg13g2_a21oi_1 _1728_ (.A1(_0228_),
    .A2(_0229_),
    .Y(_0024_),
    .B1(net227));
 sg13g2_nand2b_1 _1729_ (.Y(_0230_),
    .B(state_q_1_),
    .A_N(_0227_));
 sg13g2_inv_1 _1730_ (.Y(_0231_),
    .A(state_q_1_));
 sg13g2_o21ai_1 _1731_ (.B1(\state_q_0__$_NOT__A_Y ),
    .Y(_0232_),
    .A1(state_q_0_),
    .A2(_0223_));
 sg13g2_nor2b_1 _1732_ (.A(state_q_2_),
    .B_N(_0232_),
    .Y(_0233_));
 sg13g2_nand4_1 _1733_ (.B(_0340_),
    .C(_0227_),
    .A(_0231_),
    .Y(_0234_),
    .D(_0233_));
 sg13g2_a21oi_1 _1734_ (.A1(_0230_),
    .A2(_0234_),
    .Y(_0025_),
    .B1(net227));
 sg13g2_nand2b_1 _1735_ (.Y(_0235_),
    .B(state_q_2_),
    .A_N(_0227_));
 sg13g2_nand3_1 _1736_ (.B(dmi_req_33_),
    .C(_0227_),
    .A(_0340_),
    .Y(_0236_));
 sg13g2_a21oi_1 _1737_ (.A1(_0235_),
    .A2(_0236_),
    .Y(_0026_),
    .B1(net227));
 sg13g2_nand2b_1 _1738_ (.Y(tdo_oe_o_reg_D),
    .B(_0220_),
    .A_N(net155));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[0]_reg_4  (.L_HI(net4));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/_4__3  (.L_HI(net3));
 sg13g2_dfrbp_2 address_q_0__reg (.RESET_B(net373),
    .D(_0027_),
    .Q(address_q_0_),
    .Q_N(_0801_),
    .CLK(net426));
 sg13g2_dfrbp_1 address_q_1__reg (.CLK(net426),
    .RESET_B(net374),
    .D(_0028_),
    .Q_N(_0800_),
    .Q(address_q_1_));
 sg13g2_dfrbp_2 address_q_2__reg (.RESET_B(net377),
    .D(_0029_),
    .Q(address_q_2_),
    .Q_N(_0799_),
    .CLK(net431));
 sg13g2_dfrbp_1 address_q_3__reg (.CLK(net427),
    .RESET_B(net374),
    .D(_0030_),
    .Q_N(_0798_),
    .Q(address_q_3_));
 sg13g2_dfrbp_1 address_q_4__reg (.CLK(net427),
    .RESET_B(net374),
    .D(_0031_),
    .Q_N(_0797_),
    .Q(address_q_4_));
 sg13g2_dfrbp_1 address_q_5__reg (.CLK(net432),
    .RESET_B(net377),
    .D(_0032_),
    .Q_N(_0796_),
    .Q(address_q_5_));
 sg13g2_dfrbp_1 address_q_6__reg (.CLK(net432),
    .RESET_B(net377),
    .D(_0033_),
    .Q_N(_0795_),
    .Q(address_q_6_));
 sg13g2_dfrbp_2 data_q_0__reg (.RESET_B(net364),
    .D(_0034_),
    .Q(data_q_0_),
    .Q_N(_0794_),
    .CLK(net414));
 sg13g2_dfrbp_2 data_q_10__reg (.RESET_B(net364),
    .D(_0035_),
    .Q(data_q_10_),
    .Q_N(_0793_),
    .CLK(net415));
 sg13g2_dfrbp_2 data_q_11__reg (.RESET_B(net358),
    .D(_0036_),
    .Q(data_q_11_),
    .Q_N(_0792_),
    .CLK(net415));
 sg13g2_dfrbp_2 data_q_12__reg (.RESET_B(net361),
    .D(_0037_),
    .Q(data_q_12_),
    .Q_N(_0791_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_13__reg (.RESET_B(net368),
    .D(_0038_),
    .Q(data_q_13_),
    .Q_N(_0790_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_14__reg (.RESET_B(net368),
    .D(_0039_),
    .Q(data_q_14_),
    .Q_N(_0789_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_15__reg (.RESET_B(net368),
    .D(_0040_),
    .Q(data_q_15_),
    .Q_N(_0788_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_16__reg (.RESET_B(net370),
    .D(_0041_),
    .Q(data_q_16_),
    .Q_N(_0787_),
    .CLK(net421));
 sg13g2_dfrbp_2 data_q_17__reg (.RESET_B(net370),
    .D(_0042_),
    .Q(data_q_17_),
    .Q_N(_0786_),
    .CLK(net421));
 sg13g2_dfrbp_2 data_q_18__reg (.RESET_B(net369),
    .D(_0043_),
    .Q(data_q_18_),
    .Q_N(_0785_),
    .CLK(net420));
 sg13g2_dfrbp_2 data_q_19__reg (.RESET_B(net365),
    .D(_0044_),
    .Q(data_q_19_),
    .Q_N(_0784_),
    .CLK(net417));
 sg13g2_dfrbp_2 data_q_1__reg (.RESET_B(net373),
    .D(_0045_),
    .Q(data_q_1_),
    .Q_N(_0783_),
    .CLK(net426));
 sg13g2_dfrbp_2 data_q_20__reg (.RESET_B(net365),
    .D(_0046_),
    .Q(data_q_20_),
    .Q_N(_0782_),
    .CLK(net417));
 sg13g2_dfrbp_2 data_q_21__reg (.RESET_B(net369),
    .D(_0047_),
    .Q(data_q_21_),
    .Q_N(_0781_),
    .CLK(net420));
 sg13g2_dfrbp_2 data_q_22__reg (.RESET_B(net370),
    .D(_0048_),
    .Q(data_q_22_),
    .Q_N(_0780_),
    .CLK(net421));
 sg13g2_dfrbp_2 data_q_23__reg (.RESET_B(net373),
    .D(_0049_),
    .Q(data_q_23_),
    .Q_N(_0779_),
    .CLK(net426));
 sg13g2_dfrbp_2 data_q_24__reg (.RESET_B(net373),
    .D(_0050_),
    .Q(data_q_24_),
    .Q_N(_0778_),
    .CLK(net426));
 sg13g2_dfrbp_2 data_q_25__reg (.RESET_B(net376),
    .D(_0051_),
    .Q(data_q_25_),
    .Q_N(_0777_),
    .CLK(net431));
 sg13g2_dfrbp_2 data_q_26__reg (.RESET_B(net370),
    .D(_0052_),
    .Q(data_q_26_),
    .Q_N(_0776_),
    .CLK(net422));
 sg13g2_dfrbp_2 data_q_27__reg (.RESET_B(net376),
    .D(_0053_),
    .Q(data_q_27_),
    .Q_N(_0775_),
    .CLK(net431));
 sg13g2_dfrbp_2 data_q_28__reg (.RESET_B(net370),
    .D(_0054_),
    .Q(data_q_28_),
    .Q_N(_0774_),
    .CLK(net422));
 sg13g2_dfrbp_2 data_q_29__reg (.RESET_B(net371),
    .D(_0055_),
    .Q(data_q_29_),
    .Q_N(_0773_),
    .CLK(net421));
 sg13g2_dfrbp_2 data_q_2__reg (.RESET_B(net376),
    .D(_0056_),
    .Q(data_q_2_),
    .Q_N(_0772_),
    .CLK(net431));
 sg13g2_dfrbp_2 data_q_30__reg (.RESET_B(net365),
    .D(_0057_),
    .Q(data_q_30_),
    .Q_N(_0771_),
    .CLK(net417));
 sg13g2_dfrbp_2 data_q_31__reg (.RESET_B(net365),
    .D(_0058_),
    .Q(data_q_31_),
    .Q_N(_0770_),
    .CLK(net418));
 sg13g2_dfrbp_2 data_q_3__reg (.RESET_B(net376),
    .D(_0059_),
    .Q(data_q_3_),
    .Q_N(_0769_),
    .CLK(net431));
 sg13g2_dfrbp_2 data_q_4__reg (.RESET_B(net366),
    .D(_0060_),
    .Q(data_q_4_),
    .Q_N(_0768_),
    .CLK(net418));
 sg13g2_dfrbp_2 data_q_5__reg (.RESET_B(net365),
    .D(_0061_),
    .Q(data_q_5_),
    .Q_N(_0767_),
    .CLK(net417));
 sg13g2_dfrbp_2 data_q_6__reg (.RESET_B(net368),
    .D(_0062_),
    .Q(data_q_6_),
    .Q_N(_0766_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_7__reg (.RESET_B(net361),
    .D(_0063_),
    .Q(data_q_7_),
    .Q_N(_0765_),
    .CLK(net419));
 sg13g2_dfrbp_2 data_q_8__reg (.RESET_B(net364),
    .D(_0064_),
    .Q(data_q_8_),
    .Q_N(_0764_),
    .CLK(net413));
 sg13g2_dfrbp_2 data_q_9__reg (.RESET_B(net364),
    .D(_0065_),
    .Q(data_q_9_),
    .Q_N(_0802_),
    .CLK(net415));
 sg13g2_dfrbp_1 dmi_10__reg (.CLK(net415),
    .RESET_B(net364),
    .D(dr_d_10_),
    .Q_N(_0803_),
    .Q(dmi_10_));
 sg13g2_dfrbp_1 dmi_11__reg (.CLK(net414),
    .RESET_B(net364),
    .D(dr_d_11_),
    .Q_N(_0804_),
    .Q(dmi_11_));
 sg13g2_dfrbp_1 dmi_12__reg (.CLK(net415),
    .RESET_B(net364),
    .D(dr_d_12_),
    .Q_N(_0805_),
    .Q(dmi_12_));
 sg13g2_dfrbp_1 dmi_13__reg (.CLK(net415),
    .RESET_B(net364),
    .D(dr_d_13_),
    .Q_N(_0806_),
    .Q(dmi_13_));
 sg13g2_dfrbp_1 dmi_14__reg (.CLK(net419),
    .RESET_B(net368),
    .D(dr_d_14_),
    .Q_N(_0807_),
    .Q(dmi_14_));
 sg13g2_dfrbp_1 dmi_15__reg (.CLK(net419),
    .RESET_B(net368),
    .D(dr_d_15_),
    .Q_N(_0808_),
    .Q(dmi_15_));
 sg13g2_dfrbp_1 dmi_16__reg (.CLK(net420),
    .RESET_B(net368),
    .D(dr_d_16_),
    .Q_N(_0809_),
    .Q(dmi_16_));
 sg13g2_dfrbp_1 dmi_17__reg (.CLK(net421),
    .RESET_B(net370),
    .D(dr_d_17_),
    .Q_N(_0810_),
    .Q(dmi_17_));
 sg13g2_dfrbp_1 dmi_18__reg (.CLK(net421),
    .RESET_B(net371),
    .D(dr_d_18_),
    .Q_N(_0811_),
    .Q(dmi_18_));
 sg13g2_dfrbp_1 dmi_19__reg (.CLK(net421),
    .RESET_B(net370),
    .D(dr_d_19_),
    .Q_N(_0812_),
    .Q(dmi_19_));
 sg13g2_dfrbp_1 dmi_1__reg (.CLK(net408),
    .RESET_B(net361),
    .D(dr_d_1_),
    .Q_N(\state_q_0__reg_E_$_AND__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_NOT__Y_A_$_OR__Y_B ),
    .Q(dmi_1_));
 sg13g2_dfrbp_1 dmi_20__reg (.CLK(net420),
    .RESET_B(net369),
    .D(dr_d_20_),
    .Q_N(_0813_),
    .Q(dmi_20_));
 sg13g2_dfrbp_1 dmi_21__reg (.CLK(net416),
    .RESET_B(net365),
    .D(dr_d_21_),
    .Q_N(_0814_),
    .Q(dmi_21_));
 sg13g2_dfrbp_1 dmi_22__reg (.CLK(net416),
    .RESET_B(net367),
    .D(dr_d_22_),
    .Q_N(_0815_),
    .Q(dmi_22_));
 sg13g2_dfrbp_1 dmi_23__reg (.CLK(net416),
    .RESET_B(net367),
    .D(dr_d_23_),
    .Q_N(_0816_),
    .Q(dmi_23_));
 sg13g2_dfrbp_1 dmi_24__reg (.CLK(net417),
    .RESET_B(net370),
    .D(dr_d_24_),
    .Q_N(_0817_),
    .Q(dmi_24_));
 sg13g2_dfrbp_1 dmi_25__reg (.CLK(net418),
    .RESET_B(net366),
    .D(dr_d_25_),
    .Q_N(_0818_),
    .Q(dmi_25_));
 sg13g2_dfrbp_1 dmi_26__reg (.CLK(net418),
    .RESET_B(net373),
    .D(dr_d_26_),
    .Q_N(_0819_),
    .Q(dmi_26_));
 sg13g2_dfrbp_1 dmi_27__reg (.CLK(net422),
    .RESET_B(net376),
    .D(dr_d_27_),
    .Q_N(_0820_),
    .Q(dmi_27_));
 sg13g2_dfrbp_1 dmi_28__reg (.CLK(net422),
    .RESET_B(net371),
    .D(dr_d_28_),
    .Q_N(_0821_),
    .Q(dmi_28_));
 sg13g2_dfrbp_1 dmi_29__reg (.CLK(net422),
    .RESET_B(net376),
    .D(dr_d_29_),
    .Q_N(_0822_),
    .Q(dmi_29_));
 sg13g2_dfrbp_2 dmi_2__reg (.RESET_B(net366),
    .D(dr_d_2_),
    .Q(dmi_2_),
    .Q_N(_0823_),
    .CLK(net418));
 sg13g2_dfrbp_1 dmi_30__reg (.CLK(net422),
    .RESET_B(net371),
    .D(dr_d_30_),
    .Q_N(_0824_),
    .Q(dmi_30_));
 sg13g2_dfrbp_1 dmi_31__reg (.CLK(net421),
    .RESET_B(net371),
    .D(dr_d_31_),
    .Q_N(_0825_),
    .Q(dmi_31_));
 sg13g2_dfrbp_2 dmi_32__reg (.RESET_B(net365),
    .D(dr_d_32_),
    .Q(dmi_32_),
    .Q_N(_0826_),
    .CLK(net418));
 sg13g2_dfrbp_1 dmi_33__reg (.CLK(net417),
    .RESET_B(net366),
    .D(dr_d_33_),
    .Q_N(_0827_),
    .Q(dmi_33_));
 sg13g2_dfrbp_1 dmi_34__reg (.CLK(net426),
    .RESET_B(net373),
    .D(dr_d_34_),
    .Q_N(_0828_),
    .Q(dmi_34_));
 sg13g2_dfrbp_1 dmi_35__reg (.CLK(net427),
    .RESET_B(net373),
    .D(dr_d_35_),
    .Q_N(_0829_),
    .Q(dmi_35_));
 sg13g2_dfrbp_1 dmi_36__reg (.CLK(net432),
    .RESET_B(net377),
    .D(dr_d_36_),
    .Q_N(_0830_),
    .Q(dmi_36_));
 sg13g2_dfrbp_1 dmi_37__reg (.CLK(net427),
    .RESET_B(net374),
    .D(dr_d_37_),
    .Q_N(_0831_),
    .Q(dmi_37_));
 sg13g2_dfrbp_1 dmi_38__reg (.CLK(net427),
    .RESET_B(net374),
    .D(dr_d_38_),
    .Q_N(_0832_),
    .Q(dmi_38_));
 sg13g2_dfrbp_1 dmi_39__reg (.CLK(net432),
    .RESET_B(net377),
    .D(dr_d_39_),
    .Q_N(_0833_),
    .Q(dmi_39_));
 sg13g2_dfrbp_1 dmi_3__reg (.CLK(net426),
    .RESET_B(net374),
    .D(dr_d_3_),
    .Q_N(_0834_),
    .Q(dmi_3_));
 sg13g2_dfrbp_1 dmi_40__reg (.CLK(net431),
    .RESET_B(net376),
    .D(dr_d_40_),
    .Q_N(_0835_),
    .Q(dmi_40_));
 sg13g2_dfrbp_1 dmi_4__reg (.CLK(net431),
    .RESET_B(net374),
    .D(dr_d_4_),
    .Q_N(_0836_),
    .Q(dmi_4_));
 sg13g2_dfrbp_1 dmi_5__reg (.CLK(net426),
    .RESET_B(net373),
    .D(dr_d_5_),
    .Q_N(_0837_),
    .Q(dmi_5_));
 sg13g2_dfrbp_1 dmi_6__reg (.CLK(net417),
    .RESET_B(net366),
    .D(dr_d_6_),
    .Q_N(_0838_),
    .Q(dmi_6_));
 sg13g2_dfrbp_1 dmi_7__reg (.CLK(net417),
    .RESET_B(net365),
    .D(dr_d_7_),
    .Q_N(_0839_),
    .Q(dmi_7_));
 sg13g2_dfrbp_1 dmi_8__reg (.CLK(net415),
    .RESET_B(net368),
    .D(dr_d_8_),
    .Q_N(_0840_),
    .Q(dmi_8_));
 sg13g2_dfrbp_1 dmi_9__reg (.CLK(net415),
    .RESET_B(net358),
    .D(dr_d_9_),
    .Q_N(_0763_),
    .Q(dmi_9_));
 sg13g2_dfrbp_2 dmi_rst_no_reg (.RESET_B(net386),
    .D(_0012_),
    .Q(_0001_),
    .Q_N(dmi_rst_no),
    .CLK(clknet_5_28__leaf_clk_i));
 sg13g2_dfrbp_1 dtmcs_q_10__reg (.CLK(net404),
    .RESET_B(net358),
    .D(dtmcs_d_10_),
    .Q_N(_0841_),
    .Q(dtmcs_q_10_));
 sg13g2_dfrbp_1 dtmcs_q_11__reg (.CLK(net404),
    .RESET_B(net358),
    .D(dtmcs_d_11_),
    .Q_N(_0842_),
    .Q(dtmcs_q_11_));
 sg13g2_dfrbp_1 dtmcs_q_12__reg (.CLK(net404),
    .RESET_B(net358),
    .D(dtmcs_d_12_),
    .Q_N(_0843_),
    .Q(dtmcs_q_12_));
 sg13g2_dfrbp_1 dtmcs_q_13__reg (.CLK(net402),
    .RESET_B(net359),
    .D(dtmcs_d_13_),
    .Q_N(_0844_),
    .Q(dtmcs_q_13_));
 sg13g2_dfrbp_1 dtmcs_q_14__reg (.CLK(net403),
    .RESET_B(net355),
    .D(dtmcs_d_14_),
    .Q_N(_0845_),
    .Q(dtmcs_q_14_));
 sg13g2_dfrbp_1 dtmcs_q_15__reg (.CLK(net403),
    .RESET_B(net355),
    .D(dtmcs_d_15_),
    .Q_N(_0846_),
    .Q(dtmcs_q_15_));
 sg13g2_dfrbp_1 dtmcs_q_16__reg (.CLK(net400),
    .RESET_B(net357),
    .D(dtmcs_d_16_),
    .Q_N(_0847_),
    .Q(dtmcs_q_16_));
 sg13g2_dfrbp_1 dtmcs_q_17__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_17_),
    .Q_N(_0848_),
    .Q(dtmcs_q_17_));
 sg13g2_dfrbp_1 dtmcs_q_18__reg (.CLK(net403),
    .RESET_B(net357),
    .D(dtmcs_d_18_),
    .Q_N(_0849_),
    .Q(dtmcs_q_18_));
 sg13g2_dfrbp_1 dtmcs_q_19__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_19_),
    .Q_N(_0850_),
    .Q(dtmcs_q_19_));
 sg13g2_dfrbp_1 dtmcs_q_1__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_1_),
    .Q_N(_0851_),
    .Q(dtmcs_q_1_));
 sg13g2_dfrbp_1 dtmcs_q_20__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_20_),
    .Q_N(_0852_),
    .Q(dtmcs_q_20_));
 sg13g2_dfrbp_1 dtmcs_q_21__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_21_),
    .Q_N(_0853_),
    .Q(dtmcs_q_21_));
 sg13g2_dfrbp_1 dtmcs_q_22__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_22_),
    .Q_N(_0854_),
    .Q(dtmcs_q_22_));
 sg13g2_dfrbp_1 dtmcs_q_23__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_23_),
    .Q_N(_0855_),
    .Q(dtmcs_q_23_));
 sg13g2_dfrbp_1 dtmcs_q_24__reg (.CLK(net402),
    .RESET_B(net355),
    .D(dtmcs_d_24_),
    .Q_N(_0856_),
    .Q(dtmcs_q_24_));
 sg13g2_dfrbp_1 dtmcs_q_25__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_25_),
    .Q_N(_0857_),
    .Q(dtmcs_q_25_));
 sg13g2_dfrbp_1 dtmcs_q_26__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_26_),
    .Q_N(_0858_),
    .Q(dtmcs_q_26_));
 sg13g2_dfrbp_1 dtmcs_q_27__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_27_),
    .Q_N(_0859_),
    .Q(dtmcs_q_27_));
 sg13g2_dfrbp_1 dtmcs_q_28__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_28_),
    .Q_N(_0860_),
    .Q(dtmcs_q_28_));
 sg13g2_dfrbp_1 dtmcs_q_29__reg (.CLK(net400),
    .RESET_B(net351),
    .D(dtmcs_d_29_),
    .Q_N(_0861_),
    .Q(dtmcs_q_29_));
 sg13g2_dfrbp_1 dtmcs_q_2__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_2_),
    .Q_N(_0862_),
    .Q(dtmcs_q_2_));
 sg13g2_dfrbp_1 dtmcs_q_30__reg (.CLK(net401),
    .RESET_B(net351),
    .D(dtmcs_d_30_),
    .Q_N(_0863_),
    .Q(dtmcs_q_30_));
 sg13g2_dfrbp_1 dtmcs_q_31__reg (.CLK(net401),
    .RESET_B(net351),
    .D(dtmcs_d_31_),
    .Q_N(_0864_),
    .Q(dtmcs_q_31_));
 sg13g2_dfrbp_1 dtmcs_q_3__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_3_),
    .Q_N(_0865_),
    .Q(dtmcs_q_3_));
 sg13g2_dfrbp_1 dtmcs_q_4__reg (.CLK(net414),
    .RESET_B(net356),
    .D(dtmcs_d_4_),
    .Q_N(_0866_),
    .Q(dtmcs_q_4_));
 sg13g2_dfrbp_1 dtmcs_q_5__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_5_),
    .Q_N(_0867_),
    .Q(dtmcs_q_5_));
 sg13g2_dfrbp_1 dtmcs_q_6__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_6_),
    .Q_N(_0868_),
    .Q(dtmcs_q_6_));
 sg13g2_dfrbp_1 dtmcs_q_7__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_7_),
    .Q_N(_0869_),
    .Q(dtmcs_q_7_));
 sg13g2_dfrbp_1 dtmcs_q_8__reg (.CLK(net413),
    .RESET_B(net356),
    .D(dtmcs_d_8_),
    .Q_N(_0870_),
    .Q(dtmcs_q_8_));
 sg13g2_dfrbp_1 dtmcs_q_9__reg (.CLK(net402),
    .RESET_B(net357),
    .D(dtmcs_d_9_),
    .Q_N(_0762_),
    .Q(dtmcs_q_9_));
 sg13g2_dfrbp_1 error_q_0__reg (.CLK(net404),
    .RESET_B(net358),
    .D(_0066_),
    .Q_N(\error_q_0__$_NOT__A_Y ),
    .Q(error_q_0_));
 sg13g2_dfrbp_1 error_q_1__reg (.CLK(net405),
    .RESET_B(net358),
    .D(_0067_),
    .Q_N(\error_q_1__$_NOT__A_Y ),
    .Q(error_q_1_));
 sg13g2_dfrbp_1 \i_dmi_cdc.core_clear_pending_q_reg  (.CLK(clknet_5_28__leaf_clk_i),
    .RESET_B(net386),
    .D(\i_dmi_cdc.core_clear_pending ),
    .Q_N(\i_dmi_cdc.clear_pending_rise_edge_detect_$_AND__Y_A ),
    .Q(\i_dmi_cdc.core_clear_pending_q ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/_4_  (.A(\i_dmi_cdc.core_clear_pending ),
    .B_N(dmi_req_ready_i),
    .Y(\i_dmi_cdc.i_cdc_req/i_dst_ready_i ));
 sg13g2_nor2b_2 \i_dmi_cdc.i_cdc_req/_5_  (.A(\i_dmi_cdc.core_clear_pending ),
    .B_N(\i_dmi_cdc.i_cdc_req/s_dst_valid ),
    .Y(dmi_req_valid_o));
 sg13g2_nor2b_2 \i_dmi_cdc.i_cdc_req/_6_  (.A(\i_dmi_cdc.i_cdc_req/src_clear_pending_o ),
    .B_N(\i_dmi_cdc.i_cdc_req/s_src_ready ),
    .Y(dmi_req_ready));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/_7_  (.A(\i_dmi_cdc.i_cdc_req/src_clear_pending_o ),
    .B_N(dmi_req_valid),
    .Y(\i_dmi_cdc.i_cdc_req/i_src_valid_i ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_080_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_081_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_082_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_083_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ));
 sg13g2_buf_4 fanout205 (.X(net205),
    .A(net209));
 sg13g2_buf_2 fanout204 (.A(\i_dmi_cdc.i_cdc_resp/i_src/_036_ ),
    .X(net204));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(net204));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_087_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .A(net343));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(net204));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(\i_dmi_cdc.i_cdc_resp/i_src/_036_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_090_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_091_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_092_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_093_  (.Y(\i_dmi_cdc.i_cdc_req/s_src_clear_req ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_094_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ));
 sg13g2_buf_2 fanout200 (.A(net201),
    .X(net200));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_096_  (.A(net342),
    .B(net340),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_097_  (.B1(net344),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_098_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ),
    .B(net341),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_099_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_100_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_101_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ),
    .B(net344),
    .A_N(net341));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_102_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_103_  (.A(net341),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_104_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_105_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_106_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_107_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_108_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ),
    .A(net344),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ));
 sg13g2_or4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_109_  (.A(net344),
    .B(net342),
    .C(net340),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_110_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_111_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_112_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ),
    .A(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_113_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .A_N(net342));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_114_  (.A(net341),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ));
 sg13g2_or3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_115_  (.A(net343),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .C(net340),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_116_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_117_  (.A(\i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ),
    .B(net344),
    .C(net342),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_118_  (.B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .C1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_119_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_120_  (.A(net340),
    .B(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_121_  (.A(\i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ),
    .B(net343),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_122_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ),
    .A1(net343),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_123_  (.A(net235),
    .B(net344),
    .C(net342),
    .D(net340),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_124_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_125_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_126_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_127_  (.B1(net340),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ),
    .A1(net344),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_128_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_129_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_130_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_131_  (.A(\i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ),
    .B(net343),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_132_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B1(net342),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_133_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_134_  (.B(net343),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_135_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ),
    .A1(net235),
    .A2(net343));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_136_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_137_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_138_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_072_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_139_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_072_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_140_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(net343),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_073_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_141_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_025_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_074_ ),
    .A1(net342),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_073_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_142_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_075_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_143_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_076_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_075_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_074_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_144_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_076_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_077_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_145_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ),
    .A1(net342),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_077_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_146_  (.A(net340),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_078_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_147_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_079_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_075_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_148_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_078_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_079_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_149_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_150_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_151_  (.B1(net340),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_152_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_153_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_154_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_155_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_012_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_156_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_013_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_012_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_157_  (.Y(\i_dmi_cdc.i_cdc_req/src_clear_pending_o ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_013_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_158_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_159_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_015_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_160_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ),
    .A1(\i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_015_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_161_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_162_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_163_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_164_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ));
 sg13g2_nand2b_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_13_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_14_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_15_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_16_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_17_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_18_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_19_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_20_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_21_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_22_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_23_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_24_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_25_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_26_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/async_ack_o_reg  (.CLK(net433),
    .RESET_B(net377),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_12_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_ack ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0__reg  (.CLK(net437),
    .RESET_B(net377),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_req ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/serial_o_reg  (.CLK(net433),
    .RESET_B(net378),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__reg  (.CLK(net434),
    .RESET_B(net378),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__reg  (.CLK(net434),
    .RESET_B(net378),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_21_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_22_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_23_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/req_src_d ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_24_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_25_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_26_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_27_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_28_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_29_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_30_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_1_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_31_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_32_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_33_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_34_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_35_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_36_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_37_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_38_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_39_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_40_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_41_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_42_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_data_o[0]_reg  (.RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .CLK(net433));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_data_o[1]_reg  (.RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_20_ ),
    .CLK(net433));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_req_o_reg  (.CLK(net423),
    .RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_req ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_01_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0__reg  (.CLK(net423),
    .RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/serial_o_reg  (.CLK(net423),
    .RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__reg  (.RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .CLK(net423));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__reg  (.RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .CLK(net423));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0__reg  (.CLK(net423),
    .RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__reg  (.RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .CLK(net423));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__reg  (.RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .CLK(net424));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__reg  (.RESET_B(net372),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .CLK(net423));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__reg  (.CLK(net433),
    .RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__reg  (.CLK(net433),
    .RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(net201));
 sg13g2_buf_2 fanout198 (.A(_0548_),
    .X(net198));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_074_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .B(net336),
    .A(net338));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(net198));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_076_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_077_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .A1(net337));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_078_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_079_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_080_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_081_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_082_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_083_  (.Y(\i_dmi_cdc.i_cdc_req/s_dst_clear_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_084_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_085_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ));
 sg13g2_buf_2 fanout196 (.A(net197),
    .X(net196));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_087_  (.B1(net339),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_088_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A(net336));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_089_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_090_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_091_  (.A1(net336),
    .A2(net337),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_092_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_093_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_094_  (.A(net337),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_095_  (.A(net336),
    .B(net335),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_096_  (.A(net339),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_097_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_098_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .A1(net335),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_099_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .A(\i_dmi_cdc.i_cdc_req/s_dst_clear_ack_q ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_100_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A(net338));
 sg13g2_nand4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_101_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ),
    .D(net336));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_102_  (.A(net339),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_103_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_104_  (.A(net335),
    .B(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ));
 sg13g2_and4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_105_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net338),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_106_  (.B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ),
    .C1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_107_  (.A(net336),
    .B(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_108_  (.A(net1),
    .B(net338),
    .C(net337),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_109_  (.A1(net338),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_110_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .B(net335),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_111_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_112_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ),
    .A(net339),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_113_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_114_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A1(\i_dmi_cdc.i_cdc_req/s_dst_clear_ack_q ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_115_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_116_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_117_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_118_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net338),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_119_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ),
    .A1(net337),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_120_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_121_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_122_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ),
    .A(net338),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_123_  (.B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ),
    .C1(net335),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_124_  (.A0(net337),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_125_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net338));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_126_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ),
    .B(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ),
    .A_N(net337));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_127_  (.B1(net336),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_128_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_129_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_130_  (.A(net336),
    .B(net335),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_131_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_132_  (.A0(net335),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_133_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .A1(net335),
    .S(net339),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_134_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_135_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_136_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_137_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_138_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_139_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_140_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_141_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_142_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_143_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ),
    .Y(\i_dmi_cdc.core_clear_pending ),
    .A1(net337),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_144_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_145_  (.B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .C1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_146_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_147_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_148_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ));
 sg13g2_nand2b_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_13_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_14_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_15_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_16_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_17_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_18_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_19_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_20_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_21_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_22_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_23_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_24_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_25_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_26_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/async_ack_o_reg  (.CLK(clknet_5_15__leaf_clk_i),
    .RESET_B(net387),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_12_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_ack ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0__reg  (.CLK(clknet_5_14__leaf_clk_i),
    .RESET_B(net387),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_req ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/serial_o_reg  (.CLK(clknet_5_14__leaf_clk_i),
    .RESET_B(net387),
    .D(net446),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__reg  (.CLK(clknet_5_26__leaf_clk_i),
    .RESET_B(net387),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__reg  (.CLK(clknet_5_26__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_21_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_22_  (.B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_23_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/req_src_d ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_24_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_25_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_26_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_27_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_28_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_29_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_30_  (.A0(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_1_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_31_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_32_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_33_  (.B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .C(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_34_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_35_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_36_  (.X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_37_  (.A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_38_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_39_  (.A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_40_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_41_  (.Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ),
    .B2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_42_  (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .Y(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_data_o[0]_reg  (.CLK(clknet_5_24__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_data_o[1]_reg  (.RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_20_ ),
    .CLK(clknet_5_25__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_req_o_reg  (.CLK(clknet_5_30__leaf_clk_i),
    .RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_b2a_req ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_01_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0__reg  (.CLK(clknet_5_24__leaf_clk_i),
    .RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/async_a2b_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/serial_o_reg  (.RESET_B(net384),
    .D(net440),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_0_ ),
    .CLK(clknet_5_30__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__reg  (.RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .CLK(clknet_5_30__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__reg  (.RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .CLK(clknet_5_25__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0__reg  (.CLK(clknet_5_27__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__reg  (.CLK(clknet_5_25__leaf_clk_i),
    .RESET_B(net384),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__reg  (.RESET_B(net387),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .CLK(clknet_5_27__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__reg  (.CLK(clknet_5_27__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__reg  (.CLK(clknet_5_26__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__reg  (.CLK(clknet_5_26__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_dst/_100_  (.A(\i_dmi_cdc.i_cdc_req/s_dst_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d_$_MUX__Y_A ),
    .Y(\i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_req/i_dst/_101_  (.A2(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ),
    .A1(\i_dmi_cdc.i_cdc_req/i_dst_ready_i ),
    .B1(\i_dmi_cdc.i_cdc_req/async_ack ),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_042_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_dst/_102_  (.Y(\i_dmi_cdc.i_cdc_req/i_dst/_043_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_dst_ready_i ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_req/i_dst/_103_  (.Y(\i_dmi_cdc.i_cdc_req/i_dst/_044_ ),
    .B1(\i_dmi_cdc.i_cdc_req/i_dst/_043_ ),
    .B2(\i_dmi_cdc.i_cdc_req/async_ack ),
    .A2(\i_dmi_cdc.i_cdc_req/i_dst/_042_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d_$_MUX__Y_A ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_req/i_dst/_104_  (.A(\i_dmi_cdc.i_cdc_req/s_dst_clear_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_dst/_044_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_dst/_000_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_req/i_dst/_105_  (.Y(\i_dmi_cdc.i_cdc_req/i_dst/_045_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_req/i_dst/_106_  (.B(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ),
    .C(\i_dmi_cdc.i_cdc_req/async_ack ),
    .Y(\i_dmi_cdc.i_cdc_req/i_dst/_046_ ),
    .A_N(\i_dmi_cdc.i_cdc_req/i_dst/req_synced ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_dst/_107_  (.B1(\i_dmi_cdc.i_cdc_req/i_dst/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_dst/_047_ ),
    .A1(\i_dmi_cdc.i_cdc_req/async_ack ),
    .A2(\i_dmi_cdc.i_cdc_req/i_dst/_045_ ));
 sg13g2_buf_4 fanout195 (.X(net195),
    .A(net197));
 sg13g2_buf_2 fanout194 (.A(net198),
    .X(net194));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_110_  (.A0(dmi_req_o_0_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_0_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_111_  (.A0(dmi_req_o_10_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_10_ ),
    .S(net295),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_112_  (.A0(dmi_req_o_11_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_11_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_11_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_113_  (.A0(dmi_req_o_12_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_12_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_12_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_114_  (.A0(dmi_req_o_13_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_13_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_13_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_115_  (.A0(dmi_req_o_14_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_14_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_14_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_116_  (.A0(dmi_req_o_15_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_15_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_15_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_117_  (.A0(dmi_req_o_16_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_16_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_16_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_118_  (.A0(dmi_req_o_17_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_17_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_17_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_119_  (.A0(dmi_req_o_18_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_18_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_18_ ));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(net194));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_121_  (.A0(dmi_req_o_19_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_19_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_19_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_122_  (.A0(dmi_req_o_1_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_1_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_1_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_123_  (.A0(dmi_req_o_20_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_20_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_20_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_124_  (.A0(dmi_req_o_21_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_21_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_21_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_125_  (.A0(dmi_req_o_22_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_22_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_22_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_126_  (.A0(dmi_req_o_23_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_23_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_23_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_127_  (.A0(dmi_req_o_24_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_24_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_24_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_128_  (.A0(dmi_req_o_25_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_25_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_25_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_129_  (.A0(dmi_req_o_26_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_26_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_26_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_130_  (.A0(dmi_req_o_27_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_27_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_27_ ));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(net194));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_132_  (.A0(dmi_req_o_28_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_28_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_28_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_133_  (.A0(dmi_req_o_29_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_29_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_29_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_134_  (.A0(dmi_req_o_2_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_2_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_2_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_135_  (.A0(dmi_req_o_30_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_30_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_30_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_136_  (.A0(dmi_req_o_31_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_31_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_31_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_137_  (.A0(dmi_req_o_32_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_32_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_32_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_138_  (.A0(dmi_req_o_33_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_33_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_33_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_139_  (.A0(dmi_req_o_34_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_34_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_34_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_140_  (.A0(dmi_req_o_35_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_35_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_35_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_141_  (.A0(dmi_req_o_36_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_36_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_36_ ));
 sg13g2_buf_1 fanout191 (.A(\i_dmi_cdc.i_cdc_req/i_src/_043_ ),
    .X(net191));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_143_  (.A0(dmi_req_o_37_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_37_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_37_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_144_  (.A0(dmi_req_o_38_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_38_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_38_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_145_  (.A0(dmi_req_o_39_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_39_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_39_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_146_  (.A0(dmi_req_o_3_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_3_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_3_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_147_  (.A0(dmi_req_o_40_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_40_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_40_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_148_  (.A0(dmi_req_o_4_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_4_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_4_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_149_  (.A0(dmi_req_o_5_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_5_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_5_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_150_  (.A0(dmi_req_o_6_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_6_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_6_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_151_  (.A0(dmi_req_o_7_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_7_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_7_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_152_  (.A0(dmi_req_o_8_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_8_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_8_ ));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_154_  (.A0(dmi_req_o_9_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_9_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/data_dst_d_9_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_155_  (.A0(dmi_req_o_0_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_0_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_001_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_156_  (.A0(dmi_req_o_10_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_10_ ),
    .S(net295),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_002_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_157_  (.A0(dmi_req_o_11_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_11_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_003_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_158_  (.A0(dmi_req_o_12_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_12_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_159_  (.A0(dmi_req_o_13_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_13_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_160_  (.A0(dmi_req_o_14_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_14_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_006_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_161_  (.A0(dmi_req_o_15_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_15_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_007_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_162_  (.A0(dmi_req_o_16_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_16_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_008_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_163_  (.A0(dmi_req_o_17_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_17_ ),
    .S(net301),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_009_ ));
 sg13g2_buf_2 fanout189 (.A(net190),
    .X(net189));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_165_  (.A0(dmi_req_o_18_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_18_ ),
    .S(net301),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_010_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_166_  (.A0(dmi_req_o_19_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_19_ ),
    .S(net296),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_011_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_167_  (.A0(dmi_req_o_1_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_1_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_012_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_168_  (.A0(dmi_req_o_20_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_20_ ),
    .S(net296),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_013_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_169_  (.A0(dmi_req_o_21_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_21_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_014_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_170_  (.A0(dmi_req_o_22_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_22_ ),
    .S(net302),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_015_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_171_  (.A0(dmi_req_o_23_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_23_ ),
    .S(net290),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_016_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_172_  (.A0(dmi_req_o_24_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_24_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_017_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_173_  (.A0(dmi_req_o_25_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_25_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_018_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_174_  (.A0(dmi_req_o_26_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_26_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_019_ ));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(net190));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_176_  (.A0(dmi_req_o_27_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_27_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_020_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_177_  (.A0(dmi_req_o_28_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_28_ ),
    .S(net302),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_021_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_178_  (.A0(dmi_req_o_29_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_29_ ),
    .S(net300),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_022_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_179_  (.A0(dmi_req_o_2_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_2_ ),
    .S(net295),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_023_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_180_  (.A0(dmi_req_o_30_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_30_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_024_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_181_  (.A0(dmi_req_o_31_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_31_ ),
    .S(net294),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_025_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_182_  (.A0(dmi_req_o_32_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_32_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_026_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_183_  (.A0(dmi_req_o_33_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_33_ ),
    .S(net301),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_027_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_184_  (.A0(dmi_req_o_34_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_34_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_028_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_185_  (.A0(dmi_req_o_35_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_35_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_029_ ));
 sg13g2_buf_2 fanout187 (.A(net190),
    .X(net187));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_187_  (.A0(dmi_req_o_36_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_36_ ),
    .S(net301),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_030_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_188_  (.A0(dmi_req_o_37_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_37_ ),
    .S(net295),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_031_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_189_  (.A0(dmi_req_o_38_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_38_ ),
    .S(net292),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_032_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_190_  (.A0(dmi_req_o_39_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_39_ ),
    .S(net298),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_033_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_191_  (.A0(dmi_req_o_3_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_3_ ),
    .S(net297),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_034_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_192_  (.A0(dmi_req_o_40_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_40_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_035_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_193_  (.A0(dmi_req_o_4_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_4_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_036_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_194_  (.A0(dmi_req_o_5_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_5_ ),
    .S(net293),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_037_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_195_  (.A0(dmi_req_o_6_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_6_ ),
    .S(net299),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_038_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_196_  (.A0(dmi_req_o_7_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_7_ ),
    .S(net302),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_039_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_197_  (.A0(dmi_req_o_8_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_8_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_040_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_dst/_198_  (.A0(dmi_req_o_9_),
    .A1(\i_dmi_cdc.i_cdc_req/async_data_9_ ),
    .S(net291),
    .X(\i_dmi_cdc.i_cdc_req/i_dst/_041_ ));
 sg13g2_xor2_1 \i_dmi_cdc.i_cdc_req/i_dst/_199_  (.B(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ),
    .A(\i_dmi_cdc.i_cdc_req/async_ack ),
    .X(\i_dmi_cdc.i_cdc_req/s_dst_valid ));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[0]_reg_45  (.L_HI(net45));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/async_ack_o_reg  (.RESET_B(net386),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_000_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/ack_dst_d_$_MUX__Y_A ),
    .CLK(clknet_5_24__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[0]_reg  (.RESET_B(net4),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_001_ ),
    .Q(dmi_req_o_0_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_097_ ),
    .CLK(clknet_5_17__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[10]_reg  (.RESET_B(net5),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_002_ ),
    .Q(dmi_req_o_10_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_096_ ),
    .CLK(clknet_5_16__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[11]_reg  (.RESET_B(net6),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_003_ ),
    .Q(dmi_req_o_11_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_095_ ),
    .CLK(clknet_5_17__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[12]_reg  (.RESET_B(net7),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_004_ ),
    .Q(dmi_req_o_12_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_094_ ),
    .CLK(clknet_5_19__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[13]_reg  (.RESET_B(net8),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_005_ ),
    .Q(dmi_req_o_13_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_093_ ),
    .CLK(clknet_5_31__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[14]_reg  (.RESET_B(net9),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_006_ ),
    .Q(dmi_req_o_14_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_092_ ),
    .CLK(clknet_5_16__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[15]_reg  (.RESET_B(net10),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_007_ ),
    .Q(dmi_req_o_15_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_091_ ),
    .CLK(clknet_5_22__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[16]_reg  (.RESET_B(net11),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_008_ ),
    .Q(dmi_req_o_16_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_090_ ),
    .CLK(clknet_5_20__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[17]_reg  (.RESET_B(net12),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_009_ ),
    .Q(dmi_req_o_17_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_089_ ),
    .CLK(clknet_5_29__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[18]_reg  (.RESET_B(net13),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_010_ ),
    .Q(dmi_req_o_18_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_088_ ),
    .CLK(clknet_5_29__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[19]_reg  (.RESET_B(net14),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_011_ ),
    .Q(dmi_req_o_19_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_087_ ),
    .CLK(clknet_5_20__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[1]_reg  (.RESET_B(net15),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_012_ ),
    .Q(dmi_req_o_1_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_086_ ),
    .CLK(clknet_5_22__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[20]_reg  (.RESET_B(net16),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_013_ ),
    .Q(dmi_req_o_20_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_085_ ),
    .CLK(clknet_5_20__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[21]_reg  (.RESET_B(net17),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_014_ ),
    .Q(dmi_req_o_21_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_084_ ),
    .CLK(clknet_5_18__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[22]_reg  (.RESET_B(net18),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_015_ ),
    .Q(dmi_req_o_22_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_083_ ),
    .CLK(clknet_5_29__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[23]_reg  (.RESET_B(net19),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_016_ ),
    .Q(dmi_req_o_23_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_082_ ),
    .CLK(clknet_5_23__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[24]_reg  (.RESET_B(net20),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_017_ ),
    .Q(dmi_req_o_24_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_081_ ),
    .CLK(clknet_5_21__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[25]_reg  (.RESET_B(net21),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_018_ ),
    .Q(dmi_req_o_25_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_080_ ),
    .CLK(clknet_5_17__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[26]_reg  (.RESET_B(net22),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_019_ ),
    .Q(dmi_req_o_26_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_079_ ),
    .CLK(clknet_5_20__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[27]_reg  (.RESET_B(net23),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_020_ ),
    .Q(dmi_req_o_27_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_078_ ),
    .CLK(clknet_5_19__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[28]_reg  (.RESET_B(net24),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_021_ ),
    .Q(dmi_req_o_28_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_077_ ),
    .CLK(clknet_5_28__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[29]_reg  (.RESET_B(net25),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_022_ ),
    .Q(dmi_req_o_29_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_076_ ),
    .CLK(clknet_5_31__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[2]_reg  (.RESET_B(net26),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_023_ ),
    .Q(dmi_req_o_2_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_075_ ),
    .CLK(clknet_5_16__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[30]_reg  (.RESET_B(net27),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_024_ ),
    .Q(dmi_req_o_30_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_074_ ),
    .CLK(clknet_5_22__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[31]_reg  (.RESET_B(net28),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_025_ ),
    .Q(dmi_req_o_31_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_073_ ),
    .CLK(clknet_5_22__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[32]_reg  (.RESET_B(net29),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_026_ ),
    .Q(dmi_req_o_32_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_072_ ),
    .CLK(clknet_5_18__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[33]_reg  (.RESET_B(net30),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_027_ ),
    .Q(dmi_req_o_33_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_071_ ),
    .CLK(clknet_5_31__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[34]_reg  (.RESET_B(net31),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_028_ ),
    .Q(dmi_req_o_34_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_070_ ),
    .CLK(clknet_5_23__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[35]_reg  (.RESET_B(net32),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_029_ ),
    .Q(dmi_req_o_35_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_069_ ),
    .CLK(clknet_5_23__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[36]_reg  (.RESET_B(net33),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_030_ ),
    .Q(dmi_req_o_36_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_068_ ),
    .CLK(clknet_5_29__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[37]_reg  (.RESET_B(net34),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_031_ ),
    .Q(dmi_req_o_37_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_067_ ),
    .CLK(clknet_5_17__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[38]_reg  (.RESET_B(net35),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_032_ ),
    .Q(dmi_req_o_38_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_066_ ),
    .CLK(clknet_5_23__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[39]_reg  (.RESET_B(net36),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_033_ ),
    .Q(dmi_req_o_39_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_065_ ),
    .CLK(clknet_5_19__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[3]_reg  (.RESET_B(net37),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_034_ ),
    .Q(dmi_req_o_3_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_064_ ),
    .CLK(clknet_5_19__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[40]_reg  (.RESET_B(net38),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_035_ ),
    .Q(dmi_req_o_40_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_063_ ),
    .CLK(clknet_5_18__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[4]_reg  (.RESET_B(net39),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_036_ ),
    .Q(dmi_req_o_4_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_062_ ),
    .CLK(clknet_5_21__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[5]_reg  (.RESET_B(net40),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_037_ ),
    .Q(dmi_req_o_5_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_061_ ),
    .CLK(clknet_5_16__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[6]_reg  (.RESET_B(net41),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_038_ ),
    .Q(dmi_req_o_6_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_060_ ),
    .CLK(clknet_5_18__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[7]_reg  (.RESET_B(net42),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_039_ ),
    .Q(dmi_req_o_7_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_059_ ),
    .CLK(clknet_5_30__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[8]_reg  (.RESET_B(net43),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_040_ ),
    .Q(dmi_req_o_8_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_058_ ),
    .CLK(clknet_5_21__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/data_o[9]_reg  (.RESET_B(net44),
    .D(\i_dmi_cdc.i_cdc_req/i_dst/_041_ ),
    .Q(dmi_req_o_9_),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_098_ ),
    .CLK(clknet_5_21__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_0__reg  (.CLK(clknet_5_15__leaf_clk_i),
    .RESET_B(net386),
    .D(\i_dmi_cdc.i_cdc_req/async_req ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_1__reg  (.CLK(clknet_5_15__leaf_clk_i),
    .RESET_B(net386),
    .D(net442),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/_2_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_dst/i_sync/serial_o_reg  (.CLK(clknet_5_24__leaf_clk_i),
    .RESET_B(net386),
    .D(net439),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_dst/req_synced ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1_reg  (.RESET_B(net386),
    .D(net441),
    .Q(\i_dmi_cdc.i_cdc_req/i_dst/req_synced_q1 ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_dst/_057_ ),
    .CLK(clknet_5_28__leaf_clk_i));
 sg13g2_xnor2_1 \i_dmi_cdc.i_cdc_req/i_src/_099_  (.Y(\i_dmi_cdc.i_cdc_req/s_src_ready ),
    .A(\i_dmi_cdc.i_cdc_req/async_req ),
    .B(\i_dmi_cdc.i_cdc_req/i_src/ack_synced ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_src/_100_  (.A(\i_dmi_cdc.i_cdc_req/s_src_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_src_valid_i ),
    .Y(\i_dmi_cdc.i_cdc_req/i_src/_042_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_req/i_src/_101_  (.A(\i_dmi_cdc.i_cdc_req/s_src_ready ),
    .B(\i_dmi_cdc.i_cdc_req/i_src/_042_ ),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_043_ ));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(net190));
 sg13g2_buf_2 fanout185 (.A(net191),
    .X(net185));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_104_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_0_ ),
    .A1(data_q_0_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_000_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_105_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_10_ ),
    .A1(data_q_10_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_001_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_106_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_11_ ),
    .A1(data_q_11_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_002_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_107_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_12_ ),
    .A1(data_q_12_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_003_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_108_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_13_ ),
    .A1(data_q_13_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_109_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_14_ ),
    .A1(data_q_14_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_110_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_15_ ),
    .A1(data_q_15_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_006_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_111_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_16_ ),
    .A1(data_q_16_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_007_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_112_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_17_ ),
    .A1(data_q_17_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_008_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_113_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_18_ ),
    .A1(data_q_18_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_009_ ));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(net191));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_115_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_19_ ),
    .A1(data_q_19_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_010_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_116_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_1_ ),
    .A1(data_q_1_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_011_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_117_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_20_ ),
    .A1(data_q_20_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_012_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_118_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_21_ ),
    .A1(data_q_21_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_013_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_119_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_22_ ),
    .A1(data_q_22_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_014_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_120_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_23_ ),
    .A1(data_q_23_),
    .S(net176),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_015_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_121_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_24_ ),
    .A1(data_q_24_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_016_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_122_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_25_ ),
    .A1(data_q_25_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_017_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_123_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_26_ ),
    .A1(data_q_26_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_018_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_124_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_27_ ),
    .A1(data_q_27_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_019_ ));
 sg13g2_buf_2 fanout183 (.A(net191),
    .X(net183));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_126_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_28_ ),
    .A1(data_q_28_),
    .S(net185),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_020_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_127_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_29_ ),
    .A1(data_q_29_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_021_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_128_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_2_ ),
    .A1(data_q_2_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_022_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_129_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_30_ ),
    .A1(data_q_30_),
    .S(net181),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_023_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_130_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_31_ ),
    .A1(data_q_31_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_024_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_131_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_32_ ),
    .A1(dmi_req_32_),
    .S(net187),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_025_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_132_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_33_ ),
    .A1(dmi_req_33_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_026_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_133_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_34_ ),
    .A1(address_q_0_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_027_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_134_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_35_ ),
    .A1(address_q_1_),
    .S(net176),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_028_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_135_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_36_ ),
    .A1(address_q_2_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_029_ ));
 sg13g2_buf_4 fanout182 (.X(net182),
    .A(net183));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_137_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_37_ ),
    .A1(address_q_3_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_030_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_138_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_38_ ),
    .A1(address_q_4_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_031_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_139_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_39_ ),
    .A1(address_q_5_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_032_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_140_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_3_ ),
    .A1(data_q_3_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_033_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_141_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_40_ ),
    .A1(address_q_6_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_034_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_142_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_4_ ),
    .A1(data_q_4_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_035_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_143_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_5_ ),
    .A1(data_q_5_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_036_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_144_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_6_ ),
    .A1(data_q_6_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_037_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_145_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_7_ ),
    .A1(data_q_7_),
    .S(net185),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_038_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_146_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_8_ ),
    .A1(data_q_8_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_039_ ));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_148_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_9_ ),
    .A1(data_q_9_),
    .S(net177),
    .X(\i_dmi_cdc.i_cdc_req/i_src/_040_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_req/i_src/_149_  (.A(\i_dmi_cdc.i_cdc_req/s_src_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_req/i_src/req_src_d_$_MUX__Y_A ),
    .Y(\i_dmi_cdc.i_cdc_req/i_src/req_src_d ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_src/_150_  (.A1(\i_dmi_cdc.i_cdc_req/i_src/req_src_d_$_MUX__Y_A ),
    .A2(\i_dmi_cdc.i_cdc_req/i_src_valid_i ),
    .Y(\i_dmi_cdc.i_cdc_req/i_src/_050_ ),
    .B1(\i_dmi_cdc.i_cdc_req/async_req ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_req/i_src/_151_  (.X(\i_dmi_cdc.i_cdc_req/i_src/_051_ ),
    .B(\i_dmi_cdc.i_cdc_req/i_src/_050_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_src/ack_synced ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_req/i_src/_152_  (.Y(\i_dmi_cdc.i_cdc_req/i_src/_052_ ),
    .A(\i_dmi_cdc.i_cdc_req/i_src_valid_i ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_req/i_src/_153_  (.B1(\i_dmi_cdc.i_cdc_req/async_req ),
    .Y(\i_dmi_cdc.i_cdc_req/i_src/_053_ ),
    .A1(\i_dmi_cdc.i_cdc_req/i_src/req_src_d_$_MUX__Y_A ),
    .A2(\i_dmi_cdc.i_cdc_req/i_src/_052_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_req/i_src/_154_  (.A1(\i_dmi_cdc.i_cdc_req/i_src/_051_ ),
    .A2(\i_dmi_cdc.i_cdc_req/i_src/_053_ ),
    .Y(\i_dmi_cdc.i_cdc_req/i_src/_041_ ),
    .B1(\i_dmi_cdc.i_cdc_req/s_src_clear_req ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_155_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_0_ ),
    .A1(data_q_0_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_156_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_10_ ),
    .A1(data_q_10_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_157_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_11_ ),
    .A1(data_q_11_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_11_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_158_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_12_ ),
    .A1(data_q_12_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_12_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_159_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_13_ ),
    .A1(data_q_13_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_13_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_160_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_14_ ),
    .A1(data_q_14_),
    .S(net187),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_14_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_161_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_15_ ),
    .A1(data_q_15_),
    .S(net179),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_15_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_162_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_16_ ),
    .A1(data_q_16_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_16_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_163_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_17_ ),
    .A1(data_q_17_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_17_ ));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(net182));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_165_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_18_ ),
    .A1(data_q_18_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_18_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_166_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_19_ ),
    .A1(data_q_19_),
    .S(net179),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_19_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_167_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_1_ ),
    .A1(data_q_1_),
    .S(net183),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_1_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_168_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_20_ ),
    .A1(data_q_20_),
    .S(net182),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_20_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_169_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_21_ ),
    .A1(data_q_21_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_21_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_170_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_22_ ),
    .A1(data_q_22_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_22_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_171_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_23_ ),
    .A1(data_q_23_),
    .S(net176),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_23_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_172_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_24_ ),
    .A1(data_q_24_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_24_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_173_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_25_ ),
    .A1(data_q_25_),
    .S(net187),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_25_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_174_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_26_ ),
    .A1(data_q_26_),
    .S(net181),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_26_ ));
 sg13g2_buf_2 fanout179 (.A(net183),
    .X(net179));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_176_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_27_ ),
    .A1(data_q_27_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_27_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_177_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_28_ ),
    .A1(data_q_28_),
    .S(net185),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_28_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_178_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_29_ ),
    .A1(data_q_29_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_29_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_179_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_2_ ),
    .A1(data_q_2_),
    .S(net183),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_2_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_180_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_30_ ),
    .A1(data_q_30_),
    .S(net181),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_30_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_181_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_31_ ),
    .A1(data_q_31_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_31_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_182_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_32_ ),
    .A1(dmi_req_32_),
    .S(net187),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_32_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_183_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_33_ ),
    .A1(dmi_req_33_),
    .S(net189),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_33_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_184_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_34_ ),
    .A1(address_q_0_),
    .S(net181),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_34_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_185_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_35_ ),
    .A1(address_q_1_),
    .S(net176),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_35_ ));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(net179));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_187_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_36_ ),
    .A1(address_q_2_),
    .S(net188),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_36_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_188_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_37_ ),
    .A1(address_q_3_),
    .S(net178),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_37_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_189_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_38_ ),
    .A1(address_q_4_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_38_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_190_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_39_ ),
    .A1(address_q_5_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_39_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_191_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_3_ ),
    .A1(data_q_3_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_3_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_192_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_40_ ),
    .A1(address_q_6_),
    .S(net184),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_40_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_193_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_4_ ),
    .A1(data_q_4_),
    .S(net175),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_4_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_194_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_5_ ),
    .A1(data_q_5_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_5_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_195_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_6_ ),
    .A1(data_q_6_),
    .S(net186),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_6_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_196_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_7_ ),
    .A1(data_q_7_),
    .S(net185),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_7_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_197_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_8_ ),
    .A1(data_q_8_),
    .S(net180),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_8_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_req/i_src/_198_  (.A0(\i_dmi_cdc.i_cdc_req/async_data_9_ ),
    .A1(data_q_9_),
    .S(net177),
    .X(\i_dmi_cdc.i_cdc_req/i_src/data_src_d_9_ ));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[0]_reg_86  (.L_HI(net86));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[0]_reg  (.RESET_B(net45),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_000_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_097_ ),
    .CLK(net430));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[10]_reg  (.CLK(net429),
    .RESET_B(net46),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_096_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_10_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[11]_reg  (.CLK(net429),
    .RESET_B(net47),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_002_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_095_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_11_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[12]_reg  (.CLK(net436),
    .RESET_B(net48),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_003_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_094_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_12_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[13]_reg  (.CLK(net437),
    .RESET_B(net49),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_004_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_093_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_13_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[14]_reg  (.CLK(net435),
    .RESET_B(net50),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_092_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_14_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[15]_reg  (.CLK(net428),
    .RESET_B(net51),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_091_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_15_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[16]_reg  (.CLK(net428),
    .RESET_B(net52),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_007_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_090_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_16_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[17]_reg  (.CLK(net437),
    .RESET_B(net53),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_008_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_089_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_17_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[18]_reg  (.CLK(net435),
    .RESET_B(net54),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_009_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_088_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_18_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[19]_reg  (.CLK(net428),
    .RESET_B(net55),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_010_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_087_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_19_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[1]_reg  (.CLK(net429),
    .RESET_B(net56),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_011_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_086_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[20]_reg  (.CLK(net429),
    .RESET_B(net57),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_012_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_085_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_20_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[21]_reg  (.CLK(net435),
    .RESET_B(net58),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_013_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_084_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_21_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[22]_reg  (.CLK(net435),
    .RESET_B(net59),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_014_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_083_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_22_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[23]_reg  (.CLK(net428),
    .RESET_B(net60),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_015_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_082_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_23_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[24]_reg  (.CLK(net428),
    .RESET_B(net61),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_016_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_081_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_24_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[25]_reg  (.CLK(net435),
    .RESET_B(net62),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_017_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_080_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_25_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[26]_reg  (.CLK(net429),
    .RESET_B(net63),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_018_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_079_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_26_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[27]_reg  (.CLK(net436),
    .RESET_B(net64),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_019_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_078_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_27_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[28]_reg  (.CLK(net436),
    .RESET_B(net65),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_020_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_077_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_28_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[29]_reg  (.CLK(net437),
    .RESET_B(net66),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_021_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_076_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_29_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[2]_reg  (.CLK(net429),
    .RESET_B(net67),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_022_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_075_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_2_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[30]_reg  (.CLK(net427),
    .RESET_B(net68),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_023_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_074_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_30_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[31]_reg  (.CLK(net430),
    .RESET_B(net69),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_024_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_073_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_31_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[32]_reg  (.CLK(net435),
    .RESET_B(net70),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_025_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_072_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_32_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[33]_reg  (.CLK(net437),
    .RESET_B(net71),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_026_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_071_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_33_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[34]_reg  (.CLK(net429),
    .RESET_B(net72),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_027_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_070_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_34_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[35]_reg  (.CLK(net428),
    .RESET_B(net73),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_028_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_069_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_35_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[36]_reg  (.CLK(net435),
    .RESET_B(net74),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_029_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_068_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_36_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[37]_reg  (.CLK(net430),
    .RESET_B(net75),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_030_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_067_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_37_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[38]_reg  (.CLK(net430),
    .RESET_B(net76),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_031_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_066_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_38_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[39]_reg  (.CLK(net436),
    .RESET_B(net77),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_032_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_065_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_39_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[3]_reg  (.CLK(net435),
    .RESET_B(net78),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_033_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_064_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_3_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[40]_reg  (.CLK(net436),
    .RESET_B(net79),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_034_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_063_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_40_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[4]_reg  (.CLK(net428),
    .RESET_B(net80),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_035_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_062_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_4_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[5]_reg  (.CLK(net429),
    .RESET_B(net81),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_036_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_061_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_5_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[6]_reg  (.CLK(net436),
    .RESET_B(net82),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_037_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_060_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_6_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[7]_reg  (.CLK(net437),
    .RESET_B(net83),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_038_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_059_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_7_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[8]_reg  (.CLK(net430),
    .RESET_B(net84),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_039_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_058_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_8_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_data_o[9]_reg  (.CLK(net428),
    .RESET_B(net85),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_040_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/_057_ ),
    .Q(\i_dmi_cdc.i_cdc_req/async_data_9_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/async_req_o_reg  (.CLK(net431),
    .RESET_B(net376),
    .D(\i_dmi_cdc.i_cdc_req/i_src/_041_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/req_src_d_$_MUX__Y_A ),
    .Q(\i_dmi_cdc.i_cdc_req/async_req ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_0__reg  (.CLK(net432),
    .RESET_B(net378),
    .D(\i_dmi_cdc.i_cdc_req/async_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_1__reg  (.CLK(net432),
    .RESET_B(net378),
    .D(\i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/i_sync/_2_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/i_src/i_sync/serial_o_reg  (.CLK(net432),
    .RESET_B(net377),
    .D(\i_dmi_cdc.i_cdc_req/i_src/i_sync/reg_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_req/i_src/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_req/i_src/ack_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/s_dst_clear_ack_q_reg  (.CLK(clknet_5_27__leaf_clk_i),
    .RESET_B(net385),
    .D(\i_dmi_cdc.i_cdc_req/s_dst_clear_req ),
    .Q_N(\i_dmi_cdc.i_cdc_req/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_req/s_dst_clear_ack_q ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q_reg  (.RESET_B(net384),
    .D(\i_dmi_cdc.core_clear_pending ),
    .Q(\i_dmi_cdc.i_cdc_req/s_dst_isolate_ack_q ),
    .Q_N(\i_dmi_cdc.i_cdc_req/_2_ ),
    .CLK(clknet_5_25__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_req/s_src_clear_ack_q_reg  (.CLK(net433),
    .RESET_B(net375),
    .D(\i_dmi_cdc.i_cdc_req/s_src_clear_req ),
    .Q_N(\i_dmi_cdc.i_cdc_req/_3_ ),
    .Q(\i_dmi_cdc.i_cdc_req/s_src_clear_ack_q ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q_reg  (.RESET_B(net379),
    .D(\i_dmi_cdc.i_cdc_req/src_clear_pending_o ),
    .Q(\i_dmi_cdc.i_cdc_req/s_src_isolate_ack_q ),
    .Q_N(\i_dmi_cdc.i_cdc_req/_0_ ),
    .CLK(net433));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/_4_  (.A(\i_dmi_cdc.i_cdc_resp/dst_clear_pending_o ),
    .B_N(net3),
    .Y(\i_dmi_cdc.i_cdc_resp/i_dst_ready_i ));
 sg13g2_nor2b_2 \i_dmi_cdc.i_cdc_resp/_5_  (.A(\i_dmi_cdc.i_cdc_resp/dst_clear_pending_o ),
    .B_N(\i_dmi_cdc.i_cdc_resp/s_dst_valid ),
    .Y(dmi_resp_valid));
 sg13g2_nor2b_2 \i_dmi_cdc.i_cdc_resp/_6_  (.A(\i_dmi_cdc.i_cdc_resp/src_clear_pending_o ),
    .B_N(\i_dmi_cdc.i_cdc_resp/s_src_ready ),
    .Y(dmi_resp_ready_o));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/_7_  (.A(\i_dmi_cdc.i_cdc_resp/src_clear_pending_o ),
    .B_N(dmi_resp_valid_i),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src_valid_i ));
 sg13g2_buf_2 fanout177 (.A(net179),
    .X(net177));
 sg13g2_buf_2 fanout176 (.A(net177),
    .X(net176));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_074_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .A(net333));
 sg13g2_buf_4 fanout175 (.X(net175),
    .A(net177));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_076_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_077_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_078_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_079_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_080_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_081_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_020_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_082_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_022_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_021_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_083_  (.Y(\i_dmi_cdc.i_cdc_resp/s_src_clear_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_022_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_084_  (.A(net331),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_023_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_085_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ));
 sg13g2_buf_2 fanout174 (.A(tms_i),
    .X(net174));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_087_  (.B1(net334),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_026_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_023_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_088_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_027_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .A(net331));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_089_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_027_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_026_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_090_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_091_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .A2(net332),
    .A1(net331));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_092_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_026_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ),
    .A1(net332),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_093_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_029_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_094_  (.A(net332),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_095_  (.A(net331),
    .B(net330),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_032_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_096_  (.A(net333),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_097_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_033_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_031_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_032_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_098_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .A1(net330),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_030_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_099_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ),
    .A(\i_dmi_cdc.i_cdc_resp/s_src_clear_ack_q ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_100_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ),
    .A(net333));
 sg13g2_nand4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_101_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ),
    .D(net331));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_102_  (.A(net334),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_103_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_038_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_104_  (.A(net330),
    .B(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ));
 sg13g2_and4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_105_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(net333),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_106_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ),
    .C1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_041_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_037_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_107_  (.A(net331),
    .B(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_108_  (.A(net2),
    .B(net333),
    .C(net332),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_109_  (.A1(net333),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_043_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_044_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_110_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .B(net330),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_111_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_045_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_112_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_040_ ),
    .A(net333),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_113_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_034_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_048_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_114_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ),
    .B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_036_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/s_src_clear_ack_q ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_115_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_050_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_116_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_051_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_117_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_042_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_118_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(net334),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_119_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_014_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ),
    .A1(net332),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_053_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_120_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_054_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_121_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_122_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_024_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_056_ ),
    .A(net334),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_123_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_057_ ),
    .C1(net330),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_055_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_028_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_039_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_124_  (.A0(net332),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_058_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_125_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ),
    .B(net333));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_126_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ),
    .B(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ),
    .A_N(net332));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_127_  (.B1(net331),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_060_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_128_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_046_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_017_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_129_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_062_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_130_  (.A(net331),
    .B(net330),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_059_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_131_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_047_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_049_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_132_  (.A0(net330),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_063_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_064_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_133_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .A1(net330),
    .S(net334),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_134_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_065_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_135_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_066_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_136_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_137_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_138_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_019_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_069_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_139_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_140_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_141_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_070_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_007_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_142_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_032_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_068_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_008_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_143_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_009_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/src_clear_pending_o ),
    .A1(net332),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_067_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_144_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_145_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .C1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_071_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_010_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_018_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_146_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_147_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_148_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_011_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ));
 sg13g2_nand2b_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_13_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_14_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_15_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_16_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_04_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_17_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_18_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_19_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_06_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_05_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_20_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_ack ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_21_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_07_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_08_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_22_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_23_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_09_ ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_24_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_03_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_25_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_11_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_10_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_26_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_02_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/async_ack_o_reg  (.CLK(clknet_5_11__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/ack_dst_d ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_12_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_ack ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0__reg  (.CLK(clknet_5_11__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_req ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/serial_o_reg  (.CLK(clknet_5_11__leaf_clk_i),
    .RESET_B(net383),
    .D(net445),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/req_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__reg  (.CLK(clknet_5_11__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__reg  (.CLK(clknet_5_10__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/_01_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/state_q_1_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_21_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_22_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_23_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/req_src_d ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_24_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_08_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_25_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_26_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_27_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_09_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_28_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_29_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_0_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_30_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/data_src_d_1_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_31_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_ack ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_32_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_33_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_34_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_12_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_11_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_35_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_36_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_07_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_37_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_13_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_15_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_38_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_39_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_phase_transition_req ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_40_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_41_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_17_ ),
    .B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_18_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_16_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_42_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_19_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_data_o[0]_reg  (.CLK(clknet_5_14__leaf_clk_i),
    .RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_03_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_00_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_data_o[1]_reg  (.RESET_B(net388),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_04_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_20_ ),
    .CLK(clknet_5_14__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/async_req_o_reg  (.CLK(clknet_5_13__leaf_clk_i),
    .RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_02_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_req ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_01_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0__reg  (.CLK(clknet_5_13__leaf_clk_i),
    .RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/serial_o_reg  (.RESET_B(net381),
    .D(net447),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/ack_synced ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/_0_ ),
    .CLK(clknet_5_13__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__reg  (.RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_05_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .CLK(clknet_5_12__leaf_clk_i));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__reg  (.RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/_06_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .CLK(clknet_5_13__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0__reg  (.CLK(clknet_5_10__leaf_clk_i),
    .RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_000_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__reg  (.CLK(clknet_5_10__leaf_clk_i),
    .RESET_B(net382),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_002_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__reg  (.RESET_B(net382),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_003_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2__$_NOT__A_Y ),
    .CLK(clknet_5_10__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__reg  (.CLK(clknet_5_12__leaf_clk_i),
    .RESET_B(net381),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_004_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__reg  (.CLK(clknet_5_12__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__reg  (.CLK(clknet_5_12__leaf_clk_i),
    .RESET_B(net383),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_phase_q_1_ ));
 sg13g2_buf_1 fanout173 (.A(_0319_),
    .X(net173));
 sg13g2_buf_2 fanout172 (.A(_0319_),
    .X(net172));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_074_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .B(net326),
    .A(net328));
 sg13g2_buf_2 fanout171 (.A(net172),
    .X(net171));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_076_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .A(net325));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_077_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .A1(net327));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_078_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_079_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_080_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_081_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_020_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_082_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_021_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_083_  (.Y(\i_dmi_cdc.i_cdc_resp/s_dst_clear_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_022_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_084_  (.A(net326),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_085_  (.A(net327),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ));
 sg13g2_buf_2 fanout170 (.A(net172),
    .X(net170));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_087_  (.B1(net328),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_023_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_088_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A(net326));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_089_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_027_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .B1(net325),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_090_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_091_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .A2(net327),
    .A1(net326));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_092_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_026_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ),
    .A1(net327),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_093_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_029_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_094_  (.A(net327),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_095_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_096_  (.A(net328),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_097_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_033_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_031_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_098_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .A1(net325),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_030_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_099_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .A(\i_dmi_cdc.i_cdc_resp/s_dst_clear_ack_q ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_100_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A(net328));
 sg13g2_nand4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_101_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ),
    .D(net326));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_102_  (.A(net329),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_103_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_038_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_104_  (.A(net325),
    .B(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ));
 sg13g2_and4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_105_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net328),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_106_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ),
    .C1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_041_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_037_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_107_  (.A(net326),
    .B(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_108_  (.A(net221),
    .B(net329),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_109_  (.A1(net329),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_043_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_044_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_110_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_111_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_045_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_112_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_040_ ),
    .A(net328),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_113_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_034_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_048_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_114_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_036_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/s_dst_clear_ack_q ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_115_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_050_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_116_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_051_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_117_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_042_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_118_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net328),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_119_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_014_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ),
    .A1(net327),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_053_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_120_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_054_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_121_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ));
 sg13g2_nand3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_122_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_024_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_056_ ),
    .A(net328),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_123_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_057_ ),
    .C1(net325),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_055_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_028_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_039_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_124_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_058_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_125_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ),
    .B(net329));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_126_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ),
    .B(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ),
    .A_N(net327));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_127_  (.B1(net326),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_060_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_128_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_061_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_046_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_017_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_129_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_062_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_052_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ));
 sg13g2_nor4_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_130_  (.A(net326),
    .B(net325),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_059_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_131_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_047_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_049_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_132_  (.A0(net325),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_063_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_064_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_133_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .A1(net325),
    .S(net329),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_134_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_016_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_065_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_135_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_066_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_136_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_137_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_138_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_019_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_069_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_139_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ));
 sg13g2_nor3_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_140_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_141_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_070_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_007_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_142_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_032_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_068_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_008_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_143_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_009_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/dst_clear_pending_o ),
    .A1(net327),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_067_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_144_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ));
 sg13g2_a221oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_145_  (.B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .C1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_071_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_010_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_035_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_018_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_146_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_147_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_148_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_011_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ));
 sg13g2_nand2b_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_13_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_14_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_15_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_16_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_04_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_17_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_18_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_19_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_06_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_05_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_20_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_ack ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ));
 sg13g2_and2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_21_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_07_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_08_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_22_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_23_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_09_ ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_24_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_03_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_25_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_11_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_10_ ));
 sg13g2_a21oi_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_26_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_req ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_02_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/async_ack_o_reg  (.CLK(net406),
    .RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/ack_dst_d ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_12_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_ack ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0__reg  (.CLK(net398),
    .RESET_B(net347),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_req ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/serial_o_reg  (.CLK(net398),
    .RESET_B(net347),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/req_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__reg  (.CLK(net406),
    .RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__reg  (.CLK(net406),
    .RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/_01_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/state_q_1_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_21_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_22_  (.B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_23_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/req_src_d ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_24_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_08_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_25_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ));
 sg13g2_nor2_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_26_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_27_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_09_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_28_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_29_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_0_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_30_  (.A0(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_clear_seq_phase_1_ ),
    .S(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_10_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/data_src_d_1_ ));
 sg13g2_nor3_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_31_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_ack ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_32_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_33_  (.B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .C(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_34_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_12_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_11_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ));
 sg13g2_nand2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_35_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_36_  (.X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_14_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_07_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_37_  (.A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_13_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_15_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_38_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_39_  (.A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_phase_transition_req ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_40_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_41_  (.Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_17_ ),
    .B2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_18_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_16_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_42_  (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_19_ ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_data_o[0]_reg  (.RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_03_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_00_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_0_ ),
    .CLK(net406));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_data_o[1]_reg  (.RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_04_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/receiver_next_phase_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_20_ ),
    .CLK(net407));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/async_req_o_reg  (.CLK(net407),
    .RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_02_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_b2a_req ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_01_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0__reg  (.CLK(net407),
    .RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/async_a2b_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/serial_o_reg  (.RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/ack_synced ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/_0_ ),
    .CLK(net407));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__reg  (.RESET_B(net363),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_05_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_0__$_NOT__A_Y ),
    .CLK(net409));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__reg  (.RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/_06_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/state_q_1__$_NOT__A_Y ),
    .CLK(net407));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0__reg  (.CLK(net408),
    .RESET_B(net360),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_000_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__reg  (.CLK(net409),
    .RESET_B(net361),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_002_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__reg  (.RESET_B(net360),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_003_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_2__$_NOT__A_Y ),
    .CLK(net408));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__reg  (.CLK(net409),
    .RESET_B(net361),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_004_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__reg  (.CLK(net408),
    .RESET_B(net360),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__reg  (.CLK(net408),
    .RESET_B(net360),
    .D(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1__$_NOT__A_Y ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/receiver_phase_q_1_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_dst/_085_  (.A(\i_dmi_cdc.i_cdc_resp/s_dst_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d_$_MUX__Y_A ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d ));
 sg13g2_a21o_1 \i_dmi_cdc.i_cdc_resp/i_dst/_086_  (.A2(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_dst_ready_i ),
    .B1(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_035_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_dst/_087_  (.Y(\i_dmi_cdc.i_cdc_resp/i_dst/_036_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_dst_ready_i ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ));
 sg13g2_a22oi_1 \i_dmi_cdc.i_cdc_resp/i_dst/_088_  (.Y(\i_dmi_cdc.i_cdc_resp/i_dst/_037_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/i_dst/_036_ ),
    .B2(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_dst/_035_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d_$_MUX__Y_A ));
 sg13g2_nor2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_089_  (.A(\i_dmi_cdc.i_cdc_resp/s_dst_clear_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_dst/_037_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_dst/_000_ ));
 sg13g2_nand2b_1 \i_dmi_cdc.i_cdc_resp/i_dst/_090_  (.Y(\i_dmi_cdc.i_cdc_resp/i_dst/_038_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ));
 sg13g2_nand3b_1 \i_dmi_cdc.i_cdc_resp/i_dst/_091_  (.B(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ),
    .C(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_dst/_039_ ),
    .A_N(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_dst/_092_  (.B1(\i_dmi_cdc.i_cdc_resp/i_dst/_039_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_dst/_040_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_dst/_038_ ));
 sg13g2_buf_2 fanout169 (.A(net172),
    .X(net169));
 sg13g2_buf_2 fanout168 (.A(net172),
    .X(net168));
 sg13g2_buf_2 fanout167 (.A(net172),
    .X(net167));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_096_  (.A0(dmi_resp_0_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_0_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_097_  (.A0(dmi_resp_10_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_10_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_098_  (.A0(dmi_resp_11_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_11_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_11_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_099_  (.A0(dmi_resp_12_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_12_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_12_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_100_  (.A0(dmi_resp_13_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_13_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_13_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_101_  (.A0(dmi_resp_14_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_14_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_14_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_102_  (.A0(dmi_resp_15_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_15_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_15_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_103_  (.A0(dmi_resp_16_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_16_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_16_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_104_  (.A0(dmi_resp_17_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_17_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_17_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_105_  (.A0(dmi_resp_18_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_18_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_18_ ));
 sg13g2_buf_1 fanout166 (.A(_0287_),
    .X(net166));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_107_  (.A0(dmi_resp_19_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_19_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_19_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_108_  (.A0(net324),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_1_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_1_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_109_  (.A0(dmi_resp_20_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_20_ ),
    .S(net288),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_20_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_110_  (.A0(dmi_resp_21_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_21_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_21_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_111_  (.A0(dmi_resp_22_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_22_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_22_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_112_  (.A0(dmi_resp_23_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_23_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_23_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_113_  (.A0(dmi_resp_24_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_24_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_24_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_114_  (.A0(dmi_resp_25_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_25_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_25_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_115_  (.A0(dmi_resp_26_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_26_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_26_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_116_  (.A0(dmi_resp_27_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_27_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_27_ ));
 sg13g2_buf_2 fanout165 (.A(_0287_),
    .X(net165));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_118_  (.A0(dmi_resp_28_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_28_ ),
    .S(net281),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_28_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_119_  (.A0(dmi_resp_29_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_29_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_29_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_120_  (.A0(dmi_resp_2_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_2_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_2_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_121_  (.A0(dmi_resp_30_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_30_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_30_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_122_  (.A0(dmi_resp_31_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_31_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_31_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_123_  (.A0(dmi_resp_32_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_32_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_32_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_124_  (.A0(dmi_resp_33_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_33_ ),
    .S(net281),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_33_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_125_  (.A0(dmi_resp_3_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_3_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_3_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_126_  (.A0(dmi_resp_4_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_4_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_4_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_127_  (.A0(dmi_resp_5_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_5_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_5_ ));
 sg13g2_buf_2 fanout164 (.A(net165),
    .X(net164));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_129_  (.A0(dmi_resp_6_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_6_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_6_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_130_  (.A0(dmi_resp_7_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_7_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_7_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_131_  (.A0(dmi_resp_8_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_8_ ),
    .S(net288),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_8_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_132_  (.A0(dmi_resp_9_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_9_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/data_dst_d_9_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_133_  (.A0(dmi_resp_0_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_0_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_001_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_134_  (.A0(dmi_resp_10_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_10_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_002_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_135_  (.A0(dmi_resp_11_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_11_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_003_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_136_  (.A0(dmi_resp_12_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_12_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_137_  (.A0(dmi_resp_13_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_13_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_138_  (.A0(dmi_resp_14_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_14_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_006_ ));
 sg13g2_buf_2 fanout163 (.A(net165),
    .X(net163));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_140_  (.A0(dmi_resp_15_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_15_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_007_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_141_  (.A0(dmi_resp_16_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_16_ ),
    .S(net281),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_008_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_142_  (.A0(dmi_resp_17_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_17_ ),
    .S(net288),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_009_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_143_  (.A0(dmi_resp_18_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_18_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_010_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_144_  (.A0(dmi_resp_19_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_19_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_011_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_145_  (.A0(net324),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_1_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_012_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_146_  (.A0(dmi_resp_20_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_20_ ),
    .S(net288),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_013_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_147_  (.A0(dmi_resp_21_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_21_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_014_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_148_  (.A0(dmi_resp_22_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_22_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_015_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_149_  (.A0(dmi_resp_23_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_23_ ),
    .S(net282),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_016_ ));
 sg13g2_buf_2 fanout162 (.A(net166),
    .X(net162));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_151_  (.A0(dmi_resp_24_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_24_ ),
    .S(net283),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_017_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_152_  (.A0(dmi_resp_25_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_25_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_018_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_153_  (.A0(dmi_resp_26_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_26_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_019_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_154_  (.A0(dmi_resp_27_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_27_ ),
    .S(net283),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_020_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_155_  (.A0(dmi_resp_28_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_28_ ),
    .S(net281),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_021_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_156_  (.A0(dmi_resp_29_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_29_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_022_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_157_  (.A0(dmi_resp_2_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_2_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_023_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_158_  (.A0(dmi_resp_30_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_30_ ),
    .S(net284),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_024_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_159_  (.A0(dmi_resp_31_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_31_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_025_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_160_  (.A0(dmi_resp_32_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_32_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_026_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_161_  (.A0(dmi_resp_33_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_33_ ),
    .S(net280),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_027_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_162_  (.A0(dmi_resp_3_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_3_ ),
    .S(net285),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_028_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_163_  (.A0(dmi_resp_4_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_4_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_029_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_164_  (.A0(dmi_resp_5_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_5_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_030_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_165_  (.A0(dmi_resp_6_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_6_ ),
    .S(net279),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_031_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_166_  (.A0(dmi_resp_7_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_7_ ),
    .S(net278),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_032_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_167_  (.A0(dmi_resp_8_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_8_ ),
    .S(net287),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_033_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_168_  (.A0(dmi_resp_9_),
    .A1(\i_dmi_cdc.i_cdc_resp/async_data_9_ ),
    .S(net286),
    .X(\i_dmi_cdc.i_cdc_resp/i_dst/_034_ ));
 sg13g2_xor2_1 \i_dmi_cdc.i_cdc_resp/i_dst/_169_  (.B(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ),
    .A(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .X(\i_dmi_cdc.i_cdc_resp/s_dst_valid ));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[0]_reg_120  (.L_HI(net120));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/async_ack_o_reg  (.RESET_B(net349),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_000_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/ack_dst_d_$_MUX__Y_A ),
    .CLK(net406));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[0]_reg  (.RESET_B(net86),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_001_ ),
    .Q(dmi_resp_0_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_082_ ),
    .CLK(net393));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[10]_reg  (.RESET_B(net87),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_002_ ),
    .Q(dmi_resp_10_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_081_ ),
    .CLK(net389));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[11]_reg  (.RESET_B(net88),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_003_ ),
    .Q(dmi_resp_11_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_080_ ),
    .CLK(net392));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[12]_reg  (.RESET_B(net89),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_004_ ),
    .Q(dmi_resp_12_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_079_ ),
    .CLK(net393));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[13]_reg  (.RESET_B(net90),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_005_ ),
    .Q(dmi_resp_13_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_078_ ),
    .CLK(net392));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[14]_reg  (.RESET_B(net91),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_006_ ),
    .Q(dmi_resp_14_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_077_ ),
    .CLK(net394));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[15]_reg  (.RESET_B(net92),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_007_ ),
    .Q(dmi_resp_15_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_076_ ),
    .CLK(net394));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[16]_reg  (.CLK(net393),
    .RESET_B(net93),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_008_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_075_ ),
    .Q(dmi_resp_16_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[17]_reg  (.CLK(net394),
    .RESET_B(net94),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_009_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_074_ ),
    .Q(dmi_resp_17_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[18]_reg  (.CLK(net389),
    .RESET_B(net95),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_010_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_073_ ),
    .Q(dmi_resp_18_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[19]_reg  (.RESET_B(net96),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_011_ ),
    .Q(dmi_resp_19_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_072_ ),
    .CLK(net390));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[1]_reg  (.CLK(net392),
    .RESET_B(net97),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_012_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_071_ ),
    .Q(dmi_resp_1_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[20]_reg  (.CLK(net394),
    .RESET_B(net98),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_013_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_070_ ),
    .Q(dmi_resp_20_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[21]_reg  (.CLK(net390),
    .RESET_B(net99),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_014_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_069_ ),
    .Q(dmi_resp_21_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[22]_reg  (.RESET_B(net100),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_015_ ),
    .Q(dmi_resp_22_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_068_ ),
    .CLK(net390));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[23]_reg  (.CLK(net393),
    .RESET_B(net101),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_016_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_067_ ),
    .Q(dmi_resp_23_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[24]_reg  (.RESET_B(net102),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_017_ ),
    .Q(dmi_resp_24_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_066_ ),
    .CLK(net393));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[25]_reg  (.RESET_B(net103),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_018_ ),
    .Q(dmi_resp_25_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_065_ ),
    .CLK(net392));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[26]_reg  (.RESET_B(net104),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_019_ ),
    .Q(dmi_resp_26_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_064_ ),
    .CLK(net389));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[27]_reg  (.CLK(net395),
    .RESET_B(net105),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_020_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_063_ ),
    .Q(dmi_resp_27_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[28]_reg  (.RESET_B(net106),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_021_ ),
    .Q(dmi_resp_28_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_062_ ),
    .CLK(net393));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[29]_reg  (.CLK(net394),
    .RESET_B(net107),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_022_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_061_ ),
    .Q(dmi_resp_29_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[2]_reg  (.RESET_B(net108),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_023_ ),
    .Q(dmi_resp_2_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_060_ ),
    .CLK(net389));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[30]_reg  (.CLK(net390),
    .RESET_B(net109),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_024_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_059_ ),
    .Q(dmi_resp_30_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[31]_reg  (.CLK(net393),
    .RESET_B(net110),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_025_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_058_ ),
    .Q(dmi_resp_31_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[32]_reg  (.RESET_B(net111),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_026_ ),
    .Q(dmi_resp_32_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_057_ ),
    .CLK(net392));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[33]_reg  (.RESET_B(net112),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_027_ ),
    .Q(dmi_resp_33_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_056_ ),
    .CLK(net393));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[3]_reg  (.CLK(net389),
    .RESET_B(net113),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_028_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_055_ ),
    .Q(dmi_resp_3_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[4]_reg  (.CLK(net394),
    .RESET_B(net114),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_029_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_054_ ),
    .Q(dmi_resp_4_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[5]_reg  (.CLK(net392),
    .RESET_B(net115),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_030_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_053_ ),
    .Q(dmi_resp_5_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[6]_reg  (.CLK(net392),
    .RESET_B(net116),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_031_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_052_ ),
    .Q(dmi_resp_6_));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[7]_reg  (.RESET_B(net117),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_032_ ),
    .Q(dmi_resp_7_),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_051_ ),
    .CLK(net392));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[8]_reg  (.CLK(net394),
    .RESET_B(net118),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_033_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_050_ ),
    .Q(dmi_resp_8_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/data_o[9]_reg  (.CLK(net390),
    .RESET_B(net119),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/_034_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_083_ ),
    .Q(dmi_resp_9_));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_0__reg  (.CLK(net394),
    .RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/async_req ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_1__reg  (.CLK(net395),
    .RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_0_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_2_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_dst/i_sync/serial_o_reg  (.CLK(net395),
    .RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/reg_q_1_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1_reg  (.RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_dst/req_synced_q1 ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_dst/_049_ ),
    .CLK(net406));
 sg13g2_xnor2_1 \i_dmi_cdc.i_cdc_resp/i_src/_084_  (.Y(\i_dmi_cdc.i_cdc_resp/s_src_ready ),
    .A(\i_dmi_cdc.i_cdc_resp/async_req ),
    .B(\i_dmi_cdc.i_cdc_resp/i_src/ack_synced ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_src/_085_  (.A(\i_dmi_cdc.i_cdc_resp/s_src_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_src_valid_i ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src/_035_ ));
 sg13g2_and2_2 \i_dmi_cdc.i_cdc_resp/i_src/_086_  (.A(\i_dmi_cdc.i_cdc_resp/s_src_ready ),
    .B(\i_dmi_cdc.i_cdc_resp/i_src/_035_ ),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_036_ ));
 sg13g2_buf_2 fanout161 (.A(net166),
    .X(net161));
 sg13g2_buf_2 fanout160 (.A(net166),
    .X(net160));
 sg13g2_buf_2 fanout159 (.A(net165),
    .X(net159));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_090_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_0_ ),
    .A1(dmi_resp_i_0_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_000_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_091_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_10_ ),
    .A1(dmi_resp_i_10_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_001_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_092_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_11_ ),
    .A1(dmi_resp_i_11_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_002_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_093_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_12_ ),
    .A1(dmi_resp_i_12_),
    .S(net204),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_003_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_094_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_13_ ),
    .A1(dmi_resp_i_13_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_004_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_095_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_14_ ),
    .A1(dmi_resp_i_14_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_005_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_096_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_15_ ),
    .A1(dmi_resp_i_15_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_006_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_097_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_16_ ),
    .A1(dmi_resp_i_16_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_007_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_098_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_17_ ),
    .A1(dmi_resp_i_17_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_008_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_099_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_18_ ),
    .A1(dmi_resp_i_18_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_009_ ));
 sg13g2_buf_2 fanout158 (.A(net165),
    .X(net158));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_101_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_19_ ),
    .A1(dmi_resp_i_19_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_010_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_102_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_1_ ),
    .A1(dmi_resp_i_1_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_011_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_103_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_20_ ),
    .A1(dmi_resp_i_20_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_012_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_104_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_21_ ),
    .A1(dmi_resp_i_21_),
    .S(net206),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_013_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_105_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_22_ ),
    .A1(dmi_resp_i_22_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_014_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_106_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_23_ ),
    .A1(dmi_resp_i_23_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_015_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_107_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_24_ ),
    .A1(dmi_resp_i_24_),
    .S(net204),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_016_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_108_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_25_ ),
    .A1(dmi_resp_i_25_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_017_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_109_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_26_ ),
    .A1(dmi_resp_i_26_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_018_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_110_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_27_ ),
    .A1(dmi_resp_i_27_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_019_ ));
 sg13g2_buf_4 fanout157 (.X(net157),
    .A(net165));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_112_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_28_ ),
    .A1(dmi_resp_i_28_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_020_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_113_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_29_ ),
    .A1(dmi_resp_i_29_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_021_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_114_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_2_ ),
    .A1(dmi_resp_i_2_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_022_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_115_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_30_ ),
    .A1(dmi_resp_i_30_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_023_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_116_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_31_ ),
    .A1(dmi_resp_i_31_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_024_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_117_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_32_ ),
    .A1(dmi_resp_i_32_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_025_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_118_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_33_ ),
    .A1(dmi_resp_i_33_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_026_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_119_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_3_ ),
    .A1(dmi_resp_i_3_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_027_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_120_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_4_ ),
    .A1(dmi_resp_i_4_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_028_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_121_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_5_ ),
    .A1(dmi_resp_i_5_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_029_ ));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(net165));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_123_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_6_ ),
    .A1(dmi_resp_i_6_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_030_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_124_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_7_ ),
    .A1(dmi_resp_i_7_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_031_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_125_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_8_ ),
    .A1(dmi_resp_i_8_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_032_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_126_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_9_ ),
    .A1(dmi_resp_i_9_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/_033_ ));
 sg13g2_nor2b_1 \i_dmi_cdc.i_cdc_resp/i_src/_127_  (.A(\i_dmi_cdc.i_cdc_resp/s_src_clear_req ),
    .B_N(\i_dmi_cdc.i_cdc_resp/i_src/req_src_d_$_MUX__Y_A ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src/req_src_d ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_src/_128_  (.A1(\i_dmi_cdc.i_cdc_resp/i_src/req_src_d_$_MUX__Y_A ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_src_valid_i ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src/_043_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/async_req ));
 sg13g2_or2_1 \i_dmi_cdc.i_cdc_resp/i_src/_129_  (.X(\i_dmi_cdc.i_cdc_resp/i_src/_044_ ),
    .B(\i_dmi_cdc.i_cdc_resp/i_src/_043_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_src/ack_synced ));
 sg13g2_inv_1 \i_dmi_cdc.i_cdc_resp/i_src/_130_  (.Y(\i_dmi_cdc.i_cdc_resp/i_src/_045_ ),
    .A(\i_dmi_cdc.i_cdc_resp/i_src_valid_i ));
 sg13g2_o21ai_1 \i_dmi_cdc.i_cdc_resp/i_src/_131_  (.B1(\i_dmi_cdc.i_cdc_resp/async_req ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src/_046_ ),
    .A1(\i_dmi_cdc.i_cdc_resp/i_src/req_src_d_$_MUX__Y_A ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_src/_045_ ));
 sg13g2_a21oi_1 \i_dmi_cdc.i_cdc_resp/i_src/_132_  (.A1(\i_dmi_cdc.i_cdc_resp/i_src/_044_ ),
    .A2(\i_dmi_cdc.i_cdc_resp/i_src/_046_ ),
    .Y(\i_dmi_cdc.i_cdc_resp/i_src/_034_ ),
    .B1(\i_dmi_cdc.i_cdc_resp/s_src_clear_req ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_133_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_0_ ),
    .A1(dmi_resp_i_0_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_0_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_134_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_10_ ),
    .A1(dmi_resp_i_10_),
    .S(net206),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_10_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_135_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_11_ ),
    .A1(dmi_resp_i_11_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_11_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_136_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_12_ ),
    .A1(dmi_resp_i_12_),
    .S(net204),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_12_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_137_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_13_ ),
    .A1(dmi_resp_i_13_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_13_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_138_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_14_ ),
    .A1(dmi_resp_i_14_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_14_ ));
 sg13g2_buf_2 fanout155 (.A(net165),
    .X(net155));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_140_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_15_ ),
    .A1(dmi_resp_i_15_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_15_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_141_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_16_ ),
    .A1(dmi_resp_i_16_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_16_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_142_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_17_ ),
    .A1(dmi_resp_i_17_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_17_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_143_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_18_ ),
    .A1(dmi_resp_i_18_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_18_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_144_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_19_ ),
    .A1(dmi_resp_i_19_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_19_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_145_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_1_ ),
    .A1(dmi_resp_i_1_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_1_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_146_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_20_ ),
    .A1(dmi_resp_i_20_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_20_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_147_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_21_ ),
    .A1(dmi_resp_i_21_),
    .S(net206),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_21_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_148_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_22_ ),
    .A1(dmi_resp_i_22_),
    .S(net206),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_22_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_149_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_23_ ),
    .A1(dmi_resp_i_23_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_23_ ));
 sg13g2_buf_2 fanout154 (.A(net165),
    .X(net154));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_151_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_24_ ),
    .A1(dmi_resp_i_24_),
    .S(net204),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_24_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_152_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_25_ ),
    .A1(dmi_resp_i_25_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_25_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_153_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_26_ ),
    .A1(dmi_resp_i_26_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_26_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_154_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_27_ ),
    .A1(dmi_resp_i_27_),
    .S(net207),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_27_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_155_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_28_ ),
    .A1(dmi_resp_i_28_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_28_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_156_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_29_ ),
    .A1(dmi_resp_i_29_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_29_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_157_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_2_ ),
    .A1(dmi_resp_i_2_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_2_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_158_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_30_ ),
    .A1(dmi_resp_i_30_),
    .S(net205),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_30_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_159_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_31_ ),
    .A1(dmi_resp_i_31_),
    .S(net202),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_31_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_160_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_32_ ),
    .A1(dmi_resp_i_32_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_32_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_161_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_33_ ),
    .A1(dmi_resp_i_33_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_33_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_162_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_3_ ),
    .A1(dmi_resp_i_3_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_3_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_163_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_4_ ),
    .A1(dmi_resp_i_4_),
    .S(net203),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_4_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_164_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_5_ ),
    .A1(dmi_resp_i_5_),
    .S(net201),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_5_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_165_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_6_ ),
    .A1(dmi_resp_i_6_),
    .S(net200),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_6_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_166_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_7_ ),
    .A1(dmi_resp_i_7_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_7_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_167_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_8_ ),
    .A1(dmi_resp_i_8_),
    .S(net208),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_8_ ));
 sg13g2_mux2_1 \i_dmi_cdc.i_cdc_resp/i_src/_168_  (.A0(\i_dmi_cdc.i_cdc_resp/async_data_9_ ),
    .A1(dmi_resp_i_9_),
    .S(net199),
    .X(\i_dmi_cdc.i_cdc_resp/i_src/data_src_d_9_ ));
 sg13g2_buf_2 fanout283 (.A(net289),
    .X(net283));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[0]_reg  (.CLK(clknet_5_1__leaf_clk_i),
    .RESET_B(net120),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_000_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_082_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[10]_reg  (.CLK(clknet_5_5__leaf_clk_i),
    .RESET_B(net121),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_001_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_081_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_10_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[11]_reg  (.CLK(clknet_5_0__leaf_clk_i),
    .RESET_B(net122),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_002_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_080_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_11_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[12]_reg  (.CLK(clknet_5_3__leaf_clk_i),
    .RESET_B(net123),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_003_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_079_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_12_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[13]_reg  (.CLK(clknet_5_4__leaf_clk_i),
    .RESET_B(net124),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_004_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_078_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_13_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[14]_reg  (.CLK(clknet_5_0__leaf_clk_i),
    .RESET_B(net125),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_005_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_077_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_14_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[15]_reg  (.CLK(clknet_5_6__leaf_clk_i),
    .RESET_B(net126),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_006_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_076_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_15_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[16]_reg  (.CLK(clknet_5_2__leaf_clk_i),
    .RESET_B(net127),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_007_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_075_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_16_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[17]_reg  (.CLK(clknet_5_8__leaf_clk_i),
    .RESET_B(net128),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_008_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_074_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_17_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[18]_reg  (.CLK(clknet_5_7__leaf_clk_i),
    .RESET_B(net129),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_009_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_073_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_18_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[19]_reg  (.CLK(clknet_5_1__leaf_clk_i),
    .RESET_B(net130),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_010_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_072_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_19_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[1]_reg  (.CLK(clknet_5_1__leaf_clk_i),
    .RESET_B(net131),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_011_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_071_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[20]_reg  (.CLK(clknet_5_8__leaf_clk_i),
    .RESET_B(net132),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_012_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_070_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_20_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[21]_reg  (.CLK(clknet_5_7__leaf_clk_i),
    .RESET_B(net133),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_013_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_069_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_21_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[22]_reg  (.CLK(clknet_5_5__leaf_clk_i),
    .RESET_B(net134),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_014_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_068_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_22_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[23]_reg  (.CLK(clknet_5_6__leaf_clk_i),
    .RESET_B(net135),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_015_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_067_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_23_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[24]_reg  (.CLK(clknet_5_3__leaf_clk_i),
    .RESET_B(net136),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_016_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_066_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_24_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[25]_reg  (.CLK(clknet_5_5__leaf_clk_i),
    .RESET_B(net137),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_017_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_065_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_25_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[26]_reg  (.CLK(clknet_5_6__leaf_clk_i),
    .RESET_B(net138),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_018_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_064_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_26_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[27]_reg  (.CLK(clknet_5_3__leaf_clk_i),
    .RESET_B(net139),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_019_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_063_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_27_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[28]_reg  (.CLK(clknet_5_2__leaf_clk_i),
    .RESET_B(net140),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_020_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_062_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_28_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[29]_reg  (.CLK(clknet_5_7__leaf_clk_i),
    .RESET_B(net141),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_021_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_061_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_29_ ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[2]_reg  (.RESET_B(net142),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_022_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_2_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_060_ ),
    .CLK(clknet_5_4__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[30]_reg  (.CLK(clknet_5_5__leaf_clk_i),
    .RESET_B(net143),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_023_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_059_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_30_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[31]_reg  (.CLK(clknet_5_3__leaf_clk_i),
    .RESET_B(net144),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_024_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_058_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_31_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[32]_reg  (.CLK(clknet_5_0__leaf_clk_i),
    .RESET_B(net145),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_025_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_057_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_32_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[33]_reg  (.CLK(clknet_5_2__leaf_clk_i),
    .RESET_B(net146),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_026_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_056_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_33_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[3]_reg  (.CLK(clknet_5_7__leaf_clk_i),
    .RESET_B(net147),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_027_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_055_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_3_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[4]_reg  (.CLK(clknet_5_2__leaf_clk_i),
    .RESET_B(net148),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_028_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_054_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_4_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[5]_reg  (.CLK(clknet_5_1__leaf_clk_i),
    .RESET_B(net149),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_029_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_053_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_5_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[6]_reg  (.CLK(clknet_5_0__leaf_clk_i),
    .RESET_B(net150),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_030_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_052_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_6_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[7]_reg  (.CLK(clknet_5_4__leaf_clk_i),
    .RESET_B(net151),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_031_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_051_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_7_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[8]_reg  (.CLK(clknet_5_6__leaf_clk_i),
    .RESET_B(net152),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_032_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_050_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_8_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[9]_reg  (.CLK(clknet_5_4__leaf_clk_i),
    .RESET_B(net153),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_033_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/_049_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_data_9_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/async_req_o_reg  (.CLK(clknet_5_9__leaf_clk_i),
    .RESET_B(net382),
    .D(\i_dmi_cdc.i_cdc_resp/i_src/_034_ ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/req_src_d_$_MUX__Y_A ),
    .Q(\i_dmi_cdc.i_cdc_resp/async_req ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_0__reg  (.CLK(clknet_5_8__leaf_clk_i),
    .RESET_B(net382),
    .D(\i_dmi_cdc.i_cdc_resp/async_ack ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_1__reg  (.CLK(clknet_5_8__leaf_clk_i),
    .RESET_B(net382),
    .D(net443),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/_2_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/i_src/i_sync/serial_o_reg  (.CLK(clknet_5_9__leaf_clk_i),
    .RESET_B(net382),
    .D(net444),
    .Q_N(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/_0_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/i_src/ack_synced ));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/s_dst_clear_ack_q_reg  (.CLK(net406),
    .RESET_B(net350),
    .D(\i_dmi_cdc.i_cdc_resp/s_dst_clear_req ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/_1_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/s_dst_clear_ack_q ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q_reg  (.RESET_B(net360),
    .D(\i_dmi_cdc.i_cdc_resp/dst_clear_pending_o ),
    .Q(\i_dmi_cdc.i_cdc_resp/s_dst_isolate_ack_q ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/_2_ ),
    .CLK(net408));
 sg13g2_dfrbp_1 \i_dmi_cdc.i_cdc_resp/s_src_clear_ack_q_reg  (.CLK(clknet_5_9__leaf_clk_i),
    .RESET_B(net382),
    .D(\i_dmi_cdc.i_cdc_resp/s_src_clear_req ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/_3_ ),
    .Q(\i_dmi_cdc.i_cdc_resp/s_src_clear_ack_q ));
 sg13g2_dfrbp_2 \i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q_reg  (.RESET_B(net388),
    .D(\i_dmi_cdc.i_cdc_resp/src_clear_pending_o ),
    .Q(\i_dmi_cdc.i_cdc_resp/s_src_isolate_ack_q ),
    .Q_N(\i_dmi_cdc.i_cdc_resp/_0_ ),
    .CLK(clknet_5_9__leaf_clk_i));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.bypass_q_reg  (.CLK(net404),
    .RESET_B(net353),
    .D(\i_dmi_jtag_tap.bypass_d ),
    .Q_N(_0871_),
    .Q(\i_dmi_jtag_tap.bypass_q ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.dmi_tdo_i_reg  (.CLK(net405),
    .RESET_B(net361),
    .D(dr_d_0_),
    .Q_N(\state_d_1__$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_AND__Y_A_$_OR__Y_A ),
    .Q(dmi_0_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.dtmcs_tdo_i_reg  (.CLK(net405),
    .RESET_B(net359),
    .D(dtmcs_d_0_),
    .Q_N(_0761_),
    .Q(dtmcs_q_0_));
 sg13g2_mux2_1 \i_dmi_jtag_tap.i_dft_tck_mux/i_mux  (.A0(\i_dmi_jtag_tap.tck_ni ),
    .A1(net409),
    .S(testmode_i),
    .X(\i_dmi_jtag_tap.tck_n ));
 sg13g2_inv_1 \i_dmi_jtag_tap.i_tck_inv/i_inv  (.Y(\i_dmi_jtag_tap.tck_ni ),
    .A(net410));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_0__reg  (.CLK(net401),
    .RESET_B(net354),
    .D(_0013_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_0_ ),
    .Q(_0002_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_10__reg  (.CLK(net396),
    .RESET_B(net346),
    .D(_0014_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_10_ ),
    .Q(_0003_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_11__reg  (.CLK(net396),
    .RESET_B(net345),
    .D(_0015_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_11_ ),
    .Q(_0004_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_12__reg  (.CLK(net396),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_12_ ),
    .Q_N(_0872_),
    .Q(\i_dmi_jtag_tap.idcode_q_12_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_13__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_13_ ),
    .Q_N(_0873_),
    .Q(\i_dmi_jtag_tap.idcode_q_13_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_14__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_14_ ),
    .Q_N(_0874_),
    .Q(\i_dmi_jtag_tap.idcode_q_14_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_15__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_15_ ),
    .Q_N(_0875_),
    .Q(\i_dmi_jtag_tap.idcode_q_15_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_16__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_16_ ),
    .Q_N(_0876_),
    .Q(\i_dmi_jtag_tap.idcode_q_16_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_17__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_17_ ),
    .Q_N(_0877_),
    .Q(\i_dmi_jtag_tap.idcode_q_17_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_18__reg  (.CLK(net391),
    .RESET_B(net345),
    .D(\i_dmi_jtag_tap.idcode_d_18_ ),
    .Q_N(_0878_),
    .Q(\i_dmi_jtag_tap.idcode_q_18_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_19__reg  (.CLK(net391),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_19_ ),
    .Q_N(_0760_),
    .Q(\i_dmi_jtag_tap.idcode_q_19_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_1__reg  (.CLK(net401),
    .RESET_B(net352),
    .D(_0016_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_1_ ),
    .Q(_0005_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_20__reg  (.CLK(net389),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_20_ ),
    .Q_N(_0879_),
    .Q(\i_dmi_jtag_tap.idcode_q_20_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_21__reg  (.CLK(net398),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_21_ ),
    .Q_N(_0880_),
    .Q(\i_dmi_jtag_tap.idcode_q_21_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_22__reg  (.CLK(net389),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_22_ ),
    .Q_N(_0881_),
    .Q(\i_dmi_jtag_tap.idcode_q_22_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_23__reg  (.CLK(net389),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_23_ ),
    .Q_N(_0882_),
    .Q(\i_dmi_jtag_tap.idcode_q_23_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_24__reg  (.CLK(net398),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_24_ ),
    .Q_N(_0883_),
    .Q(\i_dmi_jtag_tap.idcode_q_24_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_25__reg  (.CLK(net398),
    .RESET_B(net347),
    .D(\i_dmi_jtag_tap.idcode_d_25_ ),
    .Q_N(_0884_),
    .Q(\i_dmi_jtag_tap.idcode_q_25_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_26__reg  (.CLK(net396),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_26_ ),
    .Q_N(_0885_),
    .Q(\i_dmi_jtag_tap.idcode_q_26_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_27__reg  (.CLK(net396),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_27_ ),
    .Q_N(_0886_),
    .Q(\i_dmi_jtag_tap.idcode_q_27_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_28__reg  (.CLK(net396),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_28_ ),
    .Q_N(_0887_),
    .Q(\i_dmi_jtag_tap.idcode_q_28_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_29__reg  (.CLK(net397),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_29_ ),
    .Q_N(_0888_),
    .Q(\i_dmi_jtag_tap.idcode_q_29_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_2__reg  (.CLK(net397),
    .RESET_B(net352),
    .D(\i_dmi_jtag_tap.idcode_d_2_ ),
    .Q_N(_0889_),
    .Q(\i_dmi_jtag_tap.idcode_q_2_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_30__reg  (.CLK(net397),
    .RESET_B(net346),
    .D(\i_dmi_jtag_tap.idcode_d_30_ ),
    .Q_N(_0890_),
    .Q(\i_dmi_jtag_tap.idcode_q_30_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_31__reg  (.CLK(net398),
    .RESET_B(net348),
    .D(\i_dmi_jtag_tap.idcode_d_31_ ),
    .Q_N(_0891_),
    .Q(\i_dmi_jtag_tap.idcode_q_31_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_3__reg  (.CLK(net397),
    .RESET_B(net352),
    .D(\i_dmi_jtag_tap.idcode_d_3_ ),
    .Q_N(_0759_),
    .Q(\i_dmi_jtag_tap.idcode_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_4__reg  (.CLK(net400),
    .RESET_B(net352),
    .D(_0017_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_4_ ),
    .Q(_0006_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_5__reg  (.CLK(net397),
    .RESET_B(net352),
    .D(_0018_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_5_ ),
    .Q(_0007_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_6__reg  (.CLK(net397),
    .RESET_B(net352),
    .D(\i_dmi_jtag_tap.idcode_d_6_ ),
    .Q_N(_0758_),
    .Q(\i_dmi_jtag_tap.idcode_q_6_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_7__reg  (.CLK(net397),
    .RESET_B(net352),
    .D(_0019_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_7_ ),
    .Q(_0008_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_8__reg  (.CLK(net396),
    .RESET_B(net348),
    .D(_0020_),
    .Q_N(\i_dmi_jtag_tap.idcode_q_8_ ),
    .Q(_0009_));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.idcode_q_9__reg  (.CLK(net396),
    .RESET_B(net348),
    .D(\i_dmi_jtag_tap.idcode_d_9_ ),
    .Q_N(_0757_),
    .Q(\i_dmi_jtag_tap.idcode_q_9_ ));
 sg13g2_dfrbp_2 \i_dmi_jtag_tap.jtag_ir_q_0__reg  (.RESET_B(net353),
    .D(_0068_),
    .Q(_0010_),
    .Q_N(\i_dmi_jtag_tap.jtag_ir_q_0_ ),
    .CLK(net404));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_q_1__reg  (.CLK(net399),
    .RESET_B(net353),
    .D(_0069_),
    .Q_N(_0756_),
    .Q(\i_dmi_jtag_tap.jtag_ir_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_q_2__reg  (.CLK(net399),
    .RESET_B(net353),
    .D(_0070_),
    .Q_N(_0755_),
    .Q(\i_dmi_jtag_tap.jtag_ir_q_2_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_q_3__reg  (.CLK(net399),
    .RESET_B(net353),
    .D(_0071_),
    .Q_N(_0754_),
    .Q(\i_dmi_jtag_tap.jtag_ir_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_q_4__reg  (.CLK(net399),
    .RESET_B(net353),
    .D(_0072_),
    .Q_N(\i_dmi_jtag_tap.jtag_ir_q_4__$_NOT__A_Y ),
    .Q(\i_dmi_jtag_tap.jtag_ir_q_4_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_shift_q_0__reg  (.CLK(net404),
    .RESET_B(net354),
    .D(_0073_),
    .Q_N(_0753_),
    .Q(\i_dmi_jtag_tap.jtag_ir_shift_q_0_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_shift_q_1__reg  (.CLK(net399),
    .RESET_B(net353),
    .D(_0074_),
    .Q_N(_0752_),
    .Q(\i_dmi_jtag_tap.jtag_ir_shift_q_1_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_shift_q_2__reg  (.CLK(net398),
    .RESET_B(net348),
    .D(_0021_),
    .Q_N(_0751_),
    .Q(\i_dmi_jtag_tap.jtag_ir_shift_q_2_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_shift_q_3__reg  (.CLK(net398),
    .RESET_B(net348),
    .D(_0022_),
    .Q_N(_0750_),
    .Q(\i_dmi_jtag_tap.jtag_ir_shift_q_3_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.jtag_ir_shift_q_4__reg  (.CLK(net399),
    .RESET_B(net348),
    .D(_0023_),
    .Q_N(_0749_),
    .Q(\i_dmi_jtag_tap.jtag_ir_shift_q_4_ ));
 sg13g2_dfrbp_1 \i_dmi_jtag_tap.tap_state_q_0__reg  (.CLK(net406),
    .RESET_B(net360),
    .D(_0011_),
    .Q_N(\i_dmi_jtag_tap.tap_state_q_0_ ),
    .Q(_0000_));
 sg13g2_dfrbp_2 \i_dmi_jtag_tap.tap_state_q_1__reg  (.RESET_B(net360),
    .D(\i_dmi_jtag_tap.tap_state_d_1_ ),
    .Q(\i_dmi_jtag_tap.tap_state_q_1_ ),
    .Q_N(\i_dmi_jtag_tap.tap_state_q_1__$_NOT__A_Y ),
    .CLK(net408));
 sg13g2_dfrbp_2 \i_dmi_jtag_tap.tap_state_q_2__reg  (.RESET_B(net360),
    .D(\i_dmi_jtag_tap.tap_state_d_2_ ),
    .Q(\i_dmi_jtag_tap.tap_state_q_2_ ),
    .Q_N(\i_dmi_jtag_tap.tap_state_q_2__$_NOT__A_Y ),
    .CLK(net408));
 sg13g2_dfrbp_2 \i_dmi_jtag_tap.tap_state_q_3__reg  (.RESET_B(net353),
    .D(\i_dmi_jtag_tap.tap_state_d_3_ ),
    .Q(\i_dmi_jtag_tap.tap_state_q_3_ ),
    .Q_N(\i_dmi_jtag_tap.tap_state_q_3__$_NOT__A_Y ),
    .CLK(net404));
 sg13g2_dfrbp_2 state_q_0__reg (.RESET_B(net361),
    .D(_0024_),
    .Q(state_q_0_),
    .Q_N(\state_q_0__$_NOT__A_Y ),
    .CLK(net409));
 sg13g2_dfrbp_2 state_q_1__reg (.RESET_B(net362),
    .D(_0025_),
    .Q(state_q_1_),
    .Q_N(\state_q_1__$_NOT__A_Y ),
    .CLK(net409));
 sg13g2_dfrbp_2 state_q_2__reg (.RESET_B(net362),
    .D(_0026_),
    .Q(state_q_2_),
    .Q_N(\state_q_0__$_OR__A_Y_$_OR__A_1_B ),
    .CLK(net409));
 sg13g2_dfrbp_2 td_o_reg (.RESET_B(net358),
    .D(\i_dmi_jtag_tap.tdo_mux ),
    .Q(td_o),
    .Q_N(_0892_),
    .CLK(\i_dmi_jtag_tap.tck_n ));
 sg13g2_dfrbp_2 tdo_oe_o_reg (.RESET_B(net362),
    .D(tdo_oe_o_reg_D),
    .Q(tdo_oe_o),
    .Q_N(_0748_),
    .CLK(\i_dmi_jtag_tap.tck_n ));
 sg13g2_tielo \i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/_108__1  (.L_LO(net1));
 sg13g2_tielo \i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/_108__2  (.L_LO(net2));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[10]_reg_5  (.L_HI(net5));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[11]_reg_6  (.L_HI(net6));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[12]_reg_7  (.L_HI(net7));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[13]_reg_8  (.L_HI(net8));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[14]_reg_9  (.L_HI(net9));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[15]_reg_10  (.L_HI(net10));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[16]_reg_11  (.L_HI(net11));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[17]_reg_12  (.L_HI(net12));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[18]_reg_13  (.L_HI(net13));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[19]_reg_14  (.L_HI(net14));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[1]_reg_15  (.L_HI(net15));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[20]_reg_16  (.L_HI(net16));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[21]_reg_17  (.L_HI(net17));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[22]_reg_18  (.L_HI(net18));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[23]_reg_19  (.L_HI(net19));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[24]_reg_20  (.L_HI(net20));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[25]_reg_21  (.L_HI(net21));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[26]_reg_22  (.L_HI(net22));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[27]_reg_23  (.L_HI(net23));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[28]_reg_24  (.L_HI(net24));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[29]_reg_25  (.L_HI(net25));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[2]_reg_26  (.L_HI(net26));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[30]_reg_27  (.L_HI(net27));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[31]_reg_28  (.L_HI(net28));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[32]_reg_29  (.L_HI(net29));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[33]_reg_30  (.L_HI(net30));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[34]_reg_31  (.L_HI(net31));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[35]_reg_32  (.L_HI(net32));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[36]_reg_33  (.L_HI(net33));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[37]_reg_34  (.L_HI(net34));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[38]_reg_35  (.L_HI(net35));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[39]_reg_36  (.L_HI(net36));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[3]_reg_37  (.L_HI(net37));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[40]_reg_38  (.L_HI(net38));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[4]_reg_39  (.L_HI(net39));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[5]_reg_40  (.L_HI(net40));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[6]_reg_41  (.L_HI(net41));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[7]_reg_42  (.L_HI(net42));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[8]_reg_43  (.L_HI(net43));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_dst/data_o[9]_reg_44  (.L_HI(net44));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[10]_reg_46  (.L_HI(net46));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[11]_reg_47  (.L_HI(net47));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[12]_reg_48  (.L_HI(net48));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[13]_reg_49  (.L_HI(net49));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[14]_reg_50  (.L_HI(net50));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[15]_reg_51  (.L_HI(net51));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[16]_reg_52  (.L_HI(net52));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[17]_reg_53  (.L_HI(net53));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[18]_reg_54  (.L_HI(net54));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[19]_reg_55  (.L_HI(net55));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[1]_reg_56  (.L_HI(net56));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[20]_reg_57  (.L_HI(net57));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[21]_reg_58  (.L_HI(net58));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[22]_reg_59  (.L_HI(net59));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[23]_reg_60  (.L_HI(net60));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[24]_reg_61  (.L_HI(net61));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[25]_reg_62  (.L_HI(net62));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[26]_reg_63  (.L_HI(net63));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[27]_reg_64  (.L_HI(net64));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[28]_reg_65  (.L_HI(net65));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[29]_reg_66  (.L_HI(net66));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[2]_reg_67  (.L_HI(net67));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[30]_reg_68  (.L_HI(net68));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[31]_reg_69  (.L_HI(net69));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[32]_reg_70  (.L_HI(net70));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[33]_reg_71  (.L_HI(net71));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[34]_reg_72  (.L_HI(net72));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[35]_reg_73  (.L_HI(net73));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[36]_reg_74  (.L_HI(net74));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[37]_reg_75  (.L_HI(net75));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[38]_reg_76  (.L_HI(net76));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[39]_reg_77  (.L_HI(net77));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[3]_reg_78  (.L_HI(net78));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[40]_reg_79  (.L_HI(net79));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[4]_reg_80  (.L_HI(net80));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[5]_reg_81  (.L_HI(net81));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[6]_reg_82  (.L_HI(net82));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[7]_reg_83  (.L_HI(net83));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[8]_reg_84  (.L_HI(net84));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_req/i_src/async_data_o[9]_reg_85  (.L_HI(net85));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[10]_reg_87  (.L_HI(net87));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[11]_reg_88  (.L_HI(net88));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[12]_reg_89  (.L_HI(net89));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[13]_reg_90  (.L_HI(net90));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[14]_reg_91  (.L_HI(net91));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[15]_reg_92  (.L_HI(net92));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[16]_reg_93  (.L_HI(net93));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[17]_reg_94  (.L_HI(net94));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[18]_reg_95  (.L_HI(net95));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[19]_reg_96  (.L_HI(net96));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[1]_reg_97  (.L_HI(net97));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[20]_reg_98  (.L_HI(net98));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[21]_reg_99  (.L_HI(net99));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[22]_reg_100  (.L_HI(net100));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[23]_reg_101  (.L_HI(net101));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[24]_reg_102  (.L_HI(net102));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[25]_reg_103  (.L_HI(net103));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[26]_reg_104  (.L_HI(net104));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[27]_reg_105  (.L_HI(net105));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[28]_reg_106  (.L_HI(net106));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[29]_reg_107  (.L_HI(net107));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[2]_reg_108  (.L_HI(net108));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[30]_reg_109  (.L_HI(net109));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[31]_reg_110  (.L_HI(net110));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[32]_reg_111  (.L_HI(net111));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[33]_reg_112  (.L_HI(net112));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[3]_reg_113  (.L_HI(net113));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[4]_reg_114  (.L_HI(net114));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[5]_reg_115  (.L_HI(net115));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[6]_reg_116  (.L_HI(net116));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[7]_reg_117  (.L_HI(net117));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[8]_reg_118  (.L_HI(net118));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_dst/data_o[9]_reg_119  (.L_HI(net119));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[10]_reg_121  (.L_HI(net121));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[11]_reg_122  (.L_HI(net122));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[12]_reg_123  (.L_HI(net123));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[13]_reg_124  (.L_HI(net124));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[14]_reg_125  (.L_HI(net125));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[15]_reg_126  (.L_HI(net126));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[16]_reg_127  (.L_HI(net127));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[17]_reg_128  (.L_HI(net128));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[18]_reg_129  (.L_HI(net129));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[19]_reg_130  (.L_HI(net130));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[1]_reg_131  (.L_HI(net131));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[20]_reg_132  (.L_HI(net132));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[21]_reg_133  (.L_HI(net133));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[22]_reg_134  (.L_HI(net134));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[23]_reg_135  (.L_HI(net135));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[24]_reg_136  (.L_HI(net136));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[25]_reg_137  (.L_HI(net137));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[26]_reg_138  (.L_HI(net138));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[27]_reg_139  (.L_HI(net139));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[28]_reg_140  (.L_HI(net140));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[29]_reg_141  (.L_HI(net141));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[2]_reg_142  (.L_HI(net142));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[30]_reg_143  (.L_HI(net143));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[31]_reg_144  (.L_HI(net144));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[32]_reg_145  (.L_HI(net145));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[33]_reg_146  (.L_HI(net146));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[3]_reg_147  (.L_HI(net147));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[4]_reg_148  (.L_HI(net148));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[5]_reg_149  (.L_HI(net149));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[6]_reg_150  (.L_HI(net150));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[7]_reg_151  (.L_HI(net151));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[8]_reg_152  (.L_HI(net152));
 sg13g2_tiehi \i_dmi_cdc.i_cdc_resp/i_src/async_data_o[9]_reg_153  (.L_HI(net153));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(net285));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(net286));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(net289));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(net289));
 sg13g2_buf_2 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_1 fanout289 (.A(\i_dmi_cdc.i_cdc_resp/i_dst/_040_ ),
    .X(net289));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(net296));
 sg13g2_buf_4 fanout291 (.X(net291),
    .A(net296));
 sg13g2_buf_4 fanout292 (.X(net292),
    .A(net293));
 sg13g2_buf_2 fanout293 (.A(net296),
    .X(net293));
 sg13g2_buf_4 fanout294 (.X(net294),
    .A(net295));
 sg13g2_buf_2 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(\i_dmi_cdc.i_cdc_req/i_dst/_047_ ),
    .X(net296));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(net302));
 sg13g2_buf_4 fanout298 (.X(net298),
    .A(net299));
 sg13g2_buf_4 fanout299 (.X(net299),
    .A(net302));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(net302));
 sg13g2_buf_2 fanout301 (.A(net302),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(\i_dmi_cdc.i_cdc_req/i_dst/_047_ ),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(net306),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(net306),
    .X(net304));
 sg13g2_buf_1 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(net309),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(net309),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(net309),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_0552_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_0394_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_0394_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_0347_),
    .X(net312));
 sg13g2_buf_1 fanout313 (.A(_0347_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(\i_dmi_jtag_tap.tap_state_q_3__$_NOT__A_Y ),
    .X(net314));
 sg13g2_buf_1 fanout315 (.A(\i_dmi_jtag_tap.tap_state_q_3__$_NOT__A_Y ),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(\i_dmi_jtag_tap.tap_state_q_2_ ),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(\i_dmi_jtag_tap.tap_state_q_1__$_NOT__A_Y ),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net320),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_1 fanout320 (.A(\i_dmi_jtag_tap.tap_state_q_0_ ),
    .X(net320));
 sg13g2_buf_2 fanout321 (.A(net323),
    .X(net321));
 sg13g2_buf_1 fanout322 (.A(net323),
    .X(net322));
 sg13g2_buf_2 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(dmi_resp_1_),
    .X(net324));
 sg13g2_buf_2 fanout325 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ),
    .X(net325));
 sg13g2_buf_2 fanout326 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .X(net326));
 sg13g2_buf_2 fanout327 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(net329),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_3_ ),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1__$_NOT__A_Y ),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .X(net332));
 sg13g2_buf_2 fanout333 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .X(net333));
 sg13g2_buf_1 fanout334 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_3_ ),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1__$_NOT__A_Y ),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_1_ ),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ),
    .X(net338));
 sg13g2_buf_1 fanout339 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/initiator_state_q_0_ ),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .X(net340));
 sg13g2_buf_1 fanout341 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_2_ ),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_1_ ),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/initiator_state_q_0_ ),
    .X(net344));
 sg13g2_buf_4 fanout345 (.X(net345),
    .A(net346));
 sg13g2_buf_4 fanout346 (.X(net346),
    .A(net348));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(net348));
 sg13g2_buf_4 fanout348 (.X(net348),
    .A(net363));
 sg13g2_buf_4 fanout349 (.X(net349),
    .A(net350));
 sg13g2_buf_4 fanout350 (.X(net350),
    .A(net363));
 sg13g2_buf_4 fanout351 (.X(net351),
    .A(net352));
 sg13g2_buf_4 fanout352 (.X(net352),
    .A(net354));
 sg13g2_buf_4 fanout353 (.X(net353),
    .A(net354));
 sg13g2_buf_2 fanout354 (.A(net362),
    .X(net354));
 sg13g2_buf_4 fanout355 (.X(net355),
    .A(net357));
 sg13g2_buf_4 fanout356 (.X(net356),
    .A(net357));
 sg13g2_buf_2 fanout357 (.A(net359),
    .X(net357));
 sg13g2_buf_4 fanout358 (.X(net358),
    .A(net359));
 sg13g2_buf_2 fanout359 (.A(net362),
    .X(net359));
 sg13g2_buf_4 fanout360 (.X(net360),
    .A(net361));
 sg13g2_buf_4 fanout361 (.X(net361),
    .A(net362));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(net363));
 sg13g2_buf_2 fanout363 (.A(trst_ni),
    .X(net363));
 sg13g2_buf_4 fanout364 (.X(net364),
    .A(net367));
 sg13g2_buf_4 fanout365 (.X(net365),
    .A(net367));
 sg13g2_buf_2 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(net380),
    .X(net367));
 sg13g2_buf_4 fanout368 (.X(net368),
    .A(net369));
 sg13g2_buf_2 fanout369 (.A(net380),
    .X(net369));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(net372));
 sg13g2_buf_2 fanout371 (.A(net372),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(net380));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(net374));
 sg13g2_buf_4 fanout374 (.X(net374),
    .A(net380));
 sg13g2_buf_4 fanout375 (.X(net375),
    .A(net379));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(net379));
 sg13g2_buf_4 fanout377 (.X(net377),
    .A(net379));
 sg13g2_buf_2 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(trst_ni),
    .X(net380));
 sg13g2_buf_4 fanout381 (.X(net381),
    .A(net382));
 sg13g2_buf_4 fanout382 (.X(net382),
    .A(net383));
 sg13g2_buf_4 fanout383 (.X(net383),
    .A(net388));
 sg13g2_buf_4 fanout384 (.X(net384),
    .A(net385));
 sg13g2_buf_4 fanout385 (.X(net385),
    .A(net386));
 sg13g2_buf_4 fanout386 (.X(net386),
    .A(net387));
 sg13g2_buf_4 fanout387 (.X(net387),
    .A(net388));
 sg13g2_buf_4 fanout388 (.X(net388),
    .A(rst_ni));
 sg13g2_buf_8 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_0_0_clk_i (.X(clknet_4_0_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_1_0_clk_i (.X(clknet_4_1_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_2_0_clk_i (.X(clknet_4_2_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_3_0_clk_i (.X(clknet_4_3_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_4_0_clk_i (.X(clknet_4_4_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_5_0_clk_i (.X(clknet_4_5_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_6_0_clk_i (.X(clknet_4_6_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_7_0_clk_i (.X(clknet_4_7_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_8_0_clk_i (.X(clknet_4_8_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_9_0_clk_i (.X(clknet_4_9_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_10_0_clk_i (.X(clknet_4_10_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_11_0_clk_i (.X(clknet_4_11_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_12_0_clk_i (.X(clknet_4_12_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_13_0_clk_i (.X(clknet_4_13_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_14_0_clk_i (.X(clknet_4_14_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_16 clkbuf_4_15_0_clk_i (.X(clknet_4_15_0_clk_i),
    .A(clknet_0_clk_i));
 sg13g2_buf_8 clkbuf_5_0__f_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_0__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_1__f_clk_i (.A(clknet_4_0_0_clk_i),
    .X(clknet_5_1__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_2__f_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_2__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_3__f_clk_i (.A(clknet_4_1_0_clk_i),
    .X(clknet_5_3__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_4__f_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_4__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_5__f_clk_i (.A(clknet_4_2_0_clk_i),
    .X(clknet_5_5__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_6__f_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_6__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_7__f_clk_i (.A(clknet_4_3_0_clk_i),
    .X(clknet_5_7__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_8__f_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_8__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_9__f_clk_i (.A(clknet_4_4_0_clk_i),
    .X(clknet_5_9__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_10__f_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_10__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_11__f_clk_i (.A(clknet_4_5_0_clk_i),
    .X(clknet_5_11__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_12__f_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_12__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_13__f_clk_i (.A(clknet_4_6_0_clk_i),
    .X(clknet_5_13__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_14__f_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_14__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_15__f_clk_i (.A(clknet_4_7_0_clk_i),
    .X(clknet_5_15__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_16__f_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_16__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_17__f_clk_i (.A(clknet_4_8_0_clk_i),
    .X(clknet_5_17__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_18__f_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_18__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_19__f_clk_i (.A(clknet_4_9_0_clk_i),
    .X(clknet_5_19__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_20__f_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_20__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_21__f_clk_i (.A(clknet_4_10_0_clk_i),
    .X(clknet_5_21__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_22__f_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_22__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_23__f_clk_i (.A(clknet_4_11_0_clk_i),
    .X(clknet_5_23__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_24__f_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_24__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_25__f_clk_i (.A(clknet_4_12_0_clk_i),
    .X(clknet_5_25__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_26__f_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_26__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_27__f_clk_i (.A(clknet_4_13_0_clk_i),
    .X(clknet_5_27__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_28__f_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_28__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_29__f_clk_i (.A(clknet_4_14_0_clk_i),
    .X(clknet_5_29__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_30__f_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_30__leaf_clk_i));
 sg13g2_buf_8 clkbuf_5_31__f_clk_i (.A(clknet_4_15_0_clk_i),
    .X(clknet_5_31__leaf_clk_i));
 sg13g2_buf_2 clkload0 (.A(clknet_5_5__leaf_clk_i));
 sg13g2_buf_2 clkload1 (.A(clknet_5_8__leaf_clk_i));
 sg13g2_buf_2 clkload2 (.A(clknet_5_11__leaf_clk_i));
 sg13g2_buf_2 clkload3 (.A(clknet_5_12__leaf_clk_i));
 sg13g2_inv_1 clkload4 (.A(clknet_5_15__leaf_clk_i));
 sg13g2_buf_2 clkload5 (.A(clknet_5_24__leaf_clk_i));
 sg13g2_buf_2 clkload6 (.A(clknet_5_26__leaf_clk_i));
 sg13g2_buf_2 clkload7 (.A(clknet_5_28__leaf_clk_i));
 sg13g2_inv_1 clkload8 (.A(clknet_5_31__leaf_clk_i));
 sg13g2_buf_1 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_1 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_1 fanout391 (.A(net412),
    .X(net391));
 sg13g2_buf_1 fanout392 (.A(net412),
    .X(net392));
 sg13g2_buf_1 fanout393 (.A(net395),
    .X(net393));
 sg13g2_buf_1 fanout394 (.A(net395),
    .X(net394));
 sg13g2_buf_1 fanout395 (.A(net412),
    .X(net395));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(net411),
    .X(net397));
 sg13g2_buf_1 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_1 fanout399 (.A(net411),
    .X(net399));
 sg13g2_buf_1 fanout400 (.A(net403),
    .X(net400));
 sg13g2_buf_1 fanout401 (.A(net403),
    .X(net401));
 sg13g2_buf_1 fanout402 (.A(net403),
    .X(net402));
 sg13g2_buf_1 fanout403 (.A(net405),
    .X(net403));
 sg13g2_buf_1 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_1 fanout405 (.A(net411),
    .X(net405));
 sg13g2_buf_1 fanout406 (.A(net410),
    .X(net406));
 sg13g2_buf_1 fanout407 (.A(net410),
    .X(net407));
 sg13g2_buf_1 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_1 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_1 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_1 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_1 fanout412 (.A(tck_i),
    .X(net412));
 sg13g2_buf_1 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_1 fanout414 (.A(net416),
    .X(net414));
 sg13g2_buf_1 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_1 fanout416 (.A(net425),
    .X(net416));
 sg13g2_buf_1 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_1 fanout418 (.A(net425),
    .X(net418));
 sg13g2_buf_1 fanout419 (.A(net425),
    .X(net419));
 sg13g2_buf_1 fanout420 (.A(net425),
    .X(net420));
 sg13g2_buf_1 fanout421 (.A(net424),
    .X(net421));
 sg13g2_buf_1 fanout422 (.A(net424),
    .X(net422));
 sg13g2_buf_1 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_1 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_1 fanout425 (.A(tck_i),
    .X(net425));
 sg13g2_buf_1 fanout426 (.A(net438),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(net438),
    .X(net427));
 sg13g2_buf_1 fanout428 (.A(net430),
    .X(net428));
 sg13g2_buf_1 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_1 fanout430 (.A(net438),
    .X(net430));
 sg13g2_buf_1 fanout431 (.A(net434),
    .X(net431));
 sg13g2_buf_1 fanout432 (.A(net434),
    .X(net432));
 sg13g2_buf_1 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_1 fanout434 (.A(net438),
    .X(net434));
 sg13g2_buf_1 fanout435 (.A(net436),
    .X(net435));
 sg13g2_buf_1 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_1 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_1 fanout438 (.A(tck_i),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_1_ ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_src/i_sync/reg_q_0_ ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_dmi_cdc.i_cdc_req/i_dst/req_synced ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold442 (.A(\i_dmi_cdc.i_cdc_req/i_dst/i_sync/reg_q_0_ ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_0_ ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold444 (.A(\i_dmi_cdc.i_cdc_resp/i_src/i_sync/reg_q_1_ ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_dst/i_sync/reg_q_0_ ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_dmi_cdc.i_cdc_req/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_b/i_state_transition_cdc_dst/i_sync/reg_q_0_ ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_dmi_cdc.i_cdc_resp/i_cdc_reset_ctrlr/i_cdc_reset_ctrlr_half_a/i_state_transition_cdc_src/i_sync/reg_q_0_ ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold448 (.A(\i_dmi_cdc.clear_pending_rise_edge_detect_$_AND__Y_A ),
    .X(net448));
 sg13g2_antennanp ANTENNA_1 (.A(_0470_));
 sg13g2_antennanp ANTENNA_2 (.A(dmi_req_ready_i));
 sg13g2_antennanp ANTENNA_3 (.A(_0470_));
 sg13g2_antennanp ANTENNA_4 (.A(_0470_));
 sg13g2_antennanp ANTENNA_5 (.A(_0470_));
 sg13g2_antennanp ANTENNA_6 (.A(_0470_));
 sg13g2_fill_8 FILLER_0_0 ();
 sg13g2_fill_8 FILLER_0_8 ();
 sg13g2_fill_8 FILLER_0_16 ();
 sg13g2_fill_8 FILLER_0_24 ();
 sg13g2_fill_8 FILLER_0_32 ();
 sg13g2_fill_8 FILLER_0_40 ();
 sg13g2_fill_8 FILLER_0_48 ();
 sg13g2_fill_8 FILLER_0_56 ();
 sg13g2_fill_8 FILLER_0_64 ();
 sg13g2_fill_8 FILLER_0_72 ();
 sg13g2_fill_8 FILLER_0_80 ();
 sg13g2_fill_8 FILLER_0_88 ();
 sg13g2_fill_8 FILLER_0_96 ();
 sg13g2_fill_8 FILLER_0_104 ();
 sg13g2_fill_8 FILLER_0_112 ();
 sg13g2_fill_8 FILLER_0_120 ();
 sg13g2_fill_8 FILLER_0_128 ();
 sg13g2_fill_8 FILLER_0_136 ();
 sg13g2_fill_8 FILLER_0_144 ();
 sg13g2_fill_8 FILLER_0_152 ();
 sg13g2_fill_8 FILLER_0_160 ();
 sg13g2_fill_8 FILLER_0_168 ();
 sg13g2_fill_8 FILLER_0_176 ();
 sg13g2_fill_8 FILLER_0_184 ();
 sg13g2_fill_8 FILLER_0_192 ();
 sg13g2_fill_8 FILLER_0_200 ();
 sg13g2_fill_8 FILLER_0_208 ();
 sg13g2_fill_8 FILLER_0_216 ();
 sg13g2_fill_8 FILLER_0_224 ();
 sg13g2_fill_8 FILLER_0_232 ();
 sg13g2_fill_8 FILLER_0_240 ();
 sg13g2_fill_8 FILLER_0_248 ();
 sg13g2_fill_8 FILLER_0_256 ();
 sg13g2_fill_8 FILLER_0_264 ();
 sg13g2_fill_8 FILLER_0_272 ();
 sg13g2_fill_8 FILLER_0_280 ();
 sg13g2_fill_8 FILLER_0_288 ();
 sg13g2_fill_8 FILLER_0_296 ();
 sg13g2_fill_8 FILLER_0_304 ();
 sg13g2_fill_8 FILLER_0_312 ();
 sg13g2_fill_8 FILLER_0_320 ();
 sg13g2_fill_8 FILLER_0_328 ();
 sg13g2_fill_8 FILLER_0_336 ();
 sg13g2_fill_8 FILLER_0_344 ();
 sg13g2_fill_8 FILLER_0_352 ();
 sg13g2_fill_8 FILLER_0_360 ();
 sg13g2_fill_8 FILLER_0_368 ();
 sg13g2_fill_8 FILLER_0_376 ();
 sg13g2_fill_8 FILLER_0_384 ();
 sg13g2_fill_8 FILLER_0_392 ();
 sg13g2_fill_8 FILLER_0_400 ();
 sg13g2_fill_8 FILLER_0_408 ();
 sg13g2_fill_8 FILLER_0_416 ();
 sg13g2_fill_8 FILLER_0_424 ();
 sg13g2_fill_8 FILLER_0_432 ();
 sg13g2_fill_8 FILLER_0_440 ();
 sg13g2_fill_8 FILLER_0_448 ();
 sg13g2_fill_8 FILLER_0_456 ();
 sg13g2_fill_8 FILLER_0_464 ();
 sg13g2_fill_8 FILLER_0_472 ();
 sg13g2_fill_8 FILLER_0_480 ();
 sg13g2_fill_8 FILLER_0_488 ();
 sg13g2_fill_8 FILLER_0_496 ();
 sg13g2_fill_8 FILLER_0_504 ();
 sg13g2_fill_8 FILLER_0_512 ();
 sg13g2_fill_8 FILLER_0_520 ();
 sg13g2_fill_8 FILLER_0_528 ();
 sg13g2_fill_8 FILLER_0_536 ();
 sg13g2_fill_8 FILLER_0_544 ();
 sg13g2_fill_8 FILLER_0_552 ();
 sg13g2_fill_8 FILLER_0_560 ();
 sg13g2_fill_8 FILLER_0_568 ();
 sg13g2_fill_8 FILLER_0_576 ();
 sg13g2_fill_8 FILLER_0_584 ();
 sg13g2_fill_8 FILLER_0_592 ();
 sg13g2_fill_8 FILLER_0_600 ();
 sg13g2_fill_8 FILLER_0_608 ();
 sg13g2_fill_8 FILLER_0_616 ();
 sg13g2_fill_8 FILLER_0_624 ();
 sg13g2_fill_8 FILLER_0_632 ();
 sg13g2_fill_8 FILLER_0_640 ();
 sg13g2_fill_8 FILLER_0_648 ();
 sg13g2_fill_8 FILLER_0_656 ();
 sg13g2_fill_8 FILLER_0_664 ();
 sg13g2_fill_8 FILLER_0_672 ();
 sg13g2_fill_8 FILLER_0_680 ();
 sg13g2_fill_8 FILLER_0_688 ();
 sg13g2_fill_8 FILLER_0_696 ();
 sg13g2_fill_8 FILLER_0_704 ();
 sg13g2_fill_8 FILLER_0_712 ();
 sg13g2_fill_8 FILLER_0_720 ();
 sg13g2_fill_8 FILLER_0_728 ();
 sg13g2_fill_8 FILLER_0_736 ();
 sg13g2_fill_8 FILLER_0_744 ();
 sg13g2_fill_8 FILLER_0_752 ();
 sg13g2_fill_8 FILLER_0_760 ();
 sg13g2_fill_8 FILLER_0_768 ();
 sg13g2_fill_8 FILLER_0_776 ();
 sg13g2_fill_8 FILLER_0_784 ();
 sg13g2_fill_8 FILLER_0_792 ();
 sg13g2_fill_8 FILLER_0_800 ();
 sg13g2_fill_8 FILLER_0_808 ();
 sg13g2_fill_8 FILLER_0_816 ();
 sg13g2_fill_8 FILLER_0_824 ();
 sg13g2_fill_8 FILLER_0_832 ();
 sg13g2_fill_8 FILLER_0_840 ();
 sg13g2_fill_8 FILLER_0_848 ();
 sg13g2_fill_8 FILLER_0_856 ();
 sg13g2_fill_8 FILLER_0_864 ();
 sg13g2_fill_8 FILLER_0_872 ();
 sg13g2_fill_8 FILLER_0_880 ();
 sg13g2_fill_8 FILLER_0_888 ();
 sg13g2_fill_8 FILLER_0_896 ();
 sg13g2_fill_8 FILLER_0_904 ();
 sg13g2_fill_8 FILLER_0_912 ();
 sg13g2_fill_8 FILLER_0_920 ();
 sg13g2_fill_8 FILLER_0_928 ();
 sg13g2_fill_8 FILLER_0_936 ();
 sg13g2_fill_8 FILLER_0_944 ();
 sg13g2_fill_8 FILLER_0_952 ();
 sg13g2_fill_8 FILLER_0_960 ();
 sg13g2_fill_8 FILLER_0_968 ();
 sg13g2_fill_8 FILLER_0_976 ();
 sg13g2_fill_8 FILLER_0_984 ();
 sg13g2_fill_8 FILLER_0_992 ();
 sg13g2_fill_8 FILLER_0_1000 ();
 sg13g2_fill_8 FILLER_0_1008 ();
 sg13g2_fill_8 FILLER_0_1016 ();
 sg13g2_fill_8 FILLER_0_1024 ();
 sg13g2_fill_8 FILLER_0_1032 ();
 sg13g2_fill_8 FILLER_0_1040 ();
 sg13g2_fill_8 FILLER_0_1048 ();
 sg13g2_fill_8 FILLER_0_1056 ();
 sg13g2_fill_8 FILLER_0_1064 ();
 sg13g2_fill_8 FILLER_0_1072 ();
 sg13g2_fill_8 FILLER_0_1080 ();
 sg13g2_fill_8 FILLER_0_1088 ();
 sg13g2_fill_8 FILLER_0_1096 ();
 sg13g2_fill_8 FILLER_0_1104 ();
 sg13g2_fill_8 FILLER_0_1112 ();
 sg13g2_fill_8 FILLER_0_1120 ();
 sg13g2_fill_8 FILLER_0_1128 ();
 sg13g2_fill_8 FILLER_0_1136 ();
 sg13g2_fill_8 FILLER_1_0 ();
 sg13g2_fill_8 FILLER_1_8 ();
 sg13g2_fill_8 FILLER_1_16 ();
 sg13g2_fill_8 FILLER_1_24 ();
 sg13g2_fill_8 FILLER_1_32 ();
 sg13g2_fill_8 FILLER_1_40 ();
 sg13g2_fill_8 FILLER_1_48 ();
 sg13g2_fill_8 FILLER_1_56 ();
 sg13g2_fill_8 FILLER_1_64 ();
 sg13g2_fill_8 FILLER_1_72 ();
 sg13g2_fill_8 FILLER_1_80 ();
 sg13g2_fill_8 FILLER_1_88 ();
 sg13g2_fill_8 FILLER_1_96 ();
 sg13g2_fill_8 FILLER_1_104 ();
 sg13g2_fill_8 FILLER_1_112 ();
 sg13g2_fill_8 FILLER_1_120 ();
 sg13g2_fill_8 FILLER_1_128 ();
 sg13g2_fill_8 FILLER_1_136 ();
 sg13g2_fill_8 FILLER_1_144 ();
 sg13g2_fill_8 FILLER_1_152 ();
 sg13g2_fill_8 FILLER_1_160 ();
 sg13g2_fill_8 FILLER_1_168 ();
 sg13g2_fill_8 FILLER_1_176 ();
 sg13g2_fill_8 FILLER_1_184 ();
 sg13g2_fill_8 FILLER_1_192 ();
 sg13g2_fill_8 FILLER_1_200 ();
 sg13g2_fill_8 FILLER_1_208 ();
 sg13g2_fill_8 FILLER_1_216 ();
 sg13g2_fill_8 FILLER_1_224 ();
 sg13g2_fill_8 FILLER_1_232 ();
 sg13g2_fill_8 FILLER_1_240 ();
 sg13g2_fill_8 FILLER_1_248 ();
 sg13g2_fill_8 FILLER_1_256 ();
 sg13g2_fill_8 FILLER_1_264 ();
 sg13g2_fill_8 FILLER_1_272 ();
 sg13g2_fill_8 FILLER_1_280 ();
 sg13g2_fill_8 FILLER_1_288 ();
 sg13g2_fill_8 FILLER_1_296 ();
 sg13g2_fill_8 FILLER_1_304 ();
 sg13g2_fill_8 FILLER_1_312 ();
 sg13g2_fill_8 FILLER_1_320 ();
 sg13g2_fill_8 FILLER_1_328 ();
 sg13g2_fill_8 FILLER_1_336 ();
 sg13g2_fill_8 FILLER_1_344 ();
 sg13g2_fill_8 FILLER_1_352 ();
 sg13g2_fill_8 FILLER_1_360 ();
 sg13g2_fill_8 FILLER_1_368 ();
 sg13g2_fill_8 FILLER_1_376 ();
 sg13g2_fill_8 FILLER_1_384 ();
 sg13g2_fill_8 FILLER_1_392 ();
 sg13g2_fill_8 FILLER_1_400 ();
 sg13g2_fill_8 FILLER_1_408 ();
 sg13g2_fill_8 FILLER_1_416 ();
 sg13g2_fill_8 FILLER_1_424 ();
 sg13g2_fill_8 FILLER_1_432 ();
 sg13g2_fill_8 FILLER_1_440 ();
 sg13g2_fill_8 FILLER_1_448 ();
 sg13g2_fill_8 FILLER_1_456 ();
 sg13g2_fill_8 FILLER_1_464 ();
 sg13g2_fill_8 FILLER_1_472 ();
 sg13g2_fill_8 FILLER_1_480 ();
 sg13g2_fill_8 FILLER_1_488 ();
 sg13g2_fill_8 FILLER_1_496 ();
 sg13g2_fill_8 FILLER_1_504 ();
 sg13g2_fill_8 FILLER_1_512 ();
 sg13g2_fill_8 FILLER_1_520 ();
 sg13g2_fill_8 FILLER_1_528 ();
 sg13g2_fill_8 FILLER_1_536 ();
 sg13g2_fill_8 FILLER_1_544 ();
 sg13g2_fill_8 FILLER_1_552 ();
 sg13g2_fill_8 FILLER_1_560 ();
 sg13g2_fill_8 FILLER_1_568 ();
 sg13g2_fill_8 FILLER_1_576 ();
 sg13g2_fill_8 FILLER_1_584 ();
 sg13g2_fill_8 FILLER_1_592 ();
 sg13g2_fill_8 FILLER_1_600 ();
 sg13g2_fill_8 FILLER_1_608 ();
 sg13g2_fill_8 FILLER_1_616 ();
 sg13g2_fill_8 FILLER_1_624 ();
 sg13g2_fill_8 FILLER_1_632 ();
 sg13g2_fill_8 FILLER_1_640 ();
 sg13g2_fill_8 FILLER_1_648 ();
 sg13g2_fill_8 FILLER_1_656 ();
 sg13g2_fill_8 FILLER_1_664 ();
 sg13g2_fill_8 FILLER_1_672 ();
 sg13g2_fill_8 FILLER_1_680 ();
 sg13g2_fill_8 FILLER_1_688 ();
 sg13g2_fill_8 FILLER_1_696 ();
 sg13g2_fill_8 FILLER_1_704 ();
 sg13g2_fill_8 FILLER_1_712 ();
 sg13g2_fill_8 FILLER_1_720 ();
 sg13g2_fill_8 FILLER_1_728 ();
 sg13g2_fill_8 FILLER_1_736 ();
 sg13g2_fill_8 FILLER_1_744 ();
 sg13g2_fill_8 FILLER_1_752 ();
 sg13g2_fill_8 FILLER_1_760 ();
 sg13g2_fill_8 FILLER_1_768 ();
 sg13g2_fill_8 FILLER_1_776 ();
 sg13g2_fill_8 FILLER_1_784 ();
 sg13g2_fill_8 FILLER_1_792 ();
 sg13g2_fill_8 FILLER_1_800 ();
 sg13g2_fill_8 FILLER_1_808 ();
 sg13g2_fill_8 FILLER_1_816 ();
 sg13g2_fill_8 FILLER_1_824 ();
 sg13g2_fill_8 FILLER_1_832 ();
 sg13g2_fill_8 FILLER_1_840 ();
 sg13g2_fill_8 FILLER_1_848 ();
 sg13g2_fill_8 FILLER_1_856 ();
 sg13g2_fill_8 FILLER_1_864 ();
 sg13g2_fill_8 FILLER_1_872 ();
 sg13g2_fill_8 FILLER_1_880 ();
 sg13g2_fill_8 FILLER_1_888 ();
 sg13g2_fill_8 FILLER_1_896 ();
 sg13g2_fill_8 FILLER_1_904 ();
 sg13g2_fill_8 FILLER_1_912 ();
 sg13g2_fill_8 FILLER_1_920 ();
 sg13g2_fill_8 FILLER_1_928 ();
 sg13g2_fill_8 FILLER_1_936 ();
 sg13g2_fill_8 FILLER_1_944 ();
 sg13g2_fill_8 FILLER_1_952 ();
 sg13g2_fill_8 FILLER_1_960 ();
 sg13g2_fill_8 FILLER_1_968 ();
 sg13g2_fill_8 FILLER_1_976 ();
 sg13g2_fill_8 FILLER_1_984 ();
 sg13g2_fill_8 FILLER_1_992 ();
 sg13g2_fill_8 FILLER_1_1000 ();
 sg13g2_fill_8 FILLER_1_1008 ();
 sg13g2_fill_8 FILLER_1_1016 ();
 sg13g2_fill_8 FILLER_1_1024 ();
 sg13g2_fill_8 FILLER_1_1032 ();
 sg13g2_fill_8 FILLER_1_1040 ();
 sg13g2_fill_8 FILLER_1_1048 ();
 sg13g2_fill_8 FILLER_1_1056 ();
 sg13g2_fill_8 FILLER_1_1064 ();
 sg13g2_fill_8 FILLER_1_1072 ();
 sg13g2_fill_8 FILLER_1_1080 ();
 sg13g2_fill_8 FILLER_1_1088 ();
 sg13g2_fill_8 FILLER_1_1096 ();
 sg13g2_fill_8 FILLER_1_1104 ();
 sg13g2_fill_8 FILLER_1_1112 ();
 sg13g2_fill_8 FILLER_1_1120 ();
 sg13g2_fill_8 FILLER_1_1128 ();
 sg13g2_fill_8 FILLER_1_1136 ();
 sg13g2_fill_8 FILLER_2_0 ();
 sg13g2_fill_8 FILLER_2_8 ();
 sg13g2_fill_8 FILLER_2_16 ();
 sg13g2_fill_8 FILLER_2_24 ();
 sg13g2_fill_8 FILLER_2_32 ();
 sg13g2_fill_8 FILLER_2_40 ();
 sg13g2_fill_8 FILLER_2_48 ();
 sg13g2_fill_8 FILLER_2_56 ();
 sg13g2_fill_8 FILLER_2_64 ();
 sg13g2_fill_8 FILLER_2_72 ();
 sg13g2_fill_8 FILLER_2_80 ();
 sg13g2_fill_8 FILLER_2_88 ();
 sg13g2_fill_8 FILLER_2_96 ();
 sg13g2_fill_8 FILLER_2_104 ();
 sg13g2_fill_8 FILLER_2_112 ();
 sg13g2_fill_8 FILLER_2_120 ();
 sg13g2_fill_8 FILLER_2_128 ();
 sg13g2_fill_8 FILLER_2_136 ();
 sg13g2_fill_8 FILLER_2_144 ();
 sg13g2_fill_8 FILLER_2_152 ();
 sg13g2_fill_8 FILLER_2_160 ();
 sg13g2_fill_8 FILLER_2_168 ();
 sg13g2_fill_8 FILLER_2_176 ();
 sg13g2_fill_8 FILLER_2_184 ();
 sg13g2_fill_8 FILLER_2_192 ();
 sg13g2_fill_8 FILLER_2_200 ();
 sg13g2_fill_8 FILLER_2_208 ();
 sg13g2_fill_8 FILLER_2_216 ();
 sg13g2_fill_8 FILLER_2_224 ();
 sg13g2_fill_8 FILLER_2_232 ();
 sg13g2_fill_8 FILLER_2_240 ();
 sg13g2_fill_8 FILLER_2_248 ();
 sg13g2_fill_8 FILLER_2_256 ();
 sg13g2_fill_8 FILLER_2_264 ();
 sg13g2_fill_8 FILLER_2_272 ();
 sg13g2_fill_8 FILLER_2_280 ();
 sg13g2_fill_8 FILLER_2_288 ();
 sg13g2_fill_8 FILLER_2_296 ();
 sg13g2_fill_8 FILLER_2_304 ();
 sg13g2_fill_8 FILLER_2_312 ();
 sg13g2_fill_8 FILLER_2_320 ();
 sg13g2_fill_8 FILLER_2_328 ();
 sg13g2_fill_8 FILLER_2_336 ();
 sg13g2_fill_8 FILLER_2_344 ();
 sg13g2_fill_8 FILLER_2_352 ();
 sg13g2_fill_8 FILLER_2_360 ();
 sg13g2_fill_8 FILLER_2_368 ();
 sg13g2_fill_8 FILLER_2_376 ();
 sg13g2_fill_8 FILLER_2_384 ();
 sg13g2_fill_8 FILLER_2_392 ();
 sg13g2_fill_8 FILLER_2_400 ();
 sg13g2_fill_8 FILLER_2_408 ();
 sg13g2_fill_8 FILLER_2_416 ();
 sg13g2_fill_8 FILLER_2_424 ();
 sg13g2_fill_8 FILLER_2_432 ();
 sg13g2_fill_8 FILLER_2_440 ();
 sg13g2_fill_8 FILLER_2_448 ();
 sg13g2_fill_8 FILLER_2_456 ();
 sg13g2_fill_8 FILLER_2_464 ();
 sg13g2_fill_8 FILLER_2_472 ();
 sg13g2_fill_8 FILLER_2_480 ();
 sg13g2_fill_8 FILLER_2_488 ();
 sg13g2_fill_8 FILLER_2_496 ();
 sg13g2_fill_8 FILLER_2_504 ();
 sg13g2_fill_8 FILLER_2_512 ();
 sg13g2_fill_8 FILLER_2_520 ();
 sg13g2_fill_8 FILLER_2_528 ();
 sg13g2_fill_8 FILLER_2_536 ();
 sg13g2_fill_8 FILLER_2_544 ();
 sg13g2_fill_8 FILLER_2_552 ();
 sg13g2_fill_8 FILLER_2_560 ();
 sg13g2_fill_8 FILLER_2_568 ();
 sg13g2_fill_8 FILLER_2_576 ();
 sg13g2_fill_8 FILLER_2_584 ();
 sg13g2_fill_8 FILLER_2_592 ();
 sg13g2_fill_8 FILLER_2_600 ();
 sg13g2_fill_8 FILLER_2_608 ();
 sg13g2_fill_8 FILLER_2_616 ();
 sg13g2_fill_8 FILLER_2_624 ();
 sg13g2_fill_8 FILLER_2_632 ();
 sg13g2_fill_8 FILLER_2_640 ();
 sg13g2_fill_8 FILLER_2_648 ();
 sg13g2_fill_8 FILLER_2_656 ();
 sg13g2_fill_8 FILLER_2_664 ();
 sg13g2_fill_8 FILLER_2_672 ();
 sg13g2_fill_8 FILLER_2_680 ();
 sg13g2_fill_8 FILLER_2_688 ();
 sg13g2_fill_8 FILLER_2_696 ();
 sg13g2_fill_8 FILLER_2_704 ();
 sg13g2_fill_8 FILLER_2_712 ();
 sg13g2_fill_8 FILLER_2_720 ();
 sg13g2_fill_8 FILLER_2_728 ();
 sg13g2_fill_8 FILLER_2_736 ();
 sg13g2_fill_8 FILLER_2_744 ();
 sg13g2_fill_8 FILLER_2_752 ();
 sg13g2_fill_8 FILLER_2_760 ();
 sg13g2_fill_8 FILLER_2_768 ();
 sg13g2_fill_8 FILLER_2_776 ();
 sg13g2_fill_8 FILLER_2_784 ();
 sg13g2_fill_8 FILLER_2_792 ();
 sg13g2_fill_8 FILLER_2_800 ();
 sg13g2_fill_8 FILLER_2_808 ();
 sg13g2_fill_8 FILLER_2_816 ();
 sg13g2_fill_8 FILLER_2_824 ();
 sg13g2_fill_8 FILLER_2_832 ();
 sg13g2_fill_8 FILLER_2_840 ();
 sg13g2_fill_8 FILLER_2_848 ();
 sg13g2_fill_8 FILLER_2_856 ();
 sg13g2_fill_8 FILLER_2_864 ();
 sg13g2_fill_8 FILLER_2_872 ();
 sg13g2_fill_8 FILLER_2_880 ();
 sg13g2_fill_8 FILLER_2_888 ();
 sg13g2_fill_8 FILLER_2_896 ();
 sg13g2_fill_8 FILLER_2_904 ();
 sg13g2_fill_8 FILLER_2_912 ();
 sg13g2_fill_8 FILLER_2_920 ();
 sg13g2_fill_8 FILLER_2_928 ();
 sg13g2_fill_8 FILLER_2_936 ();
 sg13g2_fill_8 FILLER_2_944 ();
 sg13g2_fill_8 FILLER_2_952 ();
 sg13g2_fill_8 FILLER_2_960 ();
 sg13g2_fill_8 FILLER_2_968 ();
 sg13g2_fill_8 FILLER_2_976 ();
 sg13g2_fill_8 FILLER_2_984 ();
 sg13g2_fill_8 FILLER_2_992 ();
 sg13g2_fill_8 FILLER_2_1000 ();
 sg13g2_fill_8 FILLER_2_1008 ();
 sg13g2_fill_8 FILLER_2_1016 ();
 sg13g2_fill_8 FILLER_2_1024 ();
 sg13g2_fill_8 FILLER_2_1032 ();
 sg13g2_fill_8 FILLER_2_1040 ();
 sg13g2_fill_8 FILLER_2_1048 ();
 sg13g2_fill_8 FILLER_2_1056 ();
 sg13g2_fill_8 FILLER_2_1064 ();
 sg13g2_fill_8 FILLER_2_1072 ();
 sg13g2_fill_8 FILLER_2_1080 ();
 sg13g2_fill_8 FILLER_2_1088 ();
 sg13g2_fill_8 FILLER_2_1096 ();
 sg13g2_fill_8 FILLER_2_1104 ();
 sg13g2_fill_8 FILLER_2_1112 ();
 sg13g2_fill_8 FILLER_2_1120 ();
 sg13g2_fill_8 FILLER_2_1128 ();
 sg13g2_fill_8 FILLER_2_1136 ();
 sg13g2_fill_8 FILLER_3_0 ();
 sg13g2_fill_8 FILLER_3_8 ();
 sg13g2_fill_8 FILLER_3_16 ();
 sg13g2_fill_8 FILLER_3_24 ();
 sg13g2_fill_8 FILLER_3_32 ();
 sg13g2_fill_8 FILLER_3_40 ();
 sg13g2_fill_8 FILLER_3_48 ();
 sg13g2_fill_8 FILLER_3_56 ();
 sg13g2_fill_8 FILLER_3_64 ();
 sg13g2_fill_8 FILLER_3_72 ();
 sg13g2_fill_8 FILLER_3_80 ();
 sg13g2_fill_8 FILLER_3_88 ();
 sg13g2_fill_8 FILLER_3_96 ();
 sg13g2_fill_8 FILLER_3_104 ();
 sg13g2_fill_8 FILLER_3_112 ();
 sg13g2_fill_8 FILLER_3_120 ();
 sg13g2_fill_8 FILLER_3_128 ();
 sg13g2_fill_8 FILLER_3_136 ();
 sg13g2_fill_8 FILLER_3_144 ();
 sg13g2_fill_8 FILLER_3_152 ();
 sg13g2_fill_8 FILLER_3_160 ();
 sg13g2_fill_8 FILLER_3_168 ();
 sg13g2_fill_8 FILLER_3_176 ();
 sg13g2_fill_8 FILLER_3_184 ();
 sg13g2_fill_8 FILLER_3_192 ();
 sg13g2_fill_8 FILLER_3_200 ();
 sg13g2_fill_8 FILLER_3_208 ();
 sg13g2_fill_8 FILLER_3_216 ();
 sg13g2_fill_8 FILLER_3_224 ();
 sg13g2_fill_8 FILLER_3_232 ();
 sg13g2_fill_8 FILLER_3_240 ();
 sg13g2_fill_8 FILLER_3_248 ();
 sg13g2_fill_8 FILLER_3_256 ();
 sg13g2_fill_8 FILLER_3_264 ();
 sg13g2_fill_8 FILLER_3_272 ();
 sg13g2_fill_8 FILLER_3_280 ();
 sg13g2_fill_8 FILLER_3_288 ();
 sg13g2_fill_8 FILLER_3_296 ();
 sg13g2_fill_8 FILLER_3_304 ();
 sg13g2_fill_8 FILLER_3_312 ();
 sg13g2_fill_8 FILLER_3_320 ();
 sg13g2_fill_8 FILLER_3_328 ();
 sg13g2_fill_8 FILLER_3_336 ();
 sg13g2_fill_8 FILLER_3_344 ();
 sg13g2_fill_8 FILLER_3_352 ();
 sg13g2_fill_8 FILLER_3_360 ();
 sg13g2_fill_8 FILLER_3_368 ();
 sg13g2_fill_8 FILLER_3_376 ();
 sg13g2_fill_8 FILLER_3_384 ();
 sg13g2_fill_8 FILLER_3_392 ();
 sg13g2_fill_8 FILLER_3_400 ();
 sg13g2_fill_8 FILLER_3_408 ();
 sg13g2_fill_8 FILLER_3_416 ();
 sg13g2_fill_8 FILLER_3_424 ();
 sg13g2_fill_8 FILLER_3_432 ();
 sg13g2_fill_8 FILLER_3_440 ();
 sg13g2_fill_8 FILLER_3_448 ();
 sg13g2_fill_8 FILLER_3_456 ();
 sg13g2_fill_8 FILLER_3_464 ();
 sg13g2_fill_8 FILLER_3_472 ();
 sg13g2_fill_8 FILLER_3_480 ();
 sg13g2_fill_8 FILLER_3_488 ();
 sg13g2_fill_8 FILLER_3_496 ();
 sg13g2_fill_8 FILLER_3_504 ();
 sg13g2_fill_8 FILLER_3_512 ();
 sg13g2_fill_8 FILLER_3_520 ();
 sg13g2_fill_8 FILLER_3_528 ();
 sg13g2_fill_8 FILLER_3_536 ();
 sg13g2_fill_8 FILLER_3_544 ();
 sg13g2_fill_8 FILLER_3_552 ();
 sg13g2_fill_8 FILLER_3_560 ();
 sg13g2_fill_8 FILLER_3_568 ();
 sg13g2_fill_8 FILLER_3_576 ();
 sg13g2_fill_8 FILLER_3_584 ();
 sg13g2_fill_8 FILLER_3_592 ();
 sg13g2_fill_8 FILLER_3_600 ();
 sg13g2_fill_8 FILLER_3_608 ();
 sg13g2_fill_8 FILLER_3_616 ();
 sg13g2_fill_8 FILLER_3_624 ();
 sg13g2_fill_8 FILLER_3_632 ();
 sg13g2_fill_8 FILLER_3_640 ();
 sg13g2_fill_8 FILLER_3_648 ();
 sg13g2_fill_8 FILLER_3_656 ();
 sg13g2_fill_8 FILLER_3_664 ();
 sg13g2_fill_8 FILLER_3_672 ();
 sg13g2_fill_8 FILLER_3_680 ();
 sg13g2_fill_8 FILLER_3_688 ();
 sg13g2_fill_8 FILLER_3_696 ();
 sg13g2_fill_8 FILLER_3_704 ();
 sg13g2_fill_8 FILLER_3_712 ();
 sg13g2_fill_8 FILLER_3_720 ();
 sg13g2_fill_8 FILLER_3_728 ();
 sg13g2_fill_8 FILLER_3_736 ();
 sg13g2_fill_8 FILLER_3_744 ();
 sg13g2_fill_8 FILLER_3_752 ();
 sg13g2_fill_8 FILLER_3_760 ();
 sg13g2_fill_8 FILLER_3_768 ();
 sg13g2_fill_8 FILLER_3_776 ();
 sg13g2_fill_8 FILLER_3_784 ();
 sg13g2_fill_8 FILLER_3_792 ();
 sg13g2_fill_8 FILLER_3_800 ();
 sg13g2_fill_8 FILLER_3_808 ();
 sg13g2_fill_8 FILLER_3_816 ();
 sg13g2_fill_8 FILLER_3_824 ();
 sg13g2_fill_8 FILLER_3_832 ();
 sg13g2_fill_8 FILLER_3_840 ();
 sg13g2_fill_8 FILLER_3_848 ();
 sg13g2_fill_8 FILLER_3_856 ();
 sg13g2_fill_8 FILLER_3_864 ();
 sg13g2_fill_8 FILLER_3_872 ();
 sg13g2_fill_8 FILLER_3_880 ();
 sg13g2_fill_8 FILLER_3_888 ();
 sg13g2_fill_8 FILLER_3_896 ();
 sg13g2_fill_8 FILLER_3_904 ();
 sg13g2_fill_8 FILLER_3_912 ();
 sg13g2_fill_8 FILLER_3_920 ();
 sg13g2_fill_8 FILLER_3_928 ();
 sg13g2_fill_8 FILLER_3_936 ();
 sg13g2_fill_8 FILLER_3_944 ();
 sg13g2_fill_8 FILLER_3_952 ();
 sg13g2_fill_8 FILLER_3_960 ();
 sg13g2_fill_8 FILLER_3_968 ();
 sg13g2_fill_8 FILLER_3_976 ();
 sg13g2_fill_8 FILLER_3_984 ();
 sg13g2_fill_8 FILLER_3_992 ();
 sg13g2_fill_8 FILLER_3_1000 ();
 sg13g2_fill_8 FILLER_3_1008 ();
 sg13g2_fill_8 FILLER_3_1016 ();
 sg13g2_fill_8 FILLER_3_1024 ();
 sg13g2_fill_8 FILLER_3_1032 ();
 sg13g2_fill_8 FILLER_3_1040 ();
 sg13g2_fill_8 FILLER_3_1048 ();
 sg13g2_fill_8 FILLER_3_1056 ();
 sg13g2_fill_8 FILLER_3_1064 ();
 sg13g2_fill_8 FILLER_3_1072 ();
 sg13g2_fill_8 FILLER_3_1080 ();
 sg13g2_fill_8 FILLER_3_1088 ();
 sg13g2_fill_8 FILLER_3_1096 ();
 sg13g2_fill_8 FILLER_3_1104 ();
 sg13g2_fill_8 FILLER_3_1112 ();
 sg13g2_fill_8 FILLER_3_1120 ();
 sg13g2_fill_8 FILLER_3_1128 ();
 sg13g2_fill_8 FILLER_3_1136 ();
 sg13g2_fill_8 FILLER_4_0 ();
 sg13g2_fill_8 FILLER_4_8 ();
 sg13g2_fill_8 FILLER_4_16 ();
 sg13g2_fill_8 FILLER_4_24 ();
 sg13g2_fill_8 FILLER_4_32 ();
 sg13g2_fill_8 FILLER_4_40 ();
 sg13g2_fill_8 FILLER_4_48 ();
 sg13g2_fill_8 FILLER_4_56 ();
 sg13g2_fill_8 FILLER_4_64 ();
 sg13g2_fill_8 FILLER_4_72 ();
 sg13g2_fill_8 FILLER_4_80 ();
 sg13g2_fill_8 FILLER_4_88 ();
 sg13g2_fill_8 FILLER_4_96 ();
 sg13g2_fill_8 FILLER_4_104 ();
 sg13g2_fill_8 FILLER_4_112 ();
 sg13g2_fill_8 FILLER_4_120 ();
 sg13g2_fill_8 FILLER_4_128 ();
 sg13g2_fill_8 FILLER_4_136 ();
 sg13g2_fill_8 FILLER_4_144 ();
 sg13g2_fill_8 FILLER_4_152 ();
 sg13g2_fill_8 FILLER_4_160 ();
 sg13g2_fill_8 FILLER_4_168 ();
 sg13g2_fill_8 FILLER_4_176 ();
 sg13g2_fill_8 FILLER_4_184 ();
 sg13g2_fill_8 FILLER_4_192 ();
 sg13g2_fill_8 FILLER_4_200 ();
 sg13g2_fill_8 FILLER_4_208 ();
 sg13g2_fill_8 FILLER_4_216 ();
 sg13g2_fill_8 FILLER_4_224 ();
 sg13g2_fill_8 FILLER_4_232 ();
 sg13g2_fill_8 FILLER_4_240 ();
 sg13g2_fill_8 FILLER_4_248 ();
 sg13g2_fill_8 FILLER_4_256 ();
 sg13g2_fill_8 FILLER_4_264 ();
 sg13g2_fill_8 FILLER_4_272 ();
 sg13g2_fill_8 FILLER_4_280 ();
 sg13g2_fill_8 FILLER_4_288 ();
 sg13g2_fill_8 FILLER_4_296 ();
 sg13g2_fill_8 FILLER_4_304 ();
 sg13g2_fill_8 FILLER_4_312 ();
 sg13g2_fill_8 FILLER_4_320 ();
 sg13g2_fill_8 FILLER_4_328 ();
 sg13g2_fill_8 FILLER_4_336 ();
 sg13g2_fill_8 FILLER_4_344 ();
 sg13g2_fill_8 FILLER_4_352 ();
 sg13g2_fill_8 FILLER_4_360 ();
 sg13g2_fill_8 FILLER_4_368 ();
 sg13g2_fill_8 FILLER_4_376 ();
 sg13g2_fill_8 FILLER_4_384 ();
 sg13g2_fill_8 FILLER_4_392 ();
 sg13g2_fill_8 FILLER_4_400 ();
 sg13g2_fill_8 FILLER_4_408 ();
 sg13g2_fill_8 FILLER_4_416 ();
 sg13g2_fill_8 FILLER_4_424 ();
 sg13g2_fill_8 FILLER_4_432 ();
 sg13g2_fill_8 FILLER_4_440 ();
 sg13g2_fill_8 FILLER_4_448 ();
 sg13g2_fill_8 FILLER_4_456 ();
 sg13g2_fill_8 FILLER_4_464 ();
 sg13g2_fill_8 FILLER_4_472 ();
 sg13g2_fill_8 FILLER_4_480 ();
 sg13g2_fill_8 FILLER_4_488 ();
 sg13g2_fill_8 FILLER_4_496 ();
 sg13g2_fill_8 FILLER_4_504 ();
 sg13g2_fill_8 FILLER_4_512 ();
 sg13g2_fill_8 FILLER_4_520 ();
 sg13g2_fill_8 FILLER_4_528 ();
 sg13g2_fill_8 FILLER_4_536 ();
 sg13g2_fill_8 FILLER_4_544 ();
 sg13g2_fill_8 FILLER_4_552 ();
 sg13g2_fill_8 FILLER_4_560 ();
 sg13g2_fill_8 FILLER_4_568 ();
 sg13g2_fill_8 FILLER_4_576 ();
 sg13g2_fill_8 FILLER_4_584 ();
 sg13g2_fill_8 FILLER_4_592 ();
 sg13g2_fill_8 FILLER_4_600 ();
 sg13g2_fill_8 FILLER_4_608 ();
 sg13g2_fill_8 FILLER_4_616 ();
 sg13g2_fill_8 FILLER_4_624 ();
 sg13g2_fill_8 FILLER_4_632 ();
 sg13g2_fill_8 FILLER_4_640 ();
 sg13g2_fill_8 FILLER_4_648 ();
 sg13g2_fill_8 FILLER_4_656 ();
 sg13g2_fill_8 FILLER_4_664 ();
 sg13g2_fill_8 FILLER_4_672 ();
 sg13g2_fill_8 FILLER_4_680 ();
 sg13g2_fill_8 FILLER_4_688 ();
 sg13g2_fill_8 FILLER_4_696 ();
 sg13g2_fill_8 FILLER_4_704 ();
 sg13g2_fill_8 FILLER_4_712 ();
 sg13g2_fill_8 FILLER_4_720 ();
 sg13g2_fill_8 FILLER_4_728 ();
 sg13g2_fill_8 FILLER_4_736 ();
 sg13g2_fill_8 FILLER_4_744 ();
 sg13g2_fill_8 FILLER_4_752 ();
 sg13g2_fill_8 FILLER_4_760 ();
 sg13g2_fill_8 FILLER_4_768 ();
 sg13g2_fill_8 FILLER_4_776 ();
 sg13g2_fill_8 FILLER_4_784 ();
 sg13g2_fill_8 FILLER_4_792 ();
 sg13g2_fill_8 FILLER_4_800 ();
 sg13g2_fill_8 FILLER_4_808 ();
 sg13g2_fill_8 FILLER_4_816 ();
 sg13g2_fill_8 FILLER_4_824 ();
 sg13g2_fill_8 FILLER_4_832 ();
 sg13g2_fill_8 FILLER_4_840 ();
 sg13g2_fill_8 FILLER_4_848 ();
 sg13g2_fill_8 FILLER_4_856 ();
 sg13g2_fill_8 FILLER_4_864 ();
 sg13g2_fill_8 FILLER_4_872 ();
 sg13g2_fill_8 FILLER_4_880 ();
 sg13g2_fill_8 FILLER_4_888 ();
 sg13g2_fill_8 FILLER_4_896 ();
 sg13g2_fill_8 FILLER_4_904 ();
 sg13g2_fill_8 FILLER_4_912 ();
 sg13g2_fill_8 FILLER_4_920 ();
 sg13g2_fill_8 FILLER_4_928 ();
 sg13g2_fill_8 FILLER_4_936 ();
 sg13g2_fill_8 FILLER_4_944 ();
 sg13g2_fill_8 FILLER_4_952 ();
 sg13g2_fill_8 FILLER_4_960 ();
 sg13g2_fill_8 FILLER_4_968 ();
 sg13g2_fill_8 FILLER_4_976 ();
 sg13g2_fill_8 FILLER_4_984 ();
 sg13g2_fill_8 FILLER_4_992 ();
 sg13g2_fill_8 FILLER_4_1000 ();
 sg13g2_fill_8 FILLER_4_1008 ();
 sg13g2_fill_8 FILLER_4_1016 ();
 sg13g2_fill_8 FILLER_4_1024 ();
 sg13g2_fill_8 FILLER_4_1032 ();
 sg13g2_fill_8 FILLER_4_1040 ();
 sg13g2_fill_8 FILLER_4_1048 ();
 sg13g2_fill_8 FILLER_4_1056 ();
 sg13g2_fill_8 FILLER_4_1064 ();
 sg13g2_fill_8 FILLER_4_1072 ();
 sg13g2_fill_8 FILLER_4_1080 ();
 sg13g2_fill_8 FILLER_4_1088 ();
 sg13g2_fill_8 FILLER_4_1096 ();
 sg13g2_fill_8 FILLER_4_1104 ();
 sg13g2_fill_8 FILLER_4_1112 ();
 sg13g2_fill_8 FILLER_4_1120 ();
 sg13g2_fill_8 FILLER_4_1128 ();
 sg13g2_fill_8 FILLER_4_1136 ();
 sg13g2_fill_8 FILLER_5_0 ();
 sg13g2_fill_8 FILLER_5_8 ();
 sg13g2_fill_8 FILLER_5_16 ();
 sg13g2_fill_8 FILLER_5_24 ();
 sg13g2_fill_8 FILLER_5_32 ();
 sg13g2_fill_8 FILLER_5_40 ();
 sg13g2_fill_8 FILLER_5_48 ();
 sg13g2_fill_8 FILLER_5_56 ();
 sg13g2_fill_8 FILLER_5_64 ();
 sg13g2_fill_8 FILLER_5_72 ();
 sg13g2_fill_8 FILLER_5_80 ();
 sg13g2_fill_8 FILLER_5_88 ();
 sg13g2_fill_8 FILLER_5_96 ();
 sg13g2_fill_8 FILLER_5_104 ();
 sg13g2_fill_8 FILLER_5_112 ();
 sg13g2_fill_8 FILLER_5_120 ();
 sg13g2_fill_8 FILLER_5_128 ();
 sg13g2_fill_8 FILLER_5_136 ();
 sg13g2_fill_8 FILLER_5_144 ();
 sg13g2_fill_8 FILLER_5_152 ();
 sg13g2_fill_8 FILLER_5_160 ();
 sg13g2_fill_8 FILLER_5_168 ();
 sg13g2_fill_8 FILLER_5_176 ();
 sg13g2_fill_8 FILLER_5_184 ();
 sg13g2_fill_8 FILLER_5_192 ();
 sg13g2_fill_8 FILLER_5_200 ();
 sg13g2_fill_8 FILLER_5_208 ();
 sg13g2_fill_8 FILLER_5_216 ();
 sg13g2_fill_8 FILLER_5_224 ();
 sg13g2_fill_8 FILLER_5_232 ();
 sg13g2_fill_8 FILLER_5_240 ();
 sg13g2_fill_8 FILLER_5_248 ();
 sg13g2_fill_8 FILLER_5_256 ();
 sg13g2_fill_8 FILLER_5_264 ();
 sg13g2_fill_8 FILLER_5_272 ();
 sg13g2_fill_8 FILLER_5_280 ();
 sg13g2_fill_8 FILLER_5_288 ();
 sg13g2_fill_8 FILLER_5_296 ();
 sg13g2_fill_8 FILLER_5_304 ();
 sg13g2_fill_8 FILLER_5_312 ();
 sg13g2_fill_8 FILLER_5_320 ();
 sg13g2_fill_8 FILLER_5_328 ();
 sg13g2_fill_8 FILLER_5_336 ();
 sg13g2_fill_8 FILLER_5_344 ();
 sg13g2_fill_8 FILLER_5_352 ();
 sg13g2_fill_8 FILLER_5_360 ();
 sg13g2_fill_8 FILLER_5_368 ();
 sg13g2_fill_8 FILLER_5_376 ();
 sg13g2_fill_8 FILLER_5_384 ();
 sg13g2_fill_8 FILLER_5_392 ();
 sg13g2_fill_8 FILLER_5_400 ();
 sg13g2_fill_8 FILLER_5_408 ();
 sg13g2_fill_8 FILLER_5_416 ();
 sg13g2_fill_8 FILLER_5_424 ();
 sg13g2_fill_8 FILLER_5_432 ();
 sg13g2_fill_8 FILLER_5_440 ();
 sg13g2_fill_8 FILLER_5_448 ();
 sg13g2_fill_8 FILLER_5_456 ();
 sg13g2_fill_8 FILLER_5_464 ();
 sg13g2_fill_8 FILLER_5_472 ();
 sg13g2_fill_8 FILLER_5_480 ();
 sg13g2_fill_8 FILLER_5_488 ();
 sg13g2_fill_8 FILLER_5_496 ();
 sg13g2_fill_8 FILLER_5_504 ();
 sg13g2_fill_8 FILLER_5_512 ();
 sg13g2_fill_8 FILLER_5_520 ();
 sg13g2_fill_8 FILLER_5_528 ();
 sg13g2_fill_8 FILLER_5_536 ();
 sg13g2_fill_8 FILLER_5_544 ();
 sg13g2_fill_8 FILLER_5_552 ();
 sg13g2_fill_8 FILLER_5_560 ();
 sg13g2_fill_8 FILLER_5_568 ();
 sg13g2_fill_8 FILLER_5_576 ();
 sg13g2_fill_8 FILLER_5_584 ();
 sg13g2_fill_8 FILLER_5_592 ();
 sg13g2_fill_8 FILLER_5_600 ();
 sg13g2_fill_8 FILLER_5_608 ();
 sg13g2_fill_8 FILLER_5_616 ();
 sg13g2_fill_8 FILLER_5_624 ();
 sg13g2_fill_8 FILLER_5_632 ();
 sg13g2_fill_8 FILLER_5_640 ();
 sg13g2_fill_8 FILLER_5_648 ();
 sg13g2_fill_8 FILLER_5_656 ();
 sg13g2_fill_8 FILLER_5_664 ();
 sg13g2_fill_8 FILLER_5_672 ();
 sg13g2_fill_8 FILLER_5_680 ();
 sg13g2_fill_8 FILLER_5_688 ();
 sg13g2_fill_8 FILLER_5_696 ();
 sg13g2_fill_8 FILLER_5_704 ();
 sg13g2_fill_8 FILLER_5_712 ();
 sg13g2_fill_8 FILLER_5_720 ();
 sg13g2_fill_8 FILLER_5_728 ();
 sg13g2_fill_8 FILLER_5_736 ();
 sg13g2_fill_8 FILLER_5_744 ();
 sg13g2_fill_8 FILLER_5_752 ();
 sg13g2_fill_8 FILLER_5_760 ();
 sg13g2_fill_8 FILLER_5_768 ();
 sg13g2_fill_8 FILLER_5_776 ();
 sg13g2_fill_8 FILLER_5_784 ();
 sg13g2_fill_8 FILLER_5_792 ();
 sg13g2_fill_8 FILLER_5_800 ();
 sg13g2_fill_8 FILLER_5_808 ();
 sg13g2_fill_8 FILLER_5_816 ();
 sg13g2_fill_8 FILLER_5_824 ();
 sg13g2_fill_8 FILLER_5_832 ();
 sg13g2_fill_8 FILLER_5_840 ();
 sg13g2_fill_8 FILLER_5_848 ();
 sg13g2_fill_8 FILLER_5_856 ();
 sg13g2_fill_8 FILLER_5_864 ();
 sg13g2_fill_8 FILLER_5_872 ();
 sg13g2_fill_8 FILLER_5_880 ();
 sg13g2_fill_8 FILLER_5_888 ();
 sg13g2_fill_8 FILLER_5_896 ();
 sg13g2_fill_8 FILLER_5_904 ();
 sg13g2_fill_8 FILLER_5_912 ();
 sg13g2_fill_8 FILLER_5_920 ();
 sg13g2_fill_8 FILLER_5_928 ();
 sg13g2_fill_8 FILLER_5_936 ();
 sg13g2_fill_8 FILLER_5_944 ();
 sg13g2_fill_8 FILLER_5_952 ();
 sg13g2_fill_8 FILLER_5_960 ();
 sg13g2_fill_8 FILLER_5_968 ();
 sg13g2_fill_8 FILLER_5_976 ();
 sg13g2_fill_8 FILLER_5_984 ();
 sg13g2_fill_8 FILLER_5_992 ();
 sg13g2_fill_8 FILLER_5_1000 ();
 sg13g2_fill_8 FILLER_5_1008 ();
 sg13g2_fill_8 FILLER_5_1016 ();
 sg13g2_fill_8 FILLER_5_1024 ();
 sg13g2_fill_8 FILLER_5_1032 ();
 sg13g2_fill_8 FILLER_5_1040 ();
 sg13g2_fill_8 FILLER_5_1048 ();
 sg13g2_fill_8 FILLER_5_1056 ();
 sg13g2_fill_8 FILLER_5_1064 ();
 sg13g2_fill_8 FILLER_5_1072 ();
 sg13g2_fill_8 FILLER_5_1080 ();
 sg13g2_fill_8 FILLER_5_1088 ();
 sg13g2_fill_8 FILLER_5_1096 ();
 sg13g2_fill_8 FILLER_5_1104 ();
 sg13g2_fill_8 FILLER_5_1112 ();
 sg13g2_fill_8 FILLER_5_1120 ();
 sg13g2_fill_8 FILLER_5_1128 ();
 sg13g2_fill_8 FILLER_5_1136 ();
 sg13g2_fill_8 FILLER_6_0 ();
 sg13g2_fill_8 FILLER_6_8 ();
 sg13g2_fill_8 FILLER_6_16 ();
 sg13g2_fill_8 FILLER_6_24 ();
 sg13g2_fill_8 FILLER_6_32 ();
 sg13g2_fill_8 FILLER_6_40 ();
 sg13g2_fill_8 FILLER_6_48 ();
 sg13g2_fill_8 FILLER_6_56 ();
 sg13g2_fill_8 FILLER_6_64 ();
 sg13g2_fill_8 FILLER_6_72 ();
 sg13g2_fill_8 FILLER_6_80 ();
 sg13g2_fill_8 FILLER_6_88 ();
 sg13g2_fill_8 FILLER_6_96 ();
 sg13g2_fill_8 FILLER_6_104 ();
 sg13g2_fill_8 FILLER_6_112 ();
 sg13g2_fill_8 FILLER_6_120 ();
 sg13g2_fill_8 FILLER_6_128 ();
 sg13g2_fill_8 FILLER_6_136 ();
 sg13g2_fill_8 FILLER_6_144 ();
 sg13g2_fill_8 FILLER_6_152 ();
 sg13g2_fill_8 FILLER_6_160 ();
 sg13g2_fill_8 FILLER_6_168 ();
 sg13g2_fill_8 FILLER_6_176 ();
 sg13g2_fill_8 FILLER_6_184 ();
 sg13g2_fill_8 FILLER_6_192 ();
 sg13g2_fill_8 FILLER_6_200 ();
 sg13g2_fill_8 FILLER_6_208 ();
 sg13g2_fill_8 FILLER_6_216 ();
 sg13g2_fill_8 FILLER_6_224 ();
 sg13g2_fill_8 FILLER_6_232 ();
 sg13g2_fill_8 FILLER_6_240 ();
 sg13g2_fill_8 FILLER_6_248 ();
 sg13g2_fill_8 FILLER_6_256 ();
 sg13g2_fill_8 FILLER_6_264 ();
 sg13g2_fill_8 FILLER_6_272 ();
 sg13g2_fill_8 FILLER_6_280 ();
 sg13g2_fill_8 FILLER_6_288 ();
 sg13g2_fill_8 FILLER_6_296 ();
 sg13g2_fill_8 FILLER_6_304 ();
 sg13g2_fill_8 FILLER_6_312 ();
 sg13g2_fill_8 FILLER_6_320 ();
 sg13g2_fill_8 FILLER_6_328 ();
 sg13g2_fill_8 FILLER_6_336 ();
 sg13g2_fill_8 FILLER_6_344 ();
 sg13g2_fill_8 FILLER_6_352 ();
 sg13g2_fill_8 FILLER_6_360 ();
 sg13g2_fill_8 FILLER_6_368 ();
 sg13g2_fill_8 FILLER_6_376 ();
 sg13g2_fill_8 FILLER_6_384 ();
 sg13g2_fill_8 FILLER_6_392 ();
 sg13g2_fill_8 FILLER_6_400 ();
 sg13g2_fill_8 FILLER_6_408 ();
 sg13g2_fill_8 FILLER_6_416 ();
 sg13g2_fill_8 FILLER_6_424 ();
 sg13g2_fill_8 FILLER_6_432 ();
 sg13g2_fill_8 FILLER_6_440 ();
 sg13g2_fill_8 FILLER_6_448 ();
 sg13g2_fill_8 FILLER_6_456 ();
 sg13g2_fill_8 FILLER_6_464 ();
 sg13g2_fill_8 FILLER_6_472 ();
 sg13g2_fill_8 FILLER_6_480 ();
 sg13g2_fill_8 FILLER_6_488 ();
 sg13g2_fill_8 FILLER_6_496 ();
 sg13g2_fill_8 FILLER_6_504 ();
 sg13g2_fill_8 FILLER_6_512 ();
 sg13g2_fill_8 FILLER_6_520 ();
 sg13g2_fill_8 FILLER_6_528 ();
 sg13g2_fill_8 FILLER_6_536 ();
 sg13g2_fill_8 FILLER_6_544 ();
 sg13g2_fill_8 FILLER_6_552 ();
 sg13g2_fill_8 FILLER_6_560 ();
 sg13g2_fill_8 FILLER_6_568 ();
 sg13g2_fill_8 FILLER_6_576 ();
 sg13g2_fill_8 FILLER_6_584 ();
 sg13g2_fill_8 FILLER_6_592 ();
 sg13g2_fill_8 FILLER_6_600 ();
 sg13g2_fill_8 FILLER_6_608 ();
 sg13g2_fill_8 FILLER_6_616 ();
 sg13g2_fill_8 FILLER_6_624 ();
 sg13g2_fill_8 FILLER_6_632 ();
 sg13g2_fill_8 FILLER_6_640 ();
 sg13g2_fill_8 FILLER_6_648 ();
 sg13g2_fill_8 FILLER_6_656 ();
 sg13g2_fill_8 FILLER_6_664 ();
 sg13g2_fill_8 FILLER_6_672 ();
 sg13g2_fill_8 FILLER_6_680 ();
 sg13g2_fill_8 FILLER_6_688 ();
 sg13g2_fill_8 FILLER_6_696 ();
 sg13g2_fill_8 FILLER_6_704 ();
 sg13g2_fill_8 FILLER_6_712 ();
 sg13g2_fill_8 FILLER_6_720 ();
 sg13g2_fill_8 FILLER_6_728 ();
 sg13g2_fill_8 FILLER_6_736 ();
 sg13g2_fill_8 FILLER_6_744 ();
 sg13g2_fill_8 FILLER_6_752 ();
 sg13g2_fill_8 FILLER_6_760 ();
 sg13g2_fill_8 FILLER_6_768 ();
 sg13g2_fill_8 FILLER_6_776 ();
 sg13g2_fill_8 FILLER_6_784 ();
 sg13g2_fill_8 FILLER_6_792 ();
 sg13g2_fill_8 FILLER_6_800 ();
 sg13g2_fill_8 FILLER_6_808 ();
 sg13g2_fill_8 FILLER_6_816 ();
 sg13g2_fill_8 FILLER_6_824 ();
 sg13g2_fill_8 FILLER_6_832 ();
 sg13g2_fill_8 FILLER_6_840 ();
 sg13g2_fill_8 FILLER_6_848 ();
 sg13g2_fill_8 FILLER_6_856 ();
 sg13g2_fill_8 FILLER_6_864 ();
 sg13g2_fill_8 FILLER_6_872 ();
 sg13g2_fill_8 FILLER_6_880 ();
 sg13g2_fill_8 FILLER_6_888 ();
 sg13g2_fill_8 FILLER_6_896 ();
 sg13g2_fill_8 FILLER_6_904 ();
 sg13g2_fill_8 FILLER_6_912 ();
 sg13g2_fill_8 FILLER_6_920 ();
 sg13g2_fill_8 FILLER_6_928 ();
 sg13g2_fill_8 FILLER_6_936 ();
 sg13g2_fill_8 FILLER_6_944 ();
 sg13g2_fill_8 FILLER_6_952 ();
 sg13g2_fill_8 FILLER_6_960 ();
 sg13g2_fill_8 FILLER_6_968 ();
 sg13g2_fill_8 FILLER_6_976 ();
 sg13g2_fill_8 FILLER_6_984 ();
 sg13g2_fill_8 FILLER_6_992 ();
 sg13g2_fill_8 FILLER_6_1000 ();
 sg13g2_fill_8 FILLER_6_1008 ();
 sg13g2_fill_8 FILLER_6_1016 ();
 sg13g2_fill_8 FILLER_6_1024 ();
 sg13g2_fill_8 FILLER_6_1032 ();
 sg13g2_fill_8 FILLER_6_1040 ();
 sg13g2_fill_8 FILLER_6_1048 ();
 sg13g2_fill_8 FILLER_6_1056 ();
 sg13g2_fill_8 FILLER_6_1064 ();
 sg13g2_fill_8 FILLER_6_1072 ();
 sg13g2_fill_8 FILLER_6_1080 ();
 sg13g2_fill_8 FILLER_6_1088 ();
 sg13g2_fill_8 FILLER_6_1096 ();
 sg13g2_fill_8 FILLER_6_1104 ();
 sg13g2_fill_8 FILLER_6_1112 ();
 sg13g2_fill_8 FILLER_6_1120 ();
 sg13g2_fill_8 FILLER_6_1128 ();
 sg13g2_fill_8 FILLER_6_1136 ();
 sg13g2_fill_8 FILLER_7_0 ();
 sg13g2_fill_8 FILLER_7_8 ();
 sg13g2_fill_8 FILLER_7_16 ();
 sg13g2_fill_8 FILLER_7_24 ();
 sg13g2_fill_8 FILLER_7_32 ();
 sg13g2_fill_8 FILLER_7_40 ();
 sg13g2_fill_8 FILLER_7_48 ();
 sg13g2_fill_8 FILLER_7_56 ();
 sg13g2_fill_8 FILLER_7_64 ();
 sg13g2_fill_8 FILLER_7_72 ();
 sg13g2_fill_8 FILLER_7_80 ();
 sg13g2_fill_8 FILLER_7_88 ();
 sg13g2_fill_8 FILLER_7_96 ();
 sg13g2_fill_8 FILLER_7_104 ();
 sg13g2_fill_8 FILLER_7_112 ();
 sg13g2_fill_8 FILLER_7_120 ();
 sg13g2_fill_8 FILLER_7_128 ();
 sg13g2_fill_8 FILLER_7_136 ();
 sg13g2_fill_8 FILLER_7_144 ();
 sg13g2_fill_8 FILLER_7_152 ();
 sg13g2_fill_8 FILLER_7_160 ();
 sg13g2_fill_8 FILLER_7_168 ();
 sg13g2_fill_8 FILLER_7_176 ();
 sg13g2_fill_8 FILLER_7_184 ();
 sg13g2_fill_8 FILLER_7_192 ();
 sg13g2_fill_8 FILLER_7_200 ();
 sg13g2_fill_8 FILLER_7_208 ();
 sg13g2_fill_8 FILLER_7_216 ();
 sg13g2_fill_8 FILLER_7_224 ();
 sg13g2_fill_8 FILLER_7_232 ();
 sg13g2_fill_8 FILLER_7_240 ();
 sg13g2_fill_8 FILLER_7_248 ();
 sg13g2_fill_8 FILLER_7_256 ();
 sg13g2_fill_8 FILLER_7_264 ();
 sg13g2_fill_8 FILLER_7_272 ();
 sg13g2_fill_8 FILLER_7_280 ();
 sg13g2_fill_8 FILLER_7_288 ();
 sg13g2_fill_8 FILLER_7_296 ();
 sg13g2_fill_8 FILLER_7_304 ();
 sg13g2_fill_8 FILLER_7_312 ();
 sg13g2_fill_8 FILLER_7_320 ();
 sg13g2_fill_8 FILLER_7_328 ();
 sg13g2_fill_8 FILLER_7_336 ();
 sg13g2_fill_8 FILLER_7_344 ();
 sg13g2_fill_8 FILLER_7_352 ();
 sg13g2_fill_8 FILLER_7_360 ();
 sg13g2_fill_8 FILLER_7_368 ();
 sg13g2_fill_8 FILLER_7_376 ();
 sg13g2_fill_8 FILLER_7_384 ();
 sg13g2_fill_8 FILLER_7_392 ();
 sg13g2_fill_8 FILLER_7_400 ();
 sg13g2_fill_8 FILLER_7_408 ();
 sg13g2_fill_8 FILLER_7_416 ();
 sg13g2_fill_8 FILLER_7_424 ();
 sg13g2_fill_8 FILLER_7_432 ();
 sg13g2_fill_8 FILLER_7_440 ();
 sg13g2_fill_8 FILLER_7_448 ();
 sg13g2_fill_8 FILLER_7_456 ();
 sg13g2_fill_8 FILLER_7_464 ();
 sg13g2_fill_8 FILLER_7_472 ();
 sg13g2_fill_8 FILLER_7_480 ();
 sg13g2_fill_8 FILLER_7_488 ();
 sg13g2_fill_8 FILLER_7_496 ();
 sg13g2_fill_8 FILLER_7_504 ();
 sg13g2_fill_8 FILLER_7_512 ();
 sg13g2_fill_8 FILLER_7_520 ();
 sg13g2_fill_8 FILLER_7_528 ();
 sg13g2_fill_8 FILLER_7_536 ();
 sg13g2_fill_8 FILLER_7_544 ();
 sg13g2_fill_8 FILLER_7_552 ();
 sg13g2_fill_8 FILLER_7_560 ();
 sg13g2_fill_8 FILLER_7_568 ();
 sg13g2_fill_8 FILLER_7_576 ();
 sg13g2_fill_8 FILLER_7_584 ();
 sg13g2_fill_8 FILLER_7_592 ();
 sg13g2_fill_8 FILLER_7_600 ();
 sg13g2_fill_8 FILLER_7_608 ();
 sg13g2_fill_8 FILLER_7_616 ();
 sg13g2_fill_8 FILLER_7_624 ();
 sg13g2_fill_8 FILLER_7_632 ();
 sg13g2_fill_8 FILLER_7_640 ();
 sg13g2_fill_8 FILLER_7_648 ();
 sg13g2_fill_8 FILLER_7_656 ();
 sg13g2_fill_8 FILLER_7_664 ();
 sg13g2_fill_8 FILLER_7_672 ();
 sg13g2_fill_8 FILLER_7_680 ();
 sg13g2_fill_8 FILLER_7_688 ();
 sg13g2_fill_8 FILLER_7_696 ();
 sg13g2_fill_8 FILLER_7_704 ();
 sg13g2_fill_8 FILLER_7_712 ();
 sg13g2_fill_8 FILLER_7_720 ();
 sg13g2_fill_8 FILLER_7_728 ();
 sg13g2_fill_8 FILLER_7_736 ();
 sg13g2_fill_8 FILLER_7_744 ();
 sg13g2_fill_8 FILLER_7_752 ();
 sg13g2_fill_8 FILLER_7_760 ();
 sg13g2_fill_8 FILLER_7_768 ();
 sg13g2_fill_8 FILLER_7_776 ();
 sg13g2_fill_8 FILLER_7_784 ();
 sg13g2_fill_8 FILLER_7_792 ();
 sg13g2_fill_8 FILLER_7_800 ();
 sg13g2_fill_8 FILLER_7_808 ();
 sg13g2_fill_8 FILLER_7_816 ();
 sg13g2_fill_8 FILLER_7_824 ();
 sg13g2_fill_8 FILLER_7_832 ();
 sg13g2_fill_8 FILLER_7_840 ();
 sg13g2_fill_8 FILLER_7_848 ();
 sg13g2_fill_8 FILLER_7_856 ();
 sg13g2_fill_8 FILLER_7_864 ();
 sg13g2_fill_8 FILLER_7_872 ();
 sg13g2_fill_8 FILLER_7_880 ();
 sg13g2_fill_8 FILLER_7_888 ();
 sg13g2_fill_8 FILLER_7_896 ();
 sg13g2_fill_8 FILLER_7_904 ();
 sg13g2_fill_8 FILLER_7_912 ();
 sg13g2_fill_8 FILLER_7_920 ();
 sg13g2_fill_8 FILLER_7_928 ();
 sg13g2_fill_8 FILLER_7_936 ();
 sg13g2_fill_8 FILLER_7_944 ();
 sg13g2_fill_8 FILLER_7_952 ();
 sg13g2_fill_8 FILLER_7_960 ();
 sg13g2_fill_8 FILLER_7_968 ();
 sg13g2_fill_8 FILLER_7_976 ();
 sg13g2_fill_8 FILLER_7_984 ();
 sg13g2_fill_8 FILLER_7_992 ();
 sg13g2_fill_8 FILLER_7_1000 ();
 sg13g2_fill_8 FILLER_7_1008 ();
 sg13g2_fill_8 FILLER_7_1016 ();
 sg13g2_fill_8 FILLER_7_1024 ();
 sg13g2_fill_8 FILLER_7_1032 ();
 sg13g2_fill_8 FILLER_7_1040 ();
 sg13g2_fill_8 FILLER_7_1048 ();
 sg13g2_fill_8 FILLER_7_1056 ();
 sg13g2_fill_8 FILLER_7_1064 ();
 sg13g2_fill_8 FILLER_7_1072 ();
 sg13g2_fill_8 FILLER_7_1080 ();
 sg13g2_fill_8 FILLER_7_1088 ();
 sg13g2_fill_8 FILLER_7_1096 ();
 sg13g2_fill_8 FILLER_7_1104 ();
 sg13g2_fill_8 FILLER_7_1112 ();
 sg13g2_fill_8 FILLER_7_1120 ();
 sg13g2_fill_8 FILLER_7_1128 ();
 sg13g2_fill_8 FILLER_7_1136 ();
 sg13g2_fill_8 FILLER_8_0 ();
 sg13g2_fill_8 FILLER_8_8 ();
 sg13g2_fill_8 FILLER_8_16 ();
 sg13g2_fill_8 FILLER_8_24 ();
 sg13g2_fill_8 FILLER_8_32 ();
 sg13g2_fill_8 FILLER_8_40 ();
 sg13g2_fill_8 FILLER_8_48 ();
 sg13g2_fill_8 FILLER_8_56 ();
 sg13g2_fill_8 FILLER_8_64 ();
 sg13g2_fill_8 FILLER_8_72 ();
 sg13g2_fill_8 FILLER_8_80 ();
 sg13g2_fill_8 FILLER_8_88 ();
 sg13g2_fill_8 FILLER_8_96 ();
 sg13g2_fill_8 FILLER_8_104 ();
 sg13g2_fill_8 FILLER_8_112 ();
 sg13g2_fill_8 FILLER_8_120 ();
 sg13g2_fill_8 FILLER_8_128 ();
 sg13g2_fill_8 FILLER_8_136 ();
 sg13g2_fill_8 FILLER_8_144 ();
 sg13g2_fill_8 FILLER_8_152 ();
 sg13g2_fill_8 FILLER_8_160 ();
 sg13g2_fill_8 FILLER_8_168 ();
 sg13g2_fill_8 FILLER_8_176 ();
 sg13g2_fill_8 FILLER_8_184 ();
 sg13g2_fill_8 FILLER_8_192 ();
 sg13g2_fill_8 FILLER_8_200 ();
 sg13g2_fill_8 FILLER_8_208 ();
 sg13g2_fill_8 FILLER_8_216 ();
 sg13g2_fill_8 FILLER_8_224 ();
 sg13g2_fill_8 FILLER_8_232 ();
 sg13g2_fill_8 FILLER_8_240 ();
 sg13g2_fill_8 FILLER_8_248 ();
 sg13g2_fill_8 FILLER_8_256 ();
 sg13g2_fill_8 FILLER_8_264 ();
 sg13g2_fill_8 FILLER_8_272 ();
 sg13g2_fill_8 FILLER_8_280 ();
 sg13g2_fill_8 FILLER_8_288 ();
 sg13g2_fill_8 FILLER_8_296 ();
 sg13g2_fill_8 FILLER_8_304 ();
 sg13g2_fill_8 FILLER_8_312 ();
 sg13g2_fill_8 FILLER_8_320 ();
 sg13g2_fill_8 FILLER_8_328 ();
 sg13g2_fill_8 FILLER_8_336 ();
 sg13g2_fill_8 FILLER_8_344 ();
 sg13g2_fill_8 FILLER_8_352 ();
 sg13g2_fill_8 FILLER_8_360 ();
 sg13g2_fill_8 FILLER_8_368 ();
 sg13g2_fill_8 FILLER_8_376 ();
 sg13g2_fill_8 FILLER_8_384 ();
 sg13g2_fill_8 FILLER_8_392 ();
 sg13g2_fill_8 FILLER_8_400 ();
 sg13g2_fill_8 FILLER_8_408 ();
 sg13g2_fill_8 FILLER_8_416 ();
 sg13g2_fill_8 FILLER_8_424 ();
 sg13g2_fill_8 FILLER_8_432 ();
 sg13g2_fill_8 FILLER_8_440 ();
 sg13g2_fill_8 FILLER_8_448 ();
 sg13g2_fill_8 FILLER_8_456 ();
 sg13g2_fill_8 FILLER_8_464 ();
 sg13g2_fill_8 FILLER_8_472 ();
 sg13g2_fill_8 FILLER_8_480 ();
 sg13g2_fill_8 FILLER_8_488 ();
 sg13g2_fill_8 FILLER_8_496 ();
 sg13g2_fill_8 FILLER_8_504 ();
 sg13g2_fill_8 FILLER_8_512 ();
 sg13g2_fill_8 FILLER_8_520 ();
 sg13g2_fill_8 FILLER_8_528 ();
 sg13g2_fill_8 FILLER_8_536 ();
 sg13g2_fill_8 FILLER_8_544 ();
 sg13g2_fill_8 FILLER_8_552 ();
 sg13g2_fill_8 FILLER_8_560 ();
 sg13g2_fill_8 FILLER_8_568 ();
 sg13g2_fill_8 FILLER_8_576 ();
 sg13g2_fill_8 FILLER_8_584 ();
 sg13g2_fill_8 FILLER_8_592 ();
 sg13g2_fill_8 FILLER_8_600 ();
 sg13g2_fill_8 FILLER_8_608 ();
 sg13g2_fill_8 FILLER_8_616 ();
 sg13g2_fill_8 FILLER_8_624 ();
 sg13g2_fill_8 FILLER_8_632 ();
 sg13g2_fill_8 FILLER_8_640 ();
 sg13g2_fill_8 FILLER_8_648 ();
 sg13g2_fill_8 FILLER_8_656 ();
 sg13g2_fill_8 FILLER_8_664 ();
 sg13g2_fill_8 FILLER_8_672 ();
 sg13g2_fill_8 FILLER_8_680 ();
 sg13g2_fill_8 FILLER_8_688 ();
 sg13g2_fill_8 FILLER_8_696 ();
 sg13g2_fill_8 FILLER_8_704 ();
 sg13g2_fill_8 FILLER_8_712 ();
 sg13g2_fill_8 FILLER_8_720 ();
 sg13g2_fill_8 FILLER_8_728 ();
 sg13g2_fill_8 FILLER_8_736 ();
 sg13g2_fill_8 FILLER_8_744 ();
 sg13g2_fill_8 FILLER_8_752 ();
 sg13g2_fill_8 FILLER_8_760 ();
 sg13g2_fill_8 FILLER_8_768 ();
 sg13g2_fill_8 FILLER_8_776 ();
 sg13g2_fill_8 FILLER_8_784 ();
 sg13g2_fill_8 FILLER_8_792 ();
 sg13g2_fill_8 FILLER_8_800 ();
 sg13g2_fill_8 FILLER_8_808 ();
 sg13g2_fill_8 FILLER_8_816 ();
 sg13g2_fill_8 FILLER_8_824 ();
 sg13g2_fill_8 FILLER_8_832 ();
 sg13g2_fill_8 FILLER_8_840 ();
 sg13g2_fill_8 FILLER_8_848 ();
 sg13g2_fill_8 FILLER_8_856 ();
 sg13g2_fill_8 FILLER_8_864 ();
 sg13g2_fill_8 FILLER_8_872 ();
 sg13g2_fill_8 FILLER_8_880 ();
 sg13g2_fill_8 FILLER_8_888 ();
 sg13g2_fill_8 FILLER_8_896 ();
 sg13g2_fill_8 FILLER_8_904 ();
 sg13g2_fill_8 FILLER_8_912 ();
 sg13g2_fill_8 FILLER_8_920 ();
 sg13g2_fill_8 FILLER_8_928 ();
 sg13g2_fill_8 FILLER_8_936 ();
 sg13g2_fill_8 FILLER_8_944 ();
 sg13g2_fill_8 FILLER_8_952 ();
 sg13g2_fill_8 FILLER_8_960 ();
 sg13g2_fill_8 FILLER_8_968 ();
 sg13g2_fill_8 FILLER_8_976 ();
 sg13g2_fill_8 FILLER_8_984 ();
 sg13g2_fill_8 FILLER_8_992 ();
 sg13g2_fill_8 FILLER_8_1000 ();
 sg13g2_fill_8 FILLER_8_1008 ();
 sg13g2_fill_8 FILLER_8_1016 ();
 sg13g2_fill_8 FILLER_8_1024 ();
 sg13g2_fill_8 FILLER_8_1032 ();
 sg13g2_fill_8 FILLER_8_1040 ();
 sg13g2_fill_8 FILLER_8_1048 ();
 sg13g2_fill_8 FILLER_8_1056 ();
 sg13g2_fill_8 FILLER_8_1064 ();
 sg13g2_fill_8 FILLER_8_1072 ();
 sg13g2_fill_8 FILLER_8_1080 ();
 sg13g2_fill_8 FILLER_8_1088 ();
 sg13g2_fill_8 FILLER_8_1096 ();
 sg13g2_fill_8 FILLER_8_1104 ();
 sg13g2_fill_8 FILLER_8_1112 ();
 sg13g2_fill_8 FILLER_8_1120 ();
 sg13g2_fill_8 FILLER_8_1128 ();
 sg13g2_fill_8 FILLER_8_1136 ();
 sg13g2_fill_8 FILLER_9_0 ();
 sg13g2_fill_8 FILLER_9_8 ();
 sg13g2_fill_8 FILLER_9_16 ();
 sg13g2_fill_8 FILLER_9_24 ();
 sg13g2_fill_8 FILLER_9_32 ();
 sg13g2_fill_8 FILLER_9_40 ();
 sg13g2_fill_8 FILLER_9_48 ();
 sg13g2_fill_8 FILLER_9_56 ();
 sg13g2_fill_8 FILLER_9_64 ();
 sg13g2_fill_8 FILLER_9_72 ();
 sg13g2_fill_8 FILLER_9_80 ();
 sg13g2_fill_8 FILLER_9_88 ();
 sg13g2_fill_8 FILLER_9_96 ();
 sg13g2_fill_8 FILLER_9_104 ();
 sg13g2_fill_8 FILLER_9_112 ();
 sg13g2_fill_8 FILLER_9_120 ();
 sg13g2_fill_8 FILLER_9_128 ();
 sg13g2_fill_8 FILLER_9_136 ();
 sg13g2_fill_8 FILLER_9_144 ();
 sg13g2_fill_8 FILLER_9_152 ();
 sg13g2_fill_8 FILLER_9_160 ();
 sg13g2_fill_8 FILLER_9_168 ();
 sg13g2_fill_8 FILLER_9_176 ();
 sg13g2_fill_8 FILLER_9_184 ();
 sg13g2_fill_8 FILLER_9_192 ();
 sg13g2_fill_8 FILLER_9_200 ();
 sg13g2_fill_8 FILLER_9_208 ();
 sg13g2_fill_8 FILLER_9_216 ();
 sg13g2_fill_8 FILLER_9_224 ();
 sg13g2_fill_8 FILLER_9_232 ();
 sg13g2_fill_8 FILLER_9_240 ();
 sg13g2_fill_8 FILLER_9_248 ();
 sg13g2_fill_8 FILLER_9_256 ();
 sg13g2_fill_8 FILLER_9_264 ();
 sg13g2_fill_8 FILLER_9_272 ();
 sg13g2_fill_8 FILLER_9_280 ();
 sg13g2_fill_8 FILLER_9_288 ();
 sg13g2_fill_8 FILLER_9_296 ();
 sg13g2_fill_8 FILLER_9_304 ();
 sg13g2_fill_8 FILLER_9_312 ();
 sg13g2_fill_8 FILLER_9_320 ();
 sg13g2_fill_8 FILLER_9_328 ();
 sg13g2_fill_8 FILLER_9_336 ();
 sg13g2_fill_8 FILLER_9_344 ();
 sg13g2_fill_8 FILLER_9_352 ();
 sg13g2_fill_8 FILLER_9_360 ();
 sg13g2_fill_8 FILLER_9_368 ();
 sg13g2_fill_8 FILLER_9_376 ();
 sg13g2_fill_8 FILLER_9_384 ();
 sg13g2_fill_8 FILLER_9_392 ();
 sg13g2_fill_8 FILLER_9_400 ();
 sg13g2_fill_8 FILLER_9_408 ();
 sg13g2_fill_8 FILLER_9_416 ();
 sg13g2_fill_8 FILLER_9_424 ();
 sg13g2_fill_8 FILLER_9_432 ();
 sg13g2_fill_8 FILLER_9_440 ();
 sg13g2_fill_8 FILLER_9_448 ();
 sg13g2_fill_8 FILLER_9_456 ();
 sg13g2_fill_8 FILLER_9_464 ();
 sg13g2_fill_8 FILLER_9_472 ();
 sg13g2_fill_8 FILLER_9_480 ();
 sg13g2_fill_8 FILLER_9_488 ();
 sg13g2_fill_8 FILLER_9_496 ();
 sg13g2_fill_8 FILLER_9_504 ();
 sg13g2_fill_8 FILLER_9_512 ();
 sg13g2_fill_8 FILLER_9_520 ();
 sg13g2_fill_8 FILLER_9_528 ();
 sg13g2_fill_8 FILLER_9_536 ();
 sg13g2_fill_8 FILLER_9_544 ();
 sg13g2_fill_8 FILLER_9_552 ();
 sg13g2_fill_8 FILLER_9_560 ();
 sg13g2_fill_8 FILLER_9_568 ();
 sg13g2_fill_8 FILLER_9_576 ();
 sg13g2_fill_8 FILLER_9_584 ();
 sg13g2_fill_8 FILLER_9_592 ();
 sg13g2_fill_8 FILLER_9_600 ();
 sg13g2_fill_8 FILLER_9_608 ();
 sg13g2_fill_8 FILLER_9_616 ();
 sg13g2_fill_8 FILLER_9_624 ();
 sg13g2_fill_8 FILLER_9_632 ();
 sg13g2_fill_8 FILLER_9_640 ();
 sg13g2_fill_8 FILLER_9_648 ();
 sg13g2_fill_8 FILLER_9_656 ();
 sg13g2_fill_8 FILLER_9_664 ();
 sg13g2_fill_8 FILLER_9_672 ();
 sg13g2_fill_8 FILLER_9_680 ();
 sg13g2_fill_8 FILLER_9_688 ();
 sg13g2_fill_8 FILLER_9_696 ();
 sg13g2_fill_8 FILLER_9_704 ();
 sg13g2_fill_8 FILLER_9_712 ();
 sg13g2_fill_8 FILLER_9_720 ();
 sg13g2_fill_8 FILLER_9_728 ();
 sg13g2_fill_8 FILLER_9_736 ();
 sg13g2_fill_8 FILLER_9_744 ();
 sg13g2_fill_8 FILLER_9_752 ();
 sg13g2_fill_8 FILLER_9_760 ();
 sg13g2_fill_8 FILLER_9_768 ();
 sg13g2_fill_8 FILLER_9_776 ();
 sg13g2_fill_8 FILLER_9_784 ();
 sg13g2_fill_8 FILLER_9_792 ();
 sg13g2_fill_8 FILLER_9_800 ();
 sg13g2_fill_8 FILLER_9_808 ();
 sg13g2_fill_8 FILLER_9_816 ();
 sg13g2_fill_8 FILLER_9_824 ();
 sg13g2_fill_8 FILLER_9_832 ();
 sg13g2_fill_8 FILLER_9_840 ();
 sg13g2_fill_8 FILLER_9_848 ();
 sg13g2_fill_8 FILLER_9_856 ();
 sg13g2_fill_8 FILLER_9_864 ();
 sg13g2_fill_8 FILLER_9_872 ();
 sg13g2_fill_8 FILLER_9_880 ();
 sg13g2_fill_8 FILLER_9_888 ();
 sg13g2_fill_8 FILLER_9_896 ();
 sg13g2_fill_8 FILLER_9_904 ();
 sg13g2_fill_8 FILLER_9_912 ();
 sg13g2_fill_8 FILLER_9_920 ();
 sg13g2_fill_8 FILLER_9_928 ();
 sg13g2_fill_8 FILLER_9_936 ();
 sg13g2_fill_8 FILLER_9_944 ();
 sg13g2_fill_8 FILLER_9_952 ();
 sg13g2_fill_8 FILLER_9_960 ();
 sg13g2_fill_8 FILLER_9_968 ();
 sg13g2_fill_8 FILLER_9_976 ();
 sg13g2_fill_8 FILLER_9_984 ();
 sg13g2_fill_8 FILLER_9_992 ();
 sg13g2_fill_8 FILLER_9_1000 ();
 sg13g2_fill_8 FILLER_9_1008 ();
 sg13g2_fill_8 FILLER_9_1016 ();
 sg13g2_fill_8 FILLER_9_1024 ();
 sg13g2_fill_8 FILLER_9_1032 ();
 sg13g2_fill_8 FILLER_9_1040 ();
 sg13g2_fill_8 FILLER_9_1048 ();
 sg13g2_fill_8 FILLER_9_1056 ();
 sg13g2_fill_8 FILLER_9_1064 ();
 sg13g2_fill_8 FILLER_9_1072 ();
 sg13g2_fill_8 FILLER_9_1080 ();
 sg13g2_fill_8 FILLER_9_1088 ();
 sg13g2_fill_8 FILLER_9_1096 ();
 sg13g2_fill_8 FILLER_9_1104 ();
 sg13g2_fill_8 FILLER_9_1112 ();
 sg13g2_fill_8 FILLER_9_1120 ();
 sg13g2_fill_8 FILLER_9_1128 ();
 sg13g2_fill_8 FILLER_9_1136 ();
 sg13g2_fill_8 FILLER_10_0 ();
 sg13g2_fill_8 FILLER_10_8 ();
 sg13g2_fill_8 FILLER_10_16 ();
 sg13g2_fill_8 FILLER_10_24 ();
 sg13g2_fill_8 FILLER_10_32 ();
 sg13g2_fill_8 FILLER_10_40 ();
 sg13g2_fill_8 FILLER_10_48 ();
 sg13g2_fill_8 FILLER_10_56 ();
 sg13g2_fill_8 FILLER_10_64 ();
 sg13g2_fill_8 FILLER_10_72 ();
 sg13g2_fill_8 FILLER_10_80 ();
 sg13g2_fill_8 FILLER_10_88 ();
 sg13g2_fill_8 FILLER_10_96 ();
 sg13g2_fill_8 FILLER_10_104 ();
 sg13g2_fill_8 FILLER_10_112 ();
 sg13g2_fill_8 FILLER_10_120 ();
 sg13g2_fill_8 FILLER_10_128 ();
 sg13g2_fill_8 FILLER_10_136 ();
 sg13g2_fill_8 FILLER_10_144 ();
 sg13g2_fill_8 FILLER_10_152 ();
 sg13g2_fill_8 FILLER_10_160 ();
 sg13g2_fill_8 FILLER_10_168 ();
 sg13g2_fill_8 FILLER_10_176 ();
 sg13g2_fill_8 FILLER_10_184 ();
 sg13g2_fill_8 FILLER_10_192 ();
 sg13g2_fill_8 FILLER_10_200 ();
 sg13g2_fill_8 FILLER_10_208 ();
 sg13g2_fill_8 FILLER_10_216 ();
 sg13g2_fill_8 FILLER_10_224 ();
 sg13g2_fill_8 FILLER_10_232 ();
 sg13g2_fill_8 FILLER_10_240 ();
 sg13g2_fill_8 FILLER_10_248 ();
 sg13g2_fill_8 FILLER_10_256 ();
 sg13g2_fill_8 FILLER_10_264 ();
 sg13g2_fill_8 FILLER_10_272 ();
 sg13g2_fill_8 FILLER_10_280 ();
 sg13g2_fill_8 FILLER_10_288 ();
 sg13g2_fill_8 FILLER_10_296 ();
 sg13g2_fill_8 FILLER_10_304 ();
 sg13g2_fill_8 FILLER_10_312 ();
 sg13g2_fill_8 FILLER_10_320 ();
 sg13g2_fill_8 FILLER_10_328 ();
 sg13g2_fill_8 FILLER_10_336 ();
 sg13g2_fill_8 FILLER_10_344 ();
 sg13g2_fill_8 FILLER_10_352 ();
 sg13g2_fill_8 FILLER_10_360 ();
 sg13g2_fill_8 FILLER_10_368 ();
 sg13g2_fill_8 FILLER_10_376 ();
 sg13g2_fill_8 FILLER_10_384 ();
 sg13g2_fill_8 FILLER_10_392 ();
 sg13g2_fill_8 FILLER_10_400 ();
 sg13g2_fill_8 FILLER_10_408 ();
 sg13g2_fill_8 FILLER_10_416 ();
 sg13g2_fill_8 FILLER_10_424 ();
 sg13g2_fill_8 FILLER_10_432 ();
 sg13g2_fill_8 FILLER_10_440 ();
 sg13g2_fill_8 FILLER_10_448 ();
 sg13g2_fill_8 FILLER_10_456 ();
 sg13g2_fill_8 FILLER_10_464 ();
 sg13g2_fill_8 FILLER_10_472 ();
 sg13g2_fill_8 FILLER_10_480 ();
 sg13g2_fill_8 FILLER_10_488 ();
 sg13g2_fill_8 FILLER_10_496 ();
 sg13g2_fill_8 FILLER_10_504 ();
 sg13g2_fill_8 FILLER_10_512 ();
 sg13g2_fill_8 FILLER_10_520 ();
 sg13g2_fill_8 FILLER_10_528 ();
 sg13g2_fill_8 FILLER_10_536 ();
 sg13g2_fill_8 FILLER_10_544 ();
 sg13g2_fill_8 FILLER_10_552 ();
 sg13g2_fill_8 FILLER_10_560 ();
 sg13g2_fill_8 FILLER_10_568 ();
 sg13g2_fill_8 FILLER_10_576 ();
 sg13g2_fill_8 FILLER_10_584 ();
 sg13g2_fill_8 FILLER_10_592 ();
 sg13g2_fill_8 FILLER_10_600 ();
 sg13g2_fill_8 FILLER_10_608 ();
 sg13g2_fill_8 FILLER_10_616 ();
 sg13g2_fill_8 FILLER_10_624 ();
 sg13g2_fill_8 FILLER_10_632 ();
 sg13g2_fill_8 FILLER_10_640 ();
 sg13g2_fill_8 FILLER_10_648 ();
 sg13g2_fill_8 FILLER_10_656 ();
 sg13g2_fill_8 FILLER_10_664 ();
 sg13g2_fill_8 FILLER_10_672 ();
 sg13g2_fill_8 FILLER_10_680 ();
 sg13g2_fill_8 FILLER_10_688 ();
 sg13g2_fill_8 FILLER_10_696 ();
 sg13g2_fill_8 FILLER_10_704 ();
 sg13g2_fill_8 FILLER_10_712 ();
 sg13g2_fill_8 FILLER_10_720 ();
 sg13g2_fill_8 FILLER_10_728 ();
 sg13g2_fill_8 FILLER_10_736 ();
 sg13g2_fill_8 FILLER_10_744 ();
 sg13g2_fill_8 FILLER_10_752 ();
 sg13g2_fill_8 FILLER_10_760 ();
 sg13g2_fill_8 FILLER_10_768 ();
 sg13g2_fill_8 FILLER_10_776 ();
 sg13g2_fill_8 FILLER_10_784 ();
 sg13g2_fill_8 FILLER_10_792 ();
 sg13g2_fill_8 FILLER_10_800 ();
 sg13g2_fill_8 FILLER_10_808 ();
 sg13g2_fill_8 FILLER_10_816 ();
 sg13g2_fill_8 FILLER_10_824 ();
 sg13g2_fill_8 FILLER_10_832 ();
 sg13g2_fill_8 FILLER_10_840 ();
 sg13g2_fill_8 FILLER_10_848 ();
 sg13g2_fill_8 FILLER_10_856 ();
 sg13g2_fill_8 FILLER_10_864 ();
 sg13g2_fill_8 FILLER_10_872 ();
 sg13g2_fill_8 FILLER_10_880 ();
 sg13g2_fill_8 FILLER_10_888 ();
 sg13g2_fill_8 FILLER_10_896 ();
 sg13g2_fill_8 FILLER_10_904 ();
 sg13g2_fill_8 FILLER_10_912 ();
 sg13g2_fill_8 FILLER_10_920 ();
 sg13g2_fill_8 FILLER_10_928 ();
 sg13g2_fill_8 FILLER_10_936 ();
 sg13g2_fill_8 FILLER_10_944 ();
 sg13g2_fill_8 FILLER_10_952 ();
 sg13g2_fill_8 FILLER_10_960 ();
 sg13g2_fill_8 FILLER_10_968 ();
 sg13g2_fill_8 FILLER_10_976 ();
 sg13g2_fill_8 FILLER_10_984 ();
 sg13g2_fill_8 FILLER_10_992 ();
 sg13g2_fill_8 FILLER_10_1000 ();
 sg13g2_fill_8 FILLER_10_1008 ();
 sg13g2_fill_8 FILLER_10_1016 ();
 sg13g2_fill_8 FILLER_10_1024 ();
 sg13g2_fill_8 FILLER_10_1032 ();
 sg13g2_fill_8 FILLER_10_1040 ();
 sg13g2_fill_8 FILLER_10_1048 ();
 sg13g2_fill_8 FILLER_10_1056 ();
 sg13g2_fill_8 FILLER_10_1064 ();
 sg13g2_fill_8 FILLER_10_1072 ();
 sg13g2_fill_8 FILLER_10_1080 ();
 sg13g2_fill_8 FILLER_10_1088 ();
 sg13g2_fill_8 FILLER_10_1096 ();
 sg13g2_fill_8 FILLER_10_1104 ();
 sg13g2_fill_8 FILLER_10_1112 ();
 sg13g2_fill_8 FILLER_10_1120 ();
 sg13g2_fill_8 FILLER_10_1128 ();
 sg13g2_fill_8 FILLER_10_1136 ();
 sg13g2_fill_8 FILLER_11_0 ();
 sg13g2_fill_8 FILLER_11_8 ();
 sg13g2_fill_8 FILLER_11_16 ();
 sg13g2_fill_8 FILLER_11_24 ();
 sg13g2_fill_8 FILLER_11_32 ();
 sg13g2_fill_8 FILLER_11_40 ();
 sg13g2_fill_8 FILLER_11_48 ();
 sg13g2_fill_8 FILLER_11_56 ();
 sg13g2_fill_8 FILLER_11_64 ();
 sg13g2_fill_8 FILLER_11_72 ();
 sg13g2_fill_8 FILLER_11_80 ();
 sg13g2_fill_8 FILLER_11_88 ();
 sg13g2_fill_8 FILLER_11_96 ();
 sg13g2_fill_8 FILLER_11_104 ();
 sg13g2_fill_8 FILLER_11_112 ();
 sg13g2_fill_8 FILLER_11_120 ();
 sg13g2_fill_8 FILLER_11_128 ();
 sg13g2_fill_8 FILLER_11_136 ();
 sg13g2_fill_8 FILLER_11_144 ();
 sg13g2_fill_8 FILLER_11_152 ();
 sg13g2_fill_8 FILLER_11_160 ();
 sg13g2_fill_8 FILLER_11_168 ();
 sg13g2_fill_8 FILLER_11_176 ();
 sg13g2_fill_8 FILLER_11_184 ();
 sg13g2_fill_8 FILLER_11_192 ();
 sg13g2_fill_8 FILLER_11_200 ();
 sg13g2_fill_8 FILLER_11_208 ();
 sg13g2_fill_8 FILLER_11_216 ();
 sg13g2_fill_8 FILLER_11_224 ();
 sg13g2_fill_8 FILLER_11_232 ();
 sg13g2_fill_8 FILLER_11_240 ();
 sg13g2_fill_8 FILLER_11_248 ();
 sg13g2_fill_8 FILLER_11_256 ();
 sg13g2_fill_8 FILLER_11_264 ();
 sg13g2_fill_8 FILLER_11_272 ();
 sg13g2_fill_8 FILLER_11_280 ();
 sg13g2_fill_8 FILLER_11_288 ();
 sg13g2_fill_8 FILLER_11_296 ();
 sg13g2_fill_8 FILLER_11_304 ();
 sg13g2_fill_8 FILLER_11_312 ();
 sg13g2_fill_8 FILLER_11_320 ();
 sg13g2_fill_8 FILLER_11_328 ();
 sg13g2_fill_8 FILLER_11_336 ();
 sg13g2_fill_8 FILLER_11_344 ();
 sg13g2_fill_8 FILLER_11_352 ();
 sg13g2_fill_8 FILLER_11_360 ();
 sg13g2_fill_8 FILLER_11_368 ();
 sg13g2_fill_8 FILLER_11_376 ();
 sg13g2_fill_8 FILLER_11_384 ();
 sg13g2_fill_8 FILLER_11_392 ();
 sg13g2_fill_8 FILLER_11_400 ();
 sg13g2_fill_8 FILLER_11_408 ();
 sg13g2_fill_8 FILLER_11_416 ();
 sg13g2_fill_8 FILLER_11_424 ();
 sg13g2_fill_8 FILLER_11_432 ();
 sg13g2_fill_8 FILLER_11_440 ();
 sg13g2_fill_8 FILLER_11_448 ();
 sg13g2_fill_8 FILLER_11_456 ();
 sg13g2_fill_8 FILLER_11_464 ();
 sg13g2_fill_8 FILLER_11_472 ();
 sg13g2_fill_8 FILLER_11_480 ();
 sg13g2_fill_8 FILLER_11_488 ();
 sg13g2_fill_8 FILLER_11_496 ();
 sg13g2_fill_8 FILLER_11_504 ();
 sg13g2_fill_8 FILLER_11_512 ();
 sg13g2_fill_8 FILLER_11_520 ();
 sg13g2_fill_8 FILLER_11_528 ();
 sg13g2_fill_8 FILLER_11_536 ();
 sg13g2_fill_8 FILLER_11_544 ();
 sg13g2_fill_8 FILLER_11_552 ();
 sg13g2_fill_8 FILLER_11_560 ();
 sg13g2_fill_8 FILLER_11_568 ();
 sg13g2_fill_8 FILLER_11_576 ();
 sg13g2_fill_8 FILLER_11_584 ();
 sg13g2_fill_8 FILLER_11_592 ();
 sg13g2_fill_8 FILLER_11_600 ();
 sg13g2_fill_8 FILLER_11_608 ();
 sg13g2_fill_8 FILLER_11_616 ();
 sg13g2_fill_8 FILLER_11_624 ();
 sg13g2_fill_8 FILLER_11_632 ();
 sg13g2_fill_8 FILLER_11_640 ();
 sg13g2_fill_8 FILLER_11_648 ();
 sg13g2_fill_8 FILLER_11_656 ();
 sg13g2_fill_8 FILLER_11_664 ();
 sg13g2_fill_8 FILLER_11_672 ();
 sg13g2_fill_8 FILLER_11_680 ();
 sg13g2_fill_8 FILLER_11_688 ();
 sg13g2_fill_8 FILLER_11_696 ();
 sg13g2_fill_8 FILLER_11_704 ();
 sg13g2_fill_8 FILLER_11_712 ();
 sg13g2_fill_8 FILLER_11_720 ();
 sg13g2_fill_8 FILLER_11_728 ();
 sg13g2_fill_8 FILLER_11_736 ();
 sg13g2_fill_8 FILLER_11_744 ();
 sg13g2_fill_8 FILLER_11_752 ();
 sg13g2_fill_8 FILLER_11_760 ();
 sg13g2_fill_8 FILLER_11_768 ();
 sg13g2_fill_8 FILLER_11_776 ();
 sg13g2_fill_8 FILLER_11_784 ();
 sg13g2_fill_8 FILLER_11_792 ();
 sg13g2_fill_8 FILLER_11_800 ();
 sg13g2_fill_8 FILLER_11_808 ();
 sg13g2_fill_8 FILLER_11_816 ();
 sg13g2_fill_8 FILLER_11_824 ();
 sg13g2_fill_8 FILLER_11_832 ();
 sg13g2_fill_8 FILLER_11_840 ();
 sg13g2_fill_8 FILLER_11_848 ();
 sg13g2_fill_8 FILLER_11_856 ();
 sg13g2_fill_8 FILLER_11_864 ();
 sg13g2_fill_8 FILLER_11_872 ();
 sg13g2_fill_8 FILLER_11_880 ();
 sg13g2_fill_8 FILLER_11_888 ();
 sg13g2_fill_8 FILLER_11_896 ();
 sg13g2_fill_8 FILLER_11_904 ();
 sg13g2_fill_8 FILLER_11_912 ();
 sg13g2_fill_8 FILLER_11_920 ();
 sg13g2_fill_8 FILLER_11_928 ();
 sg13g2_fill_8 FILLER_11_936 ();
 sg13g2_fill_8 FILLER_11_944 ();
 sg13g2_fill_8 FILLER_11_952 ();
 sg13g2_fill_8 FILLER_11_960 ();
 sg13g2_fill_8 FILLER_11_968 ();
 sg13g2_fill_8 FILLER_11_976 ();
 sg13g2_fill_8 FILLER_11_984 ();
 sg13g2_fill_8 FILLER_11_992 ();
 sg13g2_fill_8 FILLER_11_1000 ();
 sg13g2_fill_8 FILLER_11_1008 ();
 sg13g2_fill_8 FILLER_11_1016 ();
 sg13g2_fill_8 FILLER_11_1024 ();
 sg13g2_fill_8 FILLER_11_1032 ();
 sg13g2_fill_8 FILLER_11_1040 ();
 sg13g2_fill_8 FILLER_11_1048 ();
 sg13g2_fill_8 FILLER_11_1056 ();
 sg13g2_fill_8 FILLER_11_1064 ();
 sg13g2_fill_8 FILLER_11_1072 ();
 sg13g2_fill_8 FILLER_11_1080 ();
 sg13g2_fill_8 FILLER_11_1088 ();
 sg13g2_fill_8 FILLER_11_1096 ();
 sg13g2_fill_8 FILLER_11_1104 ();
 sg13g2_fill_8 FILLER_11_1112 ();
 sg13g2_fill_8 FILLER_11_1120 ();
 sg13g2_fill_8 FILLER_11_1128 ();
 sg13g2_fill_8 FILLER_11_1136 ();
 sg13g2_fill_8 FILLER_12_0 ();
 sg13g2_fill_8 FILLER_12_8 ();
 sg13g2_fill_8 FILLER_12_16 ();
 sg13g2_fill_8 FILLER_12_24 ();
 sg13g2_fill_8 FILLER_12_32 ();
 sg13g2_fill_8 FILLER_12_40 ();
 sg13g2_fill_8 FILLER_12_48 ();
 sg13g2_fill_8 FILLER_12_56 ();
 sg13g2_fill_8 FILLER_12_64 ();
 sg13g2_fill_8 FILLER_12_72 ();
 sg13g2_fill_8 FILLER_12_80 ();
 sg13g2_fill_8 FILLER_12_88 ();
 sg13g2_fill_8 FILLER_12_96 ();
 sg13g2_fill_8 FILLER_12_104 ();
 sg13g2_fill_8 FILLER_12_112 ();
 sg13g2_fill_8 FILLER_12_120 ();
 sg13g2_fill_8 FILLER_12_128 ();
 sg13g2_fill_8 FILLER_12_136 ();
 sg13g2_fill_8 FILLER_12_144 ();
 sg13g2_fill_8 FILLER_12_152 ();
 sg13g2_fill_8 FILLER_12_160 ();
 sg13g2_fill_8 FILLER_12_168 ();
 sg13g2_fill_8 FILLER_12_176 ();
 sg13g2_fill_8 FILLER_12_184 ();
 sg13g2_fill_8 FILLER_12_192 ();
 sg13g2_fill_8 FILLER_12_200 ();
 sg13g2_fill_8 FILLER_12_208 ();
 sg13g2_fill_8 FILLER_12_216 ();
 sg13g2_fill_8 FILLER_12_224 ();
 sg13g2_fill_8 FILLER_12_232 ();
 sg13g2_fill_8 FILLER_12_240 ();
 sg13g2_fill_8 FILLER_12_248 ();
 sg13g2_fill_8 FILLER_12_256 ();
 sg13g2_fill_8 FILLER_12_264 ();
 sg13g2_fill_8 FILLER_12_272 ();
 sg13g2_fill_8 FILLER_12_280 ();
 sg13g2_fill_8 FILLER_12_288 ();
 sg13g2_fill_8 FILLER_12_296 ();
 sg13g2_fill_8 FILLER_12_304 ();
 sg13g2_fill_8 FILLER_12_312 ();
 sg13g2_fill_8 FILLER_12_320 ();
 sg13g2_fill_8 FILLER_12_328 ();
 sg13g2_fill_8 FILLER_12_336 ();
 sg13g2_fill_8 FILLER_12_344 ();
 sg13g2_fill_8 FILLER_12_352 ();
 sg13g2_fill_8 FILLER_12_360 ();
 sg13g2_fill_8 FILLER_12_368 ();
 sg13g2_fill_8 FILLER_12_376 ();
 sg13g2_fill_8 FILLER_12_384 ();
 sg13g2_fill_8 FILLER_12_392 ();
 sg13g2_fill_8 FILLER_12_400 ();
 sg13g2_fill_8 FILLER_12_408 ();
 sg13g2_fill_8 FILLER_12_416 ();
 sg13g2_fill_8 FILLER_12_424 ();
 sg13g2_fill_8 FILLER_12_432 ();
 sg13g2_fill_8 FILLER_12_440 ();
 sg13g2_fill_8 FILLER_12_448 ();
 sg13g2_fill_8 FILLER_12_456 ();
 sg13g2_fill_8 FILLER_12_464 ();
 sg13g2_fill_8 FILLER_12_472 ();
 sg13g2_fill_8 FILLER_12_480 ();
 sg13g2_fill_8 FILLER_12_488 ();
 sg13g2_fill_8 FILLER_12_496 ();
 sg13g2_fill_8 FILLER_12_504 ();
 sg13g2_fill_8 FILLER_12_512 ();
 sg13g2_fill_8 FILLER_12_520 ();
 sg13g2_fill_8 FILLER_12_528 ();
 sg13g2_fill_8 FILLER_12_536 ();
 sg13g2_fill_8 FILLER_12_544 ();
 sg13g2_fill_8 FILLER_12_552 ();
 sg13g2_fill_8 FILLER_12_560 ();
 sg13g2_fill_8 FILLER_12_568 ();
 sg13g2_fill_8 FILLER_12_576 ();
 sg13g2_fill_8 FILLER_12_584 ();
 sg13g2_fill_8 FILLER_12_592 ();
 sg13g2_fill_8 FILLER_12_600 ();
 sg13g2_fill_8 FILLER_12_608 ();
 sg13g2_fill_8 FILLER_12_616 ();
 sg13g2_fill_8 FILLER_12_624 ();
 sg13g2_fill_8 FILLER_12_632 ();
 sg13g2_fill_8 FILLER_12_640 ();
 sg13g2_fill_8 FILLER_12_648 ();
 sg13g2_fill_8 FILLER_12_656 ();
 sg13g2_fill_8 FILLER_12_664 ();
 sg13g2_fill_8 FILLER_12_672 ();
 sg13g2_fill_8 FILLER_12_680 ();
 sg13g2_fill_8 FILLER_12_688 ();
 sg13g2_fill_8 FILLER_12_696 ();
 sg13g2_fill_8 FILLER_12_704 ();
 sg13g2_fill_8 FILLER_12_712 ();
 sg13g2_fill_8 FILLER_12_720 ();
 sg13g2_fill_8 FILLER_12_728 ();
 sg13g2_fill_8 FILLER_12_736 ();
 sg13g2_fill_8 FILLER_12_744 ();
 sg13g2_fill_8 FILLER_12_752 ();
 sg13g2_fill_8 FILLER_12_760 ();
 sg13g2_fill_8 FILLER_12_768 ();
 sg13g2_fill_8 FILLER_12_776 ();
 sg13g2_fill_8 FILLER_12_784 ();
 sg13g2_fill_8 FILLER_12_792 ();
 sg13g2_fill_8 FILLER_12_800 ();
 sg13g2_fill_8 FILLER_12_808 ();
 sg13g2_fill_8 FILLER_12_816 ();
 sg13g2_fill_8 FILLER_12_824 ();
 sg13g2_fill_8 FILLER_12_832 ();
 sg13g2_fill_8 FILLER_12_840 ();
 sg13g2_fill_8 FILLER_12_848 ();
 sg13g2_fill_8 FILLER_12_856 ();
 sg13g2_fill_8 FILLER_12_864 ();
 sg13g2_fill_8 FILLER_12_872 ();
 sg13g2_fill_8 FILLER_12_880 ();
 sg13g2_fill_8 FILLER_12_888 ();
 sg13g2_fill_8 FILLER_12_896 ();
 sg13g2_fill_8 FILLER_12_904 ();
 sg13g2_fill_8 FILLER_12_912 ();
 sg13g2_fill_8 FILLER_12_920 ();
 sg13g2_fill_8 FILLER_12_928 ();
 sg13g2_fill_8 FILLER_12_936 ();
 sg13g2_fill_8 FILLER_12_944 ();
 sg13g2_fill_8 FILLER_12_952 ();
 sg13g2_fill_8 FILLER_12_960 ();
 sg13g2_fill_8 FILLER_12_968 ();
 sg13g2_fill_8 FILLER_12_976 ();
 sg13g2_fill_8 FILLER_12_984 ();
 sg13g2_fill_8 FILLER_12_992 ();
 sg13g2_fill_8 FILLER_12_1000 ();
 sg13g2_fill_8 FILLER_12_1008 ();
 sg13g2_fill_8 FILLER_12_1016 ();
 sg13g2_fill_8 FILLER_12_1024 ();
 sg13g2_fill_8 FILLER_12_1032 ();
 sg13g2_fill_8 FILLER_12_1040 ();
 sg13g2_fill_8 FILLER_12_1048 ();
 sg13g2_fill_8 FILLER_12_1056 ();
 sg13g2_fill_8 FILLER_12_1064 ();
 sg13g2_fill_8 FILLER_12_1072 ();
 sg13g2_fill_8 FILLER_12_1080 ();
 sg13g2_fill_8 FILLER_12_1088 ();
 sg13g2_fill_8 FILLER_12_1096 ();
 sg13g2_fill_8 FILLER_12_1104 ();
 sg13g2_fill_8 FILLER_12_1112 ();
 sg13g2_fill_8 FILLER_12_1120 ();
 sg13g2_fill_8 FILLER_12_1128 ();
 sg13g2_fill_8 FILLER_12_1136 ();
 sg13g2_fill_8 FILLER_13_0 ();
 sg13g2_fill_8 FILLER_13_8 ();
 sg13g2_fill_8 FILLER_13_16 ();
 sg13g2_fill_8 FILLER_13_24 ();
 sg13g2_fill_8 FILLER_13_32 ();
 sg13g2_fill_8 FILLER_13_40 ();
 sg13g2_fill_8 FILLER_13_48 ();
 sg13g2_fill_8 FILLER_13_56 ();
 sg13g2_fill_8 FILLER_13_64 ();
 sg13g2_fill_8 FILLER_13_72 ();
 sg13g2_fill_8 FILLER_13_80 ();
 sg13g2_fill_8 FILLER_13_88 ();
 sg13g2_fill_8 FILLER_13_96 ();
 sg13g2_fill_8 FILLER_13_104 ();
 sg13g2_fill_8 FILLER_13_112 ();
 sg13g2_fill_8 FILLER_13_120 ();
 sg13g2_fill_8 FILLER_13_128 ();
 sg13g2_fill_8 FILLER_13_136 ();
 sg13g2_fill_8 FILLER_13_144 ();
 sg13g2_fill_8 FILLER_13_152 ();
 sg13g2_fill_8 FILLER_13_160 ();
 sg13g2_fill_8 FILLER_13_168 ();
 sg13g2_fill_8 FILLER_13_176 ();
 sg13g2_fill_8 FILLER_13_184 ();
 sg13g2_fill_8 FILLER_13_192 ();
 sg13g2_fill_8 FILLER_13_200 ();
 sg13g2_fill_8 FILLER_13_208 ();
 sg13g2_fill_8 FILLER_13_216 ();
 sg13g2_fill_8 FILLER_13_224 ();
 sg13g2_fill_8 FILLER_13_232 ();
 sg13g2_fill_8 FILLER_13_240 ();
 sg13g2_fill_8 FILLER_13_248 ();
 sg13g2_fill_8 FILLER_13_256 ();
 sg13g2_fill_8 FILLER_13_264 ();
 sg13g2_fill_8 FILLER_13_272 ();
 sg13g2_fill_8 FILLER_13_280 ();
 sg13g2_fill_8 FILLER_13_288 ();
 sg13g2_fill_8 FILLER_13_296 ();
 sg13g2_fill_8 FILLER_13_304 ();
 sg13g2_fill_8 FILLER_13_312 ();
 sg13g2_fill_8 FILLER_13_320 ();
 sg13g2_fill_8 FILLER_13_328 ();
 sg13g2_fill_8 FILLER_13_336 ();
 sg13g2_fill_8 FILLER_13_344 ();
 sg13g2_fill_8 FILLER_13_352 ();
 sg13g2_fill_8 FILLER_13_360 ();
 sg13g2_fill_8 FILLER_13_368 ();
 sg13g2_fill_8 FILLER_13_376 ();
 sg13g2_fill_8 FILLER_13_384 ();
 sg13g2_fill_8 FILLER_13_392 ();
 sg13g2_fill_8 FILLER_13_400 ();
 sg13g2_fill_8 FILLER_13_408 ();
 sg13g2_fill_8 FILLER_13_416 ();
 sg13g2_fill_8 FILLER_13_424 ();
 sg13g2_fill_8 FILLER_13_432 ();
 sg13g2_fill_8 FILLER_13_440 ();
 sg13g2_fill_8 FILLER_13_448 ();
 sg13g2_fill_8 FILLER_13_456 ();
 sg13g2_fill_8 FILLER_13_464 ();
 sg13g2_fill_8 FILLER_13_472 ();
 sg13g2_fill_8 FILLER_13_480 ();
 sg13g2_fill_8 FILLER_13_488 ();
 sg13g2_fill_8 FILLER_13_496 ();
 sg13g2_fill_8 FILLER_13_504 ();
 sg13g2_fill_8 FILLER_13_512 ();
 sg13g2_fill_8 FILLER_13_520 ();
 sg13g2_fill_8 FILLER_13_528 ();
 sg13g2_fill_8 FILLER_13_536 ();
 sg13g2_fill_8 FILLER_13_544 ();
 sg13g2_fill_8 FILLER_13_552 ();
 sg13g2_fill_8 FILLER_13_560 ();
 sg13g2_fill_8 FILLER_13_568 ();
 sg13g2_fill_8 FILLER_13_576 ();
 sg13g2_fill_8 FILLER_13_584 ();
 sg13g2_fill_8 FILLER_13_592 ();
 sg13g2_fill_8 FILLER_13_600 ();
 sg13g2_fill_8 FILLER_13_608 ();
 sg13g2_fill_8 FILLER_13_616 ();
 sg13g2_fill_8 FILLER_13_624 ();
 sg13g2_fill_8 FILLER_13_632 ();
 sg13g2_fill_8 FILLER_13_640 ();
 sg13g2_fill_8 FILLER_13_648 ();
 sg13g2_fill_8 FILLER_13_656 ();
 sg13g2_fill_8 FILLER_13_664 ();
 sg13g2_fill_8 FILLER_13_672 ();
 sg13g2_fill_8 FILLER_13_680 ();
 sg13g2_fill_8 FILLER_13_688 ();
 sg13g2_fill_8 FILLER_13_696 ();
 sg13g2_fill_8 FILLER_13_704 ();
 sg13g2_fill_8 FILLER_13_712 ();
 sg13g2_fill_8 FILLER_13_720 ();
 sg13g2_fill_8 FILLER_13_728 ();
 sg13g2_fill_8 FILLER_13_736 ();
 sg13g2_fill_8 FILLER_13_744 ();
 sg13g2_fill_8 FILLER_13_752 ();
 sg13g2_fill_8 FILLER_13_760 ();
 sg13g2_fill_8 FILLER_13_768 ();
 sg13g2_fill_8 FILLER_13_776 ();
 sg13g2_fill_8 FILLER_13_784 ();
 sg13g2_fill_8 FILLER_13_792 ();
 sg13g2_fill_8 FILLER_13_800 ();
 sg13g2_fill_8 FILLER_13_808 ();
 sg13g2_fill_8 FILLER_13_816 ();
 sg13g2_fill_8 FILLER_13_824 ();
 sg13g2_fill_8 FILLER_13_832 ();
 sg13g2_fill_8 FILLER_13_840 ();
 sg13g2_fill_8 FILLER_13_848 ();
 sg13g2_fill_8 FILLER_13_856 ();
 sg13g2_fill_8 FILLER_13_864 ();
 sg13g2_fill_8 FILLER_13_872 ();
 sg13g2_fill_8 FILLER_13_880 ();
 sg13g2_fill_8 FILLER_13_888 ();
 sg13g2_fill_8 FILLER_13_896 ();
 sg13g2_fill_8 FILLER_13_904 ();
 sg13g2_fill_8 FILLER_13_912 ();
 sg13g2_fill_8 FILLER_13_920 ();
 sg13g2_fill_8 FILLER_13_928 ();
 sg13g2_fill_8 FILLER_13_936 ();
 sg13g2_fill_8 FILLER_13_944 ();
 sg13g2_fill_8 FILLER_13_952 ();
 sg13g2_fill_8 FILLER_13_960 ();
 sg13g2_fill_8 FILLER_13_968 ();
 sg13g2_fill_8 FILLER_13_976 ();
 sg13g2_fill_8 FILLER_13_984 ();
 sg13g2_fill_8 FILLER_13_992 ();
 sg13g2_fill_8 FILLER_13_1000 ();
 sg13g2_fill_8 FILLER_13_1008 ();
 sg13g2_fill_8 FILLER_13_1016 ();
 sg13g2_fill_8 FILLER_13_1024 ();
 sg13g2_fill_8 FILLER_13_1032 ();
 sg13g2_fill_8 FILLER_13_1040 ();
 sg13g2_fill_8 FILLER_13_1048 ();
 sg13g2_fill_8 FILLER_13_1056 ();
 sg13g2_fill_8 FILLER_13_1064 ();
 sg13g2_fill_8 FILLER_13_1072 ();
 sg13g2_fill_8 FILLER_13_1080 ();
 sg13g2_fill_8 FILLER_13_1088 ();
 sg13g2_fill_8 FILLER_13_1096 ();
 sg13g2_fill_8 FILLER_13_1104 ();
 sg13g2_fill_8 FILLER_13_1112 ();
 sg13g2_fill_8 FILLER_13_1120 ();
 sg13g2_fill_8 FILLER_13_1128 ();
 sg13g2_fill_8 FILLER_13_1136 ();
 sg13g2_fill_8 FILLER_14_0 ();
 sg13g2_fill_8 FILLER_14_8 ();
 sg13g2_fill_8 FILLER_14_16 ();
 sg13g2_fill_8 FILLER_14_24 ();
 sg13g2_fill_8 FILLER_14_32 ();
 sg13g2_fill_8 FILLER_14_40 ();
 sg13g2_fill_8 FILLER_14_48 ();
 sg13g2_fill_8 FILLER_14_56 ();
 sg13g2_fill_8 FILLER_14_64 ();
 sg13g2_fill_8 FILLER_14_72 ();
 sg13g2_fill_8 FILLER_14_80 ();
 sg13g2_fill_8 FILLER_14_88 ();
 sg13g2_fill_8 FILLER_14_96 ();
 sg13g2_fill_8 FILLER_14_104 ();
 sg13g2_fill_8 FILLER_14_112 ();
 sg13g2_fill_8 FILLER_14_120 ();
 sg13g2_fill_8 FILLER_14_128 ();
 sg13g2_fill_8 FILLER_14_136 ();
 sg13g2_fill_8 FILLER_14_144 ();
 sg13g2_fill_8 FILLER_14_152 ();
 sg13g2_fill_8 FILLER_14_160 ();
 sg13g2_fill_8 FILLER_14_168 ();
 sg13g2_fill_8 FILLER_14_176 ();
 sg13g2_fill_8 FILLER_14_184 ();
 sg13g2_fill_8 FILLER_14_192 ();
 sg13g2_fill_8 FILLER_14_200 ();
 sg13g2_fill_8 FILLER_14_208 ();
 sg13g2_fill_8 FILLER_14_216 ();
 sg13g2_fill_8 FILLER_14_224 ();
 sg13g2_fill_8 FILLER_14_232 ();
 sg13g2_fill_8 FILLER_14_240 ();
 sg13g2_fill_8 FILLER_14_248 ();
 sg13g2_fill_8 FILLER_14_256 ();
 sg13g2_fill_8 FILLER_14_264 ();
 sg13g2_fill_8 FILLER_14_272 ();
 sg13g2_fill_8 FILLER_14_280 ();
 sg13g2_fill_8 FILLER_14_288 ();
 sg13g2_fill_8 FILLER_14_296 ();
 sg13g2_fill_8 FILLER_14_304 ();
 sg13g2_fill_8 FILLER_14_312 ();
 sg13g2_fill_8 FILLER_14_320 ();
 sg13g2_fill_8 FILLER_14_328 ();
 sg13g2_fill_8 FILLER_14_336 ();
 sg13g2_fill_8 FILLER_14_344 ();
 sg13g2_fill_8 FILLER_14_352 ();
 sg13g2_fill_8 FILLER_14_360 ();
 sg13g2_fill_8 FILLER_14_368 ();
 sg13g2_fill_8 FILLER_14_376 ();
 sg13g2_fill_8 FILLER_14_384 ();
 sg13g2_fill_8 FILLER_14_392 ();
 sg13g2_fill_8 FILLER_14_400 ();
 sg13g2_fill_8 FILLER_14_408 ();
 sg13g2_fill_8 FILLER_14_416 ();
 sg13g2_fill_8 FILLER_14_424 ();
 sg13g2_fill_8 FILLER_14_432 ();
 sg13g2_fill_8 FILLER_14_440 ();
 sg13g2_fill_8 FILLER_14_448 ();
 sg13g2_fill_8 FILLER_14_456 ();
 sg13g2_fill_8 FILLER_14_464 ();
 sg13g2_fill_8 FILLER_14_472 ();
 sg13g2_fill_8 FILLER_14_480 ();
 sg13g2_fill_8 FILLER_14_488 ();
 sg13g2_fill_8 FILLER_14_496 ();
 sg13g2_fill_8 FILLER_14_504 ();
 sg13g2_fill_8 FILLER_14_512 ();
 sg13g2_fill_8 FILLER_14_520 ();
 sg13g2_fill_8 FILLER_14_528 ();
 sg13g2_fill_8 FILLER_14_536 ();
 sg13g2_fill_8 FILLER_14_544 ();
 sg13g2_fill_8 FILLER_14_552 ();
 sg13g2_fill_8 FILLER_14_560 ();
 sg13g2_fill_8 FILLER_14_568 ();
 sg13g2_fill_8 FILLER_14_576 ();
 sg13g2_fill_8 FILLER_14_584 ();
 sg13g2_fill_8 FILLER_14_592 ();
 sg13g2_fill_8 FILLER_14_600 ();
 sg13g2_fill_8 FILLER_14_608 ();
 sg13g2_fill_8 FILLER_14_616 ();
 sg13g2_fill_8 FILLER_14_624 ();
 sg13g2_fill_8 FILLER_14_632 ();
 sg13g2_fill_8 FILLER_14_640 ();
 sg13g2_fill_8 FILLER_14_648 ();
 sg13g2_fill_8 FILLER_14_656 ();
 sg13g2_fill_8 FILLER_14_664 ();
 sg13g2_fill_8 FILLER_14_672 ();
 sg13g2_fill_8 FILLER_14_680 ();
 sg13g2_fill_8 FILLER_14_688 ();
 sg13g2_fill_8 FILLER_14_696 ();
 sg13g2_fill_8 FILLER_14_704 ();
 sg13g2_fill_8 FILLER_14_712 ();
 sg13g2_fill_8 FILLER_14_720 ();
 sg13g2_fill_8 FILLER_14_728 ();
 sg13g2_fill_8 FILLER_14_736 ();
 sg13g2_fill_8 FILLER_14_744 ();
 sg13g2_fill_8 FILLER_14_752 ();
 sg13g2_fill_8 FILLER_14_760 ();
 sg13g2_fill_8 FILLER_14_768 ();
 sg13g2_fill_8 FILLER_14_776 ();
 sg13g2_fill_8 FILLER_14_784 ();
 sg13g2_fill_8 FILLER_14_792 ();
 sg13g2_fill_8 FILLER_14_800 ();
 sg13g2_fill_8 FILLER_14_808 ();
 sg13g2_fill_8 FILLER_14_816 ();
 sg13g2_fill_8 FILLER_14_824 ();
 sg13g2_fill_8 FILLER_14_832 ();
 sg13g2_fill_8 FILLER_14_840 ();
 sg13g2_fill_8 FILLER_14_848 ();
 sg13g2_fill_8 FILLER_14_856 ();
 sg13g2_fill_8 FILLER_14_864 ();
 sg13g2_fill_8 FILLER_14_872 ();
 sg13g2_fill_8 FILLER_14_880 ();
 sg13g2_fill_8 FILLER_14_888 ();
 sg13g2_fill_8 FILLER_14_896 ();
 sg13g2_fill_8 FILLER_14_904 ();
 sg13g2_fill_8 FILLER_14_912 ();
 sg13g2_fill_8 FILLER_14_920 ();
 sg13g2_fill_8 FILLER_14_928 ();
 sg13g2_fill_8 FILLER_14_936 ();
 sg13g2_fill_8 FILLER_14_944 ();
 sg13g2_fill_8 FILLER_14_952 ();
 sg13g2_fill_8 FILLER_14_960 ();
 sg13g2_fill_8 FILLER_14_968 ();
 sg13g2_fill_8 FILLER_14_976 ();
 sg13g2_fill_8 FILLER_14_984 ();
 sg13g2_fill_8 FILLER_14_992 ();
 sg13g2_fill_8 FILLER_14_1000 ();
 sg13g2_fill_8 FILLER_14_1008 ();
 sg13g2_fill_8 FILLER_14_1016 ();
 sg13g2_fill_8 FILLER_14_1024 ();
 sg13g2_fill_8 FILLER_14_1032 ();
 sg13g2_fill_8 FILLER_14_1040 ();
 sg13g2_fill_8 FILLER_14_1048 ();
 sg13g2_fill_8 FILLER_14_1056 ();
 sg13g2_fill_8 FILLER_14_1064 ();
 sg13g2_fill_8 FILLER_14_1072 ();
 sg13g2_fill_8 FILLER_14_1080 ();
 sg13g2_fill_8 FILLER_14_1088 ();
 sg13g2_fill_8 FILLER_14_1096 ();
 sg13g2_fill_8 FILLER_14_1104 ();
 sg13g2_fill_8 FILLER_14_1112 ();
 sg13g2_fill_8 FILLER_14_1120 ();
 sg13g2_fill_8 FILLER_14_1128 ();
 sg13g2_fill_8 FILLER_14_1136 ();
 sg13g2_fill_8 FILLER_15_0 ();
 sg13g2_fill_8 FILLER_15_8 ();
 sg13g2_fill_8 FILLER_15_16 ();
 sg13g2_fill_8 FILLER_15_24 ();
 sg13g2_fill_8 FILLER_15_32 ();
 sg13g2_fill_8 FILLER_15_40 ();
 sg13g2_fill_8 FILLER_15_48 ();
 sg13g2_fill_8 FILLER_15_56 ();
 sg13g2_fill_8 FILLER_15_64 ();
 sg13g2_fill_8 FILLER_15_72 ();
 sg13g2_fill_8 FILLER_15_80 ();
 sg13g2_fill_8 FILLER_15_88 ();
 sg13g2_fill_8 FILLER_15_96 ();
 sg13g2_fill_8 FILLER_15_104 ();
 sg13g2_fill_8 FILLER_15_112 ();
 sg13g2_fill_8 FILLER_15_120 ();
 sg13g2_fill_8 FILLER_15_128 ();
 sg13g2_fill_8 FILLER_15_136 ();
 sg13g2_fill_8 FILLER_15_144 ();
 sg13g2_fill_8 FILLER_15_152 ();
 sg13g2_fill_8 FILLER_15_160 ();
 sg13g2_fill_8 FILLER_15_168 ();
 sg13g2_fill_8 FILLER_15_176 ();
 sg13g2_fill_8 FILLER_15_184 ();
 sg13g2_fill_8 FILLER_15_192 ();
 sg13g2_fill_8 FILLER_15_200 ();
 sg13g2_fill_8 FILLER_15_208 ();
 sg13g2_fill_8 FILLER_15_216 ();
 sg13g2_fill_8 FILLER_15_224 ();
 sg13g2_fill_8 FILLER_15_232 ();
 sg13g2_fill_8 FILLER_15_240 ();
 sg13g2_fill_8 FILLER_15_248 ();
 sg13g2_fill_8 FILLER_15_256 ();
 sg13g2_fill_8 FILLER_15_264 ();
 sg13g2_fill_8 FILLER_15_272 ();
 sg13g2_fill_8 FILLER_15_280 ();
 sg13g2_fill_8 FILLER_15_288 ();
 sg13g2_fill_8 FILLER_15_296 ();
 sg13g2_fill_8 FILLER_15_304 ();
 sg13g2_fill_8 FILLER_15_312 ();
 sg13g2_fill_8 FILLER_15_320 ();
 sg13g2_fill_8 FILLER_15_328 ();
 sg13g2_fill_8 FILLER_15_336 ();
 sg13g2_fill_8 FILLER_15_344 ();
 sg13g2_fill_8 FILLER_15_352 ();
 sg13g2_fill_8 FILLER_15_360 ();
 sg13g2_fill_8 FILLER_15_368 ();
 sg13g2_fill_8 FILLER_15_376 ();
 sg13g2_fill_8 FILLER_15_384 ();
 sg13g2_fill_8 FILLER_15_392 ();
 sg13g2_fill_8 FILLER_15_400 ();
 sg13g2_fill_8 FILLER_15_408 ();
 sg13g2_fill_8 FILLER_15_416 ();
 sg13g2_fill_8 FILLER_15_424 ();
 sg13g2_fill_8 FILLER_15_432 ();
 sg13g2_fill_8 FILLER_15_440 ();
 sg13g2_fill_8 FILLER_15_448 ();
 sg13g2_fill_8 FILLER_15_456 ();
 sg13g2_fill_8 FILLER_15_464 ();
 sg13g2_fill_8 FILLER_15_472 ();
 sg13g2_fill_8 FILLER_15_480 ();
 sg13g2_fill_8 FILLER_15_488 ();
 sg13g2_fill_8 FILLER_15_496 ();
 sg13g2_fill_8 FILLER_15_504 ();
 sg13g2_fill_8 FILLER_15_512 ();
 sg13g2_fill_8 FILLER_15_520 ();
 sg13g2_fill_8 FILLER_15_528 ();
 sg13g2_fill_8 FILLER_15_536 ();
 sg13g2_fill_8 FILLER_15_544 ();
 sg13g2_fill_8 FILLER_15_552 ();
 sg13g2_fill_8 FILLER_15_560 ();
 sg13g2_fill_8 FILLER_15_568 ();
 sg13g2_fill_8 FILLER_15_576 ();
 sg13g2_fill_8 FILLER_15_584 ();
 sg13g2_fill_8 FILLER_15_592 ();
 sg13g2_fill_8 FILLER_15_600 ();
 sg13g2_fill_8 FILLER_15_608 ();
 sg13g2_fill_8 FILLER_15_616 ();
 sg13g2_fill_8 FILLER_15_624 ();
 sg13g2_fill_8 FILLER_15_632 ();
 sg13g2_fill_8 FILLER_15_640 ();
 sg13g2_fill_8 FILLER_15_648 ();
 sg13g2_fill_8 FILLER_15_656 ();
 sg13g2_fill_8 FILLER_15_664 ();
 sg13g2_fill_8 FILLER_15_672 ();
 sg13g2_fill_8 FILLER_15_680 ();
 sg13g2_fill_8 FILLER_15_688 ();
 sg13g2_fill_8 FILLER_15_696 ();
 sg13g2_fill_8 FILLER_15_704 ();
 sg13g2_fill_8 FILLER_15_712 ();
 sg13g2_fill_8 FILLER_15_720 ();
 sg13g2_fill_8 FILLER_15_728 ();
 sg13g2_fill_8 FILLER_15_736 ();
 sg13g2_fill_8 FILLER_15_744 ();
 sg13g2_fill_8 FILLER_15_752 ();
 sg13g2_fill_8 FILLER_15_760 ();
 sg13g2_fill_8 FILLER_15_768 ();
 sg13g2_fill_8 FILLER_15_776 ();
 sg13g2_fill_8 FILLER_15_784 ();
 sg13g2_fill_8 FILLER_15_792 ();
 sg13g2_fill_8 FILLER_15_800 ();
 sg13g2_fill_8 FILLER_15_808 ();
 sg13g2_fill_8 FILLER_15_816 ();
 sg13g2_fill_8 FILLER_15_824 ();
 sg13g2_fill_8 FILLER_15_832 ();
 sg13g2_fill_8 FILLER_15_840 ();
 sg13g2_fill_8 FILLER_15_848 ();
 sg13g2_fill_8 FILLER_15_856 ();
 sg13g2_fill_8 FILLER_15_864 ();
 sg13g2_fill_8 FILLER_15_872 ();
 sg13g2_fill_8 FILLER_15_880 ();
 sg13g2_fill_8 FILLER_15_888 ();
 sg13g2_fill_8 FILLER_15_896 ();
 sg13g2_fill_8 FILLER_15_904 ();
 sg13g2_fill_8 FILLER_15_912 ();
 sg13g2_fill_8 FILLER_15_920 ();
 sg13g2_fill_8 FILLER_15_928 ();
 sg13g2_fill_8 FILLER_15_936 ();
 sg13g2_fill_8 FILLER_15_944 ();
 sg13g2_fill_8 FILLER_15_952 ();
 sg13g2_fill_8 FILLER_15_960 ();
 sg13g2_fill_8 FILLER_15_968 ();
 sg13g2_fill_8 FILLER_15_976 ();
 sg13g2_fill_8 FILLER_15_984 ();
 sg13g2_fill_8 FILLER_15_992 ();
 sg13g2_fill_8 FILLER_15_1000 ();
 sg13g2_fill_8 FILLER_15_1008 ();
 sg13g2_fill_8 FILLER_15_1016 ();
 sg13g2_fill_8 FILLER_15_1024 ();
 sg13g2_fill_8 FILLER_15_1032 ();
 sg13g2_fill_8 FILLER_15_1040 ();
 sg13g2_fill_8 FILLER_15_1048 ();
 sg13g2_fill_8 FILLER_15_1056 ();
 sg13g2_fill_8 FILLER_15_1064 ();
 sg13g2_fill_8 FILLER_15_1072 ();
 sg13g2_fill_8 FILLER_15_1080 ();
 sg13g2_fill_8 FILLER_15_1088 ();
 sg13g2_fill_8 FILLER_15_1096 ();
 sg13g2_fill_8 FILLER_15_1104 ();
 sg13g2_fill_8 FILLER_15_1112 ();
 sg13g2_fill_8 FILLER_15_1120 ();
 sg13g2_fill_8 FILLER_15_1128 ();
 sg13g2_fill_8 FILLER_15_1136 ();
 sg13g2_fill_8 FILLER_16_0 ();
 sg13g2_fill_8 FILLER_16_8 ();
 sg13g2_fill_8 FILLER_16_16 ();
 sg13g2_fill_8 FILLER_16_24 ();
 sg13g2_fill_8 FILLER_16_32 ();
 sg13g2_fill_8 FILLER_16_40 ();
 sg13g2_fill_8 FILLER_16_48 ();
 sg13g2_fill_8 FILLER_16_56 ();
 sg13g2_fill_8 FILLER_16_64 ();
 sg13g2_fill_8 FILLER_16_72 ();
 sg13g2_fill_8 FILLER_16_80 ();
 sg13g2_fill_8 FILLER_16_88 ();
 sg13g2_fill_8 FILLER_16_96 ();
 sg13g2_fill_8 FILLER_16_104 ();
 sg13g2_fill_8 FILLER_16_112 ();
 sg13g2_fill_8 FILLER_16_120 ();
 sg13g2_fill_8 FILLER_16_128 ();
 sg13g2_fill_8 FILLER_16_136 ();
 sg13g2_fill_8 FILLER_16_144 ();
 sg13g2_fill_8 FILLER_16_152 ();
 sg13g2_fill_8 FILLER_16_160 ();
 sg13g2_fill_8 FILLER_16_168 ();
 sg13g2_fill_8 FILLER_16_176 ();
 sg13g2_fill_8 FILLER_16_184 ();
 sg13g2_fill_8 FILLER_16_192 ();
 sg13g2_fill_8 FILLER_16_200 ();
 sg13g2_fill_8 FILLER_16_208 ();
 sg13g2_fill_8 FILLER_16_216 ();
 sg13g2_fill_8 FILLER_16_224 ();
 sg13g2_fill_8 FILLER_16_232 ();
 sg13g2_fill_8 FILLER_16_240 ();
 sg13g2_fill_8 FILLER_16_248 ();
 sg13g2_fill_8 FILLER_16_256 ();
 sg13g2_fill_8 FILLER_16_264 ();
 sg13g2_fill_8 FILLER_16_272 ();
 sg13g2_fill_8 FILLER_16_280 ();
 sg13g2_fill_8 FILLER_16_288 ();
 sg13g2_fill_8 FILLER_16_296 ();
 sg13g2_fill_8 FILLER_16_304 ();
 sg13g2_fill_8 FILLER_16_312 ();
 sg13g2_fill_8 FILLER_16_320 ();
 sg13g2_fill_8 FILLER_16_328 ();
 sg13g2_fill_8 FILLER_16_336 ();
 sg13g2_fill_8 FILLER_16_344 ();
 sg13g2_fill_8 FILLER_16_352 ();
 sg13g2_fill_8 FILLER_16_360 ();
 sg13g2_fill_8 FILLER_16_368 ();
 sg13g2_fill_8 FILLER_16_376 ();
 sg13g2_fill_8 FILLER_16_384 ();
 sg13g2_fill_8 FILLER_16_392 ();
 sg13g2_fill_8 FILLER_16_400 ();
 sg13g2_fill_8 FILLER_16_408 ();
 sg13g2_fill_8 FILLER_16_416 ();
 sg13g2_fill_8 FILLER_16_424 ();
 sg13g2_fill_8 FILLER_16_432 ();
 sg13g2_fill_8 FILLER_16_440 ();
 sg13g2_fill_8 FILLER_16_448 ();
 sg13g2_fill_8 FILLER_16_456 ();
 sg13g2_fill_8 FILLER_16_464 ();
 sg13g2_fill_8 FILLER_16_472 ();
 sg13g2_fill_8 FILLER_16_480 ();
 sg13g2_fill_8 FILLER_16_488 ();
 sg13g2_fill_8 FILLER_16_496 ();
 sg13g2_fill_8 FILLER_16_504 ();
 sg13g2_fill_8 FILLER_16_512 ();
 sg13g2_fill_8 FILLER_16_520 ();
 sg13g2_fill_8 FILLER_16_528 ();
 sg13g2_fill_8 FILLER_16_536 ();
 sg13g2_fill_8 FILLER_16_544 ();
 sg13g2_fill_8 FILLER_16_552 ();
 sg13g2_fill_8 FILLER_16_560 ();
 sg13g2_fill_8 FILLER_16_568 ();
 sg13g2_fill_8 FILLER_16_576 ();
 sg13g2_fill_8 FILLER_16_584 ();
 sg13g2_fill_8 FILLER_16_592 ();
 sg13g2_fill_8 FILLER_16_600 ();
 sg13g2_fill_8 FILLER_16_608 ();
 sg13g2_fill_8 FILLER_16_616 ();
 sg13g2_fill_8 FILLER_16_624 ();
 sg13g2_fill_8 FILLER_16_632 ();
 sg13g2_fill_8 FILLER_16_640 ();
 sg13g2_fill_8 FILLER_16_648 ();
 sg13g2_fill_8 FILLER_16_656 ();
 sg13g2_fill_8 FILLER_16_664 ();
 sg13g2_fill_8 FILLER_16_672 ();
 sg13g2_fill_8 FILLER_16_680 ();
 sg13g2_fill_8 FILLER_16_688 ();
 sg13g2_fill_8 FILLER_16_696 ();
 sg13g2_fill_8 FILLER_16_704 ();
 sg13g2_fill_8 FILLER_16_712 ();
 sg13g2_fill_8 FILLER_16_720 ();
 sg13g2_fill_8 FILLER_16_728 ();
 sg13g2_fill_8 FILLER_16_736 ();
 sg13g2_fill_8 FILLER_16_744 ();
 sg13g2_fill_8 FILLER_16_752 ();
 sg13g2_fill_8 FILLER_16_760 ();
 sg13g2_fill_8 FILLER_16_768 ();
 sg13g2_fill_8 FILLER_16_776 ();
 sg13g2_fill_8 FILLER_16_784 ();
 sg13g2_fill_8 FILLER_16_792 ();
 sg13g2_fill_8 FILLER_16_800 ();
 sg13g2_fill_8 FILLER_16_808 ();
 sg13g2_fill_8 FILLER_16_816 ();
 sg13g2_fill_8 FILLER_16_824 ();
 sg13g2_fill_8 FILLER_16_832 ();
 sg13g2_fill_8 FILLER_16_840 ();
 sg13g2_fill_8 FILLER_16_848 ();
 sg13g2_fill_8 FILLER_16_856 ();
 sg13g2_fill_8 FILLER_16_864 ();
 sg13g2_fill_8 FILLER_16_872 ();
 sg13g2_fill_8 FILLER_16_880 ();
 sg13g2_fill_8 FILLER_16_888 ();
 sg13g2_fill_8 FILLER_16_896 ();
 sg13g2_fill_8 FILLER_16_904 ();
 sg13g2_fill_8 FILLER_16_912 ();
 sg13g2_fill_8 FILLER_16_920 ();
 sg13g2_fill_8 FILLER_16_928 ();
 sg13g2_fill_8 FILLER_16_936 ();
 sg13g2_fill_8 FILLER_16_944 ();
 sg13g2_fill_8 FILLER_16_952 ();
 sg13g2_fill_8 FILLER_16_960 ();
 sg13g2_fill_8 FILLER_16_968 ();
 sg13g2_fill_8 FILLER_16_976 ();
 sg13g2_fill_8 FILLER_16_984 ();
 sg13g2_fill_8 FILLER_16_992 ();
 sg13g2_fill_8 FILLER_16_1000 ();
 sg13g2_fill_8 FILLER_16_1008 ();
 sg13g2_fill_8 FILLER_16_1016 ();
 sg13g2_fill_8 FILLER_16_1024 ();
 sg13g2_fill_8 FILLER_16_1032 ();
 sg13g2_fill_8 FILLER_16_1040 ();
 sg13g2_fill_8 FILLER_16_1048 ();
 sg13g2_fill_8 FILLER_16_1056 ();
 sg13g2_fill_8 FILLER_16_1064 ();
 sg13g2_fill_8 FILLER_16_1072 ();
 sg13g2_fill_8 FILLER_16_1080 ();
 sg13g2_fill_8 FILLER_16_1088 ();
 sg13g2_fill_8 FILLER_16_1096 ();
 sg13g2_fill_8 FILLER_16_1104 ();
 sg13g2_fill_8 FILLER_16_1112 ();
 sg13g2_fill_8 FILLER_16_1120 ();
 sg13g2_fill_8 FILLER_16_1128 ();
 sg13g2_fill_8 FILLER_16_1136 ();
 sg13g2_fill_8 FILLER_17_0 ();
 sg13g2_fill_8 FILLER_17_8 ();
 sg13g2_fill_8 FILLER_17_16 ();
 sg13g2_fill_8 FILLER_17_24 ();
 sg13g2_fill_8 FILLER_17_32 ();
 sg13g2_fill_8 FILLER_17_40 ();
 sg13g2_fill_8 FILLER_17_48 ();
 sg13g2_fill_8 FILLER_17_56 ();
 sg13g2_fill_8 FILLER_17_64 ();
 sg13g2_fill_8 FILLER_17_72 ();
 sg13g2_fill_8 FILLER_17_80 ();
 sg13g2_fill_8 FILLER_17_88 ();
 sg13g2_fill_8 FILLER_17_96 ();
 sg13g2_fill_8 FILLER_17_104 ();
 sg13g2_fill_8 FILLER_17_112 ();
 sg13g2_fill_8 FILLER_17_120 ();
 sg13g2_fill_8 FILLER_17_128 ();
 sg13g2_fill_8 FILLER_17_136 ();
 sg13g2_fill_8 FILLER_17_144 ();
 sg13g2_fill_8 FILLER_17_152 ();
 sg13g2_fill_8 FILLER_17_160 ();
 sg13g2_fill_8 FILLER_17_168 ();
 sg13g2_fill_8 FILLER_17_176 ();
 sg13g2_fill_8 FILLER_17_184 ();
 sg13g2_fill_8 FILLER_17_192 ();
 sg13g2_fill_8 FILLER_17_200 ();
 sg13g2_fill_8 FILLER_17_208 ();
 sg13g2_fill_8 FILLER_17_216 ();
 sg13g2_fill_8 FILLER_17_224 ();
 sg13g2_fill_8 FILLER_17_232 ();
 sg13g2_fill_8 FILLER_17_240 ();
 sg13g2_fill_8 FILLER_17_248 ();
 sg13g2_fill_8 FILLER_17_256 ();
 sg13g2_fill_8 FILLER_17_264 ();
 sg13g2_fill_8 FILLER_17_272 ();
 sg13g2_fill_8 FILLER_17_280 ();
 sg13g2_fill_8 FILLER_17_288 ();
 sg13g2_fill_8 FILLER_17_296 ();
 sg13g2_fill_8 FILLER_17_304 ();
 sg13g2_fill_8 FILLER_17_312 ();
 sg13g2_fill_8 FILLER_17_320 ();
 sg13g2_fill_8 FILLER_17_328 ();
 sg13g2_fill_8 FILLER_17_336 ();
 sg13g2_fill_8 FILLER_17_344 ();
 sg13g2_fill_8 FILLER_17_352 ();
 sg13g2_fill_8 FILLER_17_360 ();
 sg13g2_fill_8 FILLER_17_368 ();
 sg13g2_fill_8 FILLER_17_376 ();
 sg13g2_fill_8 FILLER_17_384 ();
 sg13g2_fill_8 FILLER_17_392 ();
 sg13g2_fill_8 FILLER_17_400 ();
 sg13g2_fill_8 FILLER_17_408 ();
 sg13g2_fill_8 FILLER_17_416 ();
 sg13g2_fill_8 FILLER_17_424 ();
 sg13g2_fill_8 FILLER_17_432 ();
 sg13g2_fill_8 FILLER_17_440 ();
 sg13g2_fill_8 FILLER_17_448 ();
 sg13g2_fill_8 FILLER_17_456 ();
 sg13g2_fill_8 FILLER_17_464 ();
 sg13g2_fill_8 FILLER_17_472 ();
 sg13g2_fill_8 FILLER_17_480 ();
 sg13g2_fill_8 FILLER_17_488 ();
 sg13g2_fill_8 FILLER_17_496 ();
 sg13g2_fill_8 FILLER_17_504 ();
 sg13g2_fill_8 FILLER_17_512 ();
 sg13g2_fill_8 FILLER_17_520 ();
 sg13g2_fill_8 FILLER_17_528 ();
 sg13g2_fill_8 FILLER_17_536 ();
 sg13g2_fill_8 FILLER_17_544 ();
 sg13g2_fill_8 FILLER_17_552 ();
 sg13g2_fill_8 FILLER_17_560 ();
 sg13g2_fill_8 FILLER_17_568 ();
 sg13g2_fill_8 FILLER_17_576 ();
 sg13g2_fill_8 FILLER_17_584 ();
 sg13g2_fill_8 FILLER_17_592 ();
 sg13g2_fill_8 FILLER_17_600 ();
 sg13g2_fill_8 FILLER_17_608 ();
 sg13g2_fill_8 FILLER_17_616 ();
 sg13g2_fill_8 FILLER_17_624 ();
 sg13g2_fill_8 FILLER_17_632 ();
 sg13g2_fill_8 FILLER_17_640 ();
 sg13g2_fill_8 FILLER_17_648 ();
 sg13g2_fill_8 FILLER_17_656 ();
 sg13g2_fill_8 FILLER_17_664 ();
 sg13g2_fill_8 FILLER_17_672 ();
 sg13g2_fill_8 FILLER_17_680 ();
 sg13g2_fill_8 FILLER_17_688 ();
 sg13g2_fill_8 FILLER_17_696 ();
 sg13g2_fill_8 FILLER_17_704 ();
 sg13g2_fill_8 FILLER_17_712 ();
 sg13g2_fill_8 FILLER_17_720 ();
 sg13g2_fill_8 FILLER_17_728 ();
 sg13g2_fill_8 FILLER_17_736 ();
 sg13g2_fill_8 FILLER_17_744 ();
 sg13g2_fill_8 FILLER_17_752 ();
 sg13g2_fill_8 FILLER_17_760 ();
 sg13g2_fill_8 FILLER_17_768 ();
 sg13g2_fill_8 FILLER_17_776 ();
 sg13g2_fill_8 FILLER_17_784 ();
 sg13g2_fill_8 FILLER_17_792 ();
 sg13g2_fill_8 FILLER_17_800 ();
 sg13g2_fill_8 FILLER_17_808 ();
 sg13g2_fill_8 FILLER_17_816 ();
 sg13g2_fill_8 FILLER_17_824 ();
 sg13g2_fill_8 FILLER_17_832 ();
 sg13g2_fill_8 FILLER_17_840 ();
 sg13g2_fill_8 FILLER_17_848 ();
 sg13g2_fill_8 FILLER_17_856 ();
 sg13g2_fill_8 FILLER_17_864 ();
 sg13g2_fill_8 FILLER_17_872 ();
 sg13g2_fill_8 FILLER_17_880 ();
 sg13g2_fill_8 FILLER_17_888 ();
 sg13g2_fill_8 FILLER_17_896 ();
 sg13g2_fill_8 FILLER_17_904 ();
 sg13g2_fill_8 FILLER_17_912 ();
 sg13g2_fill_8 FILLER_17_920 ();
 sg13g2_fill_8 FILLER_17_928 ();
 sg13g2_fill_8 FILLER_17_936 ();
 sg13g2_fill_8 FILLER_17_944 ();
 sg13g2_fill_8 FILLER_17_952 ();
 sg13g2_fill_8 FILLER_17_960 ();
 sg13g2_fill_8 FILLER_17_968 ();
 sg13g2_fill_8 FILLER_17_976 ();
 sg13g2_fill_8 FILLER_17_984 ();
 sg13g2_fill_8 FILLER_17_992 ();
 sg13g2_fill_8 FILLER_17_1000 ();
 sg13g2_fill_8 FILLER_17_1008 ();
 sg13g2_fill_8 FILLER_17_1016 ();
 sg13g2_fill_8 FILLER_17_1024 ();
 sg13g2_fill_8 FILLER_17_1032 ();
 sg13g2_fill_8 FILLER_17_1040 ();
 sg13g2_fill_8 FILLER_17_1048 ();
 sg13g2_fill_8 FILLER_17_1056 ();
 sg13g2_fill_8 FILLER_17_1064 ();
 sg13g2_fill_8 FILLER_17_1072 ();
 sg13g2_fill_8 FILLER_17_1080 ();
 sg13g2_fill_8 FILLER_17_1088 ();
 sg13g2_fill_8 FILLER_17_1096 ();
 sg13g2_fill_8 FILLER_17_1104 ();
 sg13g2_fill_8 FILLER_17_1112 ();
 sg13g2_fill_8 FILLER_17_1120 ();
 sg13g2_fill_8 FILLER_17_1128 ();
 sg13g2_fill_8 FILLER_17_1136 ();
 sg13g2_fill_8 FILLER_18_0 ();
 sg13g2_fill_8 FILLER_18_8 ();
 sg13g2_fill_8 FILLER_18_16 ();
 sg13g2_fill_8 FILLER_18_24 ();
 sg13g2_fill_8 FILLER_18_32 ();
 sg13g2_fill_8 FILLER_18_40 ();
 sg13g2_fill_8 FILLER_18_48 ();
 sg13g2_fill_8 FILLER_18_56 ();
 sg13g2_fill_8 FILLER_18_64 ();
 sg13g2_fill_8 FILLER_18_72 ();
 sg13g2_fill_8 FILLER_18_80 ();
 sg13g2_fill_8 FILLER_18_88 ();
 sg13g2_fill_8 FILLER_18_96 ();
 sg13g2_fill_8 FILLER_18_104 ();
 sg13g2_fill_8 FILLER_18_112 ();
 sg13g2_fill_8 FILLER_18_120 ();
 sg13g2_fill_8 FILLER_18_128 ();
 sg13g2_fill_8 FILLER_18_136 ();
 sg13g2_fill_8 FILLER_18_144 ();
 sg13g2_fill_8 FILLER_18_152 ();
 sg13g2_fill_8 FILLER_18_160 ();
 sg13g2_fill_8 FILLER_18_168 ();
 sg13g2_fill_8 FILLER_18_176 ();
 sg13g2_fill_8 FILLER_18_184 ();
 sg13g2_fill_8 FILLER_18_192 ();
 sg13g2_fill_8 FILLER_18_200 ();
 sg13g2_fill_8 FILLER_18_208 ();
 sg13g2_fill_8 FILLER_18_216 ();
 sg13g2_fill_8 FILLER_18_224 ();
 sg13g2_fill_8 FILLER_18_232 ();
 sg13g2_fill_8 FILLER_18_240 ();
 sg13g2_fill_8 FILLER_18_248 ();
 sg13g2_fill_8 FILLER_18_256 ();
 sg13g2_fill_8 FILLER_18_264 ();
 sg13g2_fill_8 FILLER_18_272 ();
 sg13g2_fill_8 FILLER_18_280 ();
 sg13g2_fill_8 FILLER_18_288 ();
 sg13g2_fill_8 FILLER_18_296 ();
 sg13g2_fill_8 FILLER_18_304 ();
 sg13g2_fill_8 FILLER_18_312 ();
 sg13g2_fill_8 FILLER_18_320 ();
 sg13g2_fill_8 FILLER_18_328 ();
 sg13g2_fill_8 FILLER_18_336 ();
 sg13g2_fill_8 FILLER_18_344 ();
 sg13g2_fill_8 FILLER_18_352 ();
 sg13g2_fill_8 FILLER_18_360 ();
 sg13g2_fill_8 FILLER_18_368 ();
 sg13g2_fill_8 FILLER_18_376 ();
 sg13g2_fill_8 FILLER_18_384 ();
 sg13g2_fill_8 FILLER_18_392 ();
 sg13g2_fill_8 FILLER_18_400 ();
 sg13g2_fill_8 FILLER_18_408 ();
 sg13g2_fill_8 FILLER_18_416 ();
 sg13g2_fill_8 FILLER_18_424 ();
 sg13g2_fill_8 FILLER_18_432 ();
 sg13g2_fill_8 FILLER_18_440 ();
 sg13g2_fill_8 FILLER_18_448 ();
 sg13g2_fill_8 FILLER_18_456 ();
 sg13g2_fill_8 FILLER_18_464 ();
 sg13g2_fill_8 FILLER_18_472 ();
 sg13g2_fill_8 FILLER_18_480 ();
 sg13g2_fill_8 FILLER_18_488 ();
 sg13g2_fill_8 FILLER_18_496 ();
 sg13g2_fill_8 FILLER_18_504 ();
 sg13g2_fill_8 FILLER_18_512 ();
 sg13g2_fill_8 FILLER_18_520 ();
 sg13g2_fill_8 FILLER_18_528 ();
 sg13g2_fill_8 FILLER_18_536 ();
 sg13g2_fill_8 FILLER_18_544 ();
 sg13g2_fill_8 FILLER_18_552 ();
 sg13g2_fill_8 FILLER_18_560 ();
 sg13g2_fill_8 FILLER_18_568 ();
 sg13g2_fill_8 FILLER_18_576 ();
 sg13g2_fill_8 FILLER_18_584 ();
 sg13g2_fill_8 FILLER_18_592 ();
 sg13g2_fill_8 FILLER_18_600 ();
 sg13g2_fill_8 FILLER_18_608 ();
 sg13g2_fill_8 FILLER_18_616 ();
 sg13g2_fill_8 FILLER_18_624 ();
 sg13g2_fill_8 FILLER_18_632 ();
 sg13g2_fill_8 FILLER_18_640 ();
 sg13g2_fill_8 FILLER_18_648 ();
 sg13g2_fill_8 FILLER_18_656 ();
 sg13g2_fill_8 FILLER_18_664 ();
 sg13g2_fill_8 FILLER_18_672 ();
 sg13g2_fill_8 FILLER_18_680 ();
 sg13g2_fill_8 FILLER_18_688 ();
 sg13g2_fill_8 FILLER_18_696 ();
 sg13g2_fill_8 FILLER_18_704 ();
 sg13g2_fill_8 FILLER_18_712 ();
 sg13g2_fill_8 FILLER_18_720 ();
 sg13g2_fill_8 FILLER_18_728 ();
 sg13g2_fill_8 FILLER_18_736 ();
 sg13g2_fill_8 FILLER_18_744 ();
 sg13g2_fill_8 FILLER_18_752 ();
 sg13g2_fill_8 FILLER_18_760 ();
 sg13g2_fill_8 FILLER_18_768 ();
 sg13g2_fill_8 FILLER_18_776 ();
 sg13g2_fill_8 FILLER_18_784 ();
 sg13g2_fill_8 FILLER_18_792 ();
 sg13g2_fill_8 FILLER_18_800 ();
 sg13g2_fill_8 FILLER_18_808 ();
 sg13g2_fill_8 FILLER_18_816 ();
 sg13g2_fill_8 FILLER_18_824 ();
 sg13g2_fill_8 FILLER_18_832 ();
 sg13g2_fill_8 FILLER_18_840 ();
 sg13g2_fill_8 FILLER_18_848 ();
 sg13g2_fill_8 FILLER_18_856 ();
 sg13g2_fill_8 FILLER_18_864 ();
 sg13g2_fill_8 FILLER_18_872 ();
 sg13g2_fill_8 FILLER_18_880 ();
 sg13g2_fill_8 FILLER_18_888 ();
 sg13g2_fill_8 FILLER_18_896 ();
 sg13g2_fill_8 FILLER_18_904 ();
 sg13g2_fill_8 FILLER_18_912 ();
 sg13g2_fill_8 FILLER_18_920 ();
 sg13g2_fill_8 FILLER_18_928 ();
 sg13g2_fill_8 FILLER_18_936 ();
 sg13g2_fill_8 FILLER_18_944 ();
 sg13g2_fill_8 FILLER_18_952 ();
 sg13g2_fill_8 FILLER_18_960 ();
 sg13g2_fill_8 FILLER_18_968 ();
 sg13g2_fill_8 FILLER_18_976 ();
 sg13g2_fill_8 FILLER_18_984 ();
 sg13g2_fill_8 FILLER_18_992 ();
 sg13g2_fill_8 FILLER_18_1000 ();
 sg13g2_fill_8 FILLER_18_1008 ();
 sg13g2_fill_8 FILLER_18_1016 ();
 sg13g2_fill_8 FILLER_18_1024 ();
 sg13g2_fill_8 FILLER_18_1032 ();
 sg13g2_fill_8 FILLER_18_1040 ();
 sg13g2_fill_8 FILLER_18_1048 ();
 sg13g2_fill_8 FILLER_18_1056 ();
 sg13g2_fill_8 FILLER_18_1064 ();
 sg13g2_fill_8 FILLER_18_1072 ();
 sg13g2_fill_8 FILLER_18_1080 ();
 sg13g2_fill_8 FILLER_18_1088 ();
 sg13g2_fill_8 FILLER_18_1096 ();
 sg13g2_fill_8 FILLER_18_1104 ();
 sg13g2_fill_8 FILLER_18_1112 ();
 sg13g2_fill_8 FILLER_18_1120 ();
 sg13g2_fill_8 FILLER_18_1128 ();
 sg13g2_fill_8 FILLER_18_1136 ();
 sg13g2_fill_8 FILLER_19_0 ();
 sg13g2_fill_8 FILLER_19_8 ();
 sg13g2_fill_8 FILLER_19_16 ();
 sg13g2_fill_8 FILLER_19_24 ();
 sg13g2_fill_8 FILLER_19_32 ();
 sg13g2_fill_8 FILLER_19_40 ();
 sg13g2_fill_8 FILLER_19_48 ();
 sg13g2_fill_8 FILLER_19_56 ();
 sg13g2_fill_8 FILLER_19_64 ();
 sg13g2_fill_8 FILLER_19_72 ();
 sg13g2_fill_8 FILLER_19_80 ();
 sg13g2_fill_8 FILLER_19_88 ();
 sg13g2_fill_8 FILLER_19_96 ();
 sg13g2_fill_8 FILLER_19_104 ();
 sg13g2_fill_8 FILLER_19_112 ();
 sg13g2_fill_8 FILLER_19_120 ();
 sg13g2_fill_8 FILLER_19_128 ();
 sg13g2_fill_8 FILLER_19_136 ();
 sg13g2_fill_8 FILLER_19_144 ();
 sg13g2_fill_8 FILLER_19_152 ();
 sg13g2_fill_8 FILLER_19_160 ();
 sg13g2_fill_8 FILLER_19_168 ();
 sg13g2_fill_8 FILLER_19_176 ();
 sg13g2_fill_8 FILLER_19_184 ();
 sg13g2_fill_8 FILLER_19_192 ();
 sg13g2_fill_8 FILLER_19_200 ();
 sg13g2_fill_8 FILLER_19_208 ();
 sg13g2_fill_8 FILLER_19_216 ();
 sg13g2_fill_8 FILLER_19_224 ();
 sg13g2_fill_8 FILLER_19_232 ();
 sg13g2_fill_8 FILLER_19_240 ();
 sg13g2_fill_8 FILLER_19_248 ();
 sg13g2_fill_8 FILLER_19_256 ();
 sg13g2_fill_8 FILLER_19_264 ();
 sg13g2_fill_8 FILLER_19_272 ();
 sg13g2_fill_8 FILLER_19_280 ();
 sg13g2_fill_8 FILLER_19_288 ();
 sg13g2_fill_8 FILLER_19_296 ();
 sg13g2_fill_8 FILLER_19_304 ();
 sg13g2_fill_8 FILLER_19_312 ();
 sg13g2_fill_8 FILLER_19_320 ();
 sg13g2_fill_8 FILLER_19_328 ();
 sg13g2_fill_8 FILLER_19_336 ();
 sg13g2_fill_8 FILLER_19_344 ();
 sg13g2_fill_8 FILLER_19_352 ();
 sg13g2_fill_8 FILLER_19_360 ();
 sg13g2_fill_8 FILLER_19_368 ();
 sg13g2_fill_8 FILLER_19_376 ();
 sg13g2_fill_8 FILLER_19_384 ();
 sg13g2_fill_8 FILLER_19_392 ();
 sg13g2_fill_8 FILLER_19_400 ();
 sg13g2_fill_8 FILLER_19_408 ();
 sg13g2_fill_8 FILLER_19_416 ();
 sg13g2_fill_8 FILLER_19_424 ();
 sg13g2_fill_8 FILLER_19_432 ();
 sg13g2_fill_8 FILLER_19_440 ();
 sg13g2_fill_8 FILLER_19_448 ();
 sg13g2_fill_8 FILLER_19_456 ();
 sg13g2_fill_8 FILLER_19_464 ();
 sg13g2_fill_8 FILLER_19_472 ();
 sg13g2_fill_8 FILLER_19_480 ();
 sg13g2_fill_8 FILLER_19_488 ();
 sg13g2_fill_8 FILLER_19_496 ();
 sg13g2_fill_8 FILLER_19_504 ();
 sg13g2_fill_8 FILLER_19_512 ();
 sg13g2_fill_8 FILLER_19_520 ();
 sg13g2_fill_8 FILLER_19_528 ();
 sg13g2_fill_8 FILLER_19_536 ();
 sg13g2_fill_8 FILLER_19_544 ();
 sg13g2_fill_8 FILLER_19_552 ();
 sg13g2_fill_8 FILLER_19_560 ();
 sg13g2_fill_8 FILLER_19_568 ();
 sg13g2_fill_8 FILLER_19_576 ();
 sg13g2_fill_8 FILLER_19_584 ();
 sg13g2_fill_8 FILLER_19_592 ();
 sg13g2_fill_8 FILLER_19_600 ();
 sg13g2_fill_8 FILLER_19_608 ();
 sg13g2_fill_8 FILLER_19_616 ();
 sg13g2_fill_8 FILLER_19_624 ();
 sg13g2_fill_8 FILLER_19_632 ();
 sg13g2_fill_8 FILLER_19_640 ();
 sg13g2_fill_8 FILLER_19_648 ();
 sg13g2_fill_8 FILLER_19_656 ();
 sg13g2_fill_8 FILLER_19_664 ();
 sg13g2_fill_8 FILLER_19_672 ();
 sg13g2_fill_8 FILLER_19_680 ();
 sg13g2_fill_8 FILLER_19_688 ();
 sg13g2_fill_8 FILLER_19_696 ();
 sg13g2_fill_8 FILLER_19_704 ();
 sg13g2_fill_8 FILLER_19_712 ();
 sg13g2_fill_8 FILLER_19_720 ();
 sg13g2_fill_8 FILLER_19_728 ();
 sg13g2_fill_8 FILLER_19_736 ();
 sg13g2_fill_8 FILLER_19_744 ();
 sg13g2_fill_8 FILLER_19_752 ();
 sg13g2_fill_8 FILLER_19_760 ();
 sg13g2_fill_8 FILLER_19_768 ();
 sg13g2_fill_8 FILLER_19_776 ();
 sg13g2_fill_8 FILLER_19_784 ();
 sg13g2_fill_8 FILLER_19_792 ();
 sg13g2_fill_8 FILLER_19_800 ();
 sg13g2_fill_8 FILLER_19_808 ();
 sg13g2_fill_8 FILLER_19_816 ();
 sg13g2_fill_8 FILLER_19_824 ();
 sg13g2_fill_8 FILLER_19_832 ();
 sg13g2_fill_8 FILLER_19_840 ();
 sg13g2_fill_8 FILLER_19_848 ();
 sg13g2_fill_8 FILLER_19_856 ();
 sg13g2_fill_8 FILLER_19_864 ();
 sg13g2_fill_8 FILLER_19_872 ();
 sg13g2_fill_8 FILLER_19_880 ();
 sg13g2_fill_8 FILLER_19_888 ();
 sg13g2_fill_8 FILLER_19_896 ();
 sg13g2_fill_8 FILLER_19_904 ();
 sg13g2_fill_8 FILLER_19_912 ();
 sg13g2_fill_8 FILLER_19_920 ();
 sg13g2_fill_8 FILLER_19_928 ();
 sg13g2_fill_8 FILLER_19_936 ();
 sg13g2_fill_8 FILLER_19_944 ();
 sg13g2_fill_8 FILLER_19_952 ();
 sg13g2_fill_8 FILLER_19_960 ();
 sg13g2_fill_8 FILLER_19_968 ();
 sg13g2_fill_8 FILLER_19_976 ();
 sg13g2_fill_8 FILLER_19_984 ();
 sg13g2_fill_8 FILLER_19_992 ();
 sg13g2_fill_8 FILLER_19_1000 ();
 sg13g2_fill_8 FILLER_19_1008 ();
 sg13g2_fill_8 FILLER_19_1016 ();
 sg13g2_fill_8 FILLER_19_1024 ();
 sg13g2_fill_8 FILLER_19_1032 ();
 sg13g2_fill_8 FILLER_19_1040 ();
 sg13g2_fill_8 FILLER_19_1048 ();
 sg13g2_fill_8 FILLER_19_1056 ();
 sg13g2_fill_8 FILLER_19_1064 ();
 sg13g2_fill_8 FILLER_19_1072 ();
 sg13g2_fill_8 FILLER_19_1080 ();
 sg13g2_fill_8 FILLER_19_1088 ();
 sg13g2_fill_8 FILLER_19_1096 ();
 sg13g2_fill_8 FILLER_19_1104 ();
 sg13g2_fill_8 FILLER_19_1112 ();
 sg13g2_fill_8 FILLER_19_1120 ();
 sg13g2_fill_8 FILLER_19_1128 ();
 sg13g2_fill_8 FILLER_19_1136 ();
 sg13g2_fill_8 FILLER_20_0 ();
 sg13g2_fill_8 FILLER_20_8 ();
 sg13g2_fill_8 FILLER_20_16 ();
 sg13g2_fill_8 FILLER_20_24 ();
 sg13g2_fill_8 FILLER_20_32 ();
 sg13g2_fill_8 FILLER_20_40 ();
 sg13g2_fill_8 FILLER_20_48 ();
 sg13g2_fill_8 FILLER_20_56 ();
 sg13g2_fill_8 FILLER_20_64 ();
 sg13g2_fill_8 FILLER_20_72 ();
 sg13g2_fill_8 FILLER_20_80 ();
 sg13g2_fill_8 FILLER_20_88 ();
 sg13g2_fill_8 FILLER_20_96 ();
 sg13g2_fill_8 FILLER_20_104 ();
 sg13g2_fill_8 FILLER_20_112 ();
 sg13g2_fill_8 FILLER_20_120 ();
 sg13g2_fill_8 FILLER_20_128 ();
 sg13g2_fill_8 FILLER_20_136 ();
 sg13g2_fill_8 FILLER_20_144 ();
 sg13g2_fill_8 FILLER_20_152 ();
 sg13g2_fill_8 FILLER_20_160 ();
 sg13g2_fill_8 FILLER_20_168 ();
 sg13g2_fill_8 FILLER_20_176 ();
 sg13g2_fill_8 FILLER_20_184 ();
 sg13g2_fill_8 FILLER_20_192 ();
 sg13g2_fill_8 FILLER_20_200 ();
 sg13g2_fill_8 FILLER_20_208 ();
 sg13g2_fill_8 FILLER_20_216 ();
 sg13g2_fill_8 FILLER_20_224 ();
 sg13g2_fill_8 FILLER_20_232 ();
 sg13g2_fill_8 FILLER_20_240 ();
 sg13g2_fill_8 FILLER_20_248 ();
 sg13g2_fill_8 FILLER_20_256 ();
 sg13g2_fill_8 FILLER_20_264 ();
 sg13g2_fill_8 FILLER_20_272 ();
 sg13g2_fill_8 FILLER_20_280 ();
 sg13g2_fill_8 FILLER_20_288 ();
 sg13g2_fill_8 FILLER_20_296 ();
 sg13g2_fill_8 FILLER_20_304 ();
 sg13g2_fill_8 FILLER_20_312 ();
 sg13g2_fill_8 FILLER_20_320 ();
 sg13g2_fill_8 FILLER_20_328 ();
 sg13g2_fill_8 FILLER_20_336 ();
 sg13g2_fill_8 FILLER_20_344 ();
 sg13g2_fill_8 FILLER_20_352 ();
 sg13g2_fill_8 FILLER_20_360 ();
 sg13g2_fill_8 FILLER_20_368 ();
 sg13g2_fill_8 FILLER_20_376 ();
 sg13g2_fill_8 FILLER_20_384 ();
 sg13g2_fill_8 FILLER_20_392 ();
 sg13g2_fill_8 FILLER_20_400 ();
 sg13g2_fill_8 FILLER_20_408 ();
 sg13g2_fill_8 FILLER_20_416 ();
 sg13g2_fill_8 FILLER_20_424 ();
 sg13g2_fill_8 FILLER_20_432 ();
 sg13g2_fill_8 FILLER_20_440 ();
 sg13g2_fill_8 FILLER_20_448 ();
 sg13g2_fill_8 FILLER_20_456 ();
 sg13g2_fill_8 FILLER_20_464 ();
 sg13g2_fill_8 FILLER_20_472 ();
 sg13g2_fill_8 FILLER_20_480 ();
 sg13g2_fill_8 FILLER_20_488 ();
 sg13g2_fill_8 FILLER_20_496 ();
 sg13g2_fill_8 FILLER_20_504 ();
 sg13g2_fill_8 FILLER_20_512 ();
 sg13g2_fill_8 FILLER_20_520 ();
 sg13g2_fill_8 FILLER_20_528 ();
 sg13g2_fill_8 FILLER_20_536 ();
 sg13g2_fill_8 FILLER_20_544 ();
 sg13g2_fill_8 FILLER_20_552 ();
 sg13g2_fill_8 FILLER_20_560 ();
 sg13g2_fill_8 FILLER_20_568 ();
 sg13g2_fill_8 FILLER_20_576 ();
 sg13g2_fill_8 FILLER_20_584 ();
 sg13g2_fill_8 FILLER_20_592 ();
 sg13g2_fill_8 FILLER_20_600 ();
 sg13g2_fill_8 FILLER_20_608 ();
 sg13g2_fill_8 FILLER_20_616 ();
 sg13g2_fill_8 FILLER_20_624 ();
 sg13g2_fill_8 FILLER_20_632 ();
 sg13g2_fill_8 FILLER_20_640 ();
 sg13g2_fill_8 FILLER_20_648 ();
 sg13g2_fill_8 FILLER_20_656 ();
 sg13g2_fill_8 FILLER_20_664 ();
 sg13g2_fill_8 FILLER_20_672 ();
 sg13g2_fill_8 FILLER_20_680 ();
 sg13g2_fill_8 FILLER_20_688 ();
 sg13g2_fill_8 FILLER_20_696 ();
 sg13g2_fill_8 FILLER_20_704 ();
 sg13g2_fill_8 FILLER_20_712 ();
 sg13g2_fill_8 FILLER_20_720 ();
 sg13g2_fill_8 FILLER_20_728 ();
 sg13g2_fill_8 FILLER_20_736 ();
 sg13g2_fill_8 FILLER_20_744 ();
 sg13g2_fill_8 FILLER_20_752 ();
 sg13g2_fill_8 FILLER_20_760 ();
 sg13g2_fill_8 FILLER_20_768 ();
 sg13g2_fill_8 FILLER_20_776 ();
 sg13g2_fill_8 FILLER_20_784 ();
 sg13g2_fill_8 FILLER_20_792 ();
 sg13g2_fill_8 FILLER_20_800 ();
 sg13g2_fill_8 FILLER_20_808 ();
 sg13g2_fill_8 FILLER_20_816 ();
 sg13g2_fill_8 FILLER_20_824 ();
 sg13g2_fill_8 FILLER_20_832 ();
 sg13g2_fill_8 FILLER_20_840 ();
 sg13g2_fill_8 FILLER_20_848 ();
 sg13g2_fill_8 FILLER_20_856 ();
 sg13g2_fill_8 FILLER_20_864 ();
 sg13g2_fill_8 FILLER_20_872 ();
 sg13g2_fill_8 FILLER_20_880 ();
 sg13g2_fill_8 FILLER_20_888 ();
 sg13g2_fill_8 FILLER_20_896 ();
 sg13g2_fill_8 FILLER_20_904 ();
 sg13g2_fill_8 FILLER_20_912 ();
 sg13g2_fill_8 FILLER_20_920 ();
 sg13g2_fill_8 FILLER_20_928 ();
 sg13g2_fill_8 FILLER_20_936 ();
 sg13g2_fill_8 FILLER_20_944 ();
 sg13g2_fill_8 FILLER_20_952 ();
 sg13g2_fill_8 FILLER_20_960 ();
 sg13g2_fill_8 FILLER_20_968 ();
 sg13g2_fill_8 FILLER_20_976 ();
 sg13g2_fill_8 FILLER_20_984 ();
 sg13g2_fill_8 FILLER_20_992 ();
 sg13g2_fill_8 FILLER_20_1000 ();
 sg13g2_fill_8 FILLER_20_1008 ();
 sg13g2_fill_8 FILLER_20_1016 ();
 sg13g2_fill_8 FILLER_20_1024 ();
 sg13g2_fill_8 FILLER_20_1032 ();
 sg13g2_fill_8 FILLER_20_1040 ();
 sg13g2_fill_8 FILLER_20_1048 ();
 sg13g2_fill_8 FILLER_20_1056 ();
 sg13g2_fill_8 FILLER_20_1064 ();
 sg13g2_fill_8 FILLER_20_1072 ();
 sg13g2_fill_8 FILLER_20_1080 ();
 sg13g2_fill_8 FILLER_20_1088 ();
 sg13g2_fill_8 FILLER_20_1096 ();
 sg13g2_fill_8 FILLER_20_1104 ();
 sg13g2_fill_8 FILLER_20_1112 ();
 sg13g2_fill_8 FILLER_20_1120 ();
 sg13g2_fill_8 FILLER_20_1128 ();
 sg13g2_fill_8 FILLER_20_1136 ();
 sg13g2_fill_8 FILLER_21_0 ();
 sg13g2_fill_8 FILLER_21_8 ();
 sg13g2_fill_8 FILLER_21_16 ();
 sg13g2_fill_8 FILLER_21_24 ();
 sg13g2_fill_8 FILLER_21_32 ();
 sg13g2_fill_8 FILLER_21_40 ();
 sg13g2_fill_8 FILLER_21_48 ();
 sg13g2_fill_8 FILLER_21_56 ();
 sg13g2_fill_8 FILLER_21_64 ();
 sg13g2_fill_8 FILLER_21_72 ();
 sg13g2_fill_8 FILLER_21_80 ();
 sg13g2_fill_8 FILLER_21_88 ();
 sg13g2_fill_8 FILLER_21_96 ();
 sg13g2_fill_8 FILLER_21_104 ();
 sg13g2_fill_8 FILLER_21_112 ();
 sg13g2_fill_8 FILLER_21_120 ();
 sg13g2_fill_8 FILLER_21_128 ();
 sg13g2_fill_8 FILLER_21_136 ();
 sg13g2_fill_8 FILLER_21_144 ();
 sg13g2_fill_8 FILLER_21_152 ();
 sg13g2_fill_8 FILLER_21_160 ();
 sg13g2_fill_8 FILLER_21_168 ();
 sg13g2_fill_8 FILLER_21_176 ();
 sg13g2_fill_8 FILLER_21_184 ();
 sg13g2_fill_8 FILLER_21_192 ();
 sg13g2_fill_8 FILLER_21_200 ();
 sg13g2_fill_8 FILLER_21_208 ();
 sg13g2_fill_8 FILLER_21_216 ();
 sg13g2_fill_8 FILLER_21_224 ();
 sg13g2_fill_8 FILLER_21_232 ();
 sg13g2_fill_8 FILLER_21_240 ();
 sg13g2_fill_8 FILLER_21_248 ();
 sg13g2_fill_8 FILLER_21_256 ();
 sg13g2_fill_8 FILLER_21_264 ();
 sg13g2_fill_8 FILLER_21_272 ();
 sg13g2_fill_8 FILLER_21_280 ();
 sg13g2_fill_8 FILLER_21_288 ();
 sg13g2_fill_8 FILLER_21_296 ();
 sg13g2_fill_8 FILLER_21_304 ();
 sg13g2_fill_8 FILLER_21_312 ();
 sg13g2_fill_8 FILLER_21_320 ();
 sg13g2_fill_8 FILLER_21_328 ();
 sg13g2_fill_8 FILLER_21_336 ();
 sg13g2_fill_8 FILLER_21_344 ();
 sg13g2_fill_8 FILLER_21_352 ();
 sg13g2_fill_8 FILLER_21_360 ();
 sg13g2_fill_8 FILLER_21_368 ();
 sg13g2_fill_8 FILLER_21_376 ();
 sg13g2_fill_8 FILLER_21_384 ();
 sg13g2_fill_8 FILLER_21_392 ();
 sg13g2_fill_8 FILLER_21_400 ();
 sg13g2_fill_8 FILLER_21_408 ();
 sg13g2_fill_8 FILLER_21_416 ();
 sg13g2_fill_8 FILLER_21_424 ();
 sg13g2_fill_8 FILLER_21_432 ();
 sg13g2_fill_8 FILLER_21_440 ();
 sg13g2_fill_8 FILLER_21_448 ();
 sg13g2_fill_8 FILLER_21_456 ();
 sg13g2_fill_8 FILLER_21_464 ();
 sg13g2_fill_8 FILLER_21_472 ();
 sg13g2_fill_8 FILLER_21_480 ();
 sg13g2_fill_8 FILLER_21_488 ();
 sg13g2_fill_8 FILLER_21_496 ();
 sg13g2_fill_8 FILLER_21_504 ();
 sg13g2_fill_8 FILLER_21_512 ();
 sg13g2_fill_8 FILLER_21_520 ();
 sg13g2_fill_8 FILLER_21_528 ();
 sg13g2_fill_8 FILLER_21_536 ();
 sg13g2_fill_8 FILLER_21_544 ();
 sg13g2_fill_8 FILLER_21_552 ();
 sg13g2_fill_8 FILLER_21_560 ();
 sg13g2_fill_8 FILLER_21_568 ();
 sg13g2_fill_8 FILLER_21_576 ();
 sg13g2_fill_8 FILLER_21_584 ();
 sg13g2_fill_8 FILLER_21_592 ();
 sg13g2_fill_8 FILLER_21_600 ();
 sg13g2_fill_8 FILLER_21_608 ();
 sg13g2_fill_8 FILLER_21_616 ();
 sg13g2_fill_8 FILLER_21_624 ();
 sg13g2_fill_8 FILLER_21_632 ();
 sg13g2_fill_8 FILLER_21_640 ();
 sg13g2_fill_8 FILLER_21_648 ();
 sg13g2_fill_8 FILLER_21_656 ();
 sg13g2_fill_8 FILLER_21_664 ();
 sg13g2_fill_8 FILLER_21_672 ();
 sg13g2_fill_8 FILLER_21_680 ();
 sg13g2_fill_8 FILLER_21_688 ();
 sg13g2_fill_8 FILLER_21_696 ();
 sg13g2_fill_8 FILLER_21_704 ();
 sg13g2_fill_8 FILLER_21_712 ();
 sg13g2_fill_8 FILLER_21_720 ();
 sg13g2_fill_8 FILLER_21_728 ();
 sg13g2_fill_8 FILLER_21_736 ();
 sg13g2_fill_8 FILLER_21_744 ();
 sg13g2_fill_8 FILLER_21_752 ();
 sg13g2_fill_8 FILLER_21_760 ();
 sg13g2_fill_8 FILLER_21_768 ();
 sg13g2_fill_8 FILLER_21_776 ();
 sg13g2_fill_8 FILLER_21_784 ();
 sg13g2_fill_8 FILLER_21_792 ();
 sg13g2_fill_8 FILLER_21_800 ();
 sg13g2_fill_8 FILLER_21_808 ();
 sg13g2_fill_8 FILLER_21_816 ();
 sg13g2_fill_8 FILLER_21_824 ();
 sg13g2_fill_8 FILLER_21_832 ();
 sg13g2_fill_8 FILLER_21_840 ();
 sg13g2_fill_8 FILLER_21_848 ();
 sg13g2_fill_8 FILLER_21_856 ();
 sg13g2_fill_8 FILLER_21_864 ();
 sg13g2_fill_8 FILLER_21_872 ();
 sg13g2_fill_8 FILLER_21_880 ();
 sg13g2_fill_8 FILLER_21_888 ();
 sg13g2_fill_8 FILLER_21_896 ();
 sg13g2_fill_8 FILLER_21_904 ();
 sg13g2_fill_8 FILLER_21_912 ();
 sg13g2_fill_8 FILLER_21_920 ();
 sg13g2_fill_8 FILLER_21_928 ();
 sg13g2_fill_8 FILLER_21_936 ();
 sg13g2_fill_8 FILLER_21_944 ();
 sg13g2_fill_8 FILLER_21_952 ();
 sg13g2_fill_8 FILLER_21_960 ();
 sg13g2_fill_8 FILLER_21_968 ();
 sg13g2_fill_8 FILLER_21_976 ();
 sg13g2_fill_8 FILLER_21_984 ();
 sg13g2_fill_8 FILLER_21_992 ();
 sg13g2_fill_8 FILLER_21_1000 ();
 sg13g2_fill_8 FILLER_21_1008 ();
 sg13g2_fill_8 FILLER_21_1016 ();
 sg13g2_fill_8 FILLER_21_1024 ();
 sg13g2_fill_8 FILLER_21_1032 ();
 sg13g2_fill_8 FILLER_21_1040 ();
 sg13g2_fill_8 FILLER_21_1048 ();
 sg13g2_fill_8 FILLER_21_1056 ();
 sg13g2_fill_8 FILLER_21_1064 ();
 sg13g2_fill_8 FILLER_21_1072 ();
 sg13g2_fill_8 FILLER_21_1080 ();
 sg13g2_fill_8 FILLER_21_1088 ();
 sg13g2_fill_8 FILLER_21_1096 ();
 sg13g2_fill_8 FILLER_21_1104 ();
 sg13g2_fill_8 FILLER_21_1112 ();
 sg13g2_fill_8 FILLER_21_1120 ();
 sg13g2_fill_8 FILLER_21_1128 ();
 sg13g2_fill_8 FILLER_21_1136 ();
 sg13g2_fill_8 FILLER_22_0 ();
 sg13g2_fill_8 FILLER_22_8 ();
 sg13g2_fill_8 FILLER_22_16 ();
 sg13g2_fill_8 FILLER_22_24 ();
 sg13g2_fill_8 FILLER_22_32 ();
 sg13g2_fill_8 FILLER_22_40 ();
 sg13g2_fill_8 FILLER_22_48 ();
 sg13g2_fill_8 FILLER_22_56 ();
 sg13g2_fill_8 FILLER_22_64 ();
 sg13g2_fill_8 FILLER_22_72 ();
 sg13g2_fill_8 FILLER_22_80 ();
 sg13g2_fill_8 FILLER_22_88 ();
 sg13g2_fill_8 FILLER_22_96 ();
 sg13g2_fill_8 FILLER_22_104 ();
 sg13g2_fill_8 FILLER_22_112 ();
 sg13g2_fill_8 FILLER_22_120 ();
 sg13g2_fill_8 FILLER_22_128 ();
 sg13g2_fill_8 FILLER_22_136 ();
 sg13g2_fill_8 FILLER_22_144 ();
 sg13g2_fill_8 FILLER_22_152 ();
 sg13g2_fill_8 FILLER_22_160 ();
 sg13g2_fill_8 FILLER_22_168 ();
 sg13g2_fill_8 FILLER_22_176 ();
 sg13g2_fill_8 FILLER_22_184 ();
 sg13g2_fill_8 FILLER_22_192 ();
 sg13g2_fill_8 FILLER_22_200 ();
 sg13g2_fill_8 FILLER_22_208 ();
 sg13g2_fill_8 FILLER_22_216 ();
 sg13g2_fill_8 FILLER_22_224 ();
 sg13g2_fill_8 FILLER_22_232 ();
 sg13g2_fill_8 FILLER_22_240 ();
 sg13g2_fill_8 FILLER_22_248 ();
 sg13g2_fill_8 FILLER_22_256 ();
 sg13g2_fill_8 FILLER_22_264 ();
 sg13g2_fill_8 FILLER_22_272 ();
 sg13g2_fill_8 FILLER_22_280 ();
 sg13g2_fill_8 FILLER_22_288 ();
 sg13g2_fill_8 FILLER_22_296 ();
 sg13g2_fill_8 FILLER_22_304 ();
 sg13g2_fill_8 FILLER_22_312 ();
 sg13g2_fill_8 FILLER_22_320 ();
 sg13g2_fill_8 FILLER_22_328 ();
 sg13g2_fill_8 FILLER_22_336 ();
 sg13g2_fill_8 FILLER_22_344 ();
 sg13g2_fill_8 FILLER_22_352 ();
 sg13g2_fill_8 FILLER_22_360 ();
 sg13g2_fill_8 FILLER_22_368 ();
 sg13g2_fill_8 FILLER_22_376 ();
 sg13g2_fill_8 FILLER_22_384 ();
 sg13g2_fill_8 FILLER_22_392 ();
 sg13g2_fill_8 FILLER_22_400 ();
 sg13g2_fill_8 FILLER_22_408 ();
 sg13g2_fill_8 FILLER_22_416 ();
 sg13g2_fill_8 FILLER_22_424 ();
 sg13g2_fill_8 FILLER_22_432 ();
 sg13g2_fill_8 FILLER_22_440 ();
 sg13g2_fill_8 FILLER_22_448 ();
 sg13g2_fill_8 FILLER_22_456 ();
 sg13g2_fill_8 FILLER_22_464 ();
 sg13g2_fill_8 FILLER_22_472 ();
 sg13g2_fill_8 FILLER_22_480 ();
 sg13g2_fill_8 FILLER_22_488 ();
 sg13g2_fill_8 FILLER_22_496 ();
 sg13g2_fill_8 FILLER_22_504 ();
 sg13g2_fill_8 FILLER_22_512 ();
 sg13g2_fill_8 FILLER_22_520 ();
 sg13g2_fill_8 FILLER_22_528 ();
 sg13g2_fill_8 FILLER_22_536 ();
 sg13g2_fill_8 FILLER_22_544 ();
 sg13g2_fill_8 FILLER_22_552 ();
 sg13g2_fill_8 FILLER_22_560 ();
 sg13g2_fill_8 FILLER_22_568 ();
 sg13g2_fill_8 FILLER_22_576 ();
 sg13g2_fill_8 FILLER_22_584 ();
 sg13g2_fill_8 FILLER_22_592 ();
 sg13g2_fill_8 FILLER_22_600 ();
 sg13g2_fill_8 FILLER_22_608 ();
 sg13g2_fill_8 FILLER_22_616 ();
 sg13g2_fill_8 FILLER_22_624 ();
 sg13g2_fill_8 FILLER_22_632 ();
 sg13g2_fill_8 FILLER_22_640 ();
 sg13g2_fill_8 FILLER_22_648 ();
 sg13g2_fill_8 FILLER_22_656 ();
 sg13g2_fill_8 FILLER_22_664 ();
 sg13g2_fill_8 FILLER_22_672 ();
 sg13g2_fill_8 FILLER_22_680 ();
 sg13g2_fill_8 FILLER_22_688 ();
 sg13g2_fill_8 FILLER_22_696 ();
 sg13g2_fill_8 FILLER_22_704 ();
 sg13g2_fill_8 FILLER_22_712 ();
 sg13g2_fill_8 FILLER_22_720 ();
 sg13g2_fill_8 FILLER_22_728 ();
 sg13g2_fill_8 FILLER_22_736 ();
 sg13g2_fill_8 FILLER_22_744 ();
 sg13g2_fill_8 FILLER_22_752 ();
 sg13g2_fill_8 FILLER_22_760 ();
 sg13g2_fill_8 FILLER_22_768 ();
 sg13g2_fill_8 FILLER_22_776 ();
 sg13g2_fill_8 FILLER_22_784 ();
 sg13g2_fill_8 FILLER_22_792 ();
 sg13g2_fill_8 FILLER_22_800 ();
 sg13g2_fill_8 FILLER_22_808 ();
 sg13g2_fill_8 FILLER_22_816 ();
 sg13g2_fill_8 FILLER_22_824 ();
 sg13g2_fill_8 FILLER_22_832 ();
 sg13g2_fill_8 FILLER_22_840 ();
 sg13g2_fill_8 FILLER_22_848 ();
 sg13g2_fill_8 FILLER_22_856 ();
 sg13g2_fill_8 FILLER_22_864 ();
 sg13g2_fill_8 FILLER_22_872 ();
 sg13g2_fill_8 FILLER_22_880 ();
 sg13g2_fill_8 FILLER_22_888 ();
 sg13g2_fill_8 FILLER_22_896 ();
 sg13g2_fill_8 FILLER_22_904 ();
 sg13g2_fill_8 FILLER_22_912 ();
 sg13g2_fill_8 FILLER_22_920 ();
 sg13g2_fill_8 FILLER_22_928 ();
 sg13g2_fill_8 FILLER_22_936 ();
 sg13g2_fill_8 FILLER_22_944 ();
 sg13g2_fill_8 FILLER_22_952 ();
 sg13g2_fill_8 FILLER_22_960 ();
 sg13g2_fill_8 FILLER_22_968 ();
 sg13g2_fill_8 FILLER_22_976 ();
 sg13g2_fill_8 FILLER_22_984 ();
 sg13g2_fill_8 FILLER_22_992 ();
 sg13g2_fill_8 FILLER_22_1000 ();
 sg13g2_fill_8 FILLER_22_1008 ();
 sg13g2_fill_8 FILLER_22_1016 ();
 sg13g2_fill_8 FILLER_22_1024 ();
 sg13g2_fill_8 FILLER_22_1032 ();
 sg13g2_fill_8 FILLER_22_1040 ();
 sg13g2_fill_8 FILLER_22_1048 ();
 sg13g2_fill_8 FILLER_22_1056 ();
 sg13g2_fill_8 FILLER_22_1064 ();
 sg13g2_fill_8 FILLER_22_1072 ();
 sg13g2_fill_8 FILLER_22_1080 ();
 sg13g2_fill_8 FILLER_22_1088 ();
 sg13g2_fill_8 FILLER_22_1096 ();
 sg13g2_fill_8 FILLER_22_1104 ();
 sg13g2_fill_8 FILLER_22_1112 ();
 sg13g2_fill_8 FILLER_22_1120 ();
 sg13g2_fill_8 FILLER_22_1128 ();
 sg13g2_fill_8 FILLER_22_1136 ();
 sg13g2_fill_8 FILLER_23_0 ();
 sg13g2_fill_8 FILLER_23_8 ();
 sg13g2_fill_8 FILLER_23_16 ();
 sg13g2_fill_8 FILLER_23_24 ();
 sg13g2_fill_8 FILLER_23_32 ();
 sg13g2_fill_8 FILLER_23_40 ();
 sg13g2_fill_8 FILLER_23_48 ();
 sg13g2_fill_8 FILLER_23_56 ();
 sg13g2_fill_8 FILLER_23_64 ();
 sg13g2_fill_8 FILLER_23_72 ();
 sg13g2_fill_8 FILLER_23_80 ();
 sg13g2_fill_8 FILLER_23_88 ();
 sg13g2_fill_8 FILLER_23_96 ();
 sg13g2_fill_8 FILLER_23_104 ();
 sg13g2_fill_8 FILLER_23_112 ();
 sg13g2_fill_8 FILLER_23_120 ();
 sg13g2_fill_8 FILLER_23_128 ();
 sg13g2_fill_8 FILLER_23_136 ();
 sg13g2_fill_8 FILLER_23_144 ();
 sg13g2_fill_8 FILLER_23_152 ();
 sg13g2_fill_8 FILLER_23_160 ();
 sg13g2_fill_8 FILLER_23_168 ();
 sg13g2_fill_8 FILLER_23_176 ();
 sg13g2_fill_8 FILLER_23_184 ();
 sg13g2_fill_8 FILLER_23_192 ();
 sg13g2_fill_8 FILLER_23_200 ();
 sg13g2_fill_8 FILLER_23_208 ();
 sg13g2_fill_8 FILLER_23_216 ();
 sg13g2_fill_8 FILLER_23_224 ();
 sg13g2_fill_8 FILLER_23_232 ();
 sg13g2_fill_8 FILLER_23_240 ();
 sg13g2_fill_8 FILLER_23_248 ();
 sg13g2_fill_8 FILLER_23_256 ();
 sg13g2_fill_8 FILLER_23_264 ();
 sg13g2_fill_8 FILLER_23_272 ();
 sg13g2_fill_8 FILLER_23_280 ();
 sg13g2_fill_8 FILLER_23_288 ();
 sg13g2_fill_8 FILLER_23_296 ();
 sg13g2_fill_8 FILLER_23_304 ();
 sg13g2_fill_8 FILLER_23_312 ();
 sg13g2_fill_8 FILLER_23_320 ();
 sg13g2_fill_8 FILLER_23_328 ();
 sg13g2_fill_8 FILLER_23_336 ();
 sg13g2_fill_8 FILLER_23_344 ();
 sg13g2_fill_8 FILLER_23_352 ();
 sg13g2_fill_8 FILLER_23_360 ();
 sg13g2_fill_8 FILLER_23_368 ();
 sg13g2_fill_8 FILLER_23_376 ();
 sg13g2_fill_8 FILLER_23_384 ();
 sg13g2_fill_8 FILLER_23_392 ();
 sg13g2_fill_8 FILLER_23_400 ();
 sg13g2_fill_8 FILLER_23_408 ();
 sg13g2_fill_8 FILLER_23_416 ();
 sg13g2_fill_8 FILLER_23_424 ();
 sg13g2_fill_8 FILLER_23_432 ();
 sg13g2_fill_8 FILLER_23_440 ();
 sg13g2_fill_8 FILLER_23_448 ();
 sg13g2_fill_8 FILLER_23_456 ();
 sg13g2_fill_8 FILLER_23_464 ();
 sg13g2_fill_8 FILLER_23_472 ();
 sg13g2_fill_8 FILLER_23_480 ();
 sg13g2_fill_8 FILLER_23_488 ();
 sg13g2_fill_8 FILLER_23_496 ();
 sg13g2_fill_8 FILLER_23_504 ();
 sg13g2_fill_8 FILLER_23_512 ();
 sg13g2_fill_8 FILLER_23_520 ();
 sg13g2_fill_8 FILLER_23_528 ();
 sg13g2_fill_8 FILLER_23_536 ();
 sg13g2_fill_8 FILLER_23_544 ();
 sg13g2_fill_8 FILLER_23_552 ();
 sg13g2_fill_8 FILLER_23_560 ();
 sg13g2_fill_8 FILLER_23_568 ();
 sg13g2_fill_8 FILLER_23_576 ();
 sg13g2_fill_8 FILLER_23_584 ();
 sg13g2_fill_8 FILLER_23_592 ();
 sg13g2_fill_8 FILLER_23_600 ();
 sg13g2_fill_8 FILLER_23_608 ();
 sg13g2_fill_8 FILLER_23_616 ();
 sg13g2_fill_8 FILLER_23_624 ();
 sg13g2_fill_8 FILLER_23_632 ();
 sg13g2_fill_8 FILLER_23_640 ();
 sg13g2_fill_8 FILLER_23_648 ();
 sg13g2_fill_8 FILLER_23_656 ();
 sg13g2_fill_8 FILLER_23_664 ();
 sg13g2_fill_8 FILLER_23_672 ();
 sg13g2_fill_8 FILLER_23_680 ();
 sg13g2_fill_8 FILLER_23_688 ();
 sg13g2_fill_8 FILLER_23_696 ();
 sg13g2_fill_8 FILLER_23_704 ();
 sg13g2_fill_8 FILLER_23_712 ();
 sg13g2_fill_8 FILLER_23_720 ();
 sg13g2_fill_8 FILLER_23_728 ();
 sg13g2_fill_8 FILLER_23_736 ();
 sg13g2_fill_8 FILLER_23_744 ();
 sg13g2_fill_8 FILLER_23_752 ();
 sg13g2_fill_8 FILLER_23_760 ();
 sg13g2_fill_8 FILLER_23_768 ();
 sg13g2_fill_8 FILLER_23_776 ();
 sg13g2_fill_8 FILLER_23_784 ();
 sg13g2_fill_8 FILLER_23_792 ();
 sg13g2_fill_8 FILLER_23_800 ();
 sg13g2_fill_8 FILLER_23_808 ();
 sg13g2_fill_8 FILLER_23_816 ();
 sg13g2_fill_8 FILLER_23_824 ();
 sg13g2_fill_8 FILLER_23_832 ();
 sg13g2_fill_8 FILLER_23_840 ();
 sg13g2_fill_8 FILLER_23_848 ();
 sg13g2_fill_8 FILLER_23_856 ();
 sg13g2_fill_8 FILLER_23_864 ();
 sg13g2_fill_8 FILLER_23_872 ();
 sg13g2_fill_8 FILLER_23_880 ();
 sg13g2_fill_8 FILLER_23_888 ();
 sg13g2_fill_8 FILLER_23_896 ();
 sg13g2_fill_8 FILLER_23_904 ();
 sg13g2_fill_8 FILLER_23_912 ();
 sg13g2_fill_8 FILLER_23_920 ();
 sg13g2_fill_8 FILLER_23_928 ();
 sg13g2_fill_8 FILLER_23_936 ();
 sg13g2_fill_8 FILLER_23_944 ();
 sg13g2_fill_8 FILLER_23_952 ();
 sg13g2_fill_8 FILLER_23_960 ();
 sg13g2_fill_8 FILLER_23_968 ();
 sg13g2_fill_8 FILLER_23_976 ();
 sg13g2_fill_8 FILLER_23_984 ();
 sg13g2_fill_8 FILLER_23_992 ();
 sg13g2_fill_8 FILLER_23_1000 ();
 sg13g2_fill_8 FILLER_23_1008 ();
 sg13g2_fill_8 FILLER_23_1016 ();
 sg13g2_fill_8 FILLER_23_1024 ();
 sg13g2_fill_8 FILLER_23_1032 ();
 sg13g2_fill_8 FILLER_23_1040 ();
 sg13g2_fill_8 FILLER_23_1048 ();
 sg13g2_fill_8 FILLER_23_1056 ();
 sg13g2_fill_8 FILLER_23_1064 ();
 sg13g2_fill_8 FILLER_23_1072 ();
 sg13g2_fill_8 FILLER_23_1080 ();
 sg13g2_fill_8 FILLER_23_1088 ();
 sg13g2_fill_8 FILLER_23_1096 ();
 sg13g2_fill_8 FILLER_23_1104 ();
 sg13g2_fill_8 FILLER_23_1112 ();
 sg13g2_fill_8 FILLER_23_1120 ();
 sg13g2_fill_8 FILLER_23_1128 ();
 sg13g2_fill_8 FILLER_23_1136 ();
 sg13g2_fill_8 FILLER_24_0 ();
 sg13g2_fill_8 FILLER_24_8 ();
 sg13g2_fill_8 FILLER_24_16 ();
 sg13g2_fill_8 FILLER_24_24 ();
 sg13g2_fill_8 FILLER_24_32 ();
 sg13g2_fill_8 FILLER_24_40 ();
 sg13g2_fill_8 FILLER_24_48 ();
 sg13g2_fill_8 FILLER_24_56 ();
 sg13g2_fill_8 FILLER_24_64 ();
 sg13g2_fill_8 FILLER_24_72 ();
 sg13g2_fill_8 FILLER_24_80 ();
 sg13g2_fill_8 FILLER_24_88 ();
 sg13g2_fill_8 FILLER_24_96 ();
 sg13g2_fill_8 FILLER_24_104 ();
 sg13g2_fill_8 FILLER_24_112 ();
 sg13g2_fill_8 FILLER_24_120 ();
 sg13g2_fill_8 FILLER_24_128 ();
 sg13g2_fill_8 FILLER_24_136 ();
 sg13g2_fill_8 FILLER_24_144 ();
 sg13g2_fill_8 FILLER_24_152 ();
 sg13g2_fill_8 FILLER_24_160 ();
 sg13g2_fill_8 FILLER_24_168 ();
 sg13g2_fill_8 FILLER_24_176 ();
 sg13g2_fill_8 FILLER_24_184 ();
 sg13g2_fill_8 FILLER_24_192 ();
 sg13g2_fill_8 FILLER_24_200 ();
 sg13g2_fill_8 FILLER_24_208 ();
 sg13g2_fill_8 FILLER_24_216 ();
 sg13g2_fill_8 FILLER_24_224 ();
 sg13g2_fill_8 FILLER_24_232 ();
 sg13g2_fill_8 FILLER_24_240 ();
 sg13g2_fill_8 FILLER_24_248 ();
 sg13g2_fill_8 FILLER_24_256 ();
 sg13g2_fill_8 FILLER_24_264 ();
 sg13g2_fill_8 FILLER_24_272 ();
 sg13g2_fill_8 FILLER_24_280 ();
 sg13g2_fill_8 FILLER_24_288 ();
 sg13g2_fill_8 FILLER_24_296 ();
 sg13g2_fill_8 FILLER_24_304 ();
 sg13g2_fill_8 FILLER_24_312 ();
 sg13g2_fill_8 FILLER_24_320 ();
 sg13g2_fill_8 FILLER_24_328 ();
 sg13g2_fill_8 FILLER_24_336 ();
 sg13g2_fill_8 FILLER_24_344 ();
 sg13g2_fill_8 FILLER_24_352 ();
 sg13g2_fill_8 FILLER_24_360 ();
 sg13g2_fill_8 FILLER_24_368 ();
 sg13g2_fill_8 FILLER_24_376 ();
 sg13g2_fill_8 FILLER_24_384 ();
 sg13g2_fill_8 FILLER_24_392 ();
 sg13g2_fill_8 FILLER_24_400 ();
 sg13g2_fill_8 FILLER_24_408 ();
 sg13g2_fill_8 FILLER_24_416 ();
 sg13g2_fill_8 FILLER_24_424 ();
 sg13g2_fill_8 FILLER_24_432 ();
 sg13g2_fill_8 FILLER_24_440 ();
 sg13g2_fill_8 FILLER_24_448 ();
 sg13g2_fill_8 FILLER_24_456 ();
 sg13g2_fill_8 FILLER_24_464 ();
 sg13g2_fill_8 FILLER_24_472 ();
 sg13g2_fill_8 FILLER_24_480 ();
 sg13g2_fill_8 FILLER_24_488 ();
 sg13g2_fill_8 FILLER_24_496 ();
 sg13g2_fill_8 FILLER_24_504 ();
 sg13g2_fill_8 FILLER_24_512 ();
 sg13g2_fill_8 FILLER_24_520 ();
 sg13g2_fill_8 FILLER_24_528 ();
 sg13g2_fill_8 FILLER_24_536 ();
 sg13g2_fill_8 FILLER_24_544 ();
 sg13g2_fill_8 FILLER_24_552 ();
 sg13g2_fill_8 FILLER_24_560 ();
 sg13g2_fill_8 FILLER_24_568 ();
 sg13g2_fill_8 FILLER_24_576 ();
 sg13g2_fill_8 FILLER_24_584 ();
 sg13g2_fill_8 FILLER_24_592 ();
 sg13g2_fill_8 FILLER_24_600 ();
 sg13g2_fill_8 FILLER_24_608 ();
 sg13g2_fill_8 FILLER_24_616 ();
 sg13g2_fill_8 FILLER_24_624 ();
 sg13g2_fill_8 FILLER_24_632 ();
 sg13g2_fill_8 FILLER_24_640 ();
 sg13g2_fill_8 FILLER_24_648 ();
 sg13g2_fill_8 FILLER_24_656 ();
 sg13g2_fill_8 FILLER_24_664 ();
 sg13g2_fill_8 FILLER_24_672 ();
 sg13g2_fill_8 FILLER_24_680 ();
 sg13g2_fill_8 FILLER_24_688 ();
 sg13g2_fill_8 FILLER_24_696 ();
 sg13g2_fill_8 FILLER_24_704 ();
 sg13g2_fill_8 FILLER_24_712 ();
 sg13g2_fill_8 FILLER_24_720 ();
 sg13g2_fill_8 FILLER_24_728 ();
 sg13g2_fill_8 FILLER_24_736 ();
 sg13g2_fill_8 FILLER_24_744 ();
 sg13g2_fill_8 FILLER_24_752 ();
 sg13g2_fill_8 FILLER_24_760 ();
 sg13g2_fill_8 FILLER_24_768 ();
 sg13g2_fill_8 FILLER_24_776 ();
 sg13g2_fill_8 FILLER_24_784 ();
 sg13g2_fill_8 FILLER_24_792 ();
 sg13g2_fill_8 FILLER_24_800 ();
 sg13g2_fill_8 FILLER_24_808 ();
 sg13g2_fill_8 FILLER_24_816 ();
 sg13g2_fill_8 FILLER_24_824 ();
 sg13g2_fill_8 FILLER_24_832 ();
 sg13g2_fill_8 FILLER_24_840 ();
 sg13g2_fill_8 FILLER_24_848 ();
 sg13g2_fill_8 FILLER_24_856 ();
 sg13g2_fill_8 FILLER_24_864 ();
 sg13g2_fill_8 FILLER_24_872 ();
 sg13g2_fill_8 FILLER_24_880 ();
 sg13g2_fill_8 FILLER_24_888 ();
 sg13g2_fill_8 FILLER_24_896 ();
 sg13g2_fill_8 FILLER_24_904 ();
 sg13g2_fill_8 FILLER_24_912 ();
 sg13g2_fill_8 FILLER_24_920 ();
 sg13g2_fill_8 FILLER_24_928 ();
 sg13g2_fill_8 FILLER_24_936 ();
 sg13g2_fill_8 FILLER_24_944 ();
 sg13g2_fill_8 FILLER_24_952 ();
 sg13g2_fill_8 FILLER_24_960 ();
 sg13g2_fill_8 FILLER_24_968 ();
 sg13g2_fill_8 FILLER_24_976 ();
 sg13g2_fill_8 FILLER_24_984 ();
 sg13g2_fill_8 FILLER_24_992 ();
 sg13g2_fill_8 FILLER_24_1000 ();
 sg13g2_fill_8 FILLER_24_1008 ();
 sg13g2_fill_8 FILLER_24_1016 ();
 sg13g2_fill_8 FILLER_24_1024 ();
 sg13g2_fill_8 FILLER_24_1032 ();
 sg13g2_fill_8 FILLER_24_1040 ();
 sg13g2_fill_8 FILLER_24_1048 ();
 sg13g2_fill_8 FILLER_24_1056 ();
 sg13g2_fill_8 FILLER_24_1064 ();
 sg13g2_fill_8 FILLER_24_1072 ();
 sg13g2_fill_8 FILLER_24_1080 ();
 sg13g2_fill_8 FILLER_24_1088 ();
 sg13g2_fill_8 FILLER_24_1096 ();
 sg13g2_fill_8 FILLER_24_1104 ();
 sg13g2_fill_8 FILLER_24_1112 ();
 sg13g2_fill_8 FILLER_24_1120 ();
 sg13g2_fill_8 FILLER_24_1128 ();
 sg13g2_fill_8 FILLER_24_1136 ();
 sg13g2_fill_8 FILLER_25_0 ();
 sg13g2_fill_8 FILLER_25_8 ();
 sg13g2_fill_8 FILLER_25_16 ();
 sg13g2_fill_8 FILLER_25_24 ();
 sg13g2_fill_8 FILLER_25_32 ();
 sg13g2_fill_8 FILLER_25_40 ();
 sg13g2_fill_8 FILLER_25_48 ();
 sg13g2_fill_8 FILLER_25_56 ();
 sg13g2_fill_8 FILLER_25_64 ();
 sg13g2_fill_8 FILLER_25_72 ();
 sg13g2_fill_8 FILLER_25_80 ();
 sg13g2_fill_8 FILLER_25_88 ();
 sg13g2_fill_8 FILLER_25_96 ();
 sg13g2_fill_8 FILLER_25_104 ();
 sg13g2_fill_8 FILLER_25_112 ();
 sg13g2_fill_8 FILLER_25_120 ();
 sg13g2_fill_8 FILLER_25_128 ();
 sg13g2_fill_8 FILLER_25_136 ();
 sg13g2_fill_8 FILLER_25_144 ();
 sg13g2_fill_8 FILLER_25_152 ();
 sg13g2_fill_8 FILLER_25_160 ();
 sg13g2_fill_8 FILLER_25_168 ();
 sg13g2_fill_8 FILLER_25_176 ();
 sg13g2_fill_8 FILLER_25_184 ();
 sg13g2_fill_8 FILLER_25_192 ();
 sg13g2_fill_8 FILLER_25_200 ();
 sg13g2_fill_8 FILLER_25_208 ();
 sg13g2_fill_8 FILLER_25_216 ();
 sg13g2_fill_8 FILLER_25_224 ();
 sg13g2_fill_8 FILLER_25_232 ();
 sg13g2_fill_8 FILLER_25_240 ();
 sg13g2_fill_8 FILLER_25_248 ();
 sg13g2_fill_8 FILLER_25_256 ();
 sg13g2_fill_8 FILLER_25_264 ();
 sg13g2_fill_8 FILLER_25_272 ();
 sg13g2_fill_8 FILLER_25_280 ();
 sg13g2_fill_8 FILLER_25_288 ();
 sg13g2_fill_8 FILLER_25_296 ();
 sg13g2_fill_8 FILLER_25_304 ();
 sg13g2_fill_8 FILLER_25_312 ();
 sg13g2_fill_8 FILLER_25_320 ();
 sg13g2_fill_8 FILLER_25_328 ();
 sg13g2_fill_8 FILLER_25_336 ();
 sg13g2_fill_8 FILLER_25_344 ();
 sg13g2_fill_8 FILLER_25_352 ();
 sg13g2_fill_8 FILLER_25_360 ();
 sg13g2_fill_8 FILLER_25_368 ();
 sg13g2_fill_8 FILLER_25_376 ();
 sg13g2_fill_8 FILLER_25_384 ();
 sg13g2_fill_8 FILLER_25_392 ();
 sg13g2_fill_8 FILLER_25_400 ();
 sg13g2_fill_8 FILLER_25_408 ();
 sg13g2_fill_8 FILLER_25_416 ();
 sg13g2_fill_8 FILLER_25_424 ();
 sg13g2_fill_8 FILLER_25_432 ();
 sg13g2_fill_8 FILLER_25_440 ();
 sg13g2_fill_8 FILLER_25_448 ();
 sg13g2_fill_8 FILLER_25_456 ();
 sg13g2_fill_8 FILLER_25_464 ();
 sg13g2_fill_8 FILLER_25_472 ();
 sg13g2_fill_8 FILLER_25_480 ();
 sg13g2_fill_8 FILLER_25_488 ();
 sg13g2_fill_8 FILLER_25_496 ();
 sg13g2_fill_8 FILLER_25_504 ();
 sg13g2_fill_8 FILLER_25_512 ();
 sg13g2_fill_8 FILLER_25_520 ();
 sg13g2_fill_8 FILLER_25_528 ();
 sg13g2_fill_8 FILLER_25_536 ();
 sg13g2_fill_8 FILLER_25_544 ();
 sg13g2_fill_8 FILLER_25_552 ();
 sg13g2_fill_8 FILLER_25_560 ();
 sg13g2_fill_8 FILLER_25_568 ();
 sg13g2_fill_8 FILLER_25_576 ();
 sg13g2_fill_8 FILLER_25_584 ();
 sg13g2_fill_8 FILLER_25_592 ();
 sg13g2_fill_8 FILLER_25_600 ();
 sg13g2_fill_8 FILLER_25_608 ();
 sg13g2_fill_8 FILLER_25_616 ();
 sg13g2_fill_8 FILLER_25_624 ();
 sg13g2_fill_8 FILLER_25_632 ();
 sg13g2_fill_8 FILLER_25_640 ();
 sg13g2_fill_8 FILLER_25_648 ();
 sg13g2_fill_8 FILLER_25_656 ();
 sg13g2_fill_8 FILLER_25_664 ();
 sg13g2_fill_8 FILLER_25_672 ();
 sg13g2_fill_8 FILLER_25_680 ();
 sg13g2_fill_8 FILLER_25_688 ();
 sg13g2_fill_8 FILLER_25_696 ();
 sg13g2_fill_8 FILLER_25_704 ();
 sg13g2_fill_8 FILLER_25_712 ();
 sg13g2_fill_8 FILLER_25_720 ();
 sg13g2_fill_8 FILLER_25_728 ();
 sg13g2_fill_8 FILLER_25_736 ();
 sg13g2_fill_8 FILLER_25_744 ();
 sg13g2_fill_8 FILLER_25_752 ();
 sg13g2_fill_8 FILLER_25_760 ();
 sg13g2_fill_8 FILLER_25_768 ();
 sg13g2_fill_8 FILLER_25_776 ();
 sg13g2_fill_8 FILLER_25_784 ();
 sg13g2_fill_8 FILLER_25_792 ();
 sg13g2_fill_8 FILLER_25_800 ();
 sg13g2_fill_8 FILLER_25_808 ();
 sg13g2_fill_8 FILLER_25_816 ();
 sg13g2_fill_8 FILLER_25_824 ();
 sg13g2_fill_8 FILLER_25_832 ();
 sg13g2_fill_8 FILLER_25_840 ();
 sg13g2_fill_8 FILLER_25_848 ();
 sg13g2_fill_8 FILLER_25_856 ();
 sg13g2_fill_8 FILLER_25_864 ();
 sg13g2_fill_8 FILLER_25_872 ();
 sg13g2_fill_8 FILLER_25_880 ();
 sg13g2_fill_8 FILLER_25_888 ();
 sg13g2_fill_8 FILLER_25_896 ();
 sg13g2_fill_8 FILLER_25_904 ();
 sg13g2_fill_8 FILLER_25_912 ();
 sg13g2_fill_8 FILLER_25_920 ();
 sg13g2_fill_8 FILLER_25_928 ();
 sg13g2_fill_8 FILLER_25_936 ();
 sg13g2_fill_8 FILLER_25_944 ();
 sg13g2_fill_8 FILLER_25_952 ();
 sg13g2_fill_8 FILLER_25_960 ();
 sg13g2_fill_8 FILLER_25_968 ();
 sg13g2_fill_8 FILLER_25_976 ();
 sg13g2_fill_8 FILLER_25_984 ();
 sg13g2_fill_8 FILLER_25_992 ();
 sg13g2_fill_8 FILLER_25_1000 ();
 sg13g2_fill_8 FILLER_25_1008 ();
 sg13g2_fill_8 FILLER_25_1016 ();
 sg13g2_fill_8 FILLER_25_1024 ();
 sg13g2_fill_8 FILLER_25_1032 ();
 sg13g2_fill_8 FILLER_25_1040 ();
 sg13g2_fill_8 FILLER_25_1048 ();
 sg13g2_fill_8 FILLER_25_1056 ();
 sg13g2_fill_8 FILLER_25_1064 ();
 sg13g2_fill_8 FILLER_25_1072 ();
 sg13g2_fill_8 FILLER_25_1080 ();
 sg13g2_fill_8 FILLER_25_1088 ();
 sg13g2_fill_8 FILLER_25_1096 ();
 sg13g2_fill_8 FILLER_25_1104 ();
 sg13g2_fill_8 FILLER_25_1112 ();
 sg13g2_fill_8 FILLER_25_1120 ();
 sg13g2_fill_8 FILLER_25_1128 ();
 sg13g2_fill_8 FILLER_25_1136 ();
 sg13g2_fill_8 FILLER_26_0 ();
 sg13g2_fill_8 FILLER_26_8 ();
 sg13g2_fill_8 FILLER_26_16 ();
 sg13g2_fill_8 FILLER_26_24 ();
 sg13g2_fill_8 FILLER_26_32 ();
 sg13g2_fill_8 FILLER_26_40 ();
 sg13g2_fill_8 FILLER_26_48 ();
 sg13g2_fill_8 FILLER_26_56 ();
 sg13g2_fill_8 FILLER_26_64 ();
 sg13g2_fill_8 FILLER_26_72 ();
 sg13g2_fill_8 FILLER_26_80 ();
 sg13g2_fill_8 FILLER_26_88 ();
 sg13g2_fill_8 FILLER_26_96 ();
 sg13g2_fill_8 FILLER_26_104 ();
 sg13g2_fill_8 FILLER_26_112 ();
 sg13g2_fill_8 FILLER_26_120 ();
 sg13g2_fill_8 FILLER_26_128 ();
 sg13g2_fill_8 FILLER_26_136 ();
 sg13g2_fill_8 FILLER_26_144 ();
 sg13g2_fill_8 FILLER_26_152 ();
 sg13g2_fill_8 FILLER_26_160 ();
 sg13g2_fill_8 FILLER_26_168 ();
 sg13g2_fill_8 FILLER_26_176 ();
 sg13g2_fill_8 FILLER_26_184 ();
 sg13g2_fill_8 FILLER_26_192 ();
 sg13g2_fill_8 FILLER_26_200 ();
 sg13g2_fill_8 FILLER_26_208 ();
 sg13g2_fill_8 FILLER_26_216 ();
 sg13g2_fill_8 FILLER_26_224 ();
 sg13g2_fill_8 FILLER_26_232 ();
 sg13g2_fill_8 FILLER_26_240 ();
 sg13g2_fill_8 FILLER_26_248 ();
 sg13g2_fill_8 FILLER_26_256 ();
 sg13g2_fill_8 FILLER_26_264 ();
 sg13g2_fill_8 FILLER_26_272 ();
 sg13g2_fill_8 FILLER_26_280 ();
 sg13g2_fill_8 FILLER_26_288 ();
 sg13g2_fill_8 FILLER_26_296 ();
 sg13g2_fill_8 FILLER_26_304 ();
 sg13g2_fill_8 FILLER_26_312 ();
 sg13g2_fill_8 FILLER_26_320 ();
 sg13g2_fill_8 FILLER_26_328 ();
 sg13g2_fill_8 FILLER_26_336 ();
 sg13g2_fill_8 FILLER_26_344 ();
 sg13g2_fill_8 FILLER_26_352 ();
 sg13g2_fill_8 FILLER_26_360 ();
 sg13g2_fill_8 FILLER_26_368 ();
 sg13g2_fill_8 FILLER_26_376 ();
 sg13g2_fill_8 FILLER_26_384 ();
 sg13g2_fill_8 FILLER_26_392 ();
 sg13g2_fill_8 FILLER_26_400 ();
 sg13g2_fill_8 FILLER_26_408 ();
 sg13g2_fill_8 FILLER_26_416 ();
 sg13g2_fill_8 FILLER_26_424 ();
 sg13g2_fill_8 FILLER_26_432 ();
 sg13g2_fill_8 FILLER_26_440 ();
 sg13g2_fill_8 FILLER_26_448 ();
 sg13g2_fill_8 FILLER_26_456 ();
 sg13g2_fill_8 FILLER_26_464 ();
 sg13g2_fill_8 FILLER_26_472 ();
 sg13g2_fill_8 FILLER_26_480 ();
 sg13g2_fill_8 FILLER_26_488 ();
 sg13g2_fill_8 FILLER_26_496 ();
 sg13g2_fill_8 FILLER_26_504 ();
 sg13g2_fill_8 FILLER_26_512 ();
 sg13g2_fill_8 FILLER_26_520 ();
 sg13g2_fill_8 FILLER_26_528 ();
 sg13g2_fill_8 FILLER_26_536 ();
 sg13g2_fill_8 FILLER_26_544 ();
 sg13g2_fill_8 FILLER_26_552 ();
 sg13g2_fill_8 FILLER_26_560 ();
 sg13g2_fill_8 FILLER_26_568 ();
 sg13g2_fill_8 FILLER_26_576 ();
 sg13g2_fill_8 FILLER_26_584 ();
 sg13g2_fill_8 FILLER_26_592 ();
 sg13g2_fill_8 FILLER_26_600 ();
 sg13g2_fill_8 FILLER_26_608 ();
 sg13g2_fill_8 FILLER_26_616 ();
 sg13g2_fill_8 FILLER_26_624 ();
 sg13g2_fill_8 FILLER_26_632 ();
 sg13g2_fill_8 FILLER_26_640 ();
 sg13g2_fill_8 FILLER_26_648 ();
 sg13g2_fill_8 FILLER_26_656 ();
 sg13g2_fill_8 FILLER_26_664 ();
 sg13g2_fill_8 FILLER_26_672 ();
 sg13g2_fill_8 FILLER_26_680 ();
 sg13g2_fill_8 FILLER_26_688 ();
 sg13g2_fill_8 FILLER_26_696 ();
 sg13g2_fill_8 FILLER_26_704 ();
 sg13g2_fill_8 FILLER_26_712 ();
 sg13g2_fill_8 FILLER_26_720 ();
 sg13g2_fill_8 FILLER_26_728 ();
 sg13g2_fill_8 FILLER_26_736 ();
 sg13g2_fill_8 FILLER_26_744 ();
 sg13g2_fill_8 FILLER_26_752 ();
 sg13g2_fill_8 FILLER_26_760 ();
 sg13g2_fill_8 FILLER_26_768 ();
 sg13g2_fill_8 FILLER_26_776 ();
 sg13g2_fill_8 FILLER_26_784 ();
 sg13g2_fill_8 FILLER_26_792 ();
 sg13g2_fill_8 FILLER_26_800 ();
 sg13g2_fill_8 FILLER_26_808 ();
 sg13g2_fill_8 FILLER_26_816 ();
 sg13g2_fill_8 FILLER_26_824 ();
 sg13g2_fill_8 FILLER_26_832 ();
 sg13g2_fill_8 FILLER_26_840 ();
 sg13g2_fill_8 FILLER_26_848 ();
 sg13g2_fill_8 FILLER_26_856 ();
 sg13g2_fill_8 FILLER_26_864 ();
 sg13g2_fill_8 FILLER_26_872 ();
 sg13g2_fill_8 FILLER_26_880 ();
 sg13g2_fill_8 FILLER_26_888 ();
 sg13g2_fill_8 FILLER_26_896 ();
 sg13g2_fill_8 FILLER_26_904 ();
 sg13g2_fill_8 FILLER_26_912 ();
 sg13g2_fill_8 FILLER_26_920 ();
 sg13g2_fill_8 FILLER_26_928 ();
 sg13g2_fill_8 FILLER_26_936 ();
 sg13g2_fill_8 FILLER_26_944 ();
 sg13g2_fill_8 FILLER_26_952 ();
 sg13g2_fill_8 FILLER_26_960 ();
 sg13g2_fill_8 FILLER_26_968 ();
 sg13g2_fill_8 FILLER_26_976 ();
 sg13g2_fill_8 FILLER_26_984 ();
 sg13g2_fill_8 FILLER_26_992 ();
 sg13g2_fill_8 FILLER_26_1000 ();
 sg13g2_fill_8 FILLER_26_1008 ();
 sg13g2_fill_8 FILLER_26_1016 ();
 sg13g2_fill_8 FILLER_26_1024 ();
 sg13g2_fill_8 FILLER_26_1032 ();
 sg13g2_fill_8 FILLER_26_1040 ();
 sg13g2_fill_8 FILLER_26_1048 ();
 sg13g2_fill_8 FILLER_26_1056 ();
 sg13g2_fill_8 FILLER_26_1064 ();
 sg13g2_fill_8 FILLER_26_1072 ();
 sg13g2_fill_8 FILLER_26_1080 ();
 sg13g2_fill_8 FILLER_26_1088 ();
 sg13g2_fill_8 FILLER_26_1096 ();
 sg13g2_fill_8 FILLER_26_1104 ();
 sg13g2_fill_8 FILLER_26_1112 ();
 sg13g2_fill_8 FILLER_26_1120 ();
 sg13g2_fill_8 FILLER_26_1128 ();
 sg13g2_fill_8 FILLER_26_1136 ();
 sg13g2_fill_8 FILLER_27_0 ();
 sg13g2_fill_8 FILLER_27_8 ();
 sg13g2_fill_8 FILLER_27_16 ();
 sg13g2_fill_8 FILLER_27_24 ();
 sg13g2_fill_8 FILLER_27_32 ();
 sg13g2_fill_8 FILLER_27_40 ();
 sg13g2_fill_8 FILLER_27_48 ();
 sg13g2_fill_8 FILLER_27_56 ();
 sg13g2_fill_8 FILLER_27_64 ();
 sg13g2_fill_8 FILLER_27_72 ();
 sg13g2_fill_8 FILLER_27_80 ();
 sg13g2_fill_8 FILLER_27_88 ();
 sg13g2_fill_8 FILLER_27_96 ();
 sg13g2_fill_8 FILLER_27_104 ();
 sg13g2_fill_8 FILLER_27_112 ();
 sg13g2_fill_8 FILLER_27_120 ();
 sg13g2_fill_8 FILLER_27_128 ();
 sg13g2_fill_8 FILLER_27_136 ();
 sg13g2_fill_8 FILLER_27_144 ();
 sg13g2_fill_8 FILLER_27_152 ();
 sg13g2_fill_8 FILLER_27_160 ();
 sg13g2_fill_8 FILLER_27_168 ();
 sg13g2_fill_8 FILLER_27_176 ();
 sg13g2_fill_8 FILLER_27_184 ();
 sg13g2_fill_8 FILLER_27_192 ();
 sg13g2_fill_8 FILLER_27_200 ();
 sg13g2_fill_8 FILLER_27_208 ();
 sg13g2_fill_8 FILLER_27_216 ();
 sg13g2_fill_8 FILLER_27_224 ();
 sg13g2_fill_8 FILLER_27_232 ();
 sg13g2_fill_8 FILLER_27_240 ();
 sg13g2_fill_8 FILLER_27_248 ();
 sg13g2_fill_8 FILLER_27_256 ();
 sg13g2_fill_8 FILLER_27_264 ();
 sg13g2_fill_8 FILLER_27_272 ();
 sg13g2_fill_8 FILLER_27_280 ();
 sg13g2_fill_8 FILLER_27_288 ();
 sg13g2_fill_8 FILLER_27_296 ();
 sg13g2_fill_8 FILLER_27_304 ();
 sg13g2_fill_8 FILLER_27_312 ();
 sg13g2_fill_8 FILLER_27_320 ();
 sg13g2_fill_8 FILLER_27_328 ();
 sg13g2_fill_8 FILLER_27_336 ();
 sg13g2_fill_8 FILLER_27_344 ();
 sg13g2_fill_8 FILLER_27_352 ();
 sg13g2_fill_8 FILLER_27_360 ();
 sg13g2_fill_8 FILLER_27_368 ();
 sg13g2_fill_8 FILLER_27_376 ();
 sg13g2_fill_8 FILLER_27_384 ();
 sg13g2_fill_8 FILLER_27_392 ();
 sg13g2_fill_8 FILLER_27_400 ();
 sg13g2_fill_8 FILLER_27_408 ();
 sg13g2_fill_8 FILLER_27_416 ();
 sg13g2_fill_8 FILLER_27_424 ();
 sg13g2_fill_8 FILLER_27_432 ();
 sg13g2_fill_8 FILLER_27_440 ();
 sg13g2_fill_8 FILLER_27_448 ();
 sg13g2_fill_8 FILLER_27_456 ();
 sg13g2_fill_8 FILLER_27_464 ();
 sg13g2_fill_8 FILLER_27_472 ();
 sg13g2_fill_8 FILLER_27_480 ();
 sg13g2_fill_8 FILLER_27_488 ();
 sg13g2_fill_8 FILLER_27_496 ();
 sg13g2_fill_8 FILLER_27_504 ();
 sg13g2_fill_8 FILLER_27_512 ();
 sg13g2_fill_8 FILLER_27_520 ();
 sg13g2_fill_8 FILLER_27_528 ();
 sg13g2_fill_8 FILLER_27_536 ();
 sg13g2_fill_8 FILLER_27_544 ();
 sg13g2_fill_8 FILLER_27_552 ();
 sg13g2_fill_8 FILLER_27_560 ();
 sg13g2_fill_8 FILLER_27_568 ();
 sg13g2_fill_8 FILLER_27_576 ();
 sg13g2_fill_8 FILLER_27_584 ();
 sg13g2_fill_8 FILLER_27_592 ();
 sg13g2_fill_8 FILLER_27_600 ();
 sg13g2_fill_8 FILLER_27_608 ();
 sg13g2_fill_8 FILLER_27_616 ();
 sg13g2_fill_8 FILLER_27_624 ();
 sg13g2_fill_8 FILLER_27_632 ();
 sg13g2_fill_8 FILLER_27_640 ();
 sg13g2_fill_8 FILLER_27_648 ();
 sg13g2_fill_8 FILLER_27_656 ();
 sg13g2_fill_8 FILLER_27_664 ();
 sg13g2_fill_8 FILLER_27_672 ();
 sg13g2_fill_8 FILLER_27_680 ();
 sg13g2_fill_8 FILLER_27_688 ();
 sg13g2_fill_8 FILLER_27_696 ();
 sg13g2_fill_8 FILLER_27_704 ();
 sg13g2_fill_8 FILLER_27_712 ();
 sg13g2_fill_8 FILLER_27_720 ();
 sg13g2_fill_8 FILLER_27_728 ();
 sg13g2_fill_8 FILLER_27_736 ();
 sg13g2_fill_8 FILLER_27_744 ();
 sg13g2_fill_8 FILLER_27_752 ();
 sg13g2_fill_8 FILLER_27_760 ();
 sg13g2_fill_8 FILLER_27_768 ();
 sg13g2_fill_8 FILLER_27_776 ();
 sg13g2_fill_8 FILLER_27_784 ();
 sg13g2_fill_8 FILLER_27_792 ();
 sg13g2_fill_8 FILLER_27_800 ();
 sg13g2_fill_8 FILLER_27_808 ();
 sg13g2_fill_8 FILLER_27_816 ();
 sg13g2_fill_8 FILLER_27_824 ();
 sg13g2_fill_8 FILLER_27_832 ();
 sg13g2_fill_8 FILLER_27_840 ();
 sg13g2_fill_8 FILLER_27_848 ();
 sg13g2_fill_8 FILLER_27_856 ();
 sg13g2_fill_8 FILLER_27_864 ();
 sg13g2_fill_8 FILLER_27_872 ();
 sg13g2_fill_8 FILLER_27_880 ();
 sg13g2_fill_8 FILLER_27_888 ();
 sg13g2_fill_8 FILLER_27_896 ();
 sg13g2_fill_8 FILLER_27_904 ();
 sg13g2_fill_8 FILLER_27_912 ();
 sg13g2_fill_8 FILLER_27_920 ();
 sg13g2_fill_8 FILLER_27_928 ();
 sg13g2_fill_8 FILLER_27_936 ();
 sg13g2_fill_8 FILLER_27_944 ();
 sg13g2_fill_8 FILLER_27_952 ();
 sg13g2_fill_8 FILLER_27_960 ();
 sg13g2_fill_8 FILLER_27_968 ();
 sg13g2_fill_8 FILLER_27_976 ();
 sg13g2_fill_8 FILLER_27_984 ();
 sg13g2_fill_8 FILLER_27_992 ();
 sg13g2_fill_8 FILLER_27_1000 ();
 sg13g2_fill_8 FILLER_27_1008 ();
 sg13g2_fill_8 FILLER_27_1016 ();
 sg13g2_fill_8 FILLER_27_1024 ();
 sg13g2_fill_8 FILLER_27_1032 ();
 sg13g2_fill_8 FILLER_27_1040 ();
 sg13g2_fill_8 FILLER_27_1048 ();
 sg13g2_fill_8 FILLER_27_1056 ();
 sg13g2_fill_8 FILLER_27_1064 ();
 sg13g2_fill_8 FILLER_27_1072 ();
 sg13g2_fill_8 FILLER_27_1080 ();
 sg13g2_fill_8 FILLER_27_1088 ();
 sg13g2_fill_8 FILLER_27_1096 ();
 sg13g2_fill_8 FILLER_27_1104 ();
 sg13g2_fill_8 FILLER_27_1112 ();
 sg13g2_fill_8 FILLER_27_1120 ();
 sg13g2_fill_8 FILLER_27_1128 ();
 sg13g2_fill_8 FILLER_27_1136 ();
 sg13g2_fill_8 FILLER_28_0 ();
 sg13g2_fill_8 FILLER_28_8 ();
 sg13g2_fill_8 FILLER_28_16 ();
 sg13g2_fill_8 FILLER_28_24 ();
 sg13g2_fill_8 FILLER_28_32 ();
 sg13g2_fill_8 FILLER_28_40 ();
 sg13g2_fill_8 FILLER_28_48 ();
 sg13g2_fill_8 FILLER_28_56 ();
 sg13g2_fill_8 FILLER_28_64 ();
 sg13g2_fill_8 FILLER_28_72 ();
 sg13g2_fill_8 FILLER_28_80 ();
 sg13g2_fill_8 FILLER_28_88 ();
 sg13g2_fill_8 FILLER_28_96 ();
 sg13g2_fill_8 FILLER_28_104 ();
 sg13g2_fill_8 FILLER_28_112 ();
 sg13g2_fill_8 FILLER_28_120 ();
 sg13g2_fill_8 FILLER_28_128 ();
 sg13g2_fill_8 FILLER_28_136 ();
 sg13g2_fill_8 FILLER_28_144 ();
 sg13g2_fill_8 FILLER_28_152 ();
 sg13g2_fill_8 FILLER_28_160 ();
 sg13g2_fill_8 FILLER_28_168 ();
 sg13g2_fill_8 FILLER_28_176 ();
 sg13g2_fill_8 FILLER_28_184 ();
 sg13g2_fill_8 FILLER_28_192 ();
 sg13g2_fill_8 FILLER_28_200 ();
 sg13g2_fill_8 FILLER_28_208 ();
 sg13g2_fill_8 FILLER_28_216 ();
 sg13g2_fill_8 FILLER_28_224 ();
 sg13g2_fill_8 FILLER_28_232 ();
 sg13g2_fill_8 FILLER_28_240 ();
 sg13g2_fill_8 FILLER_28_248 ();
 sg13g2_fill_8 FILLER_28_256 ();
 sg13g2_fill_8 FILLER_28_264 ();
 sg13g2_fill_8 FILLER_28_272 ();
 sg13g2_fill_8 FILLER_28_280 ();
 sg13g2_fill_8 FILLER_28_288 ();
 sg13g2_fill_8 FILLER_28_296 ();
 sg13g2_fill_8 FILLER_28_304 ();
 sg13g2_fill_8 FILLER_28_312 ();
 sg13g2_fill_8 FILLER_28_320 ();
 sg13g2_fill_8 FILLER_28_328 ();
 sg13g2_fill_8 FILLER_28_336 ();
 sg13g2_fill_8 FILLER_28_344 ();
 sg13g2_fill_8 FILLER_28_352 ();
 sg13g2_fill_8 FILLER_28_360 ();
 sg13g2_fill_8 FILLER_28_368 ();
 sg13g2_fill_8 FILLER_28_376 ();
 sg13g2_fill_8 FILLER_28_384 ();
 sg13g2_fill_8 FILLER_28_392 ();
 sg13g2_fill_8 FILLER_28_400 ();
 sg13g2_fill_8 FILLER_28_408 ();
 sg13g2_fill_8 FILLER_28_416 ();
 sg13g2_fill_8 FILLER_28_424 ();
 sg13g2_fill_8 FILLER_28_432 ();
 sg13g2_fill_8 FILLER_28_440 ();
 sg13g2_fill_8 FILLER_28_448 ();
 sg13g2_fill_8 FILLER_28_456 ();
 sg13g2_fill_8 FILLER_28_464 ();
 sg13g2_fill_8 FILLER_28_472 ();
 sg13g2_fill_8 FILLER_28_480 ();
 sg13g2_fill_8 FILLER_28_488 ();
 sg13g2_fill_8 FILLER_28_496 ();
 sg13g2_fill_8 FILLER_28_504 ();
 sg13g2_fill_8 FILLER_28_512 ();
 sg13g2_fill_8 FILLER_28_520 ();
 sg13g2_fill_8 FILLER_28_528 ();
 sg13g2_fill_8 FILLER_28_536 ();
 sg13g2_fill_8 FILLER_28_544 ();
 sg13g2_fill_8 FILLER_28_552 ();
 sg13g2_fill_8 FILLER_28_560 ();
 sg13g2_fill_8 FILLER_28_568 ();
 sg13g2_fill_8 FILLER_28_576 ();
 sg13g2_fill_8 FILLER_28_584 ();
 sg13g2_fill_8 FILLER_28_592 ();
 sg13g2_fill_8 FILLER_28_600 ();
 sg13g2_fill_8 FILLER_28_608 ();
 sg13g2_fill_8 FILLER_28_616 ();
 sg13g2_fill_8 FILLER_28_624 ();
 sg13g2_fill_8 FILLER_28_632 ();
 sg13g2_fill_8 FILLER_28_640 ();
 sg13g2_fill_8 FILLER_28_648 ();
 sg13g2_fill_8 FILLER_28_656 ();
 sg13g2_fill_8 FILLER_28_664 ();
 sg13g2_fill_8 FILLER_28_672 ();
 sg13g2_fill_8 FILLER_28_680 ();
 sg13g2_fill_8 FILLER_28_688 ();
 sg13g2_fill_8 FILLER_28_696 ();
 sg13g2_fill_8 FILLER_28_704 ();
 sg13g2_fill_8 FILLER_28_712 ();
 sg13g2_fill_8 FILLER_28_720 ();
 sg13g2_fill_8 FILLER_28_728 ();
 sg13g2_fill_8 FILLER_28_736 ();
 sg13g2_fill_8 FILLER_28_744 ();
 sg13g2_fill_8 FILLER_28_752 ();
 sg13g2_fill_8 FILLER_28_760 ();
 sg13g2_fill_8 FILLER_28_768 ();
 sg13g2_fill_8 FILLER_28_776 ();
 sg13g2_fill_8 FILLER_28_784 ();
 sg13g2_fill_8 FILLER_28_792 ();
 sg13g2_fill_8 FILLER_28_800 ();
 sg13g2_fill_8 FILLER_28_808 ();
 sg13g2_fill_8 FILLER_28_816 ();
 sg13g2_fill_8 FILLER_28_824 ();
 sg13g2_fill_8 FILLER_28_832 ();
 sg13g2_fill_8 FILLER_28_840 ();
 sg13g2_fill_8 FILLER_28_848 ();
 sg13g2_fill_8 FILLER_28_856 ();
 sg13g2_fill_8 FILLER_28_864 ();
 sg13g2_fill_8 FILLER_28_872 ();
 sg13g2_fill_8 FILLER_28_880 ();
 sg13g2_fill_8 FILLER_28_888 ();
 sg13g2_fill_8 FILLER_28_896 ();
 sg13g2_fill_8 FILLER_28_904 ();
 sg13g2_fill_8 FILLER_28_912 ();
 sg13g2_fill_8 FILLER_28_920 ();
 sg13g2_fill_8 FILLER_28_928 ();
 sg13g2_fill_8 FILLER_28_936 ();
 sg13g2_fill_8 FILLER_28_944 ();
 sg13g2_fill_8 FILLER_28_952 ();
 sg13g2_fill_8 FILLER_28_960 ();
 sg13g2_fill_8 FILLER_28_968 ();
 sg13g2_fill_8 FILLER_28_976 ();
 sg13g2_fill_8 FILLER_28_984 ();
 sg13g2_fill_8 FILLER_28_992 ();
 sg13g2_fill_8 FILLER_28_1000 ();
 sg13g2_fill_8 FILLER_28_1008 ();
 sg13g2_fill_8 FILLER_28_1016 ();
 sg13g2_fill_8 FILLER_28_1024 ();
 sg13g2_fill_8 FILLER_28_1032 ();
 sg13g2_fill_8 FILLER_28_1040 ();
 sg13g2_fill_8 FILLER_28_1048 ();
 sg13g2_fill_8 FILLER_28_1056 ();
 sg13g2_fill_8 FILLER_28_1064 ();
 sg13g2_fill_8 FILLER_28_1072 ();
 sg13g2_fill_8 FILLER_28_1080 ();
 sg13g2_fill_8 FILLER_28_1088 ();
 sg13g2_fill_8 FILLER_28_1096 ();
 sg13g2_fill_8 FILLER_28_1104 ();
 sg13g2_fill_8 FILLER_28_1112 ();
 sg13g2_fill_8 FILLER_28_1120 ();
 sg13g2_fill_8 FILLER_28_1128 ();
 sg13g2_fill_8 FILLER_28_1136 ();
 sg13g2_fill_8 FILLER_29_0 ();
 sg13g2_fill_8 FILLER_29_8 ();
 sg13g2_fill_8 FILLER_29_16 ();
 sg13g2_fill_8 FILLER_29_24 ();
 sg13g2_fill_8 FILLER_29_32 ();
 sg13g2_fill_8 FILLER_29_40 ();
 sg13g2_fill_8 FILLER_29_48 ();
 sg13g2_fill_8 FILLER_29_56 ();
 sg13g2_fill_8 FILLER_29_64 ();
 sg13g2_fill_8 FILLER_29_72 ();
 sg13g2_fill_8 FILLER_29_80 ();
 sg13g2_fill_8 FILLER_29_88 ();
 sg13g2_fill_8 FILLER_29_96 ();
 sg13g2_fill_8 FILLER_29_104 ();
 sg13g2_fill_8 FILLER_29_112 ();
 sg13g2_fill_8 FILLER_29_120 ();
 sg13g2_fill_8 FILLER_29_128 ();
 sg13g2_fill_8 FILLER_29_136 ();
 sg13g2_fill_8 FILLER_29_144 ();
 sg13g2_fill_8 FILLER_29_152 ();
 sg13g2_fill_8 FILLER_29_160 ();
 sg13g2_fill_8 FILLER_29_168 ();
 sg13g2_fill_8 FILLER_29_176 ();
 sg13g2_fill_8 FILLER_29_184 ();
 sg13g2_fill_8 FILLER_29_192 ();
 sg13g2_fill_8 FILLER_29_200 ();
 sg13g2_fill_8 FILLER_29_208 ();
 sg13g2_fill_8 FILLER_29_216 ();
 sg13g2_fill_8 FILLER_29_224 ();
 sg13g2_fill_8 FILLER_29_232 ();
 sg13g2_fill_8 FILLER_29_240 ();
 sg13g2_fill_8 FILLER_29_248 ();
 sg13g2_fill_8 FILLER_29_256 ();
 sg13g2_fill_8 FILLER_29_264 ();
 sg13g2_fill_8 FILLER_29_272 ();
 sg13g2_fill_8 FILLER_29_280 ();
 sg13g2_fill_8 FILLER_29_288 ();
 sg13g2_fill_8 FILLER_29_296 ();
 sg13g2_fill_8 FILLER_29_304 ();
 sg13g2_fill_8 FILLER_29_312 ();
 sg13g2_fill_8 FILLER_29_320 ();
 sg13g2_fill_8 FILLER_29_328 ();
 sg13g2_fill_8 FILLER_29_336 ();
 sg13g2_fill_8 FILLER_29_344 ();
 sg13g2_fill_8 FILLER_29_352 ();
 sg13g2_fill_8 FILLER_29_360 ();
 sg13g2_fill_8 FILLER_29_368 ();
 sg13g2_fill_8 FILLER_29_376 ();
 sg13g2_fill_8 FILLER_29_384 ();
 sg13g2_fill_8 FILLER_29_392 ();
 sg13g2_fill_8 FILLER_29_400 ();
 sg13g2_fill_8 FILLER_29_408 ();
 sg13g2_fill_8 FILLER_29_416 ();
 sg13g2_fill_8 FILLER_29_424 ();
 sg13g2_fill_8 FILLER_29_432 ();
 sg13g2_fill_8 FILLER_29_440 ();
 sg13g2_fill_8 FILLER_29_448 ();
 sg13g2_fill_8 FILLER_29_456 ();
 sg13g2_fill_8 FILLER_29_464 ();
 sg13g2_fill_8 FILLER_29_472 ();
 sg13g2_fill_8 FILLER_29_480 ();
 sg13g2_fill_8 FILLER_29_488 ();
 sg13g2_fill_8 FILLER_29_496 ();
 sg13g2_fill_8 FILLER_29_504 ();
 sg13g2_fill_8 FILLER_29_512 ();
 sg13g2_fill_8 FILLER_29_520 ();
 sg13g2_fill_8 FILLER_29_528 ();
 sg13g2_fill_8 FILLER_29_536 ();
 sg13g2_fill_8 FILLER_29_544 ();
 sg13g2_fill_8 FILLER_29_552 ();
 sg13g2_fill_8 FILLER_29_560 ();
 sg13g2_fill_8 FILLER_29_568 ();
 sg13g2_fill_8 FILLER_29_576 ();
 sg13g2_fill_8 FILLER_29_584 ();
 sg13g2_fill_8 FILLER_29_592 ();
 sg13g2_fill_8 FILLER_29_600 ();
 sg13g2_fill_8 FILLER_29_608 ();
 sg13g2_fill_8 FILLER_29_616 ();
 sg13g2_fill_8 FILLER_29_624 ();
 sg13g2_fill_8 FILLER_29_632 ();
 sg13g2_fill_8 FILLER_29_640 ();
 sg13g2_fill_8 FILLER_29_648 ();
 sg13g2_fill_8 FILLER_29_656 ();
 sg13g2_fill_8 FILLER_29_664 ();
 sg13g2_fill_8 FILLER_29_672 ();
 sg13g2_fill_8 FILLER_29_680 ();
 sg13g2_fill_8 FILLER_29_688 ();
 sg13g2_fill_8 FILLER_29_696 ();
 sg13g2_fill_8 FILLER_29_704 ();
 sg13g2_fill_8 FILLER_29_712 ();
 sg13g2_fill_8 FILLER_29_720 ();
 sg13g2_fill_8 FILLER_29_728 ();
 sg13g2_fill_8 FILLER_29_736 ();
 sg13g2_fill_8 FILLER_29_744 ();
 sg13g2_fill_8 FILLER_29_752 ();
 sg13g2_fill_8 FILLER_29_760 ();
 sg13g2_fill_8 FILLER_29_768 ();
 sg13g2_fill_8 FILLER_29_776 ();
 sg13g2_fill_8 FILLER_29_784 ();
 sg13g2_fill_8 FILLER_29_792 ();
 sg13g2_fill_8 FILLER_29_800 ();
 sg13g2_fill_8 FILLER_29_808 ();
 sg13g2_fill_8 FILLER_29_816 ();
 sg13g2_fill_8 FILLER_29_824 ();
 sg13g2_fill_8 FILLER_29_832 ();
 sg13g2_fill_8 FILLER_29_840 ();
 sg13g2_fill_8 FILLER_29_848 ();
 sg13g2_fill_8 FILLER_29_856 ();
 sg13g2_fill_8 FILLER_29_864 ();
 sg13g2_fill_8 FILLER_29_872 ();
 sg13g2_fill_8 FILLER_29_880 ();
 sg13g2_fill_8 FILLER_29_888 ();
 sg13g2_fill_8 FILLER_29_896 ();
 sg13g2_fill_8 FILLER_29_904 ();
 sg13g2_fill_8 FILLER_29_912 ();
 sg13g2_fill_8 FILLER_29_920 ();
 sg13g2_fill_8 FILLER_29_928 ();
 sg13g2_fill_8 FILLER_29_936 ();
 sg13g2_fill_8 FILLER_29_944 ();
 sg13g2_fill_8 FILLER_29_952 ();
 sg13g2_fill_8 FILLER_29_960 ();
 sg13g2_fill_8 FILLER_29_968 ();
 sg13g2_fill_8 FILLER_29_976 ();
 sg13g2_fill_8 FILLER_29_984 ();
 sg13g2_fill_8 FILLER_29_992 ();
 sg13g2_fill_8 FILLER_29_1000 ();
 sg13g2_fill_8 FILLER_29_1008 ();
 sg13g2_fill_8 FILLER_29_1016 ();
 sg13g2_fill_8 FILLER_29_1024 ();
 sg13g2_fill_8 FILLER_29_1032 ();
 sg13g2_fill_8 FILLER_29_1040 ();
 sg13g2_fill_8 FILLER_29_1048 ();
 sg13g2_fill_8 FILLER_29_1056 ();
 sg13g2_fill_8 FILLER_29_1064 ();
 sg13g2_fill_8 FILLER_29_1072 ();
 sg13g2_fill_8 FILLER_29_1080 ();
 sg13g2_fill_8 FILLER_29_1088 ();
 sg13g2_fill_8 FILLER_29_1096 ();
 sg13g2_fill_8 FILLER_29_1104 ();
 sg13g2_fill_8 FILLER_29_1112 ();
 sg13g2_fill_8 FILLER_29_1120 ();
 sg13g2_fill_8 FILLER_29_1128 ();
 sg13g2_fill_8 FILLER_29_1136 ();
 sg13g2_fill_8 FILLER_30_0 ();
 sg13g2_fill_8 FILLER_30_8 ();
 sg13g2_fill_8 FILLER_30_16 ();
 sg13g2_fill_8 FILLER_30_24 ();
 sg13g2_fill_8 FILLER_30_32 ();
 sg13g2_fill_8 FILLER_30_40 ();
 sg13g2_fill_8 FILLER_30_48 ();
 sg13g2_fill_8 FILLER_30_56 ();
 sg13g2_fill_8 FILLER_30_64 ();
 sg13g2_fill_8 FILLER_30_72 ();
 sg13g2_fill_8 FILLER_30_80 ();
 sg13g2_fill_8 FILLER_30_88 ();
 sg13g2_fill_8 FILLER_30_96 ();
 sg13g2_fill_8 FILLER_30_104 ();
 sg13g2_fill_8 FILLER_30_112 ();
 sg13g2_fill_8 FILLER_30_120 ();
 sg13g2_fill_8 FILLER_30_128 ();
 sg13g2_fill_8 FILLER_30_136 ();
 sg13g2_fill_8 FILLER_30_144 ();
 sg13g2_fill_8 FILLER_30_152 ();
 sg13g2_fill_8 FILLER_30_160 ();
 sg13g2_fill_8 FILLER_30_168 ();
 sg13g2_fill_8 FILLER_30_176 ();
 sg13g2_fill_8 FILLER_30_184 ();
 sg13g2_fill_8 FILLER_30_192 ();
 sg13g2_fill_8 FILLER_30_200 ();
 sg13g2_fill_8 FILLER_30_208 ();
 sg13g2_fill_8 FILLER_30_216 ();
 sg13g2_fill_8 FILLER_30_224 ();
 sg13g2_fill_8 FILLER_30_232 ();
 sg13g2_fill_8 FILLER_30_240 ();
 sg13g2_fill_8 FILLER_30_248 ();
 sg13g2_fill_8 FILLER_30_256 ();
 sg13g2_fill_8 FILLER_30_264 ();
 sg13g2_fill_8 FILLER_30_272 ();
 sg13g2_fill_8 FILLER_30_280 ();
 sg13g2_fill_8 FILLER_30_288 ();
 sg13g2_fill_8 FILLER_30_296 ();
 sg13g2_fill_8 FILLER_30_304 ();
 sg13g2_fill_8 FILLER_30_312 ();
 sg13g2_fill_8 FILLER_30_320 ();
 sg13g2_fill_8 FILLER_30_328 ();
 sg13g2_fill_8 FILLER_30_336 ();
 sg13g2_fill_8 FILLER_30_344 ();
 sg13g2_fill_8 FILLER_30_352 ();
 sg13g2_fill_8 FILLER_30_360 ();
 sg13g2_fill_8 FILLER_30_368 ();
 sg13g2_fill_8 FILLER_30_376 ();
 sg13g2_fill_8 FILLER_30_384 ();
 sg13g2_fill_8 FILLER_30_392 ();
 sg13g2_fill_8 FILLER_30_400 ();
 sg13g2_fill_8 FILLER_30_408 ();
 sg13g2_fill_8 FILLER_30_416 ();
 sg13g2_fill_8 FILLER_30_424 ();
 sg13g2_fill_8 FILLER_30_432 ();
 sg13g2_fill_8 FILLER_30_440 ();
 sg13g2_fill_8 FILLER_30_448 ();
 sg13g2_fill_8 FILLER_30_456 ();
 sg13g2_fill_8 FILLER_30_464 ();
 sg13g2_fill_8 FILLER_30_472 ();
 sg13g2_fill_8 FILLER_30_480 ();
 sg13g2_fill_8 FILLER_30_488 ();
 sg13g2_fill_8 FILLER_30_496 ();
 sg13g2_fill_8 FILLER_30_504 ();
 sg13g2_fill_8 FILLER_30_512 ();
 sg13g2_fill_8 FILLER_30_520 ();
 sg13g2_fill_8 FILLER_30_528 ();
 sg13g2_fill_8 FILLER_30_536 ();
 sg13g2_fill_8 FILLER_30_544 ();
 sg13g2_fill_8 FILLER_30_552 ();
 sg13g2_fill_8 FILLER_30_560 ();
 sg13g2_fill_8 FILLER_30_568 ();
 sg13g2_fill_8 FILLER_30_576 ();
 sg13g2_fill_8 FILLER_30_584 ();
 sg13g2_fill_8 FILLER_30_592 ();
 sg13g2_fill_8 FILLER_30_600 ();
 sg13g2_fill_8 FILLER_30_608 ();
 sg13g2_fill_8 FILLER_30_616 ();
 sg13g2_fill_8 FILLER_30_624 ();
 sg13g2_fill_8 FILLER_30_632 ();
 sg13g2_fill_8 FILLER_30_640 ();
 sg13g2_fill_8 FILLER_30_648 ();
 sg13g2_fill_8 FILLER_30_656 ();
 sg13g2_fill_8 FILLER_30_664 ();
 sg13g2_fill_8 FILLER_30_672 ();
 sg13g2_fill_8 FILLER_30_680 ();
 sg13g2_fill_8 FILLER_30_688 ();
 sg13g2_fill_8 FILLER_30_696 ();
 sg13g2_fill_8 FILLER_30_704 ();
 sg13g2_fill_8 FILLER_30_712 ();
 sg13g2_fill_8 FILLER_30_720 ();
 sg13g2_fill_8 FILLER_30_728 ();
 sg13g2_fill_8 FILLER_30_736 ();
 sg13g2_fill_8 FILLER_30_744 ();
 sg13g2_fill_8 FILLER_30_752 ();
 sg13g2_fill_8 FILLER_30_760 ();
 sg13g2_fill_8 FILLER_30_768 ();
 sg13g2_fill_8 FILLER_30_776 ();
 sg13g2_fill_8 FILLER_30_784 ();
 sg13g2_fill_8 FILLER_30_792 ();
 sg13g2_fill_8 FILLER_30_800 ();
 sg13g2_fill_8 FILLER_30_808 ();
 sg13g2_fill_8 FILLER_30_816 ();
 sg13g2_fill_8 FILLER_30_824 ();
 sg13g2_fill_8 FILLER_30_832 ();
 sg13g2_fill_8 FILLER_30_840 ();
 sg13g2_fill_8 FILLER_30_848 ();
 sg13g2_fill_8 FILLER_30_856 ();
 sg13g2_fill_8 FILLER_30_864 ();
 sg13g2_fill_8 FILLER_30_872 ();
 sg13g2_fill_8 FILLER_30_880 ();
 sg13g2_fill_8 FILLER_30_888 ();
 sg13g2_fill_8 FILLER_30_896 ();
 sg13g2_fill_8 FILLER_30_904 ();
 sg13g2_fill_8 FILLER_30_912 ();
 sg13g2_fill_8 FILLER_30_920 ();
 sg13g2_fill_8 FILLER_30_928 ();
 sg13g2_fill_8 FILLER_30_936 ();
 sg13g2_fill_8 FILLER_30_944 ();
 sg13g2_fill_8 FILLER_30_952 ();
 sg13g2_fill_8 FILLER_30_960 ();
 sg13g2_fill_8 FILLER_30_968 ();
 sg13g2_fill_8 FILLER_30_976 ();
 sg13g2_fill_8 FILLER_30_984 ();
 sg13g2_fill_8 FILLER_30_992 ();
 sg13g2_fill_8 FILLER_30_1000 ();
 sg13g2_fill_8 FILLER_30_1008 ();
 sg13g2_fill_8 FILLER_30_1016 ();
 sg13g2_fill_8 FILLER_30_1024 ();
 sg13g2_fill_8 FILLER_30_1032 ();
 sg13g2_fill_8 FILLER_30_1040 ();
 sg13g2_fill_8 FILLER_30_1048 ();
 sg13g2_fill_8 FILLER_30_1056 ();
 sg13g2_fill_8 FILLER_30_1064 ();
 sg13g2_fill_8 FILLER_30_1072 ();
 sg13g2_fill_8 FILLER_30_1080 ();
 sg13g2_fill_8 FILLER_30_1088 ();
 sg13g2_fill_8 FILLER_30_1096 ();
 sg13g2_fill_8 FILLER_30_1104 ();
 sg13g2_fill_8 FILLER_30_1112 ();
 sg13g2_fill_8 FILLER_30_1120 ();
 sg13g2_fill_8 FILLER_30_1128 ();
 sg13g2_fill_8 FILLER_30_1136 ();
 sg13g2_fill_8 FILLER_31_0 ();
 sg13g2_fill_8 FILLER_31_8 ();
 sg13g2_fill_8 FILLER_31_16 ();
 sg13g2_fill_8 FILLER_31_24 ();
 sg13g2_fill_8 FILLER_31_32 ();
 sg13g2_fill_8 FILLER_31_40 ();
 sg13g2_fill_8 FILLER_31_48 ();
 sg13g2_fill_8 FILLER_31_56 ();
 sg13g2_fill_8 FILLER_31_64 ();
 sg13g2_fill_8 FILLER_31_72 ();
 sg13g2_fill_8 FILLER_31_80 ();
 sg13g2_fill_8 FILLER_31_88 ();
 sg13g2_fill_8 FILLER_31_96 ();
 sg13g2_fill_8 FILLER_31_104 ();
 sg13g2_fill_8 FILLER_31_112 ();
 sg13g2_fill_8 FILLER_31_120 ();
 sg13g2_fill_8 FILLER_31_128 ();
 sg13g2_fill_8 FILLER_31_136 ();
 sg13g2_fill_8 FILLER_31_144 ();
 sg13g2_fill_8 FILLER_31_152 ();
 sg13g2_fill_8 FILLER_31_160 ();
 sg13g2_fill_8 FILLER_31_168 ();
 sg13g2_fill_8 FILLER_31_176 ();
 sg13g2_fill_8 FILLER_31_184 ();
 sg13g2_fill_8 FILLER_31_192 ();
 sg13g2_fill_8 FILLER_31_200 ();
 sg13g2_fill_8 FILLER_31_208 ();
 sg13g2_fill_8 FILLER_31_216 ();
 sg13g2_fill_8 FILLER_31_224 ();
 sg13g2_fill_8 FILLER_31_232 ();
 sg13g2_fill_8 FILLER_31_240 ();
 sg13g2_fill_8 FILLER_31_248 ();
 sg13g2_fill_8 FILLER_31_256 ();
 sg13g2_fill_8 FILLER_31_264 ();
 sg13g2_fill_8 FILLER_31_272 ();
 sg13g2_fill_8 FILLER_31_280 ();
 sg13g2_fill_8 FILLER_31_288 ();
 sg13g2_fill_8 FILLER_31_296 ();
 sg13g2_fill_8 FILLER_31_304 ();
 sg13g2_fill_8 FILLER_31_312 ();
 sg13g2_fill_8 FILLER_31_320 ();
 sg13g2_fill_8 FILLER_31_328 ();
 sg13g2_fill_8 FILLER_31_336 ();
 sg13g2_fill_8 FILLER_31_344 ();
 sg13g2_fill_8 FILLER_31_352 ();
 sg13g2_fill_8 FILLER_31_360 ();
 sg13g2_fill_8 FILLER_31_368 ();
 sg13g2_fill_8 FILLER_31_376 ();
 sg13g2_fill_8 FILLER_31_384 ();
 sg13g2_fill_8 FILLER_31_392 ();
 sg13g2_fill_8 FILLER_31_400 ();
 sg13g2_fill_8 FILLER_31_408 ();
 sg13g2_fill_8 FILLER_31_416 ();
 sg13g2_fill_8 FILLER_31_424 ();
 sg13g2_fill_8 FILLER_31_432 ();
 sg13g2_fill_8 FILLER_31_440 ();
 sg13g2_fill_8 FILLER_31_448 ();
 sg13g2_fill_8 FILLER_31_456 ();
 sg13g2_fill_8 FILLER_31_464 ();
 sg13g2_fill_8 FILLER_31_472 ();
 sg13g2_fill_8 FILLER_31_480 ();
 sg13g2_fill_8 FILLER_31_488 ();
 sg13g2_fill_8 FILLER_31_496 ();
 sg13g2_fill_8 FILLER_31_504 ();
 sg13g2_fill_8 FILLER_31_512 ();
 sg13g2_fill_8 FILLER_31_520 ();
 sg13g2_fill_8 FILLER_31_528 ();
 sg13g2_fill_8 FILLER_31_536 ();
 sg13g2_fill_8 FILLER_31_544 ();
 sg13g2_fill_8 FILLER_31_552 ();
 sg13g2_fill_8 FILLER_31_560 ();
 sg13g2_fill_8 FILLER_31_568 ();
 sg13g2_fill_8 FILLER_31_576 ();
 sg13g2_fill_8 FILLER_31_584 ();
 sg13g2_fill_8 FILLER_31_592 ();
 sg13g2_fill_8 FILLER_31_600 ();
 sg13g2_fill_8 FILLER_31_608 ();
 sg13g2_fill_8 FILLER_31_616 ();
 sg13g2_fill_8 FILLER_31_624 ();
 sg13g2_fill_8 FILLER_31_632 ();
 sg13g2_fill_8 FILLER_31_640 ();
 sg13g2_fill_8 FILLER_31_648 ();
 sg13g2_fill_8 FILLER_31_656 ();
 sg13g2_fill_8 FILLER_31_664 ();
 sg13g2_fill_8 FILLER_31_672 ();
 sg13g2_fill_8 FILLER_31_680 ();
 sg13g2_fill_8 FILLER_31_688 ();
 sg13g2_fill_8 FILLER_31_696 ();
 sg13g2_fill_8 FILLER_31_704 ();
 sg13g2_fill_8 FILLER_31_712 ();
 sg13g2_fill_8 FILLER_31_720 ();
 sg13g2_fill_8 FILLER_31_728 ();
 sg13g2_fill_8 FILLER_31_736 ();
 sg13g2_fill_8 FILLER_31_744 ();
 sg13g2_fill_8 FILLER_31_752 ();
 sg13g2_fill_8 FILLER_31_760 ();
 sg13g2_fill_8 FILLER_31_768 ();
 sg13g2_fill_8 FILLER_31_776 ();
 sg13g2_fill_8 FILLER_31_784 ();
 sg13g2_fill_8 FILLER_31_792 ();
 sg13g2_fill_8 FILLER_31_800 ();
 sg13g2_fill_8 FILLER_31_808 ();
 sg13g2_fill_8 FILLER_31_816 ();
 sg13g2_fill_8 FILLER_31_824 ();
 sg13g2_fill_8 FILLER_31_832 ();
 sg13g2_fill_8 FILLER_31_840 ();
 sg13g2_fill_8 FILLER_31_848 ();
 sg13g2_fill_8 FILLER_31_856 ();
 sg13g2_fill_8 FILLER_31_864 ();
 sg13g2_fill_8 FILLER_31_872 ();
 sg13g2_fill_8 FILLER_31_880 ();
 sg13g2_fill_8 FILLER_31_888 ();
 sg13g2_fill_8 FILLER_31_896 ();
 sg13g2_fill_8 FILLER_31_904 ();
 sg13g2_fill_8 FILLER_31_912 ();
 sg13g2_fill_8 FILLER_31_920 ();
 sg13g2_fill_8 FILLER_31_928 ();
 sg13g2_fill_8 FILLER_31_936 ();
 sg13g2_fill_8 FILLER_31_944 ();
 sg13g2_fill_8 FILLER_31_952 ();
 sg13g2_fill_8 FILLER_31_960 ();
 sg13g2_fill_8 FILLER_31_968 ();
 sg13g2_fill_8 FILLER_31_976 ();
 sg13g2_fill_8 FILLER_31_984 ();
 sg13g2_fill_8 FILLER_31_992 ();
 sg13g2_fill_8 FILLER_31_1000 ();
 sg13g2_fill_8 FILLER_31_1008 ();
 sg13g2_fill_8 FILLER_31_1016 ();
 sg13g2_fill_8 FILLER_31_1024 ();
 sg13g2_fill_8 FILLER_31_1032 ();
 sg13g2_fill_8 FILLER_31_1040 ();
 sg13g2_fill_8 FILLER_31_1048 ();
 sg13g2_fill_8 FILLER_31_1056 ();
 sg13g2_fill_8 FILLER_31_1064 ();
 sg13g2_fill_8 FILLER_31_1072 ();
 sg13g2_fill_8 FILLER_31_1080 ();
 sg13g2_fill_8 FILLER_31_1088 ();
 sg13g2_fill_8 FILLER_31_1096 ();
 sg13g2_fill_8 FILLER_31_1104 ();
 sg13g2_fill_8 FILLER_31_1112 ();
 sg13g2_fill_8 FILLER_31_1120 ();
 sg13g2_fill_8 FILLER_31_1128 ();
 sg13g2_fill_8 FILLER_31_1136 ();
 sg13g2_fill_8 FILLER_32_0 ();
 sg13g2_fill_8 FILLER_32_8 ();
 sg13g2_fill_8 FILLER_32_16 ();
 sg13g2_fill_8 FILLER_32_24 ();
 sg13g2_fill_8 FILLER_32_32 ();
 sg13g2_fill_8 FILLER_32_40 ();
 sg13g2_fill_8 FILLER_32_48 ();
 sg13g2_fill_8 FILLER_32_56 ();
 sg13g2_fill_8 FILLER_32_64 ();
 sg13g2_fill_8 FILLER_32_72 ();
 sg13g2_fill_8 FILLER_32_80 ();
 sg13g2_fill_8 FILLER_32_88 ();
 sg13g2_fill_8 FILLER_32_96 ();
 sg13g2_fill_8 FILLER_32_104 ();
 sg13g2_fill_8 FILLER_32_112 ();
 sg13g2_fill_8 FILLER_32_120 ();
 sg13g2_fill_8 FILLER_32_128 ();
 sg13g2_fill_8 FILLER_32_136 ();
 sg13g2_fill_8 FILLER_32_144 ();
 sg13g2_fill_8 FILLER_32_152 ();
 sg13g2_fill_8 FILLER_32_160 ();
 sg13g2_fill_8 FILLER_32_168 ();
 sg13g2_fill_8 FILLER_32_176 ();
 sg13g2_fill_8 FILLER_32_184 ();
 sg13g2_fill_8 FILLER_32_192 ();
 sg13g2_fill_8 FILLER_32_200 ();
 sg13g2_fill_8 FILLER_32_208 ();
 sg13g2_fill_8 FILLER_32_216 ();
 sg13g2_fill_8 FILLER_32_224 ();
 sg13g2_fill_8 FILLER_32_232 ();
 sg13g2_fill_8 FILLER_32_240 ();
 sg13g2_fill_8 FILLER_32_248 ();
 sg13g2_fill_8 FILLER_32_256 ();
 sg13g2_fill_8 FILLER_32_264 ();
 sg13g2_fill_8 FILLER_32_272 ();
 sg13g2_fill_8 FILLER_32_280 ();
 sg13g2_fill_8 FILLER_32_288 ();
 sg13g2_fill_8 FILLER_32_296 ();
 sg13g2_fill_8 FILLER_32_304 ();
 sg13g2_fill_8 FILLER_32_312 ();
 sg13g2_fill_8 FILLER_32_320 ();
 sg13g2_fill_8 FILLER_32_328 ();
 sg13g2_fill_8 FILLER_32_336 ();
 sg13g2_fill_8 FILLER_32_344 ();
 sg13g2_fill_8 FILLER_32_352 ();
 sg13g2_fill_8 FILLER_32_360 ();
 sg13g2_fill_8 FILLER_32_368 ();
 sg13g2_fill_8 FILLER_32_376 ();
 sg13g2_fill_8 FILLER_32_384 ();
 sg13g2_fill_8 FILLER_32_392 ();
 sg13g2_fill_8 FILLER_32_400 ();
 sg13g2_fill_8 FILLER_32_408 ();
 sg13g2_fill_8 FILLER_32_416 ();
 sg13g2_fill_8 FILLER_32_424 ();
 sg13g2_fill_8 FILLER_32_432 ();
 sg13g2_fill_8 FILLER_32_440 ();
 sg13g2_fill_8 FILLER_32_448 ();
 sg13g2_fill_8 FILLER_32_456 ();
 sg13g2_fill_8 FILLER_32_464 ();
 sg13g2_fill_8 FILLER_32_472 ();
 sg13g2_fill_8 FILLER_32_480 ();
 sg13g2_fill_8 FILLER_32_488 ();
 sg13g2_fill_8 FILLER_32_496 ();
 sg13g2_fill_8 FILLER_32_504 ();
 sg13g2_fill_8 FILLER_32_512 ();
 sg13g2_fill_8 FILLER_32_520 ();
 sg13g2_fill_8 FILLER_32_528 ();
 sg13g2_fill_8 FILLER_32_536 ();
 sg13g2_fill_8 FILLER_32_544 ();
 sg13g2_fill_8 FILLER_32_552 ();
 sg13g2_fill_8 FILLER_32_560 ();
 sg13g2_fill_8 FILLER_32_568 ();
 sg13g2_fill_8 FILLER_32_576 ();
 sg13g2_fill_8 FILLER_32_584 ();
 sg13g2_fill_8 FILLER_32_592 ();
 sg13g2_fill_8 FILLER_32_600 ();
 sg13g2_fill_8 FILLER_32_608 ();
 sg13g2_fill_8 FILLER_32_616 ();
 sg13g2_fill_8 FILLER_32_624 ();
 sg13g2_fill_8 FILLER_32_632 ();
 sg13g2_fill_8 FILLER_32_640 ();
 sg13g2_fill_8 FILLER_32_648 ();
 sg13g2_fill_8 FILLER_32_656 ();
 sg13g2_fill_8 FILLER_32_664 ();
 sg13g2_fill_8 FILLER_32_672 ();
 sg13g2_fill_8 FILLER_32_680 ();
 sg13g2_fill_8 FILLER_32_688 ();
 sg13g2_fill_8 FILLER_32_696 ();
 sg13g2_fill_8 FILLER_32_704 ();
 sg13g2_fill_8 FILLER_32_712 ();
 sg13g2_fill_8 FILLER_32_720 ();
 sg13g2_fill_8 FILLER_32_728 ();
 sg13g2_fill_8 FILLER_32_736 ();
 sg13g2_fill_8 FILLER_32_744 ();
 sg13g2_fill_8 FILLER_32_752 ();
 sg13g2_fill_8 FILLER_32_760 ();
 sg13g2_fill_8 FILLER_32_768 ();
 sg13g2_fill_8 FILLER_32_776 ();
 sg13g2_fill_8 FILLER_32_784 ();
 sg13g2_fill_8 FILLER_32_792 ();
 sg13g2_fill_8 FILLER_32_800 ();
 sg13g2_fill_8 FILLER_32_808 ();
 sg13g2_fill_8 FILLER_32_816 ();
 sg13g2_fill_8 FILLER_32_824 ();
 sg13g2_fill_8 FILLER_32_832 ();
 sg13g2_fill_8 FILLER_32_840 ();
 sg13g2_fill_8 FILLER_32_848 ();
 sg13g2_fill_8 FILLER_32_856 ();
 sg13g2_fill_8 FILLER_32_864 ();
 sg13g2_fill_8 FILLER_32_872 ();
 sg13g2_fill_8 FILLER_32_880 ();
 sg13g2_fill_8 FILLER_32_888 ();
 sg13g2_fill_8 FILLER_32_896 ();
 sg13g2_fill_8 FILLER_32_904 ();
 sg13g2_fill_8 FILLER_32_912 ();
 sg13g2_fill_8 FILLER_32_920 ();
 sg13g2_fill_8 FILLER_32_928 ();
 sg13g2_fill_8 FILLER_32_936 ();
 sg13g2_fill_8 FILLER_32_944 ();
 sg13g2_fill_8 FILLER_32_952 ();
 sg13g2_fill_8 FILLER_32_960 ();
 sg13g2_fill_8 FILLER_32_968 ();
 sg13g2_fill_8 FILLER_32_976 ();
 sg13g2_fill_8 FILLER_32_984 ();
 sg13g2_fill_8 FILLER_32_992 ();
 sg13g2_fill_8 FILLER_32_1000 ();
 sg13g2_fill_8 FILLER_32_1008 ();
 sg13g2_fill_8 FILLER_32_1016 ();
 sg13g2_fill_8 FILLER_32_1024 ();
 sg13g2_fill_8 FILLER_32_1032 ();
 sg13g2_fill_8 FILLER_32_1040 ();
 sg13g2_fill_8 FILLER_32_1048 ();
 sg13g2_fill_8 FILLER_32_1056 ();
 sg13g2_fill_8 FILLER_32_1064 ();
 sg13g2_fill_8 FILLER_32_1072 ();
 sg13g2_fill_8 FILLER_32_1080 ();
 sg13g2_fill_8 FILLER_32_1088 ();
 sg13g2_fill_8 FILLER_32_1096 ();
 sg13g2_fill_8 FILLER_32_1104 ();
 sg13g2_fill_8 FILLER_32_1112 ();
 sg13g2_fill_8 FILLER_32_1120 ();
 sg13g2_fill_8 FILLER_32_1128 ();
 sg13g2_fill_8 FILLER_32_1136 ();
 sg13g2_fill_8 FILLER_33_0 ();
 sg13g2_fill_8 FILLER_33_8 ();
 sg13g2_fill_8 FILLER_33_16 ();
 sg13g2_fill_8 FILLER_33_24 ();
 sg13g2_fill_8 FILLER_33_32 ();
 sg13g2_fill_8 FILLER_33_40 ();
 sg13g2_fill_8 FILLER_33_48 ();
 sg13g2_fill_8 FILLER_33_56 ();
 sg13g2_fill_8 FILLER_33_64 ();
 sg13g2_fill_8 FILLER_33_72 ();
 sg13g2_fill_8 FILLER_33_80 ();
 sg13g2_fill_8 FILLER_33_88 ();
 sg13g2_fill_8 FILLER_33_96 ();
 sg13g2_fill_8 FILLER_33_104 ();
 sg13g2_fill_8 FILLER_33_112 ();
 sg13g2_fill_8 FILLER_33_120 ();
 sg13g2_fill_8 FILLER_33_128 ();
 sg13g2_fill_8 FILLER_33_136 ();
 sg13g2_fill_8 FILLER_33_144 ();
 sg13g2_fill_8 FILLER_33_152 ();
 sg13g2_fill_8 FILLER_33_160 ();
 sg13g2_fill_8 FILLER_33_168 ();
 sg13g2_fill_8 FILLER_33_176 ();
 sg13g2_fill_8 FILLER_33_184 ();
 sg13g2_fill_8 FILLER_33_192 ();
 sg13g2_fill_8 FILLER_33_200 ();
 sg13g2_fill_8 FILLER_33_208 ();
 sg13g2_fill_8 FILLER_33_216 ();
 sg13g2_fill_8 FILLER_33_224 ();
 sg13g2_fill_8 FILLER_33_232 ();
 sg13g2_fill_8 FILLER_33_240 ();
 sg13g2_fill_8 FILLER_33_248 ();
 sg13g2_fill_8 FILLER_33_256 ();
 sg13g2_fill_8 FILLER_33_264 ();
 sg13g2_fill_8 FILLER_33_272 ();
 sg13g2_fill_8 FILLER_33_280 ();
 sg13g2_fill_8 FILLER_33_288 ();
 sg13g2_fill_8 FILLER_33_296 ();
 sg13g2_fill_8 FILLER_33_304 ();
 sg13g2_fill_8 FILLER_33_312 ();
 sg13g2_fill_8 FILLER_33_320 ();
 sg13g2_fill_8 FILLER_33_328 ();
 sg13g2_fill_8 FILLER_33_336 ();
 sg13g2_fill_8 FILLER_33_344 ();
 sg13g2_fill_8 FILLER_33_352 ();
 sg13g2_fill_8 FILLER_33_360 ();
 sg13g2_fill_8 FILLER_33_368 ();
 sg13g2_fill_8 FILLER_33_376 ();
 sg13g2_fill_8 FILLER_33_384 ();
 sg13g2_fill_8 FILLER_33_392 ();
 sg13g2_fill_8 FILLER_33_400 ();
 sg13g2_fill_8 FILLER_33_408 ();
 sg13g2_fill_8 FILLER_33_416 ();
 sg13g2_fill_8 FILLER_33_424 ();
 sg13g2_fill_8 FILLER_33_432 ();
 sg13g2_fill_8 FILLER_33_440 ();
 sg13g2_fill_8 FILLER_33_448 ();
 sg13g2_fill_8 FILLER_33_456 ();
 sg13g2_fill_8 FILLER_33_464 ();
 sg13g2_fill_8 FILLER_33_472 ();
 sg13g2_fill_8 FILLER_33_480 ();
 sg13g2_fill_8 FILLER_33_488 ();
 sg13g2_fill_8 FILLER_33_496 ();
 sg13g2_fill_8 FILLER_33_504 ();
 sg13g2_fill_8 FILLER_33_512 ();
 sg13g2_fill_8 FILLER_33_520 ();
 sg13g2_fill_8 FILLER_33_528 ();
 sg13g2_fill_8 FILLER_33_536 ();
 sg13g2_fill_8 FILLER_33_544 ();
 sg13g2_fill_8 FILLER_33_552 ();
 sg13g2_fill_8 FILLER_33_560 ();
 sg13g2_fill_8 FILLER_33_568 ();
 sg13g2_fill_8 FILLER_33_576 ();
 sg13g2_fill_8 FILLER_33_584 ();
 sg13g2_fill_8 FILLER_33_592 ();
 sg13g2_fill_8 FILLER_33_600 ();
 sg13g2_fill_8 FILLER_33_608 ();
 sg13g2_fill_8 FILLER_33_616 ();
 sg13g2_fill_8 FILLER_33_624 ();
 sg13g2_fill_8 FILLER_33_632 ();
 sg13g2_fill_8 FILLER_33_640 ();
 sg13g2_fill_8 FILLER_33_648 ();
 sg13g2_fill_8 FILLER_33_656 ();
 sg13g2_fill_8 FILLER_33_664 ();
 sg13g2_fill_8 FILLER_33_672 ();
 sg13g2_fill_8 FILLER_33_680 ();
 sg13g2_fill_8 FILLER_33_688 ();
 sg13g2_fill_8 FILLER_33_696 ();
 sg13g2_fill_8 FILLER_33_704 ();
 sg13g2_fill_8 FILLER_33_712 ();
 sg13g2_fill_8 FILLER_33_720 ();
 sg13g2_fill_8 FILLER_33_728 ();
 sg13g2_fill_8 FILLER_33_736 ();
 sg13g2_fill_8 FILLER_33_744 ();
 sg13g2_fill_8 FILLER_33_752 ();
 sg13g2_fill_8 FILLER_33_760 ();
 sg13g2_fill_8 FILLER_33_768 ();
 sg13g2_fill_8 FILLER_33_776 ();
 sg13g2_fill_8 FILLER_33_784 ();
 sg13g2_fill_8 FILLER_33_792 ();
 sg13g2_fill_8 FILLER_33_800 ();
 sg13g2_fill_8 FILLER_33_808 ();
 sg13g2_fill_8 FILLER_33_816 ();
 sg13g2_fill_8 FILLER_33_824 ();
 sg13g2_fill_8 FILLER_33_832 ();
 sg13g2_fill_8 FILLER_33_840 ();
 sg13g2_fill_8 FILLER_33_848 ();
 sg13g2_fill_8 FILLER_33_856 ();
 sg13g2_fill_8 FILLER_33_864 ();
 sg13g2_fill_8 FILLER_33_872 ();
 sg13g2_fill_8 FILLER_33_880 ();
 sg13g2_fill_8 FILLER_33_888 ();
 sg13g2_fill_8 FILLER_33_896 ();
 sg13g2_fill_8 FILLER_33_904 ();
 sg13g2_fill_8 FILLER_33_912 ();
 sg13g2_fill_8 FILLER_33_920 ();
 sg13g2_fill_8 FILLER_33_928 ();
 sg13g2_fill_8 FILLER_33_936 ();
 sg13g2_fill_8 FILLER_33_944 ();
 sg13g2_fill_8 FILLER_33_952 ();
 sg13g2_fill_8 FILLER_33_960 ();
 sg13g2_fill_8 FILLER_33_968 ();
 sg13g2_fill_8 FILLER_33_976 ();
 sg13g2_fill_8 FILLER_33_984 ();
 sg13g2_fill_8 FILLER_33_992 ();
 sg13g2_fill_8 FILLER_33_1000 ();
 sg13g2_fill_8 FILLER_33_1008 ();
 sg13g2_fill_8 FILLER_33_1016 ();
 sg13g2_fill_8 FILLER_33_1024 ();
 sg13g2_fill_8 FILLER_33_1032 ();
 sg13g2_fill_8 FILLER_33_1040 ();
 sg13g2_fill_8 FILLER_33_1048 ();
 sg13g2_fill_8 FILLER_33_1056 ();
 sg13g2_fill_8 FILLER_33_1064 ();
 sg13g2_fill_8 FILLER_33_1072 ();
 sg13g2_fill_8 FILLER_33_1080 ();
 sg13g2_fill_8 FILLER_33_1088 ();
 sg13g2_fill_8 FILLER_33_1096 ();
 sg13g2_fill_8 FILLER_33_1104 ();
 sg13g2_fill_8 FILLER_33_1112 ();
 sg13g2_fill_8 FILLER_33_1120 ();
 sg13g2_fill_8 FILLER_33_1128 ();
 sg13g2_fill_8 FILLER_33_1136 ();
 sg13g2_fill_8 FILLER_34_0 ();
 sg13g2_fill_8 FILLER_34_8 ();
 sg13g2_fill_8 FILLER_34_16 ();
 sg13g2_fill_8 FILLER_34_24 ();
 sg13g2_fill_8 FILLER_34_32 ();
 sg13g2_fill_8 FILLER_34_40 ();
 sg13g2_fill_8 FILLER_34_48 ();
 sg13g2_fill_8 FILLER_34_56 ();
 sg13g2_fill_8 FILLER_34_64 ();
 sg13g2_fill_8 FILLER_34_72 ();
 sg13g2_fill_8 FILLER_34_80 ();
 sg13g2_fill_8 FILLER_34_88 ();
 sg13g2_fill_8 FILLER_34_96 ();
 sg13g2_fill_8 FILLER_34_104 ();
 sg13g2_fill_8 FILLER_34_112 ();
 sg13g2_fill_8 FILLER_34_120 ();
 sg13g2_fill_8 FILLER_34_128 ();
 sg13g2_fill_8 FILLER_34_136 ();
 sg13g2_fill_8 FILLER_34_144 ();
 sg13g2_fill_8 FILLER_34_152 ();
 sg13g2_fill_8 FILLER_34_160 ();
 sg13g2_fill_8 FILLER_34_168 ();
 sg13g2_fill_8 FILLER_34_176 ();
 sg13g2_fill_8 FILLER_34_184 ();
 sg13g2_fill_8 FILLER_34_192 ();
 sg13g2_fill_8 FILLER_34_200 ();
 sg13g2_fill_8 FILLER_34_208 ();
 sg13g2_fill_8 FILLER_34_216 ();
 sg13g2_fill_8 FILLER_34_224 ();
 sg13g2_fill_8 FILLER_34_232 ();
 sg13g2_fill_8 FILLER_34_240 ();
 sg13g2_fill_8 FILLER_34_248 ();
 sg13g2_fill_8 FILLER_34_256 ();
 sg13g2_fill_8 FILLER_34_264 ();
 sg13g2_fill_8 FILLER_34_272 ();
 sg13g2_fill_8 FILLER_34_280 ();
 sg13g2_fill_8 FILLER_34_288 ();
 sg13g2_fill_8 FILLER_34_296 ();
 sg13g2_fill_8 FILLER_34_304 ();
 sg13g2_fill_8 FILLER_34_312 ();
 sg13g2_fill_8 FILLER_34_320 ();
 sg13g2_fill_8 FILLER_34_328 ();
 sg13g2_fill_8 FILLER_34_336 ();
 sg13g2_fill_8 FILLER_34_344 ();
 sg13g2_fill_8 FILLER_34_352 ();
 sg13g2_fill_8 FILLER_34_360 ();
 sg13g2_fill_8 FILLER_34_368 ();
 sg13g2_fill_8 FILLER_34_376 ();
 sg13g2_fill_8 FILLER_34_384 ();
 sg13g2_fill_8 FILLER_34_392 ();
 sg13g2_fill_8 FILLER_34_400 ();
 sg13g2_fill_8 FILLER_34_408 ();
 sg13g2_fill_8 FILLER_34_416 ();
 sg13g2_fill_8 FILLER_34_424 ();
 sg13g2_fill_8 FILLER_34_432 ();
 sg13g2_fill_8 FILLER_34_440 ();
 sg13g2_fill_8 FILLER_34_448 ();
 sg13g2_fill_8 FILLER_34_456 ();
 sg13g2_fill_8 FILLER_34_464 ();
 sg13g2_fill_8 FILLER_34_472 ();
 sg13g2_fill_8 FILLER_34_480 ();
 sg13g2_fill_8 FILLER_34_488 ();
 sg13g2_fill_8 FILLER_34_496 ();
 sg13g2_fill_8 FILLER_34_504 ();
 sg13g2_fill_8 FILLER_34_512 ();
 sg13g2_fill_8 FILLER_34_520 ();
 sg13g2_fill_8 FILLER_34_528 ();
 sg13g2_fill_8 FILLER_34_536 ();
 sg13g2_fill_8 FILLER_34_544 ();
 sg13g2_fill_8 FILLER_34_552 ();
 sg13g2_fill_8 FILLER_34_560 ();
 sg13g2_fill_8 FILLER_34_568 ();
 sg13g2_fill_8 FILLER_34_576 ();
 sg13g2_fill_8 FILLER_34_584 ();
 sg13g2_fill_8 FILLER_34_592 ();
 sg13g2_fill_8 FILLER_34_600 ();
 sg13g2_fill_8 FILLER_34_608 ();
 sg13g2_fill_8 FILLER_34_616 ();
 sg13g2_fill_8 FILLER_34_624 ();
 sg13g2_fill_8 FILLER_34_632 ();
 sg13g2_fill_8 FILLER_34_640 ();
 sg13g2_fill_8 FILLER_34_648 ();
 sg13g2_fill_8 FILLER_34_656 ();
 sg13g2_fill_8 FILLER_34_664 ();
 sg13g2_fill_8 FILLER_34_672 ();
 sg13g2_fill_8 FILLER_34_680 ();
 sg13g2_fill_8 FILLER_34_688 ();
 sg13g2_fill_8 FILLER_34_696 ();
 sg13g2_fill_8 FILLER_34_704 ();
 sg13g2_fill_8 FILLER_34_712 ();
 sg13g2_fill_8 FILLER_34_720 ();
 sg13g2_fill_8 FILLER_34_728 ();
 sg13g2_fill_8 FILLER_34_736 ();
 sg13g2_fill_8 FILLER_34_744 ();
 sg13g2_fill_8 FILLER_34_752 ();
 sg13g2_fill_8 FILLER_34_760 ();
 sg13g2_fill_8 FILLER_34_768 ();
 sg13g2_fill_8 FILLER_34_776 ();
 sg13g2_fill_8 FILLER_34_784 ();
 sg13g2_fill_8 FILLER_34_792 ();
 sg13g2_fill_8 FILLER_34_800 ();
 sg13g2_fill_8 FILLER_34_808 ();
 sg13g2_fill_8 FILLER_34_816 ();
 sg13g2_fill_8 FILLER_34_824 ();
 sg13g2_fill_8 FILLER_34_832 ();
 sg13g2_fill_8 FILLER_34_840 ();
 sg13g2_fill_8 FILLER_34_848 ();
 sg13g2_fill_8 FILLER_34_856 ();
 sg13g2_fill_8 FILLER_34_864 ();
 sg13g2_fill_8 FILLER_34_872 ();
 sg13g2_fill_8 FILLER_34_880 ();
 sg13g2_fill_8 FILLER_34_888 ();
 sg13g2_fill_8 FILLER_34_896 ();
 sg13g2_fill_8 FILLER_34_904 ();
 sg13g2_fill_8 FILLER_34_912 ();
 sg13g2_fill_8 FILLER_34_920 ();
 sg13g2_fill_8 FILLER_34_928 ();
 sg13g2_fill_8 FILLER_34_936 ();
 sg13g2_fill_8 FILLER_34_944 ();
 sg13g2_fill_8 FILLER_34_952 ();
 sg13g2_fill_8 FILLER_34_960 ();
 sg13g2_fill_8 FILLER_34_968 ();
 sg13g2_fill_8 FILLER_34_976 ();
 sg13g2_fill_8 FILLER_34_984 ();
 sg13g2_fill_8 FILLER_34_992 ();
 sg13g2_fill_8 FILLER_34_1000 ();
 sg13g2_fill_8 FILLER_34_1008 ();
 sg13g2_fill_8 FILLER_34_1016 ();
 sg13g2_fill_8 FILLER_34_1024 ();
 sg13g2_fill_8 FILLER_34_1032 ();
 sg13g2_fill_8 FILLER_34_1040 ();
 sg13g2_fill_8 FILLER_34_1048 ();
 sg13g2_fill_8 FILLER_34_1056 ();
 sg13g2_fill_8 FILLER_34_1064 ();
 sg13g2_fill_8 FILLER_34_1072 ();
 sg13g2_fill_8 FILLER_34_1080 ();
 sg13g2_fill_8 FILLER_34_1088 ();
 sg13g2_fill_8 FILLER_34_1096 ();
 sg13g2_fill_8 FILLER_34_1104 ();
 sg13g2_fill_8 FILLER_34_1112 ();
 sg13g2_fill_8 FILLER_34_1120 ();
 sg13g2_fill_8 FILLER_34_1128 ();
 sg13g2_fill_8 FILLER_34_1136 ();
 sg13g2_fill_8 FILLER_35_0 ();
 sg13g2_fill_8 FILLER_35_8 ();
 sg13g2_fill_8 FILLER_35_16 ();
 sg13g2_fill_8 FILLER_35_24 ();
 sg13g2_fill_8 FILLER_35_32 ();
 sg13g2_fill_8 FILLER_35_40 ();
 sg13g2_fill_8 FILLER_35_48 ();
 sg13g2_fill_8 FILLER_35_56 ();
 sg13g2_fill_8 FILLER_35_64 ();
 sg13g2_fill_8 FILLER_35_72 ();
 sg13g2_fill_8 FILLER_35_80 ();
 sg13g2_fill_8 FILLER_35_88 ();
 sg13g2_fill_8 FILLER_35_96 ();
 sg13g2_fill_8 FILLER_35_104 ();
 sg13g2_fill_8 FILLER_35_112 ();
 sg13g2_fill_8 FILLER_35_120 ();
 sg13g2_fill_8 FILLER_35_128 ();
 sg13g2_fill_8 FILLER_35_136 ();
 sg13g2_fill_8 FILLER_35_144 ();
 sg13g2_fill_8 FILLER_35_152 ();
 sg13g2_fill_8 FILLER_35_160 ();
 sg13g2_fill_8 FILLER_35_168 ();
 sg13g2_fill_8 FILLER_35_176 ();
 sg13g2_fill_8 FILLER_35_184 ();
 sg13g2_fill_8 FILLER_35_192 ();
 sg13g2_fill_8 FILLER_35_200 ();
 sg13g2_fill_8 FILLER_35_208 ();
 sg13g2_fill_8 FILLER_35_216 ();
 sg13g2_fill_8 FILLER_35_224 ();
 sg13g2_fill_8 FILLER_35_232 ();
 sg13g2_fill_8 FILLER_35_240 ();
 sg13g2_fill_8 FILLER_35_248 ();
 sg13g2_fill_8 FILLER_35_256 ();
 sg13g2_fill_8 FILLER_35_264 ();
 sg13g2_fill_8 FILLER_35_272 ();
 sg13g2_fill_8 FILLER_35_280 ();
 sg13g2_fill_8 FILLER_35_288 ();
 sg13g2_fill_8 FILLER_35_296 ();
 sg13g2_fill_8 FILLER_35_304 ();
 sg13g2_fill_8 FILLER_35_312 ();
 sg13g2_fill_8 FILLER_35_320 ();
 sg13g2_fill_8 FILLER_35_328 ();
 sg13g2_fill_8 FILLER_35_336 ();
 sg13g2_fill_8 FILLER_35_344 ();
 sg13g2_fill_8 FILLER_35_352 ();
 sg13g2_fill_8 FILLER_35_360 ();
 sg13g2_fill_8 FILLER_35_368 ();
 sg13g2_fill_8 FILLER_35_376 ();
 sg13g2_fill_8 FILLER_35_384 ();
 sg13g2_fill_8 FILLER_35_392 ();
 sg13g2_fill_8 FILLER_35_400 ();
 sg13g2_fill_8 FILLER_35_408 ();
 sg13g2_fill_8 FILLER_35_416 ();
 sg13g2_fill_8 FILLER_35_424 ();
 sg13g2_fill_8 FILLER_35_432 ();
 sg13g2_fill_8 FILLER_35_440 ();
 sg13g2_fill_8 FILLER_35_448 ();
 sg13g2_fill_8 FILLER_35_456 ();
 sg13g2_fill_8 FILLER_35_464 ();
 sg13g2_fill_8 FILLER_35_472 ();
 sg13g2_fill_8 FILLER_35_480 ();
 sg13g2_fill_8 FILLER_35_488 ();
 sg13g2_fill_8 FILLER_35_496 ();
 sg13g2_fill_8 FILLER_35_504 ();
 sg13g2_fill_8 FILLER_35_512 ();
 sg13g2_fill_8 FILLER_35_520 ();
 sg13g2_fill_8 FILLER_35_528 ();
 sg13g2_fill_8 FILLER_35_536 ();
 sg13g2_fill_8 FILLER_35_544 ();
 sg13g2_fill_8 FILLER_35_552 ();
 sg13g2_fill_8 FILLER_35_560 ();
 sg13g2_fill_8 FILLER_35_568 ();
 sg13g2_fill_8 FILLER_35_576 ();
 sg13g2_fill_8 FILLER_35_584 ();
 sg13g2_fill_8 FILLER_35_592 ();
 sg13g2_fill_8 FILLER_35_600 ();
 sg13g2_fill_8 FILLER_35_608 ();
 sg13g2_fill_8 FILLER_35_616 ();
 sg13g2_fill_8 FILLER_35_624 ();
 sg13g2_fill_8 FILLER_35_632 ();
 sg13g2_fill_8 FILLER_35_640 ();
 sg13g2_fill_8 FILLER_35_648 ();
 sg13g2_fill_8 FILLER_35_656 ();
 sg13g2_fill_8 FILLER_35_664 ();
 sg13g2_fill_8 FILLER_35_672 ();
 sg13g2_fill_8 FILLER_35_680 ();
 sg13g2_fill_8 FILLER_35_688 ();
 sg13g2_fill_8 FILLER_35_696 ();
 sg13g2_fill_8 FILLER_35_704 ();
 sg13g2_fill_8 FILLER_35_712 ();
 sg13g2_fill_8 FILLER_35_720 ();
 sg13g2_fill_8 FILLER_35_728 ();
 sg13g2_fill_8 FILLER_35_736 ();
 sg13g2_fill_8 FILLER_35_744 ();
 sg13g2_fill_8 FILLER_35_752 ();
 sg13g2_fill_8 FILLER_35_760 ();
 sg13g2_fill_8 FILLER_35_768 ();
 sg13g2_fill_8 FILLER_35_776 ();
 sg13g2_fill_8 FILLER_35_784 ();
 sg13g2_fill_8 FILLER_35_792 ();
 sg13g2_fill_8 FILLER_35_800 ();
 sg13g2_fill_8 FILLER_35_808 ();
 sg13g2_fill_8 FILLER_35_816 ();
 sg13g2_fill_8 FILLER_35_824 ();
 sg13g2_fill_8 FILLER_35_832 ();
 sg13g2_fill_8 FILLER_35_840 ();
 sg13g2_fill_8 FILLER_35_848 ();
 sg13g2_fill_8 FILLER_35_856 ();
 sg13g2_fill_8 FILLER_35_864 ();
 sg13g2_fill_8 FILLER_35_872 ();
 sg13g2_fill_8 FILLER_35_880 ();
 sg13g2_fill_8 FILLER_35_888 ();
 sg13g2_fill_8 FILLER_35_896 ();
 sg13g2_fill_8 FILLER_35_904 ();
 sg13g2_fill_8 FILLER_35_912 ();
 sg13g2_fill_8 FILLER_35_920 ();
 sg13g2_fill_8 FILLER_35_928 ();
 sg13g2_fill_8 FILLER_35_936 ();
 sg13g2_fill_8 FILLER_35_944 ();
 sg13g2_fill_8 FILLER_35_952 ();
 sg13g2_fill_8 FILLER_35_960 ();
 sg13g2_fill_8 FILLER_35_968 ();
 sg13g2_fill_8 FILLER_35_976 ();
 sg13g2_fill_8 FILLER_35_984 ();
 sg13g2_fill_8 FILLER_35_992 ();
 sg13g2_fill_8 FILLER_35_1000 ();
 sg13g2_fill_8 FILLER_35_1008 ();
 sg13g2_fill_8 FILLER_35_1016 ();
 sg13g2_fill_8 FILLER_35_1024 ();
 sg13g2_fill_8 FILLER_35_1032 ();
 sg13g2_fill_8 FILLER_35_1040 ();
 sg13g2_fill_8 FILLER_35_1048 ();
 sg13g2_fill_8 FILLER_35_1056 ();
 sg13g2_fill_8 FILLER_35_1064 ();
 sg13g2_fill_8 FILLER_35_1072 ();
 sg13g2_fill_8 FILLER_35_1080 ();
 sg13g2_fill_8 FILLER_35_1088 ();
 sg13g2_fill_8 FILLER_35_1096 ();
 sg13g2_fill_8 FILLER_35_1104 ();
 sg13g2_fill_8 FILLER_35_1112 ();
 sg13g2_fill_8 FILLER_35_1120 ();
 sg13g2_fill_8 FILLER_35_1128 ();
 sg13g2_fill_8 FILLER_35_1136 ();
 sg13g2_fill_8 FILLER_36_0 ();
 sg13g2_fill_8 FILLER_36_8 ();
 sg13g2_fill_8 FILLER_36_16 ();
 sg13g2_fill_8 FILLER_36_24 ();
 sg13g2_fill_8 FILLER_36_32 ();
 sg13g2_fill_8 FILLER_36_40 ();
 sg13g2_fill_8 FILLER_36_48 ();
 sg13g2_fill_8 FILLER_36_56 ();
 sg13g2_fill_8 FILLER_36_64 ();
 sg13g2_fill_8 FILLER_36_72 ();
 sg13g2_fill_8 FILLER_36_80 ();
 sg13g2_fill_8 FILLER_36_88 ();
 sg13g2_fill_8 FILLER_36_96 ();
 sg13g2_fill_8 FILLER_36_104 ();
 sg13g2_fill_8 FILLER_36_112 ();
 sg13g2_fill_8 FILLER_36_120 ();
 sg13g2_fill_8 FILLER_36_128 ();
 sg13g2_fill_8 FILLER_36_136 ();
 sg13g2_fill_8 FILLER_36_144 ();
 sg13g2_fill_8 FILLER_36_152 ();
 sg13g2_fill_8 FILLER_36_160 ();
 sg13g2_fill_8 FILLER_36_168 ();
 sg13g2_fill_8 FILLER_36_176 ();
 sg13g2_fill_8 FILLER_36_184 ();
 sg13g2_fill_8 FILLER_36_192 ();
 sg13g2_fill_8 FILLER_36_200 ();
 sg13g2_fill_8 FILLER_36_208 ();
 sg13g2_fill_8 FILLER_36_216 ();
 sg13g2_fill_8 FILLER_36_224 ();
 sg13g2_fill_8 FILLER_36_232 ();
 sg13g2_fill_8 FILLER_36_240 ();
 sg13g2_fill_8 FILLER_36_248 ();
 sg13g2_fill_8 FILLER_36_256 ();
 sg13g2_fill_8 FILLER_36_264 ();
 sg13g2_fill_8 FILLER_36_272 ();
 sg13g2_fill_8 FILLER_36_280 ();
 sg13g2_fill_8 FILLER_36_288 ();
 sg13g2_fill_8 FILLER_36_296 ();
 sg13g2_fill_8 FILLER_36_304 ();
 sg13g2_fill_8 FILLER_36_312 ();
 sg13g2_fill_8 FILLER_36_320 ();
 sg13g2_fill_8 FILLER_36_328 ();
 sg13g2_fill_8 FILLER_36_336 ();
 sg13g2_fill_8 FILLER_36_344 ();
 sg13g2_fill_8 FILLER_36_352 ();
 sg13g2_fill_8 FILLER_36_360 ();
 sg13g2_fill_8 FILLER_36_368 ();
 sg13g2_fill_8 FILLER_36_376 ();
 sg13g2_fill_8 FILLER_36_384 ();
 sg13g2_fill_8 FILLER_36_392 ();
 sg13g2_fill_8 FILLER_36_400 ();
 sg13g2_fill_8 FILLER_36_408 ();
 sg13g2_fill_8 FILLER_36_416 ();
 sg13g2_fill_8 FILLER_36_424 ();
 sg13g2_fill_8 FILLER_36_432 ();
 sg13g2_fill_8 FILLER_36_440 ();
 sg13g2_fill_8 FILLER_36_448 ();
 sg13g2_fill_8 FILLER_36_456 ();
 sg13g2_fill_8 FILLER_36_464 ();
 sg13g2_fill_8 FILLER_36_472 ();
 sg13g2_fill_8 FILLER_36_480 ();
 sg13g2_fill_8 FILLER_36_488 ();
 sg13g2_fill_8 FILLER_36_496 ();
 sg13g2_fill_8 FILLER_36_504 ();
 sg13g2_fill_8 FILLER_36_512 ();
 sg13g2_fill_8 FILLER_36_520 ();
 sg13g2_fill_8 FILLER_36_528 ();
 sg13g2_fill_8 FILLER_36_536 ();
 sg13g2_fill_8 FILLER_36_544 ();
 sg13g2_fill_8 FILLER_36_552 ();
 sg13g2_fill_8 FILLER_36_560 ();
 sg13g2_fill_8 FILLER_36_568 ();
 sg13g2_fill_8 FILLER_36_576 ();
 sg13g2_fill_8 FILLER_36_584 ();
 sg13g2_fill_8 FILLER_36_592 ();
 sg13g2_fill_8 FILLER_36_600 ();
 sg13g2_fill_8 FILLER_36_608 ();
 sg13g2_fill_8 FILLER_36_616 ();
 sg13g2_fill_8 FILLER_36_624 ();
 sg13g2_fill_8 FILLER_36_632 ();
 sg13g2_fill_8 FILLER_36_640 ();
 sg13g2_fill_8 FILLER_36_648 ();
 sg13g2_fill_8 FILLER_36_656 ();
 sg13g2_fill_8 FILLER_36_664 ();
 sg13g2_fill_8 FILLER_36_672 ();
 sg13g2_fill_8 FILLER_36_680 ();
 sg13g2_fill_8 FILLER_36_688 ();
 sg13g2_fill_8 FILLER_36_696 ();
 sg13g2_fill_8 FILLER_36_704 ();
 sg13g2_fill_8 FILLER_36_712 ();
 sg13g2_fill_8 FILLER_36_720 ();
 sg13g2_fill_8 FILLER_36_728 ();
 sg13g2_fill_8 FILLER_36_736 ();
 sg13g2_fill_8 FILLER_36_744 ();
 sg13g2_fill_8 FILLER_36_752 ();
 sg13g2_fill_8 FILLER_36_760 ();
 sg13g2_fill_8 FILLER_36_768 ();
 sg13g2_fill_8 FILLER_36_776 ();
 sg13g2_fill_8 FILLER_36_784 ();
 sg13g2_fill_8 FILLER_36_792 ();
 sg13g2_fill_8 FILLER_36_800 ();
 sg13g2_fill_8 FILLER_36_808 ();
 sg13g2_fill_8 FILLER_36_816 ();
 sg13g2_fill_8 FILLER_36_824 ();
 sg13g2_fill_8 FILLER_36_832 ();
 sg13g2_fill_8 FILLER_36_840 ();
 sg13g2_fill_8 FILLER_36_848 ();
 sg13g2_fill_8 FILLER_36_856 ();
 sg13g2_fill_8 FILLER_36_864 ();
 sg13g2_fill_8 FILLER_36_872 ();
 sg13g2_fill_8 FILLER_36_880 ();
 sg13g2_fill_8 FILLER_36_888 ();
 sg13g2_fill_8 FILLER_36_896 ();
 sg13g2_fill_8 FILLER_36_904 ();
 sg13g2_fill_8 FILLER_36_912 ();
 sg13g2_fill_8 FILLER_36_920 ();
 sg13g2_fill_8 FILLER_36_928 ();
 sg13g2_fill_8 FILLER_36_936 ();
 sg13g2_fill_8 FILLER_36_944 ();
 sg13g2_fill_8 FILLER_36_952 ();
 sg13g2_fill_8 FILLER_36_960 ();
 sg13g2_fill_8 FILLER_36_968 ();
 sg13g2_fill_8 FILLER_36_976 ();
 sg13g2_fill_8 FILLER_36_984 ();
 sg13g2_fill_8 FILLER_36_992 ();
 sg13g2_fill_8 FILLER_36_1000 ();
 sg13g2_fill_8 FILLER_36_1008 ();
 sg13g2_fill_8 FILLER_36_1016 ();
 sg13g2_fill_8 FILLER_36_1024 ();
 sg13g2_fill_8 FILLER_36_1032 ();
 sg13g2_fill_8 FILLER_36_1040 ();
 sg13g2_fill_8 FILLER_36_1048 ();
 sg13g2_fill_8 FILLER_36_1056 ();
 sg13g2_fill_8 FILLER_36_1064 ();
 sg13g2_fill_8 FILLER_36_1072 ();
 sg13g2_fill_8 FILLER_36_1080 ();
 sg13g2_fill_8 FILLER_36_1088 ();
 sg13g2_fill_8 FILLER_36_1096 ();
 sg13g2_fill_8 FILLER_36_1104 ();
 sg13g2_fill_8 FILLER_36_1112 ();
 sg13g2_fill_8 FILLER_36_1120 ();
 sg13g2_fill_8 FILLER_36_1128 ();
 sg13g2_fill_8 FILLER_36_1136 ();
 sg13g2_fill_8 FILLER_37_0 ();
 sg13g2_fill_8 FILLER_37_8 ();
 sg13g2_fill_8 FILLER_37_16 ();
 sg13g2_fill_8 FILLER_37_24 ();
 sg13g2_fill_8 FILLER_37_32 ();
 sg13g2_fill_8 FILLER_37_40 ();
 sg13g2_fill_8 FILLER_37_48 ();
 sg13g2_fill_8 FILLER_37_56 ();
 sg13g2_fill_8 FILLER_37_64 ();
 sg13g2_fill_8 FILLER_37_72 ();
 sg13g2_fill_8 FILLER_37_80 ();
 sg13g2_fill_8 FILLER_37_88 ();
 sg13g2_fill_8 FILLER_37_96 ();
 sg13g2_fill_8 FILLER_37_104 ();
 sg13g2_fill_8 FILLER_37_112 ();
 sg13g2_fill_8 FILLER_37_120 ();
 sg13g2_fill_8 FILLER_37_128 ();
 sg13g2_fill_8 FILLER_37_136 ();
 sg13g2_fill_8 FILLER_37_144 ();
 sg13g2_fill_8 FILLER_37_152 ();
 sg13g2_fill_8 FILLER_37_160 ();
 sg13g2_fill_8 FILLER_37_168 ();
 sg13g2_fill_8 FILLER_37_176 ();
 sg13g2_fill_8 FILLER_37_184 ();
 sg13g2_fill_8 FILLER_37_192 ();
 sg13g2_fill_8 FILLER_37_200 ();
 sg13g2_fill_8 FILLER_37_208 ();
 sg13g2_fill_8 FILLER_37_216 ();
 sg13g2_fill_8 FILLER_37_224 ();
 sg13g2_fill_8 FILLER_37_232 ();
 sg13g2_fill_8 FILLER_37_240 ();
 sg13g2_fill_8 FILLER_37_248 ();
 sg13g2_fill_8 FILLER_37_256 ();
 sg13g2_fill_8 FILLER_37_264 ();
 sg13g2_fill_8 FILLER_37_272 ();
 sg13g2_fill_8 FILLER_37_280 ();
 sg13g2_fill_8 FILLER_37_288 ();
 sg13g2_fill_8 FILLER_37_296 ();
 sg13g2_fill_8 FILLER_37_304 ();
 sg13g2_fill_8 FILLER_37_312 ();
 sg13g2_fill_8 FILLER_37_320 ();
 sg13g2_fill_8 FILLER_37_328 ();
 sg13g2_fill_8 FILLER_37_336 ();
 sg13g2_fill_8 FILLER_37_344 ();
 sg13g2_fill_8 FILLER_37_352 ();
 sg13g2_fill_8 FILLER_37_360 ();
 sg13g2_fill_8 FILLER_37_368 ();
 sg13g2_fill_8 FILLER_37_376 ();
 sg13g2_fill_8 FILLER_37_384 ();
 sg13g2_fill_8 FILLER_37_392 ();
 sg13g2_fill_8 FILLER_37_400 ();
 sg13g2_fill_8 FILLER_37_408 ();
 sg13g2_fill_8 FILLER_37_416 ();
 sg13g2_fill_8 FILLER_37_424 ();
 sg13g2_fill_8 FILLER_37_432 ();
 sg13g2_fill_8 FILLER_37_440 ();
 sg13g2_fill_8 FILLER_37_448 ();
 sg13g2_fill_8 FILLER_37_456 ();
 sg13g2_fill_8 FILLER_37_464 ();
 sg13g2_fill_8 FILLER_37_472 ();
 sg13g2_fill_8 FILLER_37_480 ();
 sg13g2_fill_8 FILLER_37_488 ();
 sg13g2_fill_8 FILLER_37_496 ();
 sg13g2_fill_8 FILLER_37_504 ();
 sg13g2_fill_8 FILLER_37_512 ();
 sg13g2_fill_8 FILLER_37_520 ();
 sg13g2_fill_8 FILLER_37_528 ();
 sg13g2_fill_8 FILLER_37_536 ();
 sg13g2_fill_8 FILLER_37_544 ();
 sg13g2_fill_8 FILLER_37_552 ();
 sg13g2_fill_8 FILLER_37_560 ();
 sg13g2_fill_8 FILLER_37_568 ();
 sg13g2_fill_8 FILLER_37_576 ();
 sg13g2_fill_8 FILLER_37_584 ();
 sg13g2_fill_8 FILLER_37_592 ();
 sg13g2_fill_8 FILLER_37_600 ();
 sg13g2_fill_8 FILLER_37_608 ();
 sg13g2_fill_8 FILLER_37_616 ();
 sg13g2_fill_8 FILLER_37_624 ();
 sg13g2_fill_8 FILLER_37_632 ();
 sg13g2_fill_8 FILLER_37_640 ();
 sg13g2_fill_8 FILLER_37_648 ();
 sg13g2_fill_8 FILLER_37_656 ();
 sg13g2_fill_8 FILLER_37_664 ();
 sg13g2_fill_8 FILLER_37_672 ();
 sg13g2_fill_8 FILLER_37_680 ();
 sg13g2_fill_8 FILLER_37_688 ();
 sg13g2_fill_8 FILLER_37_696 ();
 sg13g2_fill_8 FILLER_37_704 ();
 sg13g2_fill_8 FILLER_37_712 ();
 sg13g2_fill_8 FILLER_37_720 ();
 sg13g2_fill_8 FILLER_37_728 ();
 sg13g2_fill_8 FILLER_37_736 ();
 sg13g2_fill_8 FILLER_37_744 ();
 sg13g2_fill_8 FILLER_37_752 ();
 sg13g2_fill_8 FILLER_37_760 ();
 sg13g2_fill_8 FILLER_37_768 ();
 sg13g2_fill_8 FILLER_37_776 ();
 sg13g2_fill_8 FILLER_37_784 ();
 sg13g2_fill_8 FILLER_37_792 ();
 sg13g2_fill_8 FILLER_37_800 ();
 sg13g2_fill_8 FILLER_37_808 ();
 sg13g2_fill_8 FILLER_37_816 ();
 sg13g2_fill_8 FILLER_37_824 ();
 sg13g2_fill_8 FILLER_37_832 ();
 sg13g2_fill_8 FILLER_37_840 ();
 sg13g2_fill_8 FILLER_37_848 ();
 sg13g2_fill_8 FILLER_37_856 ();
 sg13g2_fill_8 FILLER_37_864 ();
 sg13g2_fill_8 FILLER_37_872 ();
 sg13g2_fill_8 FILLER_37_880 ();
 sg13g2_fill_8 FILLER_37_888 ();
 sg13g2_fill_8 FILLER_37_896 ();
 sg13g2_fill_8 FILLER_37_904 ();
 sg13g2_fill_8 FILLER_37_912 ();
 sg13g2_fill_8 FILLER_37_920 ();
 sg13g2_fill_8 FILLER_37_928 ();
 sg13g2_fill_8 FILLER_37_936 ();
 sg13g2_fill_8 FILLER_37_944 ();
 sg13g2_fill_8 FILLER_37_952 ();
 sg13g2_fill_8 FILLER_37_960 ();
 sg13g2_fill_8 FILLER_37_968 ();
 sg13g2_fill_8 FILLER_37_976 ();
 sg13g2_fill_8 FILLER_37_984 ();
 sg13g2_fill_8 FILLER_37_992 ();
 sg13g2_fill_8 FILLER_37_1000 ();
 sg13g2_fill_8 FILLER_37_1008 ();
 sg13g2_fill_8 FILLER_37_1016 ();
 sg13g2_fill_8 FILLER_37_1024 ();
 sg13g2_fill_8 FILLER_37_1032 ();
 sg13g2_fill_8 FILLER_37_1040 ();
 sg13g2_fill_8 FILLER_37_1048 ();
 sg13g2_fill_8 FILLER_37_1056 ();
 sg13g2_fill_8 FILLER_37_1064 ();
 sg13g2_fill_8 FILLER_37_1072 ();
 sg13g2_fill_8 FILLER_37_1080 ();
 sg13g2_fill_8 FILLER_37_1088 ();
 sg13g2_fill_8 FILLER_37_1096 ();
 sg13g2_fill_8 FILLER_37_1104 ();
 sg13g2_fill_8 FILLER_37_1112 ();
 sg13g2_fill_8 FILLER_37_1120 ();
 sg13g2_fill_8 FILLER_37_1128 ();
 sg13g2_fill_8 FILLER_37_1136 ();
 sg13g2_fill_8 FILLER_38_0 ();
 sg13g2_fill_8 FILLER_38_8 ();
 sg13g2_fill_8 FILLER_38_16 ();
 sg13g2_fill_8 FILLER_38_24 ();
 sg13g2_fill_8 FILLER_38_32 ();
 sg13g2_fill_8 FILLER_38_40 ();
 sg13g2_fill_8 FILLER_38_48 ();
 sg13g2_fill_8 FILLER_38_56 ();
 sg13g2_fill_8 FILLER_38_64 ();
 sg13g2_fill_8 FILLER_38_72 ();
 sg13g2_fill_8 FILLER_38_80 ();
 sg13g2_fill_8 FILLER_38_88 ();
 sg13g2_fill_8 FILLER_38_96 ();
 sg13g2_fill_8 FILLER_38_104 ();
 sg13g2_fill_8 FILLER_38_112 ();
 sg13g2_fill_8 FILLER_38_120 ();
 sg13g2_fill_8 FILLER_38_128 ();
 sg13g2_fill_8 FILLER_38_136 ();
 sg13g2_fill_8 FILLER_38_144 ();
 sg13g2_fill_8 FILLER_38_152 ();
 sg13g2_fill_8 FILLER_38_160 ();
 sg13g2_fill_8 FILLER_38_168 ();
 sg13g2_fill_8 FILLER_38_176 ();
 sg13g2_fill_8 FILLER_38_184 ();
 sg13g2_fill_8 FILLER_38_192 ();
 sg13g2_fill_8 FILLER_38_200 ();
 sg13g2_fill_8 FILLER_38_208 ();
 sg13g2_fill_8 FILLER_38_216 ();
 sg13g2_fill_8 FILLER_38_224 ();
 sg13g2_fill_8 FILLER_38_232 ();
 sg13g2_fill_8 FILLER_38_240 ();
 sg13g2_fill_8 FILLER_38_248 ();
 sg13g2_fill_8 FILLER_38_256 ();
 sg13g2_fill_8 FILLER_38_264 ();
 sg13g2_fill_8 FILLER_38_272 ();
 sg13g2_fill_8 FILLER_38_280 ();
 sg13g2_fill_8 FILLER_38_288 ();
 sg13g2_fill_8 FILLER_38_296 ();
 sg13g2_fill_8 FILLER_38_304 ();
 sg13g2_fill_8 FILLER_38_312 ();
 sg13g2_fill_8 FILLER_38_320 ();
 sg13g2_fill_8 FILLER_38_328 ();
 sg13g2_fill_8 FILLER_38_336 ();
 sg13g2_fill_8 FILLER_38_344 ();
 sg13g2_fill_8 FILLER_38_352 ();
 sg13g2_fill_8 FILLER_38_360 ();
 sg13g2_fill_8 FILLER_38_368 ();
 sg13g2_fill_8 FILLER_38_376 ();
 sg13g2_fill_8 FILLER_38_384 ();
 sg13g2_fill_8 FILLER_38_392 ();
 sg13g2_fill_8 FILLER_38_400 ();
 sg13g2_fill_8 FILLER_38_408 ();
 sg13g2_fill_8 FILLER_38_416 ();
 sg13g2_fill_8 FILLER_38_424 ();
 sg13g2_fill_8 FILLER_38_432 ();
 sg13g2_fill_8 FILLER_38_440 ();
 sg13g2_fill_8 FILLER_38_448 ();
 sg13g2_fill_8 FILLER_38_456 ();
 sg13g2_fill_8 FILLER_38_464 ();
 sg13g2_fill_8 FILLER_38_472 ();
 sg13g2_fill_8 FILLER_38_480 ();
 sg13g2_fill_8 FILLER_38_488 ();
 sg13g2_fill_8 FILLER_38_496 ();
 sg13g2_fill_8 FILLER_38_504 ();
 sg13g2_fill_8 FILLER_38_512 ();
 sg13g2_fill_8 FILLER_38_520 ();
 sg13g2_fill_8 FILLER_38_528 ();
 sg13g2_fill_8 FILLER_38_536 ();
 sg13g2_fill_8 FILLER_38_544 ();
 sg13g2_fill_8 FILLER_38_552 ();
 sg13g2_fill_8 FILLER_38_560 ();
 sg13g2_fill_8 FILLER_38_568 ();
 sg13g2_fill_8 FILLER_38_576 ();
 sg13g2_fill_8 FILLER_38_584 ();
 sg13g2_fill_8 FILLER_38_592 ();
 sg13g2_fill_8 FILLER_38_600 ();
 sg13g2_fill_8 FILLER_38_608 ();
 sg13g2_fill_8 FILLER_38_616 ();
 sg13g2_fill_8 FILLER_38_624 ();
 sg13g2_fill_8 FILLER_38_632 ();
 sg13g2_fill_8 FILLER_38_640 ();
 sg13g2_fill_8 FILLER_38_648 ();
 sg13g2_fill_8 FILLER_38_656 ();
 sg13g2_fill_8 FILLER_38_664 ();
 sg13g2_fill_8 FILLER_38_672 ();
 sg13g2_fill_8 FILLER_38_680 ();
 sg13g2_fill_8 FILLER_38_688 ();
 sg13g2_fill_8 FILLER_38_696 ();
 sg13g2_fill_8 FILLER_38_704 ();
 sg13g2_fill_8 FILLER_38_712 ();
 sg13g2_fill_8 FILLER_38_720 ();
 sg13g2_fill_8 FILLER_38_728 ();
 sg13g2_fill_8 FILLER_38_736 ();
 sg13g2_fill_8 FILLER_38_744 ();
 sg13g2_fill_8 FILLER_38_752 ();
 sg13g2_fill_8 FILLER_38_760 ();
 sg13g2_fill_8 FILLER_38_768 ();
 sg13g2_fill_8 FILLER_38_776 ();
 sg13g2_fill_8 FILLER_38_784 ();
 sg13g2_fill_8 FILLER_38_792 ();
 sg13g2_fill_8 FILLER_38_800 ();
 sg13g2_fill_8 FILLER_38_808 ();
 sg13g2_fill_8 FILLER_38_816 ();
 sg13g2_fill_8 FILLER_38_824 ();
 sg13g2_fill_8 FILLER_38_832 ();
 sg13g2_fill_8 FILLER_38_840 ();
 sg13g2_fill_8 FILLER_38_848 ();
 sg13g2_fill_8 FILLER_38_856 ();
 sg13g2_fill_8 FILLER_38_864 ();
 sg13g2_fill_8 FILLER_38_872 ();
 sg13g2_fill_8 FILLER_38_880 ();
 sg13g2_fill_8 FILLER_38_888 ();
 sg13g2_fill_8 FILLER_38_896 ();
 sg13g2_fill_8 FILLER_38_904 ();
 sg13g2_fill_8 FILLER_38_912 ();
 sg13g2_fill_8 FILLER_38_920 ();
 sg13g2_fill_8 FILLER_38_928 ();
 sg13g2_fill_8 FILLER_38_936 ();
 sg13g2_fill_8 FILLER_38_944 ();
 sg13g2_fill_8 FILLER_38_952 ();
 sg13g2_fill_8 FILLER_38_960 ();
 sg13g2_fill_8 FILLER_38_968 ();
 sg13g2_fill_8 FILLER_38_976 ();
 sg13g2_fill_8 FILLER_38_984 ();
 sg13g2_fill_8 FILLER_38_992 ();
 sg13g2_fill_8 FILLER_38_1000 ();
 sg13g2_fill_8 FILLER_38_1008 ();
 sg13g2_fill_8 FILLER_38_1016 ();
 sg13g2_fill_8 FILLER_38_1024 ();
 sg13g2_fill_8 FILLER_38_1032 ();
 sg13g2_fill_8 FILLER_38_1040 ();
 sg13g2_fill_8 FILLER_38_1048 ();
 sg13g2_fill_8 FILLER_38_1056 ();
 sg13g2_fill_8 FILLER_38_1064 ();
 sg13g2_fill_8 FILLER_38_1072 ();
 sg13g2_fill_8 FILLER_38_1080 ();
 sg13g2_fill_8 FILLER_38_1088 ();
 sg13g2_fill_8 FILLER_38_1096 ();
 sg13g2_fill_8 FILLER_38_1104 ();
 sg13g2_fill_8 FILLER_38_1112 ();
 sg13g2_fill_8 FILLER_38_1120 ();
 sg13g2_fill_8 FILLER_38_1128 ();
 sg13g2_fill_8 FILLER_38_1136 ();
 sg13g2_fill_8 FILLER_39_0 ();
 sg13g2_fill_8 FILLER_39_8 ();
 sg13g2_fill_8 FILLER_39_16 ();
 sg13g2_fill_8 FILLER_39_24 ();
 sg13g2_fill_8 FILLER_39_32 ();
 sg13g2_fill_8 FILLER_39_40 ();
 sg13g2_fill_8 FILLER_39_48 ();
 sg13g2_fill_8 FILLER_39_56 ();
 sg13g2_fill_8 FILLER_39_64 ();
 sg13g2_fill_8 FILLER_39_72 ();
 sg13g2_fill_8 FILLER_39_80 ();
 sg13g2_fill_8 FILLER_39_88 ();
 sg13g2_fill_8 FILLER_39_96 ();
 sg13g2_fill_8 FILLER_39_104 ();
 sg13g2_fill_8 FILLER_39_112 ();
 sg13g2_fill_8 FILLER_39_120 ();
 sg13g2_fill_8 FILLER_39_128 ();
 sg13g2_fill_8 FILLER_39_136 ();
 sg13g2_fill_8 FILLER_39_144 ();
 sg13g2_fill_8 FILLER_39_152 ();
 sg13g2_fill_8 FILLER_39_160 ();
 sg13g2_fill_8 FILLER_39_168 ();
 sg13g2_fill_8 FILLER_39_176 ();
 sg13g2_fill_8 FILLER_39_184 ();
 sg13g2_fill_8 FILLER_39_192 ();
 sg13g2_fill_8 FILLER_39_200 ();
 sg13g2_fill_8 FILLER_39_208 ();
 sg13g2_fill_8 FILLER_39_216 ();
 sg13g2_fill_8 FILLER_39_224 ();
 sg13g2_fill_8 FILLER_39_232 ();
 sg13g2_fill_8 FILLER_39_240 ();
 sg13g2_fill_8 FILLER_39_248 ();
 sg13g2_fill_8 FILLER_39_256 ();
 sg13g2_fill_8 FILLER_39_264 ();
 sg13g2_fill_8 FILLER_39_272 ();
 sg13g2_fill_8 FILLER_39_280 ();
 sg13g2_fill_8 FILLER_39_288 ();
 sg13g2_fill_8 FILLER_39_296 ();
 sg13g2_fill_8 FILLER_39_304 ();
 sg13g2_fill_8 FILLER_39_312 ();
 sg13g2_fill_8 FILLER_39_320 ();
 sg13g2_fill_8 FILLER_39_328 ();
 sg13g2_fill_8 FILLER_39_336 ();
 sg13g2_fill_8 FILLER_39_344 ();
 sg13g2_fill_8 FILLER_39_352 ();
 sg13g2_fill_8 FILLER_39_360 ();
 sg13g2_fill_8 FILLER_39_368 ();
 sg13g2_fill_8 FILLER_39_376 ();
 sg13g2_fill_8 FILLER_39_384 ();
 sg13g2_fill_8 FILLER_39_392 ();
 sg13g2_fill_8 FILLER_39_400 ();
 sg13g2_fill_8 FILLER_39_408 ();
 sg13g2_fill_8 FILLER_39_416 ();
 sg13g2_fill_8 FILLER_39_424 ();
 sg13g2_fill_8 FILLER_39_432 ();
 sg13g2_fill_8 FILLER_39_440 ();
 sg13g2_fill_8 FILLER_39_448 ();
 sg13g2_fill_8 FILLER_39_456 ();
 sg13g2_fill_8 FILLER_39_464 ();
 sg13g2_fill_8 FILLER_39_472 ();
 sg13g2_fill_8 FILLER_39_480 ();
 sg13g2_fill_8 FILLER_39_488 ();
 sg13g2_fill_8 FILLER_39_496 ();
 sg13g2_fill_8 FILLER_39_504 ();
 sg13g2_fill_8 FILLER_39_512 ();
 sg13g2_fill_8 FILLER_39_520 ();
 sg13g2_fill_8 FILLER_39_528 ();
 sg13g2_fill_8 FILLER_39_536 ();
 sg13g2_fill_8 FILLER_39_544 ();
 sg13g2_fill_8 FILLER_39_552 ();
 sg13g2_fill_8 FILLER_39_560 ();
 sg13g2_fill_8 FILLER_39_568 ();
 sg13g2_fill_8 FILLER_39_576 ();
 sg13g2_fill_8 FILLER_39_584 ();
 sg13g2_fill_8 FILLER_39_592 ();
 sg13g2_fill_8 FILLER_39_600 ();
 sg13g2_fill_8 FILLER_39_608 ();
 sg13g2_fill_8 FILLER_39_616 ();
 sg13g2_fill_8 FILLER_39_624 ();
 sg13g2_fill_8 FILLER_39_632 ();
 sg13g2_fill_8 FILLER_39_640 ();
 sg13g2_fill_8 FILLER_39_648 ();
 sg13g2_fill_8 FILLER_39_656 ();
 sg13g2_fill_8 FILLER_39_664 ();
 sg13g2_fill_8 FILLER_39_672 ();
 sg13g2_fill_8 FILLER_39_680 ();
 sg13g2_fill_8 FILLER_39_688 ();
 sg13g2_fill_8 FILLER_39_696 ();
 sg13g2_fill_8 FILLER_39_704 ();
 sg13g2_fill_8 FILLER_39_712 ();
 sg13g2_fill_8 FILLER_39_720 ();
 sg13g2_fill_8 FILLER_39_728 ();
 sg13g2_fill_8 FILLER_39_736 ();
 sg13g2_fill_8 FILLER_39_744 ();
 sg13g2_fill_8 FILLER_39_752 ();
 sg13g2_fill_8 FILLER_39_760 ();
 sg13g2_fill_8 FILLER_39_768 ();
 sg13g2_fill_8 FILLER_39_776 ();
 sg13g2_fill_8 FILLER_39_784 ();
 sg13g2_fill_8 FILLER_39_792 ();
 sg13g2_fill_8 FILLER_39_800 ();
 sg13g2_fill_8 FILLER_39_808 ();
 sg13g2_fill_8 FILLER_39_816 ();
 sg13g2_fill_8 FILLER_39_824 ();
 sg13g2_fill_8 FILLER_39_832 ();
 sg13g2_fill_8 FILLER_39_840 ();
 sg13g2_fill_8 FILLER_39_848 ();
 sg13g2_fill_8 FILLER_39_856 ();
 sg13g2_fill_8 FILLER_39_864 ();
 sg13g2_fill_8 FILLER_39_872 ();
 sg13g2_fill_8 FILLER_39_880 ();
 sg13g2_fill_8 FILLER_39_888 ();
 sg13g2_fill_8 FILLER_39_896 ();
 sg13g2_fill_8 FILLER_39_904 ();
 sg13g2_fill_8 FILLER_39_912 ();
 sg13g2_fill_8 FILLER_39_920 ();
 sg13g2_fill_8 FILLER_39_928 ();
 sg13g2_fill_8 FILLER_39_936 ();
 sg13g2_fill_8 FILLER_39_944 ();
 sg13g2_fill_8 FILLER_39_952 ();
 sg13g2_fill_8 FILLER_39_960 ();
 sg13g2_fill_8 FILLER_39_968 ();
 sg13g2_fill_8 FILLER_39_976 ();
 sg13g2_fill_8 FILLER_39_984 ();
 sg13g2_fill_8 FILLER_39_992 ();
 sg13g2_fill_8 FILLER_39_1000 ();
 sg13g2_fill_8 FILLER_39_1008 ();
 sg13g2_fill_8 FILLER_39_1016 ();
 sg13g2_fill_8 FILLER_39_1024 ();
 sg13g2_fill_8 FILLER_39_1032 ();
 sg13g2_fill_8 FILLER_39_1040 ();
 sg13g2_fill_8 FILLER_39_1048 ();
 sg13g2_fill_8 FILLER_39_1056 ();
 sg13g2_fill_8 FILLER_39_1064 ();
 sg13g2_fill_8 FILLER_39_1072 ();
 sg13g2_fill_8 FILLER_39_1080 ();
 sg13g2_fill_8 FILLER_39_1088 ();
 sg13g2_fill_8 FILLER_39_1096 ();
 sg13g2_fill_8 FILLER_39_1104 ();
 sg13g2_fill_8 FILLER_39_1112 ();
 sg13g2_fill_8 FILLER_39_1120 ();
 sg13g2_fill_8 FILLER_39_1128 ();
 sg13g2_fill_8 FILLER_39_1136 ();
 sg13g2_fill_8 FILLER_40_0 ();
 sg13g2_fill_8 FILLER_40_8 ();
 sg13g2_fill_8 FILLER_40_16 ();
 sg13g2_fill_8 FILLER_40_24 ();
 sg13g2_fill_8 FILLER_40_32 ();
 sg13g2_fill_8 FILLER_40_40 ();
 sg13g2_fill_8 FILLER_40_48 ();
 sg13g2_fill_8 FILLER_40_56 ();
 sg13g2_fill_8 FILLER_40_64 ();
 sg13g2_fill_8 FILLER_40_72 ();
 sg13g2_fill_8 FILLER_40_80 ();
 sg13g2_fill_8 FILLER_40_88 ();
 sg13g2_fill_8 FILLER_40_96 ();
 sg13g2_fill_8 FILLER_40_104 ();
 sg13g2_fill_8 FILLER_40_112 ();
 sg13g2_fill_8 FILLER_40_120 ();
 sg13g2_fill_8 FILLER_40_128 ();
 sg13g2_fill_8 FILLER_40_136 ();
 sg13g2_fill_8 FILLER_40_144 ();
 sg13g2_fill_8 FILLER_40_152 ();
 sg13g2_fill_8 FILLER_40_160 ();
 sg13g2_fill_8 FILLER_40_168 ();
 sg13g2_fill_8 FILLER_40_176 ();
 sg13g2_fill_8 FILLER_40_184 ();
 sg13g2_fill_8 FILLER_40_192 ();
 sg13g2_fill_8 FILLER_40_200 ();
 sg13g2_fill_8 FILLER_40_208 ();
 sg13g2_fill_8 FILLER_40_216 ();
 sg13g2_fill_8 FILLER_40_224 ();
 sg13g2_fill_8 FILLER_40_232 ();
 sg13g2_fill_8 FILLER_40_240 ();
 sg13g2_fill_8 FILLER_40_248 ();
 sg13g2_fill_8 FILLER_40_256 ();
 sg13g2_fill_8 FILLER_40_264 ();
 sg13g2_fill_8 FILLER_40_272 ();
 sg13g2_fill_8 FILLER_40_280 ();
 sg13g2_fill_8 FILLER_40_288 ();
 sg13g2_fill_8 FILLER_40_296 ();
 sg13g2_fill_8 FILLER_40_304 ();
 sg13g2_fill_8 FILLER_40_312 ();
 sg13g2_fill_8 FILLER_40_320 ();
 sg13g2_fill_8 FILLER_40_328 ();
 sg13g2_fill_8 FILLER_40_336 ();
 sg13g2_fill_8 FILLER_40_344 ();
 sg13g2_fill_8 FILLER_40_352 ();
 sg13g2_fill_8 FILLER_40_360 ();
 sg13g2_fill_8 FILLER_40_368 ();
 sg13g2_fill_8 FILLER_40_376 ();
 sg13g2_fill_8 FILLER_40_384 ();
 sg13g2_fill_8 FILLER_40_392 ();
 sg13g2_fill_8 FILLER_40_400 ();
 sg13g2_fill_8 FILLER_40_408 ();
 sg13g2_fill_8 FILLER_40_416 ();
 sg13g2_fill_8 FILLER_40_424 ();
 sg13g2_fill_8 FILLER_40_432 ();
 sg13g2_fill_8 FILLER_40_440 ();
 sg13g2_fill_8 FILLER_40_448 ();
 sg13g2_fill_8 FILLER_40_456 ();
 sg13g2_fill_8 FILLER_40_464 ();
 sg13g2_fill_8 FILLER_40_472 ();
 sg13g2_fill_8 FILLER_40_480 ();
 sg13g2_fill_8 FILLER_40_488 ();
 sg13g2_fill_8 FILLER_40_496 ();
 sg13g2_fill_8 FILLER_40_504 ();
 sg13g2_fill_8 FILLER_40_512 ();
 sg13g2_fill_8 FILLER_40_520 ();
 sg13g2_fill_8 FILLER_40_528 ();
 sg13g2_fill_8 FILLER_40_536 ();
 sg13g2_fill_8 FILLER_40_544 ();
 sg13g2_fill_8 FILLER_40_552 ();
 sg13g2_fill_8 FILLER_40_560 ();
 sg13g2_fill_8 FILLER_40_568 ();
 sg13g2_fill_8 FILLER_40_576 ();
 sg13g2_fill_8 FILLER_40_584 ();
 sg13g2_fill_8 FILLER_40_592 ();
 sg13g2_fill_8 FILLER_40_600 ();
 sg13g2_fill_8 FILLER_40_608 ();
 sg13g2_fill_8 FILLER_40_616 ();
 sg13g2_fill_8 FILLER_40_624 ();
 sg13g2_fill_8 FILLER_40_632 ();
 sg13g2_fill_8 FILLER_40_640 ();
 sg13g2_fill_8 FILLER_40_648 ();
 sg13g2_fill_8 FILLER_40_656 ();
 sg13g2_fill_8 FILLER_40_664 ();
 sg13g2_fill_8 FILLER_40_672 ();
 sg13g2_fill_8 FILLER_40_680 ();
 sg13g2_fill_8 FILLER_40_688 ();
 sg13g2_fill_8 FILLER_40_696 ();
 sg13g2_fill_8 FILLER_40_704 ();
 sg13g2_fill_8 FILLER_40_712 ();
 sg13g2_fill_8 FILLER_40_720 ();
 sg13g2_fill_8 FILLER_40_728 ();
 sg13g2_fill_8 FILLER_40_736 ();
 sg13g2_fill_8 FILLER_40_744 ();
 sg13g2_fill_8 FILLER_40_752 ();
 sg13g2_fill_8 FILLER_40_760 ();
 sg13g2_fill_8 FILLER_40_768 ();
 sg13g2_fill_8 FILLER_40_776 ();
 sg13g2_fill_8 FILLER_40_784 ();
 sg13g2_fill_8 FILLER_40_792 ();
 sg13g2_fill_8 FILLER_40_800 ();
 sg13g2_fill_8 FILLER_40_808 ();
 sg13g2_fill_8 FILLER_40_816 ();
 sg13g2_fill_8 FILLER_40_824 ();
 sg13g2_fill_8 FILLER_40_832 ();
 sg13g2_fill_8 FILLER_40_840 ();
 sg13g2_fill_8 FILLER_40_848 ();
 sg13g2_fill_8 FILLER_40_856 ();
 sg13g2_fill_8 FILLER_40_864 ();
 sg13g2_fill_8 FILLER_40_872 ();
 sg13g2_fill_8 FILLER_40_880 ();
 sg13g2_fill_8 FILLER_40_888 ();
 sg13g2_fill_8 FILLER_40_896 ();
 sg13g2_fill_8 FILLER_40_904 ();
 sg13g2_fill_8 FILLER_40_912 ();
 sg13g2_fill_8 FILLER_40_920 ();
 sg13g2_fill_8 FILLER_40_928 ();
 sg13g2_fill_8 FILLER_40_936 ();
 sg13g2_fill_8 FILLER_40_944 ();
 sg13g2_fill_8 FILLER_40_952 ();
 sg13g2_fill_8 FILLER_40_960 ();
 sg13g2_fill_8 FILLER_40_968 ();
 sg13g2_fill_8 FILLER_40_976 ();
 sg13g2_fill_8 FILLER_40_984 ();
 sg13g2_fill_8 FILLER_40_992 ();
 sg13g2_fill_8 FILLER_40_1000 ();
 sg13g2_fill_8 FILLER_40_1008 ();
 sg13g2_fill_8 FILLER_40_1016 ();
 sg13g2_fill_8 FILLER_40_1024 ();
 sg13g2_fill_8 FILLER_40_1032 ();
 sg13g2_fill_8 FILLER_40_1040 ();
 sg13g2_fill_8 FILLER_40_1048 ();
 sg13g2_fill_8 FILLER_40_1056 ();
 sg13g2_fill_8 FILLER_40_1064 ();
 sg13g2_fill_8 FILLER_40_1072 ();
 sg13g2_fill_8 FILLER_40_1080 ();
 sg13g2_fill_8 FILLER_40_1088 ();
 sg13g2_fill_8 FILLER_40_1096 ();
 sg13g2_fill_8 FILLER_40_1104 ();
 sg13g2_fill_8 FILLER_40_1112 ();
 sg13g2_fill_8 FILLER_40_1120 ();
 sg13g2_fill_8 FILLER_40_1128 ();
 sg13g2_fill_8 FILLER_40_1136 ();
 sg13g2_fill_8 FILLER_41_0 ();
 sg13g2_fill_8 FILLER_41_8 ();
 sg13g2_fill_8 FILLER_41_16 ();
 sg13g2_fill_8 FILLER_41_24 ();
 sg13g2_fill_8 FILLER_41_32 ();
 sg13g2_fill_8 FILLER_41_40 ();
 sg13g2_fill_8 FILLER_41_48 ();
 sg13g2_fill_8 FILLER_41_56 ();
 sg13g2_fill_8 FILLER_41_64 ();
 sg13g2_fill_8 FILLER_41_72 ();
 sg13g2_fill_8 FILLER_41_80 ();
 sg13g2_fill_8 FILLER_41_88 ();
 sg13g2_fill_8 FILLER_41_96 ();
 sg13g2_fill_8 FILLER_41_104 ();
 sg13g2_fill_8 FILLER_41_112 ();
 sg13g2_fill_8 FILLER_41_120 ();
 sg13g2_fill_8 FILLER_41_128 ();
 sg13g2_fill_8 FILLER_41_136 ();
 sg13g2_fill_8 FILLER_41_144 ();
 sg13g2_fill_8 FILLER_41_152 ();
 sg13g2_fill_8 FILLER_41_160 ();
 sg13g2_fill_8 FILLER_41_168 ();
 sg13g2_fill_8 FILLER_41_176 ();
 sg13g2_fill_8 FILLER_41_184 ();
 sg13g2_fill_8 FILLER_41_192 ();
 sg13g2_fill_8 FILLER_41_200 ();
 sg13g2_fill_8 FILLER_41_208 ();
 sg13g2_fill_8 FILLER_41_216 ();
 sg13g2_fill_8 FILLER_41_224 ();
 sg13g2_fill_8 FILLER_41_232 ();
 sg13g2_fill_8 FILLER_41_240 ();
 sg13g2_fill_8 FILLER_41_248 ();
 sg13g2_fill_8 FILLER_41_256 ();
 sg13g2_fill_8 FILLER_41_264 ();
 sg13g2_fill_8 FILLER_41_272 ();
 sg13g2_fill_8 FILLER_41_280 ();
 sg13g2_fill_8 FILLER_41_288 ();
 sg13g2_fill_8 FILLER_41_296 ();
 sg13g2_fill_8 FILLER_41_304 ();
 sg13g2_fill_8 FILLER_41_312 ();
 sg13g2_fill_8 FILLER_41_320 ();
 sg13g2_fill_8 FILLER_41_328 ();
 sg13g2_fill_8 FILLER_41_336 ();
 sg13g2_fill_8 FILLER_41_344 ();
 sg13g2_fill_8 FILLER_41_352 ();
 sg13g2_fill_8 FILLER_41_360 ();
 sg13g2_fill_8 FILLER_41_368 ();
 sg13g2_fill_8 FILLER_41_376 ();
 sg13g2_fill_8 FILLER_41_384 ();
 sg13g2_fill_8 FILLER_41_392 ();
 sg13g2_fill_8 FILLER_41_400 ();
 sg13g2_fill_8 FILLER_41_408 ();
 sg13g2_fill_8 FILLER_41_416 ();
 sg13g2_fill_8 FILLER_41_424 ();
 sg13g2_fill_8 FILLER_41_432 ();
 sg13g2_fill_8 FILLER_41_440 ();
 sg13g2_fill_8 FILLER_41_448 ();
 sg13g2_fill_8 FILLER_41_456 ();
 sg13g2_fill_8 FILLER_41_464 ();
 sg13g2_fill_8 FILLER_41_472 ();
 sg13g2_fill_8 FILLER_41_480 ();
 sg13g2_fill_8 FILLER_41_488 ();
 sg13g2_fill_8 FILLER_41_496 ();
 sg13g2_fill_8 FILLER_41_504 ();
 sg13g2_fill_8 FILLER_41_512 ();
 sg13g2_fill_8 FILLER_41_520 ();
 sg13g2_fill_8 FILLER_41_528 ();
 sg13g2_fill_8 FILLER_41_536 ();
 sg13g2_fill_8 FILLER_41_544 ();
 sg13g2_fill_8 FILLER_41_552 ();
 sg13g2_fill_8 FILLER_41_560 ();
 sg13g2_fill_8 FILLER_41_568 ();
 sg13g2_fill_8 FILLER_41_576 ();
 sg13g2_fill_8 FILLER_41_584 ();
 sg13g2_fill_8 FILLER_41_592 ();
 sg13g2_fill_8 FILLER_41_600 ();
 sg13g2_fill_8 FILLER_41_608 ();
 sg13g2_fill_8 FILLER_41_616 ();
 sg13g2_fill_8 FILLER_41_624 ();
 sg13g2_fill_8 FILLER_41_632 ();
 sg13g2_fill_8 FILLER_41_640 ();
 sg13g2_fill_8 FILLER_41_648 ();
 sg13g2_fill_8 FILLER_41_656 ();
 sg13g2_fill_8 FILLER_41_664 ();
 sg13g2_fill_8 FILLER_41_672 ();
 sg13g2_fill_8 FILLER_41_680 ();
 sg13g2_fill_8 FILLER_41_688 ();
 sg13g2_fill_8 FILLER_41_696 ();
 sg13g2_fill_8 FILLER_41_704 ();
 sg13g2_fill_8 FILLER_41_712 ();
 sg13g2_fill_8 FILLER_41_720 ();
 sg13g2_fill_8 FILLER_41_728 ();
 sg13g2_fill_8 FILLER_41_736 ();
 sg13g2_fill_8 FILLER_41_744 ();
 sg13g2_fill_8 FILLER_41_752 ();
 sg13g2_fill_8 FILLER_41_760 ();
 sg13g2_fill_8 FILLER_41_768 ();
 sg13g2_fill_8 FILLER_41_776 ();
 sg13g2_fill_8 FILLER_41_784 ();
 sg13g2_fill_8 FILLER_41_792 ();
 sg13g2_fill_8 FILLER_41_800 ();
 sg13g2_fill_8 FILLER_41_808 ();
 sg13g2_fill_8 FILLER_41_816 ();
 sg13g2_fill_8 FILLER_41_824 ();
 sg13g2_fill_8 FILLER_41_832 ();
 sg13g2_fill_8 FILLER_41_840 ();
 sg13g2_fill_8 FILLER_41_848 ();
 sg13g2_fill_8 FILLER_41_856 ();
 sg13g2_fill_8 FILLER_41_864 ();
 sg13g2_fill_8 FILLER_41_872 ();
 sg13g2_fill_8 FILLER_41_880 ();
 sg13g2_fill_8 FILLER_41_888 ();
 sg13g2_fill_8 FILLER_41_896 ();
 sg13g2_fill_8 FILLER_41_904 ();
 sg13g2_fill_8 FILLER_41_912 ();
 sg13g2_fill_8 FILLER_41_920 ();
 sg13g2_fill_8 FILLER_41_928 ();
 sg13g2_fill_8 FILLER_41_936 ();
 sg13g2_fill_8 FILLER_41_944 ();
 sg13g2_fill_8 FILLER_41_952 ();
 sg13g2_fill_8 FILLER_41_960 ();
 sg13g2_fill_8 FILLER_41_968 ();
 sg13g2_fill_8 FILLER_41_976 ();
 sg13g2_fill_8 FILLER_41_984 ();
 sg13g2_fill_8 FILLER_41_992 ();
 sg13g2_fill_8 FILLER_41_1000 ();
 sg13g2_fill_8 FILLER_41_1008 ();
 sg13g2_fill_8 FILLER_41_1016 ();
 sg13g2_fill_8 FILLER_41_1024 ();
 sg13g2_fill_8 FILLER_41_1032 ();
 sg13g2_fill_8 FILLER_41_1040 ();
 sg13g2_fill_8 FILLER_41_1048 ();
 sg13g2_fill_8 FILLER_41_1056 ();
 sg13g2_fill_8 FILLER_41_1064 ();
 sg13g2_fill_8 FILLER_41_1072 ();
 sg13g2_fill_8 FILLER_41_1080 ();
 sg13g2_fill_8 FILLER_41_1088 ();
 sg13g2_fill_8 FILLER_41_1096 ();
 sg13g2_fill_8 FILLER_41_1104 ();
 sg13g2_fill_8 FILLER_41_1112 ();
 sg13g2_fill_8 FILLER_41_1120 ();
 sg13g2_fill_8 FILLER_41_1128 ();
 sg13g2_fill_8 FILLER_41_1136 ();
 sg13g2_fill_8 FILLER_42_0 ();
 sg13g2_fill_8 FILLER_42_8 ();
 sg13g2_fill_8 FILLER_42_16 ();
 sg13g2_fill_8 FILLER_42_24 ();
 sg13g2_fill_8 FILLER_42_32 ();
 sg13g2_fill_8 FILLER_42_40 ();
 sg13g2_fill_8 FILLER_42_48 ();
 sg13g2_fill_8 FILLER_42_56 ();
 sg13g2_fill_8 FILLER_42_64 ();
 sg13g2_fill_8 FILLER_42_72 ();
 sg13g2_fill_8 FILLER_42_80 ();
 sg13g2_fill_8 FILLER_42_88 ();
 sg13g2_fill_8 FILLER_42_96 ();
 sg13g2_fill_8 FILLER_42_104 ();
 sg13g2_fill_8 FILLER_42_112 ();
 sg13g2_fill_8 FILLER_42_120 ();
 sg13g2_fill_8 FILLER_42_128 ();
 sg13g2_fill_8 FILLER_42_136 ();
 sg13g2_fill_8 FILLER_42_144 ();
 sg13g2_fill_8 FILLER_42_152 ();
 sg13g2_fill_8 FILLER_42_160 ();
 sg13g2_fill_8 FILLER_42_168 ();
 sg13g2_fill_8 FILLER_42_176 ();
 sg13g2_fill_8 FILLER_42_184 ();
 sg13g2_fill_8 FILLER_42_192 ();
 sg13g2_fill_8 FILLER_42_200 ();
 sg13g2_fill_8 FILLER_42_208 ();
 sg13g2_fill_8 FILLER_42_216 ();
 sg13g2_fill_8 FILLER_42_224 ();
 sg13g2_fill_8 FILLER_42_232 ();
 sg13g2_fill_8 FILLER_42_240 ();
 sg13g2_fill_8 FILLER_42_248 ();
 sg13g2_fill_8 FILLER_42_256 ();
 sg13g2_fill_8 FILLER_42_264 ();
 sg13g2_fill_8 FILLER_42_272 ();
 sg13g2_fill_8 FILLER_42_280 ();
 sg13g2_fill_8 FILLER_42_288 ();
 sg13g2_fill_8 FILLER_42_296 ();
 sg13g2_fill_8 FILLER_42_304 ();
 sg13g2_fill_8 FILLER_42_312 ();
 sg13g2_fill_8 FILLER_42_320 ();
 sg13g2_fill_8 FILLER_42_328 ();
 sg13g2_fill_8 FILLER_42_336 ();
 sg13g2_fill_8 FILLER_42_344 ();
 sg13g2_fill_8 FILLER_42_352 ();
 sg13g2_fill_8 FILLER_42_360 ();
 sg13g2_fill_8 FILLER_42_368 ();
 sg13g2_fill_8 FILLER_42_376 ();
 sg13g2_fill_8 FILLER_42_384 ();
 sg13g2_fill_8 FILLER_42_392 ();
 sg13g2_fill_8 FILLER_42_400 ();
 sg13g2_fill_8 FILLER_42_408 ();
 sg13g2_fill_8 FILLER_42_416 ();
 sg13g2_fill_8 FILLER_42_424 ();
 sg13g2_fill_8 FILLER_42_432 ();
 sg13g2_fill_8 FILLER_42_440 ();
 sg13g2_fill_8 FILLER_42_448 ();
 sg13g2_fill_8 FILLER_42_456 ();
 sg13g2_fill_8 FILLER_42_464 ();
 sg13g2_fill_8 FILLER_42_472 ();
 sg13g2_fill_8 FILLER_42_480 ();
 sg13g2_fill_8 FILLER_42_488 ();
 sg13g2_fill_8 FILLER_42_496 ();
 sg13g2_fill_8 FILLER_42_504 ();
 sg13g2_fill_8 FILLER_42_512 ();
 sg13g2_fill_8 FILLER_42_520 ();
 sg13g2_fill_8 FILLER_42_528 ();
 sg13g2_fill_8 FILLER_42_536 ();
 sg13g2_fill_8 FILLER_42_544 ();
 sg13g2_fill_8 FILLER_42_552 ();
 sg13g2_fill_8 FILLER_42_560 ();
 sg13g2_fill_8 FILLER_42_568 ();
 sg13g2_fill_8 FILLER_42_576 ();
 sg13g2_fill_8 FILLER_42_584 ();
 sg13g2_fill_8 FILLER_42_592 ();
 sg13g2_fill_8 FILLER_42_600 ();
 sg13g2_fill_8 FILLER_42_608 ();
 sg13g2_fill_8 FILLER_42_616 ();
 sg13g2_fill_8 FILLER_42_624 ();
 sg13g2_fill_8 FILLER_42_632 ();
 sg13g2_fill_8 FILLER_42_640 ();
 sg13g2_fill_8 FILLER_42_648 ();
 sg13g2_fill_8 FILLER_42_656 ();
 sg13g2_fill_8 FILLER_42_664 ();
 sg13g2_fill_8 FILLER_42_672 ();
 sg13g2_fill_8 FILLER_42_680 ();
 sg13g2_fill_8 FILLER_42_688 ();
 sg13g2_fill_8 FILLER_42_696 ();
 sg13g2_fill_8 FILLER_42_704 ();
 sg13g2_fill_8 FILLER_42_712 ();
 sg13g2_fill_8 FILLER_42_720 ();
 sg13g2_fill_8 FILLER_42_728 ();
 sg13g2_fill_8 FILLER_42_736 ();
 sg13g2_fill_8 FILLER_42_744 ();
 sg13g2_fill_8 FILLER_42_752 ();
 sg13g2_fill_8 FILLER_42_760 ();
 sg13g2_fill_8 FILLER_42_768 ();
 sg13g2_fill_8 FILLER_42_776 ();
 sg13g2_fill_8 FILLER_42_784 ();
 sg13g2_fill_8 FILLER_42_792 ();
 sg13g2_fill_8 FILLER_42_800 ();
 sg13g2_fill_8 FILLER_42_808 ();
 sg13g2_fill_8 FILLER_42_816 ();
 sg13g2_fill_8 FILLER_42_824 ();
 sg13g2_fill_8 FILLER_42_832 ();
 sg13g2_fill_8 FILLER_42_840 ();
 sg13g2_fill_8 FILLER_42_848 ();
 sg13g2_fill_8 FILLER_42_856 ();
 sg13g2_fill_8 FILLER_42_864 ();
 sg13g2_fill_8 FILLER_42_872 ();
 sg13g2_fill_8 FILLER_42_880 ();
 sg13g2_fill_8 FILLER_42_888 ();
 sg13g2_fill_8 FILLER_42_896 ();
 sg13g2_fill_8 FILLER_42_904 ();
 sg13g2_fill_8 FILLER_42_912 ();
 sg13g2_fill_8 FILLER_42_920 ();
 sg13g2_fill_8 FILLER_42_928 ();
 sg13g2_fill_8 FILLER_42_936 ();
 sg13g2_fill_8 FILLER_42_944 ();
 sg13g2_fill_8 FILLER_42_952 ();
 sg13g2_fill_8 FILLER_42_960 ();
 sg13g2_fill_8 FILLER_42_968 ();
 sg13g2_fill_8 FILLER_42_976 ();
 sg13g2_fill_8 FILLER_42_984 ();
 sg13g2_fill_8 FILLER_42_992 ();
 sg13g2_fill_8 FILLER_42_1000 ();
 sg13g2_fill_8 FILLER_42_1008 ();
 sg13g2_fill_8 FILLER_42_1016 ();
 sg13g2_fill_8 FILLER_42_1024 ();
 sg13g2_fill_8 FILLER_42_1032 ();
 sg13g2_fill_8 FILLER_42_1040 ();
 sg13g2_fill_8 FILLER_42_1048 ();
 sg13g2_fill_8 FILLER_42_1056 ();
 sg13g2_fill_8 FILLER_42_1064 ();
 sg13g2_fill_8 FILLER_42_1072 ();
 sg13g2_fill_8 FILLER_42_1080 ();
 sg13g2_fill_8 FILLER_42_1088 ();
 sg13g2_fill_8 FILLER_42_1096 ();
 sg13g2_fill_8 FILLER_42_1104 ();
 sg13g2_fill_8 FILLER_42_1112 ();
 sg13g2_fill_8 FILLER_42_1120 ();
 sg13g2_fill_8 FILLER_42_1128 ();
 sg13g2_fill_8 FILLER_42_1136 ();
 sg13g2_fill_8 FILLER_43_0 ();
 sg13g2_fill_8 FILLER_43_8 ();
 sg13g2_fill_8 FILLER_43_16 ();
 sg13g2_fill_8 FILLER_43_24 ();
 sg13g2_fill_8 FILLER_43_32 ();
 sg13g2_fill_8 FILLER_43_40 ();
 sg13g2_fill_8 FILLER_43_48 ();
 sg13g2_fill_8 FILLER_43_56 ();
 sg13g2_fill_8 FILLER_43_64 ();
 sg13g2_fill_8 FILLER_43_72 ();
 sg13g2_fill_8 FILLER_43_80 ();
 sg13g2_fill_8 FILLER_43_88 ();
 sg13g2_fill_8 FILLER_43_96 ();
 sg13g2_fill_8 FILLER_43_104 ();
 sg13g2_fill_8 FILLER_43_112 ();
 sg13g2_fill_8 FILLER_43_120 ();
 sg13g2_fill_8 FILLER_43_128 ();
 sg13g2_fill_8 FILLER_43_136 ();
 sg13g2_fill_8 FILLER_43_144 ();
 sg13g2_fill_8 FILLER_43_152 ();
 sg13g2_fill_8 FILLER_43_160 ();
 sg13g2_fill_8 FILLER_43_168 ();
 sg13g2_fill_8 FILLER_43_176 ();
 sg13g2_fill_8 FILLER_43_184 ();
 sg13g2_fill_8 FILLER_43_192 ();
 sg13g2_fill_8 FILLER_43_200 ();
 sg13g2_fill_8 FILLER_43_208 ();
 sg13g2_fill_8 FILLER_43_216 ();
 sg13g2_fill_8 FILLER_43_224 ();
 sg13g2_fill_8 FILLER_43_232 ();
 sg13g2_fill_8 FILLER_43_240 ();
 sg13g2_fill_8 FILLER_43_248 ();
 sg13g2_fill_8 FILLER_43_256 ();
 sg13g2_fill_8 FILLER_43_264 ();
 sg13g2_fill_8 FILLER_43_272 ();
 sg13g2_fill_8 FILLER_43_280 ();
 sg13g2_fill_8 FILLER_43_288 ();
 sg13g2_fill_8 FILLER_43_296 ();
 sg13g2_fill_8 FILLER_43_304 ();
 sg13g2_fill_8 FILLER_43_312 ();
 sg13g2_fill_8 FILLER_43_320 ();
 sg13g2_fill_8 FILLER_43_328 ();
 sg13g2_fill_8 FILLER_43_336 ();
 sg13g2_fill_8 FILLER_43_344 ();
 sg13g2_fill_8 FILLER_43_352 ();
 sg13g2_fill_8 FILLER_43_360 ();
 sg13g2_fill_8 FILLER_43_368 ();
 sg13g2_fill_8 FILLER_43_376 ();
 sg13g2_fill_8 FILLER_43_384 ();
 sg13g2_fill_8 FILLER_43_392 ();
 sg13g2_fill_8 FILLER_43_400 ();
 sg13g2_fill_8 FILLER_43_408 ();
 sg13g2_fill_8 FILLER_43_416 ();
 sg13g2_fill_8 FILLER_43_424 ();
 sg13g2_fill_8 FILLER_43_432 ();
 sg13g2_fill_8 FILLER_43_440 ();
 sg13g2_fill_8 FILLER_43_448 ();
 sg13g2_fill_8 FILLER_43_456 ();
 sg13g2_fill_8 FILLER_43_464 ();
 sg13g2_fill_8 FILLER_43_472 ();
 sg13g2_fill_8 FILLER_43_480 ();
 sg13g2_fill_8 FILLER_43_488 ();
 sg13g2_fill_8 FILLER_43_496 ();
 sg13g2_fill_8 FILLER_43_504 ();
 sg13g2_fill_8 FILLER_43_512 ();
 sg13g2_fill_8 FILLER_43_520 ();
 sg13g2_fill_8 FILLER_43_528 ();
 sg13g2_fill_8 FILLER_43_536 ();
 sg13g2_fill_8 FILLER_43_544 ();
 sg13g2_fill_8 FILLER_43_552 ();
 sg13g2_fill_8 FILLER_43_560 ();
 sg13g2_fill_8 FILLER_43_568 ();
 sg13g2_fill_8 FILLER_43_576 ();
 sg13g2_fill_8 FILLER_43_584 ();
 sg13g2_fill_8 FILLER_43_592 ();
 sg13g2_fill_8 FILLER_43_600 ();
 sg13g2_fill_8 FILLER_43_608 ();
 sg13g2_fill_8 FILLER_43_616 ();
 sg13g2_fill_8 FILLER_43_624 ();
 sg13g2_fill_8 FILLER_43_632 ();
 sg13g2_fill_8 FILLER_43_640 ();
 sg13g2_fill_8 FILLER_43_648 ();
 sg13g2_fill_8 FILLER_43_656 ();
 sg13g2_fill_8 FILLER_43_664 ();
 sg13g2_fill_8 FILLER_43_672 ();
 sg13g2_fill_8 FILLER_43_680 ();
 sg13g2_fill_8 FILLER_43_688 ();
 sg13g2_fill_8 FILLER_43_696 ();
 sg13g2_fill_8 FILLER_43_704 ();
 sg13g2_fill_8 FILLER_43_712 ();
 sg13g2_fill_8 FILLER_43_720 ();
 sg13g2_fill_8 FILLER_43_728 ();
 sg13g2_fill_8 FILLER_43_736 ();
 sg13g2_fill_8 FILLER_43_744 ();
 sg13g2_fill_8 FILLER_43_752 ();
 sg13g2_fill_8 FILLER_43_760 ();
 sg13g2_fill_8 FILLER_43_768 ();
 sg13g2_fill_8 FILLER_43_776 ();
 sg13g2_fill_8 FILLER_43_784 ();
 sg13g2_fill_8 FILLER_43_792 ();
 sg13g2_fill_8 FILLER_43_800 ();
 sg13g2_fill_8 FILLER_43_808 ();
 sg13g2_fill_8 FILLER_43_816 ();
 sg13g2_fill_8 FILLER_43_824 ();
 sg13g2_fill_8 FILLER_43_832 ();
 sg13g2_fill_8 FILLER_43_840 ();
 sg13g2_fill_8 FILLER_43_848 ();
 sg13g2_fill_8 FILLER_43_856 ();
 sg13g2_fill_8 FILLER_43_864 ();
 sg13g2_fill_8 FILLER_43_872 ();
 sg13g2_fill_8 FILLER_43_880 ();
 sg13g2_fill_8 FILLER_43_888 ();
 sg13g2_fill_8 FILLER_43_896 ();
 sg13g2_fill_8 FILLER_43_904 ();
 sg13g2_fill_8 FILLER_43_912 ();
 sg13g2_fill_8 FILLER_43_920 ();
 sg13g2_fill_8 FILLER_43_928 ();
 sg13g2_fill_8 FILLER_43_936 ();
 sg13g2_fill_8 FILLER_43_944 ();
 sg13g2_fill_8 FILLER_43_952 ();
 sg13g2_fill_8 FILLER_43_960 ();
 sg13g2_fill_8 FILLER_43_968 ();
 sg13g2_fill_8 FILLER_43_976 ();
 sg13g2_fill_8 FILLER_43_984 ();
 sg13g2_fill_8 FILLER_43_992 ();
 sg13g2_fill_8 FILLER_43_1000 ();
 sg13g2_fill_8 FILLER_43_1008 ();
 sg13g2_fill_8 FILLER_43_1016 ();
 sg13g2_fill_8 FILLER_43_1024 ();
 sg13g2_fill_8 FILLER_43_1032 ();
 sg13g2_fill_8 FILLER_43_1040 ();
 sg13g2_fill_8 FILLER_43_1048 ();
 sg13g2_fill_8 FILLER_43_1056 ();
 sg13g2_fill_8 FILLER_43_1064 ();
 sg13g2_fill_8 FILLER_43_1072 ();
 sg13g2_fill_8 FILLER_43_1080 ();
 sg13g2_fill_8 FILLER_43_1088 ();
 sg13g2_fill_8 FILLER_43_1096 ();
 sg13g2_fill_8 FILLER_43_1104 ();
 sg13g2_fill_8 FILLER_43_1112 ();
 sg13g2_fill_8 FILLER_43_1120 ();
 sg13g2_fill_8 FILLER_43_1128 ();
 sg13g2_fill_8 FILLER_43_1136 ();
 sg13g2_fill_8 FILLER_44_0 ();
 sg13g2_fill_8 FILLER_44_8 ();
 sg13g2_fill_8 FILLER_44_16 ();
 sg13g2_fill_8 FILLER_44_24 ();
 sg13g2_fill_8 FILLER_44_32 ();
 sg13g2_fill_8 FILLER_44_40 ();
 sg13g2_fill_8 FILLER_44_48 ();
 sg13g2_fill_8 FILLER_44_56 ();
 sg13g2_fill_8 FILLER_44_64 ();
 sg13g2_fill_8 FILLER_44_72 ();
 sg13g2_fill_8 FILLER_44_80 ();
 sg13g2_fill_8 FILLER_44_88 ();
 sg13g2_fill_8 FILLER_44_96 ();
 sg13g2_fill_8 FILLER_44_104 ();
 sg13g2_fill_8 FILLER_44_112 ();
 sg13g2_fill_8 FILLER_44_120 ();
 sg13g2_fill_8 FILLER_44_128 ();
 sg13g2_fill_8 FILLER_44_136 ();
 sg13g2_fill_8 FILLER_44_144 ();
 sg13g2_fill_8 FILLER_44_152 ();
 sg13g2_fill_8 FILLER_44_160 ();
 sg13g2_fill_8 FILLER_44_168 ();
 sg13g2_fill_8 FILLER_44_176 ();
 sg13g2_fill_8 FILLER_44_184 ();
 sg13g2_fill_8 FILLER_44_192 ();
 sg13g2_fill_8 FILLER_44_200 ();
 sg13g2_fill_8 FILLER_44_208 ();
 sg13g2_fill_8 FILLER_44_216 ();
 sg13g2_fill_8 FILLER_44_224 ();
 sg13g2_fill_8 FILLER_44_232 ();
 sg13g2_fill_8 FILLER_44_240 ();
 sg13g2_fill_8 FILLER_44_248 ();
 sg13g2_fill_8 FILLER_44_256 ();
 sg13g2_fill_8 FILLER_44_264 ();
 sg13g2_fill_8 FILLER_44_272 ();
 sg13g2_fill_8 FILLER_44_280 ();
 sg13g2_fill_8 FILLER_44_288 ();
 sg13g2_fill_8 FILLER_44_296 ();
 sg13g2_fill_8 FILLER_44_304 ();
 sg13g2_fill_8 FILLER_44_312 ();
 sg13g2_fill_8 FILLER_44_320 ();
 sg13g2_fill_8 FILLER_44_328 ();
 sg13g2_fill_8 FILLER_44_336 ();
 sg13g2_fill_8 FILLER_44_344 ();
 sg13g2_fill_8 FILLER_44_352 ();
 sg13g2_fill_8 FILLER_44_360 ();
 sg13g2_fill_8 FILLER_44_368 ();
 sg13g2_fill_8 FILLER_44_376 ();
 sg13g2_fill_8 FILLER_44_384 ();
 sg13g2_fill_8 FILLER_44_392 ();
 sg13g2_fill_8 FILLER_44_400 ();
 sg13g2_fill_8 FILLER_44_408 ();
 sg13g2_fill_8 FILLER_44_416 ();
 sg13g2_fill_8 FILLER_44_424 ();
 sg13g2_fill_8 FILLER_44_432 ();
 sg13g2_fill_8 FILLER_44_440 ();
 sg13g2_fill_8 FILLER_44_448 ();
 sg13g2_fill_8 FILLER_44_456 ();
 sg13g2_fill_8 FILLER_44_464 ();
 sg13g2_fill_8 FILLER_44_472 ();
 sg13g2_fill_8 FILLER_44_480 ();
 sg13g2_fill_8 FILLER_44_488 ();
 sg13g2_fill_8 FILLER_44_496 ();
 sg13g2_fill_8 FILLER_44_504 ();
 sg13g2_fill_8 FILLER_44_512 ();
 sg13g2_fill_8 FILLER_44_520 ();
 sg13g2_fill_8 FILLER_44_528 ();
 sg13g2_fill_8 FILLER_44_536 ();
 sg13g2_fill_8 FILLER_44_544 ();
 sg13g2_fill_8 FILLER_44_552 ();
 sg13g2_fill_8 FILLER_44_560 ();
 sg13g2_fill_8 FILLER_44_568 ();
 sg13g2_fill_8 FILLER_44_576 ();
 sg13g2_fill_8 FILLER_44_584 ();
 sg13g2_fill_8 FILLER_44_592 ();
 sg13g2_fill_8 FILLER_44_600 ();
 sg13g2_fill_8 FILLER_44_608 ();
 sg13g2_fill_8 FILLER_44_616 ();
 sg13g2_fill_8 FILLER_44_624 ();
 sg13g2_fill_8 FILLER_44_632 ();
 sg13g2_fill_8 FILLER_44_640 ();
 sg13g2_fill_8 FILLER_44_648 ();
 sg13g2_fill_8 FILLER_44_656 ();
 sg13g2_fill_8 FILLER_44_664 ();
 sg13g2_fill_8 FILLER_44_672 ();
 sg13g2_fill_8 FILLER_44_680 ();
 sg13g2_fill_8 FILLER_44_688 ();
 sg13g2_fill_8 FILLER_44_696 ();
 sg13g2_fill_8 FILLER_44_704 ();
 sg13g2_fill_8 FILLER_44_712 ();
 sg13g2_fill_8 FILLER_44_720 ();
 sg13g2_fill_8 FILLER_44_728 ();
 sg13g2_fill_8 FILLER_44_736 ();
 sg13g2_fill_8 FILLER_44_744 ();
 sg13g2_fill_8 FILLER_44_752 ();
 sg13g2_fill_8 FILLER_44_760 ();
 sg13g2_fill_8 FILLER_44_768 ();
 sg13g2_fill_8 FILLER_44_776 ();
 sg13g2_fill_8 FILLER_44_784 ();
 sg13g2_fill_8 FILLER_44_792 ();
 sg13g2_fill_8 FILLER_44_800 ();
 sg13g2_fill_8 FILLER_44_808 ();
 sg13g2_fill_8 FILLER_44_816 ();
 sg13g2_fill_8 FILLER_44_824 ();
 sg13g2_fill_8 FILLER_44_832 ();
 sg13g2_fill_8 FILLER_44_840 ();
 sg13g2_fill_8 FILLER_44_848 ();
 sg13g2_fill_8 FILLER_44_856 ();
 sg13g2_fill_8 FILLER_44_864 ();
 sg13g2_fill_8 FILLER_44_872 ();
 sg13g2_fill_8 FILLER_44_880 ();
 sg13g2_fill_8 FILLER_44_888 ();
 sg13g2_fill_8 FILLER_44_896 ();
 sg13g2_fill_8 FILLER_44_904 ();
 sg13g2_fill_8 FILLER_44_912 ();
 sg13g2_fill_8 FILLER_44_920 ();
 sg13g2_fill_8 FILLER_44_928 ();
 sg13g2_fill_8 FILLER_44_936 ();
 sg13g2_fill_8 FILLER_44_944 ();
 sg13g2_fill_8 FILLER_44_952 ();
 sg13g2_fill_8 FILLER_44_960 ();
 sg13g2_fill_8 FILLER_44_968 ();
 sg13g2_fill_8 FILLER_44_976 ();
 sg13g2_fill_8 FILLER_44_984 ();
 sg13g2_fill_8 FILLER_44_992 ();
 sg13g2_fill_8 FILLER_44_1000 ();
 sg13g2_fill_8 FILLER_44_1008 ();
 sg13g2_fill_8 FILLER_44_1016 ();
 sg13g2_fill_8 FILLER_44_1024 ();
 sg13g2_fill_8 FILLER_44_1032 ();
 sg13g2_fill_8 FILLER_44_1040 ();
 sg13g2_fill_8 FILLER_44_1048 ();
 sg13g2_fill_8 FILLER_44_1056 ();
 sg13g2_fill_8 FILLER_44_1064 ();
 sg13g2_fill_8 FILLER_44_1072 ();
 sg13g2_fill_8 FILLER_44_1080 ();
 sg13g2_fill_8 FILLER_44_1088 ();
 sg13g2_fill_8 FILLER_44_1096 ();
 sg13g2_fill_8 FILLER_44_1104 ();
 sg13g2_fill_8 FILLER_44_1112 ();
 sg13g2_fill_8 FILLER_44_1120 ();
 sg13g2_fill_8 FILLER_44_1128 ();
 sg13g2_fill_8 FILLER_44_1136 ();
 sg13g2_fill_8 FILLER_45_0 ();
 sg13g2_fill_8 FILLER_45_8 ();
 sg13g2_fill_8 FILLER_45_16 ();
 sg13g2_fill_8 FILLER_45_24 ();
 sg13g2_fill_8 FILLER_45_32 ();
 sg13g2_fill_8 FILLER_45_40 ();
 sg13g2_fill_8 FILLER_45_48 ();
 sg13g2_fill_8 FILLER_45_56 ();
 sg13g2_fill_8 FILLER_45_64 ();
 sg13g2_fill_8 FILLER_45_72 ();
 sg13g2_fill_8 FILLER_45_80 ();
 sg13g2_fill_8 FILLER_45_88 ();
 sg13g2_fill_8 FILLER_45_96 ();
 sg13g2_fill_8 FILLER_45_104 ();
 sg13g2_fill_8 FILLER_45_112 ();
 sg13g2_fill_8 FILLER_45_120 ();
 sg13g2_fill_8 FILLER_45_128 ();
 sg13g2_fill_8 FILLER_45_136 ();
 sg13g2_fill_8 FILLER_45_144 ();
 sg13g2_fill_8 FILLER_45_152 ();
 sg13g2_fill_8 FILLER_45_160 ();
 sg13g2_fill_8 FILLER_45_168 ();
 sg13g2_fill_8 FILLER_45_176 ();
 sg13g2_fill_8 FILLER_45_184 ();
 sg13g2_fill_8 FILLER_45_192 ();
 sg13g2_fill_8 FILLER_45_200 ();
 sg13g2_fill_8 FILLER_45_208 ();
 sg13g2_fill_8 FILLER_45_216 ();
 sg13g2_fill_8 FILLER_45_224 ();
 sg13g2_fill_8 FILLER_45_232 ();
 sg13g2_fill_8 FILLER_45_240 ();
 sg13g2_fill_8 FILLER_45_248 ();
 sg13g2_fill_8 FILLER_45_256 ();
 sg13g2_fill_8 FILLER_45_264 ();
 sg13g2_fill_8 FILLER_45_272 ();
 sg13g2_fill_8 FILLER_45_280 ();
 sg13g2_fill_8 FILLER_45_288 ();
 sg13g2_fill_8 FILLER_45_296 ();
 sg13g2_fill_8 FILLER_45_304 ();
 sg13g2_fill_8 FILLER_45_312 ();
 sg13g2_fill_8 FILLER_45_320 ();
 sg13g2_fill_8 FILLER_45_328 ();
 sg13g2_fill_8 FILLER_45_336 ();
 sg13g2_fill_8 FILLER_45_344 ();
 sg13g2_fill_8 FILLER_45_352 ();
 sg13g2_fill_8 FILLER_45_360 ();
 sg13g2_fill_8 FILLER_45_368 ();
 sg13g2_fill_8 FILLER_45_376 ();
 sg13g2_fill_8 FILLER_45_384 ();
 sg13g2_fill_8 FILLER_45_392 ();
 sg13g2_fill_8 FILLER_45_400 ();
 sg13g2_fill_8 FILLER_45_408 ();
 sg13g2_fill_8 FILLER_45_416 ();
 sg13g2_fill_8 FILLER_45_424 ();
 sg13g2_fill_8 FILLER_45_432 ();
 sg13g2_fill_8 FILLER_45_440 ();
 sg13g2_fill_8 FILLER_45_448 ();
 sg13g2_fill_8 FILLER_45_456 ();
 sg13g2_fill_8 FILLER_45_464 ();
 sg13g2_fill_4 FILLER_45_472 ();
 sg13g2_fill_2 FILLER_45_476 ();
 sg13g2_fill_4 FILLER_45_510 ();
 sg13g2_fill_4 FILLER_45_517 ();
 sg13g2_fill_2 FILLER_45_521 ();
 sg13g2_fill_1 FILLER_45_523 ();
 sg13g2_fill_8 FILLER_45_553 ();
 sg13g2_fill_8 FILLER_45_561 ();
 sg13g2_fill_8 FILLER_45_569 ();
 sg13g2_fill_8 FILLER_45_577 ();
 sg13g2_fill_8 FILLER_45_585 ();
 sg13g2_fill_8 FILLER_45_593 ();
 sg13g2_fill_8 FILLER_45_601 ();
 sg13g2_fill_8 FILLER_45_609 ();
 sg13g2_fill_8 FILLER_45_617 ();
 sg13g2_fill_8 FILLER_45_625 ();
 sg13g2_fill_8 FILLER_45_633 ();
 sg13g2_fill_8 FILLER_45_641 ();
 sg13g2_fill_8 FILLER_45_649 ();
 sg13g2_fill_8 FILLER_45_657 ();
 sg13g2_fill_8 FILLER_45_665 ();
 sg13g2_fill_8 FILLER_45_673 ();
 sg13g2_fill_8 FILLER_45_681 ();
 sg13g2_fill_8 FILLER_45_689 ();
 sg13g2_fill_8 FILLER_45_697 ();
 sg13g2_fill_8 FILLER_45_705 ();
 sg13g2_fill_8 FILLER_45_713 ();
 sg13g2_fill_8 FILLER_45_721 ();
 sg13g2_fill_8 FILLER_45_729 ();
 sg13g2_fill_8 FILLER_45_737 ();
 sg13g2_fill_8 FILLER_45_745 ();
 sg13g2_fill_8 FILLER_45_753 ();
 sg13g2_fill_8 FILLER_45_761 ();
 sg13g2_fill_8 FILLER_45_769 ();
 sg13g2_fill_8 FILLER_45_777 ();
 sg13g2_fill_8 FILLER_45_785 ();
 sg13g2_fill_8 FILLER_45_793 ();
 sg13g2_fill_8 FILLER_45_801 ();
 sg13g2_fill_8 FILLER_45_809 ();
 sg13g2_fill_8 FILLER_45_817 ();
 sg13g2_fill_8 FILLER_45_825 ();
 sg13g2_fill_8 FILLER_45_833 ();
 sg13g2_fill_8 FILLER_45_841 ();
 sg13g2_fill_8 FILLER_45_849 ();
 sg13g2_fill_8 FILLER_45_857 ();
 sg13g2_fill_8 FILLER_45_865 ();
 sg13g2_fill_8 FILLER_45_873 ();
 sg13g2_fill_8 FILLER_45_881 ();
 sg13g2_fill_8 FILLER_45_889 ();
 sg13g2_fill_8 FILLER_45_897 ();
 sg13g2_fill_8 FILLER_45_905 ();
 sg13g2_fill_8 FILLER_45_913 ();
 sg13g2_fill_8 FILLER_45_921 ();
 sg13g2_fill_8 FILLER_45_929 ();
 sg13g2_fill_8 FILLER_45_937 ();
 sg13g2_fill_8 FILLER_45_945 ();
 sg13g2_fill_8 FILLER_45_953 ();
 sg13g2_fill_8 FILLER_45_961 ();
 sg13g2_fill_8 FILLER_45_969 ();
 sg13g2_fill_8 FILLER_45_977 ();
 sg13g2_fill_8 FILLER_45_985 ();
 sg13g2_fill_8 FILLER_45_993 ();
 sg13g2_fill_8 FILLER_45_1001 ();
 sg13g2_fill_8 FILLER_45_1009 ();
 sg13g2_fill_8 FILLER_45_1017 ();
 sg13g2_fill_8 FILLER_45_1025 ();
 sg13g2_fill_8 FILLER_45_1033 ();
 sg13g2_fill_8 FILLER_45_1041 ();
 sg13g2_fill_8 FILLER_45_1049 ();
 sg13g2_fill_8 FILLER_45_1057 ();
 sg13g2_fill_8 FILLER_45_1065 ();
 sg13g2_fill_8 FILLER_45_1073 ();
 sg13g2_fill_8 FILLER_45_1081 ();
 sg13g2_fill_8 FILLER_45_1089 ();
 sg13g2_fill_8 FILLER_45_1097 ();
 sg13g2_fill_8 FILLER_45_1105 ();
 sg13g2_fill_8 FILLER_45_1113 ();
 sg13g2_fill_8 FILLER_45_1121 ();
 sg13g2_fill_8 FILLER_45_1129 ();
 sg13g2_fill_4 FILLER_45_1137 ();
 sg13g2_fill_2 FILLER_45_1141 ();
 sg13g2_fill_1 FILLER_45_1143 ();
 sg13g2_fill_8 FILLER_46_0 ();
 sg13g2_fill_8 FILLER_46_8 ();
 sg13g2_fill_8 FILLER_46_16 ();
 sg13g2_fill_8 FILLER_46_24 ();
 sg13g2_fill_8 FILLER_46_32 ();
 sg13g2_fill_8 FILLER_46_40 ();
 sg13g2_fill_8 FILLER_46_48 ();
 sg13g2_fill_8 FILLER_46_56 ();
 sg13g2_fill_8 FILLER_46_64 ();
 sg13g2_fill_8 FILLER_46_72 ();
 sg13g2_fill_8 FILLER_46_80 ();
 sg13g2_fill_8 FILLER_46_88 ();
 sg13g2_fill_8 FILLER_46_96 ();
 sg13g2_fill_8 FILLER_46_104 ();
 sg13g2_fill_8 FILLER_46_112 ();
 sg13g2_fill_8 FILLER_46_120 ();
 sg13g2_fill_8 FILLER_46_128 ();
 sg13g2_fill_8 FILLER_46_136 ();
 sg13g2_fill_8 FILLER_46_144 ();
 sg13g2_fill_8 FILLER_46_152 ();
 sg13g2_fill_8 FILLER_46_160 ();
 sg13g2_fill_8 FILLER_46_168 ();
 sg13g2_fill_8 FILLER_46_176 ();
 sg13g2_fill_8 FILLER_46_184 ();
 sg13g2_fill_8 FILLER_46_192 ();
 sg13g2_fill_8 FILLER_46_200 ();
 sg13g2_fill_8 FILLER_46_208 ();
 sg13g2_fill_8 FILLER_46_216 ();
 sg13g2_fill_8 FILLER_46_224 ();
 sg13g2_fill_8 FILLER_46_232 ();
 sg13g2_fill_8 FILLER_46_240 ();
 sg13g2_fill_8 FILLER_46_248 ();
 sg13g2_fill_8 FILLER_46_256 ();
 sg13g2_fill_8 FILLER_46_264 ();
 sg13g2_fill_8 FILLER_46_272 ();
 sg13g2_fill_8 FILLER_46_280 ();
 sg13g2_fill_8 FILLER_46_288 ();
 sg13g2_fill_8 FILLER_46_296 ();
 sg13g2_fill_8 FILLER_46_304 ();
 sg13g2_fill_8 FILLER_46_312 ();
 sg13g2_fill_8 FILLER_46_320 ();
 sg13g2_fill_2 FILLER_46_328 ();
 sg13g2_fill_8 FILLER_46_361 ();
 sg13g2_fill_8 FILLER_46_369 ();
 sg13g2_fill_8 FILLER_46_377 ();
 sg13g2_fill_8 FILLER_46_385 ();
 sg13g2_fill_8 FILLER_46_393 ();
 sg13g2_fill_8 FILLER_46_401 ();
 sg13g2_fill_8 FILLER_46_409 ();
 sg13g2_fill_8 FILLER_46_417 ();
 sg13g2_fill_8 FILLER_46_425 ();
 sg13g2_fill_8 FILLER_46_433 ();
 sg13g2_fill_8 FILLER_46_441 ();
 sg13g2_fill_8 FILLER_46_449 ();
 sg13g2_fill_8 FILLER_46_457 ();
 sg13g2_fill_8 FILLER_46_465 ();
 sg13g2_fill_4 FILLER_46_473 ();
 sg13g2_fill_2 FILLER_46_477 ();
 sg13g2_fill_4 FILLER_46_537 ();
 sg13g2_fill_8 FILLER_46_570 ();
 sg13g2_fill_8 FILLER_46_578 ();
 sg13g2_fill_8 FILLER_46_586 ();
 sg13g2_fill_8 FILLER_46_594 ();
 sg13g2_fill_8 FILLER_46_602 ();
 sg13g2_fill_8 FILLER_46_610 ();
 sg13g2_fill_8 FILLER_46_618 ();
 sg13g2_fill_8 FILLER_46_626 ();
 sg13g2_fill_8 FILLER_46_634 ();
 sg13g2_fill_8 FILLER_46_642 ();
 sg13g2_fill_8 FILLER_46_650 ();
 sg13g2_fill_8 FILLER_46_658 ();
 sg13g2_fill_8 FILLER_46_666 ();
 sg13g2_fill_8 FILLER_46_674 ();
 sg13g2_fill_8 FILLER_46_682 ();
 sg13g2_fill_8 FILLER_46_690 ();
 sg13g2_fill_8 FILLER_46_698 ();
 sg13g2_fill_8 FILLER_46_706 ();
 sg13g2_fill_8 FILLER_46_714 ();
 sg13g2_fill_8 FILLER_46_722 ();
 sg13g2_fill_8 FILLER_46_730 ();
 sg13g2_fill_8 FILLER_46_738 ();
 sg13g2_fill_8 FILLER_46_746 ();
 sg13g2_fill_8 FILLER_46_754 ();
 sg13g2_fill_8 FILLER_46_762 ();
 sg13g2_fill_8 FILLER_46_770 ();
 sg13g2_fill_8 FILLER_46_778 ();
 sg13g2_fill_8 FILLER_46_786 ();
 sg13g2_fill_8 FILLER_46_794 ();
 sg13g2_fill_8 FILLER_46_802 ();
 sg13g2_fill_8 FILLER_46_810 ();
 sg13g2_fill_8 FILLER_46_818 ();
 sg13g2_fill_8 FILLER_46_826 ();
 sg13g2_fill_8 FILLER_46_834 ();
 sg13g2_fill_8 FILLER_46_842 ();
 sg13g2_fill_8 FILLER_46_850 ();
 sg13g2_fill_8 FILLER_46_858 ();
 sg13g2_fill_8 FILLER_46_866 ();
 sg13g2_fill_8 FILLER_46_874 ();
 sg13g2_fill_8 FILLER_46_882 ();
 sg13g2_fill_8 FILLER_46_890 ();
 sg13g2_fill_8 FILLER_46_898 ();
 sg13g2_fill_8 FILLER_46_906 ();
 sg13g2_fill_8 FILLER_46_914 ();
 sg13g2_fill_8 FILLER_46_922 ();
 sg13g2_fill_8 FILLER_46_930 ();
 sg13g2_fill_8 FILLER_46_938 ();
 sg13g2_fill_8 FILLER_46_946 ();
 sg13g2_fill_8 FILLER_46_954 ();
 sg13g2_fill_8 FILLER_46_962 ();
 sg13g2_fill_8 FILLER_46_970 ();
 sg13g2_fill_8 FILLER_46_978 ();
 sg13g2_fill_8 FILLER_46_986 ();
 sg13g2_fill_8 FILLER_46_994 ();
 sg13g2_fill_8 FILLER_46_1002 ();
 sg13g2_fill_8 FILLER_46_1010 ();
 sg13g2_fill_8 FILLER_46_1018 ();
 sg13g2_fill_8 FILLER_46_1026 ();
 sg13g2_fill_8 FILLER_46_1034 ();
 sg13g2_fill_8 FILLER_46_1042 ();
 sg13g2_fill_8 FILLER_46_1050 ();
 sg13g2_fill_8 FILLER_46_1058 ();
 sg13g2_fill_8 FILLER_46_1066 ();
 sg13g2_fill_8 FILLER_46_1074 ();
 sg13g2_fill_8 FILLER_46_1082 ();
 sg13g2_fill_8 FILLER_46_1090 ();
 sg13g2_fill_8 FILLER_46_1098 ();
 sg13g2_fill_8 FILLER_46_1106 ();
 sg13g2_fill_8 FILLER_46_1114 ();
 sg13g2_fill_8 FILLER_46_1122 ();
 sg13g2_fill_8 FILLER_46_1130 ();
 sg13g2_fill_4 FILLER_46_1138 ();
 sg13g2_fill_2 FILLER_46_1142 ();
 sg13g2_fill_8 FILLER_47_0 ();
 sg13g2_fill_8 FILLER_47_8 ();
 sg13g2_fill_8 FILLER_47_16 ();
 sg13g2_fill_8 FILLER_47_24 ();
 sg13g2_fill_8 FILLER_47_32 ();
 sg13g2_fill_8 FILLER_47_40 ();
 sg13g2_fill_8 FILLER_47_48 ();
 sg13g2_fill_8 FILLER_47_56 ();
 sg13g2_fill_8 FILLER_47_64 ();
 sg13g2_fill_8 FILLER_47_72 ();
 sg13g2_fill_8 FILLER_47_80 ();
 sg13g2_fill_8 FILLER_47_88 ();
 sg13g2_fill_8 FILLER_47_96 ();
 sg13g2_fill_8 FILLER_47_104 ();
 sg13g2_fill_8 FILLER_47_112 ();
 sg13g2_fill_8 FILLER_47_120 ();
 sg13g2_fill_8 FILLER_47_128 ();
 sg13g2_fill_8 FILLER_47_136 ();
 sg13g2_fill_8 FILLER_47_144 ();
 sg13g2_fill_8 FILLER_47_152 ();
 sg13g2_fill_8 FILLER_47_160 ();
 sg13g2_fill_8 FILLER_47_168 ();
 sg13g2_fill_8 FILLER_47_176 ();
 sg13g2_fill_8 FILLER_47_184 ();
 sg13g2_fill_8 FILLER_47_192 ();
 sg13g2_fill_8 FILLER_47_200 ();
 sg13g2_fill_8 FILLER_47_208 ();
 sg13g2_fill_8 FILLER_47_216 ();
 sg13g2_fill_8 FILLER_47_224 ();
 sg13g2_fill_8 FILLER_47_232 ();
 sg13g2_fill_8 FILLER_47_240 ();
 sg13g2_fill_8 FILLER_47_248 ();
 sg13g2_fill_8 FILLER_47_256 ();
 sg13g2_fill_8 FILLER_47_264 ();
 sg13g2_fill_8 FILLER_47_272 ();
 sg13g2_fill_8 FILLER_47_280 ();
 sg13g2_fill_8 FILLER_47_288 ();
 sg13g2_fill_8 FILLER_47_296 ();
 sg13g2_fill_4 FILLER_47_304 ();
 sg13g2_fill_1 FILLER_47_308 ();
 sg13g2_fill_2 FILLER_47_339 ();
 sg13g2_fill_8 FILLER_47_372 ();
 sg13g2_fill_8 FILLER_47_380 ();
 sg13g2_fill_8 FILLER_47_388 ();
 sg13g2_fill_8 FILLER_47_396 ();
 sg13g2_fill_8 FILLER_47_404 ();
 sg13g2_fill_8 FILLER_47_412 ();
 sg13g2_fill_8 FILLER_47_420 ();
 sg13g2_fill_8 FILLER_47_428 ();
 sg13g2_fill_8 FILLER_47_436 ();
 sg13g2_fill_8 FILLER_47_444 ();
 sg13g2_fill_8 FILLER_47_452 ();
 sg13g2_fill_8 FILLER_47_460 ();
 sg13g2_fill_4 FILLER_47_468 ();
 sg13g2_fill_1 FILLER_47_472 ();
 sg13g2_fill_4 FILLER_47_511 ();
 sg13g2_fill_4 FILLER_47_521 ();
 sg13g2_fill_2 FILLER_47_525 ();
 sg13g2_fill_8 FILLER_47_533 ();
 sg13g2_fill_2 FILLER_47_541 ();
 sg13g2_fill_1 FILLER_47_543 ();
 sg13g2_fill_1 FILLER_47_576 ();
 sg13g2_fill_8 FILLER_47_603 ();
 sg13g2_fill_8 FILLER_47_611 ();
 sg13g2_fill_8 FILLER_47_619 ();
 sg13g2_fill_8 FILLER_47_627 ();
 sg13g2_fill_8 FILLER_47_635 ();
 sg13g2_fill_8 FILLER_47_643 ();
 sg13g2_fill_8 FILLER_47_651 ();
 sg13g2_fill_8 FILLER_47_659 ();
 sg13g2_fill_8 FILLER_47_667 ();
 sg13g2_fill_8 FILLER_47_675 ();
 sg13g2_fill_8 FILLER_47_683 ();
 sg13g2_fill_8 FILLER_47_691 ();
 sg13g2_fill_8 FILLER_47_699 ();
 sg13g2_fill_8 FILLER_47_707 ();
 sg13g2_fill_8 FILLER_47_715 ();
 sg13g2_fill_8 FILLER_47_723 ();
 sg13g2_fill_8 FILLER_47_731 ();
 sg13g2_fill_8 FILLER_47_739 ();
 sg13g2_fill_8 FILLER_47_747 ();
 sg13g2_fill_8 FILLER_47_755 ();
 sg13g2_fill_8 FILLER_47_763 ();
 sg13g2_fill_8 FILLER_47_771 ();
 sg13g2_fill_8 FILLER_47_779 ();
 sg13g2_fill_8 FILLER_47_787 ();
 sg13g2_fill_8 FILLER_47_795 ();
 sg13g2_fill_8 FILLER_47_803 ();
 sg13g2_fill_8 FILLER_47_811 ();
 sg13g2_fill_8 FILLER_47_819 ();
 sg13g2_fill_8 FILLER_47_827 ();
 sg13g2_fill_8 FILLER_47_835 ();
 sg13g2_fill_8 FILLER_47_843 ();
 sg13g2_fill_8 FILLER_47_851 ();
 sg13g2_fill_8 FILLER_47_859 ();
 sg13g2_fill_8 FILLER_47_867 ();
 sg13g2_fill_8 FILLER_47_875 ();
 sg13g2_fill_8 FILLER_47_883 ();
 sg13g2_fill_8 FILLER_47_891 ();
 sg13g2_fill_8 FILLER_47_899 ();
 sg13g2_fill_8 FILLER_47_907 ();
 sg13g2_fill_8 FILLER_47_915 ();
 sg13g2_fill_8 FILLER_47_923 ();
 sg13g2_fill_8 FILLER_47_931 ();
 sg13g2_fill_8 FILLER_47_939 ();
 sg13g2_fill_8 FILLER_47_947 ();
 sg13g2_fill_8 FILLER_47_955 ();
 sg13g2_fill_8 FILLER_47_963 ();
 sg13g2_fill_8 FILLER_47_971 ();
 sg13g2_fill_8 FILLER_47_979 ();
 sg13g2_fill_8 FILLER_47_987 ();
 sg13g2_fill_8 FILLER_47_995 ();
 sg13g2_fill_8 FILLER_47_1003 ();
 sg13g2_fill_8 FILLER_47_1011 ();
 sg13g2_fill_8 FILLER_47_1019 ();
 sg13g2_fill_8 FILLER_47_1027 ();
 sg13g2_fill_8 FILLER_47_1035 ();
 sg13g2_fill_8 FILLER_47_1043 ();
 sg13g2_fill_8 FILLER_47_1051 ();
 sg13g2_fill_8 FILLER_47_1059 ();
 sg13g2_fill_8 FILLER_47_1067 ();
 sg13g2_fill_8 FILLER_47_1075 ();
 sg13g2_fill_8 FILLER_47_1083 ();
 sg13g2_fill_8 FILLER_47_1091 ();
 sg13g2_fill_8 FILLER_47_1099 ();
 sg13g2_fill_8 FILLER_47_1107 ();
 sg13g2_fill_8 FILLER_47_1115 ();
 sg13g2_fill_8 FILLER_47_1123 ();
 sg13g2_fill_8 FILLER_47_1131 ();
 sg13g2_fill_4 FILLER_47_1139 ();
 sg13g2_fill_1 FILLER_47_1143 ();
 sg13g2_fill_8 FILLER_48_0 ();
 sg13g2_fill_8 FILLER_48_8 ();
 sg13g2_fill_8 FILLER_48_16 ();
 sg13g2_fill_8 FILLER_48_24 ();
 sg13g2_fill_8 FILLER_48_32 ();
 sg13g2_fill_8 FILLER_48_40 ();
 sg13g2_fill_8 FILLER_48_48 ();
 sg13g2_fill_8 FILLER_48_56 ();
 sg13g2_fill_8 FILLER_48_64 ();
 sg13g2_fill_8 FILLER_48_72 ();
 sg13g2_fill_8 FILLER_48_80 ();
 sg13g2_fill_8 FILLER_48_88 ();
 sg13g2_fill_8 FILLER_48_96 ();
 sg13g2_fill_8 FILLER_48_104 ();
 sg13g2_fill_8 FILLER_48_112 ();
 sg13g2_fill_8 FILLER_48_120 ();
 sg13g2_fill_8 FILLER_48_128 ();
 sg13g2_fill_8 FILLER_48_136 ();
 sg13g2_fill_8 FILLER_48_144 ();
 sg13g2_fill_8 FILLER_48_152 ();
 sg13g2_fill_8 FILLER_48_160 ();
 sg13g2_fill_8 FILLER_48_168 ();
 sg13g2_fill_8 FILLER_48_176 ();
 sg13g2_fill_8 FILLER_48_184 ();
 sg13g2_fill_8 FILLER_48_192 ();
 sg13g2_fill_8 FILLER_48_200 ();
 sg13g2_fill_8 FILLER_48_208 ();
 sg13g2_fill_8 FILLER_48_216 ();
 sg13g2_fill_8 FILLER_48_224 ();
 sg13g2_fill_8 FILLER_48_232 ();
 sg13g2_fill_8 FILLER_48_240 ();
 sg13g2_fill_8 FILLER_48_248 ();
 sg13g2_fill_8 FILLER_48_256 ();
 sg13g2_fill_8 FILLER_48_264 ();
 sg13g2_fill_8 FILLER_48_272 ();
 sg13g2_fill_8 FILLER_48_280 ();
 sg13g2_fill_8 FILLER_48_288 ();
 sg13g2_fill_8 FILLER_48_296 ();
 sg13g2_fill_4 FILLER_48_330 ();
 sg13g2_fill_4 FILLER_48_340 ();
 sg13g2_fill_2 FILLER_48_344 ();
 sg13g2_fill_1 FILLER_48_346 ();
 sg13g2_fill_1 FILLER_48_352 ();
 sg13g2_fill_8 FILLER_48_358 ();
 sg13g2_fill_8 FILLER_48_366 ();
 sg13g2_fill_8 FILLER_48_374 ();
 sg13g2_fill_8 FILLER_48_382 ();
 sg13g2_fill_8 FILLER_48_390 ();
 sg13g2_fill_8 FILLER_48_398 ();
 sg13g2_fill_8 FILLER_48_406 ();
 sg13g2_fill_8 FILLER_48_414 ();
 sg13g2_fill_8 FILLER_48_422 ();
 sg13g2_fill_8 FILLER_48_430 ();
 sg13g2_fill_8 FILLER_48_438 ();
 sg13g2_fill_8 FILLER_48_446 ();
 sg13g2_fill_8 FILLER_48_454 ();
 sg13g2_fill_8 FILLER_48_462 ();
 sg13g2_fill_8 FILLER_48_470 ();
 sg13g2_fill_4 FILLER_48_478 ();
 sg13g2_fill_1 FILLER_48_485 ();
 sg13g2_fill_8 FILLER_48_489 ();
 sg13g2_fill_8 FILLER_48_497 ();
 sg13g2_fill_8 FILLER_48_505 ();
 sg13g2_fill_8 FILLER_48_513 ();
 sg13g2_fill_8 FILLER_48_536 ();
 sg13g2_fill_8 FILLER_48_544 ();
 sg13g2_fill_2 FILLER_48_561 ();
 sg13g2_fill_8 FILLER_48_615 ();
 sg13g2_fill_8 FILLER_48_623 ();
 sg13g2_fill_8 FILLER_48_631 ();
 sg13g2_fill_8 FILLER_48_639 ();
 sg13g2_fill_8 FILLER_48_647 ();
 sg13g2_fill_8 FILLER_48_655 ();
 sg13g2_fill_8 FILLER_48_663 ();
 sg13g2_fill_8 FILLER_48_671 ();
 sg13g2_fill_8 FILLER_48_679 ();
 sg13g2_fill_8 FILLER_48_687 ();
 sg13g2_fill_8 FILLER_48_695 ();
 sg13g2_fill_8 FILLER_48_703 ();
 sg13g2_fill_8 FILLER_48_711 ();
 sg13g2_fill_8 FILLER_48_719 ();
 sg13g2_fill_8 FILLER_48_727 ();
 sg13g2_fill_8 FILLER_48_735 ();
 sg13g2_fill_8 FILLER_48_743 ();
 sg13g2_fill_8 FILLER_48_751 ();
 sg13g2_fill_8 FILLER_48_759 ();
 sg13g2_fill_8 FILLER_48_767 ();
 sg13g2_fill_8 FILLER_48_775 ();
 sg13g2_fill_8 FILLER_48_783 ();
 sg13g2_fill_8 FILLER_48_791 ();
 sg13g2_fill_8 FILLER_48_799 ();
 sg13g2_fill_8 FILLER_48_807 ();
 sg13g2_fill_8 FILLER_48_815 ();
 sg13g2_fill_8 FILLER_48_823 ();
 sg13g2_fill_8 FILLER_48_831 ();
 sg13g2_fill_8 FILLER_48_839 ();
 sg13g2_fill_8 FILLER_48_847 ();
 sg13g2_fill_8 FILLER_48_855 ();
 sg13g2_fill_8 FILLER_48_863 ();
 sg13g2_fill_8 FILLER_48_871 ();
 sg13g2_fill_8 FILLER_48_879 ();
 sg13g2_fill_8 FILLER_48_887 ();
 sg13g2_fill_8 FILLER_48_895 ();
 sg13g2_fill_8 FILLER_48_903 ();
 sg13g2_fill_8 FILLER_48_911 ();
 sg13g2_fill_8 FILLER_48_919 ();
 sg13g2_fill_8 FILLER_48_927 ();
 sg13g2_fill_8 FILLER_48_935 ();
 sg13g2_fill_8 FILLER_48_943 ();
 sg13g2_fill_8 FILLER_48_951 ();
 sg13g2_fill_8 FILLER_48_959 ();
 sg13g2_fill_8 FILLER_48_967 ();
 sg13g2_fill_8 FILLER_48_975 ();
 sg13g2_fill_8 FILLER_48_983 ();
 sg13g2_fill_8 FILLER_48_991 ();
 sg13g2_fill_8 FILLER_48_999 ();
 sg13g2_fill_8 FILLER_48_1007 ();
 sg13g2_fill_8 FILLER_48_1015 ();
 sg13g2_fill_8 FILLER_48_1023 ();
 sg13g2_fill_8 FILLER_48_1031 ();
 sg13g2_fill_8 FILLER_48_1039 ();
 sg13g2_fill_8 FILLER_48_1047 ();
 sg13g2_fill_8 FILLER_48_1055 ();
 sg13g2_fill_8 FILLER_48_1063 ();
 sg13g2_fill_8 FILLER_48_1071 ();
 sg13g2_fill_8 FILLER_48_1079 ();
 sg13g2_fill_8 FILLER_48_1087 ();
 sg13g2_fill_8 FILLER_48_1095 ();
 sg13g2_fill_8 FILLER_48_1103 ();
 sg13g2_fill_8 FILLER_48_1111 ();
 sg13g2_fill_8 FILLER_48_1119 ();
 sg13g2_fill_8 FILLER_48_1127 ();
 sg13g2_fill_8 FILLER_48_1135 ();
 sg13g2_fill_1 FILLER_48_1143 ();
 sg13g2_fill_8 FILLER_49_0 ();
 sg13g2_fill_8 FILLER_49_8 ();
 sg13g2_fill_8 FILLER_49_16 ();
 sg13g2_fill_8 FILLER_49_24 ();
 sg13g2_fill_8 FILLER_49_32 ();
 sg13g2_fill_8 FILLER_49_40 ();
 sg13g2_fill_8 FILLER_49_48 ();
 sg13g2_fill_8 FILLER_49_56 ();
 sg13g2_fill_8 FILLER_49_64 ();
 sg13g2_fill_8 FILLER_49_72 ();
 sg13g2_fill_8 FILLER_49_80 ();
 sg13g2_fill_8 FILLER_49_88 ();
 sg13g2_fill_8 FILLER_49_96 ();
 sg13g2_fill_8 FILLER_49_104 ();
 sg13g2_fill_8 FILLER_49_112 ();
 sg13g2_fill_8 FILLER_49_120 ();
 sg13g2_fill_8 FILLER_49_128 ();
 sg13g2_fill_8 FILLER_49_136 ();
 sg13g2_fill_8 FILLER_49_144 ();
 sg13g2_fill_8 FILLER_49_152 ();
 sg13g2_fill_8 FILLER_49_160 ();
 sg13g2_fill_8 FILLER_49_168 ();
 sg13g2_fill_8 FILLER_49_176 ();
 sg13g2_fill_8 FILLER_49_184 ();
 sg13g2_fill_8 FILLER_49_192 ();
 sg13g2_fill_8 FILLER_49_200 ();
 sg13g2_fill_8 FILLER_49_208 ();
 sg13g2_fill_8 FILLER_49_216 ();
 sg13g2_fill_8 FILLER_49_224 ();
 sg13g2_fill_8 FILLER_49_232 ();
 sg13g2_fill_8 FILLER_49_240 ();
 sg13g2_fill_8 FILLER_49_248 ();
 sg13g2_fill_8 FILLER_49_256 ();
 sg13g2_fill_8 FILLER_49_264 ();
 sg13g2_fill_8 FILLER_49_272 ();
 sg13g2_fill_8 FILLER_49_280 ();
 sg13g2_fill_8 FILLER_49_288 ();
 sg13g2_fill_8 FILLER_49_296 ();
 sg13g2_fill_8 FILLER_49_304 ();
 sg13g2_fill_2 FILLER_49_312 ();
 sg13g2_fill_1 FILLER_49_322 ();
 sg13g2_fill_8 FILLER_49_335 ();
 sg13g2_fill_8 FILLER_49_343 ();
 sg13g2_fill_2 FILLER_49_356 ();
 sg13g2_fill_1 FILLER_49_358 ();
 sg13g2_fill_2 FILLER_49_365 ();
 sg13g2_fill_4 FILLER_49_393 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_fill_1 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_405 ();
 sg13g2_fill_1 FILLER_49_407 ();
 sg13g2_fill_8 FILLER_49_434 ();
 sg13g2_fill_1 FILLER_49_442 ();
 sg13g2_fill_8 FILLER_49_448 ();
 sg13g2_fill_8 FILLER_49_456 ();
 sg13g2_fill_8 FILLER_49_464 ();
 sg13g2_fill_4 FILLER_49_472 ();
 sg13g2_fill_2 FILLER_49_476 ();
 sg13g2_fill_8 FILLER_49_509 ();
 sg13g2_fill_8 FILLER_49_543 ();
 sg13g2_fill_8 FILLER_49_551 ();
 sg13g2_fill_8 FILLER_49_559 ();
 sg13g2_fill_1 FILLER_49_567 ();
 sg13g2_fill_2 FILLER_49_577 ();
 sg13g2_fill_1 FILLER_49_579 ();
 sg13g2_fill_4 FILLER_49_598 ();
 sg13g2_fill_1 FILLER_49_602 ();
 sg13g2_fill_8 FILLER_49_609 ();
 sg13g2_fill_8 FILLER_49_617 ();
 sg13g2_fill_8 FILLER_49_625 ();
 sg13g2_fill_8 FILLER_49_633 ();
 sg13g2_fill_8 FILLER_49_641 ();
 sg13g2_fill_8 FILLER_49_649 ();
 sg13g2_fill_8 FILLER_49_657 ();
 sg13g2_fill_8 FILLER_49_665 ();
 sg13g2_fill_8 FILLER_49_673 ();
 sg13g2_fill_8 FILLER_49_681 ();
 sg13g2_fill_8 FILLER_49_689 ();
 sg13g2_fill_8 FILLER_49_697 ();
 sg13g2_fill_8 FILLER_49_705 ();
 sg13g2_fill_8 FILLER_49_713 ();
 sg13g2_fill_8 FILLER_49_721 ();
 sg13g2_fill_8 FILLER_49_729 ();
 sg13g2_fill_8 FILLER_49_737 ();
 sg13g2_fill_8 FILLER_49_745 ();
 sg13g2_fill_8 FILLER_49_753 ();
 sg13g2_fill_8 FILLER_49_761 ();
 sg13g2_fill_8 FILLER_49_769 ();
 sg13g2_fill_8 FILLER_49_777 ();
 sg13g2_fill_8 FILLER_49_785 ();
 sg13g2_fill_8 FILLER_49_793 ();
 sg13g2_fill_8 FILLER_49_801 ();
 sg13g2_fill_8 FILLER_49_809 ();
 sg13g2_fill_8 FILLER_49_817 ();
 sg13g2_fill_8 FILLER_49_825 ();
 sg13g2_fill_8 FILLER_49_833 ();
 sg13g2_fill_8 FILLER_49_841 ();
 sg13g2_fill_8 FILLER_49_849 ();
 sg13g2_fill_8 FILLER_49_857 ();
 sg13g2_fill_8 FILLER_49_865 ();
 sg13g2_fill_8 FILLER_49_873 ();
 sg13g2_fill_8 FILLER_49_881 ();
 sg13g2_fill_8 FILLER_49_889 ();
 sg13g2_fill_8 FILLER_49_897 ();
 sg13g2_fill_8 FILLER_49_905 ();
 sg13g2_fill_8 FILLER_49_913 ();
 sg13g2_fill_8 FILLER_49_921 ();
 sg13g2_fill_8 FILLER_49_929 ();
 sg13g2_fill_8 FILLER_49_937 ();
 sg13g2_fill_8 FILLER_49_945 ();
 sg13g2_fill_8 FILLER_49_953 ();
 sg13g2_fill_8 FILLER_49_961 ();
 sg13g2_fill_8 FILLER_49_969 ();
 sg13g2_fill_8 FILLER_49_977 ();
 sg13g2_fill_8 FILLER_49_985 ();
 sg13g2_fill_8 FILLER_49_993 ();
 sg13g2_fill_8 FILLER_49_1001 ();
 sg13g2_fill_8 FILLER_49_1009 ();
 sg13g2_fill_8 FILLER_49_1017 ();
 sg13g2_fill_8 FILLER_49_1025 ();
 sg13g2_fill_8 FILLER_49_1033 ();
 sg13g2_fill_8 FILLER_49_1041 ();
 sg13g2_fill_8 FILLER_49_1049 ();
 sg13g2_fill_8 FILLER_49_1057 ();
 sg13g2_fill_8 FILLER_49_1065 ();
 sg13g2_fill_8 FILLER_49_1073 ();
 sg13g2_fill_8 FILLER_49_1081 ();
 sg13g2_fill_8 FILLER_49_1089 ();
 sg13g2_fill_8 FILLER_49_1097 ();
 sg13g2_fill_8 FILLER_49_1105 ();
 sg13g2_fill_8 FILLER_49_1113 ();
 sg13g2_fill_8 FILLER_49_1121 ();
 sg13g2_fill_8 FILLER_49_1129 ();
 sg13g2_fill_4 FILLER_49_1137 ();
 sg13g2_fill_2 FILLER_49_1141 ();
 sg13g2_fill_1 FILLER_49_1143 ();
 sg13g2_fill_8 FILLER_50_0 ();
 sg13g2_fill_8 FILLER_50_8 ();
 sg13g2_fill_8 FILLER_50_16 ();
 sg13g2_fill_8 FILLER_50_24 ();
 sg13g2_fill_8 FILLER_50_32 ();
 sg13g2_fill_8 FILLER_50_40 ();
 sg13g2_fill_8 FILLER_50_48 ();
 sg13g2_fill_8 FILLER_50_56 ();
 sg13g2_fill_8 FILLER_50_64 ();
 sg13g2_fill_8 FILLER_50_72 ();
 sg13g2_fill_8 FILLER_50_80 ();
 sg13g2_fill_8 FILLER_50_88 ();
 sg13g2_fill_8 FILLER_50_96 ();
 sg13g2_fill_8 FILLER_50_104 ();
 sg13g2_fill_8 FILLER_50_112 ();
 sg13g2_fill_8 FILLER_50_120 ();
 sg13g2_fill_8 FILLER_50_128 ();
 sg13g2_fill_8 FILLER_50_136 ();
 sg13g2_fill_8 FILLER_50_144 ();
 sg13g2_fill_8 FILLER_50_152 ();
 sg13g2_fill_8 FILLER_50_160 ();
 sg13g2_fill_8 FILLER_50_168 ();
 sg13g2_fill_8 FILLER_50_176 ();
 sg13g2_fill_8 FILLER_50_184 ();
 sg13g2_fill_8 FILLER_50_192 ();
 sg13g2_fill_8 FILLER_50_200 ();
 sg13g2_fill_8 FILLER_50_208 ();
 sg13g2_fill_8 FILLER_50_216 ();
 sg13g2_fill_8 FILLER_50_224 ();
 sg13g2_fill_8 FILLER_50_232 ();
 sg13g2_fill_8 FILLER_50_240 ();
 sg13g2_fill_8 FILLER_50_248 ();
 sg13g2_fill_8 FILLER_50_256 ();
 sg13g2_fill_8 FILLER_50_264 ();
 sg13g2_fill_8 FILLER_50_272 ();
 sg13g2_fill_8 FILLER_50_280 ();
 sg13g2_fill_8 FILLER_50_288 ();
 sg13g2_fill_8 FILLER_50_296 ();
 sg13g2_fill_1 FILLER_50_304 ();
 sg13g2_fill_8 FILLER_50_331 ();
 sg13g2_fill_4 FILLER_50_339 ();
 sg13g2_fill_1 FILLER_50_343 ();
 sg13g2_fill_2 FILLER_50_375 ();
 sg13g2_fill_1 FILLER_50_413 ();
 sg13g2_fill_2 FILLER_50_440 ();
 sg13g2_fill_1 FILLER_50_442 ();
 sg13g2_fill_8 FILLER_50_469 ();
 sg13g2_fill_2 FILLER_50_477 ();
 sg13g2_fill_2 FILLER_50_516 ();
 sg13g2_fill_8 FILLER_50_544 ();
 sg13g2_fill_2 FILLER_50_552 ();
 sg13g2_fill_1 FILLER_50_554 ();
 sg13g2_fill_8 FILLER_50_571 ();
 sg13g2_fill_2 FILLER_50_579 ();
 sg13g2_fill_1 FILLER_50_581 ();
 sg13g2_fill_8 FILLER_50_614 ();
 sg13g2_fill_8 FILLER_50_622 ();
 sg13g2_fill_8 FILLER_50_630 ();
 sg13g2_fill_8 FILLER_50_638 ();
 sg13g2_fill_8 FILLER_50_646 ();
 sg13g2_fill_8 FILLER_50_654 ();
 sg13g2_fill_8 FILLER_50_662 ();
 sg13g2_fill_8 FILLER_50_670 ();
 sg13g2_fill_8 FILLER_50_678 ();
 sg13g2_fill_8 FILLER_50_686 ();
 sg13g2_fill_8 FILLER_50_694 ();
 sg13g2_fill_8 FILLER_50_702 ();
 sg13g2_fill_8 FILLER_50_710 ();
 sg13g2_fill_8 FILLER_50_718 ();
 sg13g2_fill_8 FILLER_50_726 ();
 sg13g2_fill_8 FILLER_50_734 ();
 sg13g2_fill_8 FILLER_50_742 ();
 sg13g2_fill_8 FILLER_50_750 ();
 sg13g2_fill_8 FILLER_50_758 ();
 sg13g2_fill_8 FILLER_50_766 ();
 sg13g2_fill_8 FILLER_50_774 ();
 sg13g2_fill_8 FILLER_50_782 ();
 sg13g2_fill_8 FILLER_50_790 ();
 sg13g2_fill_8 FILLER_50_798 ();
 sg13g2_fill_8 FILLER_50_806 ();
 sg13g2_fill_8 FILLER_50_814 ();
 sg13g2_fill_8 FILLER_50_822 ();
 sg13g2_fill_8 FILLER_50_830 ();
 sg13g2_fill_8 FILLER_50_838 ();
 sg13g2_fill_8 FILLER_50_846 ();
 sg13g2_fill_8 FILLER_50_854 ();
 sg13g2_fill_8 FILLER_50_862 ();
 sg13g2_fill_8 FILLER_50_870 ();
 sg13g2_fill_8 FILLER_50_878 ();
 sg13g2_fill_8 FILLER_50_886 ();
 sg13g2_fill_8 FILLER_50_894 ();
 sg13g2_fill_8 FILLER_50_902 ();
 sg13g2_fill_8 FILLER_50_910 ();
 sg13g2_fill_8 FILLER_50_918 ();
 sg13g2_fill_8 FILLER_50_926 ();
 sg13g2_fill_8 FILLER_50_934 ();
 sg13g2_fill_8 FILLER_50_942 ();
 sg13g2_fill_8 FILLER_50_950 ();
 sg13g2_fill_8 FILLER_50_958 ();
 sg13g2_fill_8 FILLER_50_966 ();
 sg13g2_fill_8 FILLER_50_974 ();
 sg13g2_fill_8 FILLER_50_982 ();
 sg13g2_fill_8 FILLER_50_990 ();
 sg13g2_fill_8 FILLER_50_998 ();
 sg13g2_fill_8 FILLER_50_1006 ();
 sg13g2_fill_8 FILLER_50_1014 ();
 sg13g2_fill_8 FILLER_50_1022 ();
 sg13g2_fill_8 FILLER_50_1030 ();
 sg13g2_fill_8 FILLER_50_1038 ();
 sg13g2_fill_8 FILLER_50_1046 ();
 sg13g2_fill_8 FILLER_50_1054 ();
 sg13g2_fill_8 FILLER_50_1062 ();
 sg13g2_fill_8 FILLER_50_1070 ();
 sg13g2_fill_8 FILLER_50_1078 ();
 sg13g2_fill_8 FILLER_50_1086 ();
 sg13g2_fill_8 FILLER_50_1094 ();
 sg13g2_fill_8 FILLER_50_1102 ();
 sg13g2_fill_8 FILLER_50_1110 ();
 sg13g2_fill_8 FILLER_50_1118 ();
 sg13g2_fill_8 FILLER_50_1126 ();
 sg13g2_fill_8 FILLER_50_1134 ();
 sg13g2_fill_2 FILLER_50_1142 ();
 sg13g2_fill_8 FILLER_51_0 ();
 sg13g2_fill_8 FILLER_51_8 ();
 sg13g2_fill_8 FILLER_51_16 ();
 sg13g2_fill_8 FILLER_51_24 ();
 sg13g2_fill_8 FILLER_51_32 ();
 sg13g2_fill_8 FILLER_51_40 ();
 sg13g2_fill_8 FILLER_51_48 ();
 sg13g2_fill_8 FILLER_51_56 ();
 sg13g2_fill_8 FILLER_51_64 ();
 sg13g2_fill_8 FILLER_51_72 ();
 sg13g2_fill_8 FILLER_51_80 ();
 sg13g2_fill_8 FILLER_51_88 ();
 sg13g2_fill_8 FILLER_51_96 ();
 sg13g2_fill_8 FILLER_51_104 ();
 sg13g2_fill_8 FILLER_51_112 ();
 sg13g2_fill_8 FILLER_51_120 ();
 sg13g2_fill_8 FILLER_51_128 ();
 sg13g2_fill_8 FILLER_51_136 ();
 sg13g2_fill_8 FILLER_51_144 ();
 sg13g2_fill_8 FILLER_51_152 ();
 sg13g2_fill_8 FILLER_51_160 ();
 sg13g2_fill_8 FILLER_51_168 ();
 sg13g2_fill_8 FILLER_51_176 ();
 sg13g2_fill_8 FILLER_51_184 ();
 sg13g2_fill_8 FILLER_51_192 ();
 sg13g2_fill_8 FILLER_51_200 ();
 sg13g2_fill_8 FILLER_51_208 ();
 sg13g2_fill_8 FILLER_51_216 ();
 sg13g2_fill_8 FILLER_51_224 ();
 sg13g2_fill_8 FILLER_51_232 ();
 sg13g2_fill_8 FILLER_51_240 ();
 sg13g2_fill_8 FILLER_51_248 ();
 sg13g2_fill_8 FILLER_51_256 ();
 sg13g2_fill_8 FILLER_51_264 ();
 sg13g2_fill_8 FILLER_51_272 ();
 sg13g2_fill_8 FILLER_51_280 ();
 sg13g2_fill_8 FILLER_51_288 ();
 sg13g2_fill_8 FILLER_51_296 ();
 sg13g2_fill_8 FILLER_51_340 ();
 sg13g2_fill_8 FILLER_51_348 ();
 sg13g2_fill_8 FILLER_51_370 ();
 sg13g2_fill_4 FILLER_51_378 ();
 sg13g2_fill_2 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_384 ();
 sg13g2_fill_4 FILLER_51_398 ();
 sg13g2_fill_2 FILLER_51_402 ();
 sg13g2_fill_1 FILLER_51_404 ();
 sg13g2_fill_4 FILLER_51_410 ();
 sg13g2_fill_2 FILLER_51_414 ();
 sg13g2_fill_2 FILLER_51_431 ();
 sg13g2_fill_4 FILLER_51_482 ();
 sg13g2_fill_1 FILLER_51_486 ();
 sg13g2_fill_8 FILLER_51_490 ();
 sg13g2_fill_8 FILLER_51_504 ();
 sg13g2_fill_4 FILLER_51_512 ();
 sg13g2_fill_1 FILLER_51_516 ();
 sg13g2_fill_1 FILLER_51_520 ();
 sg13g2_fill_8 FILLER_51_530 ();
 sg13g2_fill_8 FILLER_51_538 ();
 sg13g2_fill_2 FILLER_51_546 ();
 sg13g2_fill_1 FILLER_51_548 ();
 sg13g2_fill_8 FILLER_51_575 ();
 sg13g2_fill_4 FILLER_51_583 ();
 sg13g2_fill_1 FILLER_51_587 ();
 sg13g2_fill_8 FILLER_51_597 ();
 sg13g2_fill_8 FILLER_51_605 ();
 sg13g2_fill_8 FILLER_51_613 ();
 sg13g2_fill_8 FILLER_51_621 ();
 sg13g2_fill_8 FILLER_51_629 ();
 sg13g2_fill_8 FILLER_51_637 ();
 sg13g2_fill_8 FILLER_51_645 ();
 sg13g2_fill_8 FILLER_51_653 ();
 sg13g2_fill_8 FILLER_51_661 ();
 sg13g2_fill_8 FILLER_51_669 ();
 sg13g2_fill_8 FILLER_51_677 ();
 sg13g2_fill_8 FILLER_51_685 ();
 sg13g2_fill_8 FILLER_51_693 ();
 sg13g2_fill_8 FILLER_51_701 ();
 sg13g2_fill_8 FILLER_51_709 ();
 sg13g2_fill_8 FILLER_51_717 ();
 sg13g2_fill_8 FILLER_51_725 ();
 sg13g2_fill_8 FILLER_51_733 ();
 sg13g2_fill_8 FILLER_51_741 ();
 sg13g2_fill_8 FILLER_51_749 ();
 sg13g2_fill_8 FILLER_51_757 ();
 sg13g2_fill_8 FILLER_51_765 ();
 sg13g2_fill_8 FILLER_51_773 ();
 sg13g2_fill_8 FILLER_51_781 ();
 sg13g2_fill_8 FILLER_51_789 ();
 sg13g2_fill_8 FILLER_51_797 ();
 sg13g2_fill_8 FILLER_51_805 ();
 sg13g2_fill_8 FILLER_51_813 ();
 sg13g2_fill_8 FILLER_51_821 ();
 sg13g2_fill_8 FILLER_51_829 ();
 sg13g2_fill_8 FILLER_51_837 ();
 sg13g2_fill_8 FILLER_51_845 ();
 sg13g2_fill_8 FILLER_51_853 ();
 sg13g2_fill_8 FILLER_51_861 ();
 sg13g2_fill_8 FILLER_51_869 ();
 sg13g2_fill_8 FILLER_51_877 ();
 sg13g2_fill_8 FILLER_51_885 ();
 sg13g2_fill_8 FILLER_51_893 ();
 sg13g2_fill_8 FILLER_51_901 ();
 sg13g2_fill_8 FILLER_51_909 ();
 sg13g2_fill_8 FILLER_51_917 ();
 sg13g2_fill_8 FILLER_51_925 ();
 sg13g2_fill_8 FILLER_51_933 ();
 sg13g2_fill_8 FILLER_51_941 ();
 sg13g2_fill_8 FILLER_51_949 ();
 sg13g2_fill_8 FILLER_51_957 ();
 sg13g2_fill_8 FILLER_51_965 ();
 sg13g2_fill_8 FILLER_51_973 ();
 sg13g2_fill_8 FILLER_51_981 ();
 sg13g2_fill_8 FILLER_51_989 ();
 sg13g2_fill_8 FILLER_51_997 ();
 sg13g2_fill_8 FILLER_51_1005 ();
 sg13g2_fill_8 FILLER_51_1013 ();
 sg13g2_fill_8 FILLER_51_1021 ();
 sg13g2_fill_8 FILLER_51_1029 ();
 sg13g2_fill_8 FILLER_51_1037 ();
 sg13g2_fill_8 FILLER_51_1045 ();
 sg13g2_fill_8 FILLER_51_1053 ();
 sg13g2_fill_8 FILLER_51_1061 ();
 sg13g2_fill_8 FILLER_51_1069 ();
 sg13g2_fill_8 FILLER_51_1077 ();
 sg13g2_fill_8 FILLER_51_1085 ();
 sg13g2_fill_8 FILLER_51_1093 ();
 sg13g2_fill_8 FILLER_51_1101 ();
 sg13g2_fill_8 FILLER_51_1109 ();
 sg13g2_fill_8 FILLER_51_1117 ();
 sg13g2_fill_8 FILLER_51_1125 ();
 sg13g2_fill_8 FILLER_51_1133 ();
 sg13g2_fill_2 FILLER_51_1141 ();
 sg13g2_fill_1 FILLER_51_1143 ();
 sg13g2_fill_8 FILLER_52_0 ();
 sg13g2_fill_8 FILLER_52_8 ();
 sg13g2_fill_8 FILLER_52_16 ();
 sg13g2_fill_8 FILLER_52_24 ();
 sg13g2_fill_8 FILLER_52_32 ();
 sg13g2_fill_8 FILLER_52_40 ();
 sg13g2_fill_8 FILLER_52_48 ();
 sg13g2_fill_8 FILLER_52_56 ();
 sg13g2_fill_8 FILLER_52_64 ();
 sg13g2_fill_8 FILLER_52_72 ();
 sg13g2_fill_8 FILLER_52_80 ();
 sg13g2_fill_8 FILLER_52_88 ();
 sg13g2_fill_8 FILLER_52_96 ();
 sg13g2_fill_8 FILLER_52_104 ();
 sg13g2_fill_8 FILLER_52_112 ();
 sg13g2_fill_8 FILLER_52_120 ();
 sg13g2_fill_8 FILLER_52_128 ();
 sg13g2_fill_8 FILLER_52_136 ();
 sg13g2_fill_8 FILLER_52_144 ();
 sg13g2_fill_8 FILLER_52_152 ();
 sg13g2_fill_8 FILLER_52_160 ();
 sg13g2_fill_8 FILLER_52_168 ();
 sg13g2_fill_8 FILLER_52_176 ();
 sg13g2_fill_8 FILLER_52_184 ();
 sg13g2_fill_8 FILLER_52_192 ();
 sg13g2_fill_8 FILLER_52_200 ();
 sg13g2_fill_8 FILLER_52_208 ();
 sg13g2_fill_8 FILLER_52_216 ();
 sg13g2_fill_8 FILLER_52_224 ();
 sg13g2_fill_8 FILLER_52_232 ();
 sg13g2_fill_8 FILLER_52_240 ();
 sg13g2_fill_8 FILLER_52_248 ();
 sg13g2_fill_8 FILLER_52_256 ();
 sg13g2_fill_8 FILLER_52_264 ();
 sg13g2_fill_8 FILLER_52_272 ();
 sg13g2_fill_8 FILLER_52_280 ();
 sg13g2_fill_8 FILLER_52_288 ();
 sg13g2_fill_8 FILLER_52_296 ();
 sg13g2_fill_8 FILLER_52_304 ();
 sg13g2_fill_2 FILLER_52_312 ();
 sg13g2_fill_2 FILLER_52_322 ();
 sg13g2_fill_8 FILLER_52_330 ();
 sg13g2_fill_2 FILLER_52_338 ();
 sg13g2_fill_8 FILLER_52_348 ();
 sg13g2_fill_2 FILLER_52_356 ();
 sg13g2_fill_1 FILLER_52_358 ();
 sg13g2_fill_8 FILLER_52_368 ();
 sg13g2_fill_8 FILLER_52_376 ();
 sg13g2_fill_8 FILLER_52_384 ();
 sg13g2_fill_8 FILLER_52_392 ();
 sg13g2_fill_8 FILLER_52_400 ();
 sg13g2_fill_8 FILLER_52_408 ();
 sg13g2_fill_8 FILLER_52_416 ();
 sg13g2_fill_8 FILLER_52_424 ();
 sg13g2_fill_8 FILLER_52_432 ();
 sg13g2_fill_4 FILLER_52_440 ();
 sg13g2_fill_1 FILLER_52_444 ();
 sg13g2_fill_8 FILLER_52_459 ();
 sg13g2_fill_8 FILLER_52_467 ();
 sg13g2_fill_4 FILLER_52_475 ();
 sg13g2_fill_4 FILLER_52_505 ();
 sg13g2_fill_2 FILLER_52_509 ();
 sg13g2_fill_1 FILLER_52_511 ();
 sg13g2_fill_4 FILLER_52_538 ();
 sg13g2_fill_2 FILLER_52_542 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_fill_1 FILLER_52_554 ();
 sg13g2_fill_1 FILLER_52_558 ();
 sg13g2_fill_8 FILLER_52_576 ();
 sg13g2_fill_2 FILLER_52_584 ();
 sg13g2_fill_8 FILLER_52_612 ();
 sg13g2_fill_8 FILLER_52_620 ();
 sg13g2_fill_8 FILLER_52_628 ();
 sg13g2_fill_8 FILLER_52_636 ();
 sg13g2_fill_8 FILLER_52_644 ();
 sg13g2_fill_8 FILLER_52_652 ();
 sg13g2_fill_8 FILLER_52_660 ();
 sg13g2_fill_8 FILLER_52_668 ();
 sg13g2_fill_8 FILLER_52_676 ();
 sg13g2_fill_8 FILLER_52_684 ();
 sg13g2_fill_8 FILLER_52_692 ();
 sg13g2_fill_8 FILLER_52_700 ();
 sg13g2_fill_8 FILLER_52_708 ();
 sg13g2_fill_8 FILLER_52_716 ();
 sg13g2_fill_8 FILLER_52_724 ();
 sg13g2_fill_8 FILLER_52_732 ();
 sg13g2_fill_8 FILLER_52_740 ();
 sg13g2_fill_8 FILLER_52_748 ();
 sg13g2_fill_8 FILLER_52_756 ();
 sg13g2_fill_8 FILLER_52_764 ();
 sg13g2_fill_8 FILLER_52_772 ();
 sg13g2_fill_8 FILLER_52_780 ();
 sg13g2_fill_8 FILLER_52_788 ();
 sg13g2_fill_8 FILLER_52_796 ();
 sg13g2_fill_8 FILLER_52_804 ();
 sg13g2_fill_8 FILLER_52_812 ();
 sg13g2_fill_8 FILLER_52_820 ();
 sg13g2_fill_8 FILLER_52_828 ();
 sg13g2_fill_8 FILLER_52_836 ();
 sg13g2_fill_8 FILLER_52_844 ();
 sg13g2_fill_8 FILLER_52_852 ();
 sg13g2_fill_8 FILLER_52_860 ();
 sg13g2_fill_8 FILLER_52_868 ();
 sg13g2_fill_8 FILLER_52_876 ();
 sg13g2_fill_8 FILLER_52_884 ();
 sg13g2_fill_8 FILLER_52_892 ();
 sg13g2_fill_8 FILLER_52_900 ();
 sg13g2_fill_8 FILLER_52_908 ();
 sg13g2_fill_8 FILLER_52_916 ();
 sg13g2_fill_8 FILLER_52_924 ();
 sg13g2_fill_8 FILLER_52_932 ();
 sg13g2_fill_8 FILLER_52_940 ();
 sg13g2_fill_8 FILLER_52_948 ();
 sg13g2_fill_8 FILLER_52_956 ();
 sg13g2_fill_8 FILLER_52_964 ();
 sg13g2_fill_8 FILLER_52_972 ();
 sg13g2_fill_8 FILLER_52_980 ();
 sg13g2_fill_8 FILLER_52_988 ();
 sg13g2_fill_8 FILLER_52_996 ();
 sg13g2_fill_8 FILLER_52_1004 ();
 sg13g2_fill_8 FILLER_52_1012 ();
 sg13g2_fill_8 FILLER_52_1020 ();
 sg13g2_fill_8 FILLER_52_1028 ();
 sg13g2_fill_8 FILLER_52_1036 ();
 sg13g2_fill_8 FILLER_52_1044 ();
 sg13g2_fill_8 FILLER_52_1052 ();
 sg13g2_fill_8 FILLER_52_1060 ();
 sg13g2_fill_8 FILLER_52_1068 ();
 sg13g2_fill_8 FILLER_52_1076 ();
 sg13g2_fill_8 FILLER_52_1084 ();
 sg13g2_fill_8 FILLER_52_1092 ();
 sg13g2_fill_8 FILLER_52_1100 ();
 sg13g2_fill_8 FILLER_52_1108 ();
 sg13g2_fill_8 FILLER_52_1116 ();
 sg13g2_fill_8 FILLER_52_1124 ();
 sg13g2_fill_8 FILLER_52_1132 ();
 sg13g2_fill_4 FILLER_52_1140 ();
 sg13g2_fill_8 FILLER_53_0 ();
 sg13g2_fill_8 FILLER_53_8 ();
 sg13g2_fill_8 FILLER_53_16 ();
 sg13g2_fill_8 FILLER_53_24 ();
 sg13g2_fill_8 FILLER_53_32 ();
 sg13g2_fill_8 FILLER_53_40 ();
 sg13g2_fill_8 FILLER_53_48 ();
 sg13g2_fill_8 FILLER_53_56 ();
 sg13g2_fill_8 FILLER_53_64 ();
 sg13g2_fill_8 FILLER_53_72 ();
 sg13g2_fill_8 FILLER_53_80 ();
 sg13g2_fill_8 FILLER_53_88 ();
 sg13g2_fill_8 FILLER_53_96 ();
 sg13g2_fill_8 FILLER_53_104 ();
 sg13g2_fill_8 FILLER_53_112 ();
 sg13g2_fill_8 FILLER_53_120 ();
 sg13g2_fill_8 FILLER_53_128 ();
 sg13g2_fill_8 FILLER_53_136 ();
 sg13g2_fill_8 FILLER_53_144 ();
 sg13g2_fill_8 FILLER_53_152 ();
 sg13g2_fill_8 FILLER_53_160 ();
 sg13g2_fill_8 FILLER_53_168 ();
 sg13g2_fill_8 FILLER_53_176 ();
 sg13g2_fill_8 FILLER_53_184 ();
 sg13g2_fill_8 FILLER_53_192 ();
 sg13g2_fill_8 FILLER_53_200 ();
 sg13g2_fill_8 FILLER_53_208 ();
 sg13g2_fill_8 FILLER_53_216 ();
 sg13g2_fill_8 FILLER_53_224 ();
 sg13g2_fill_8 FILLER_53_232 ();
 sg13g2_fill_8 FILLER_53_240 ();
 sg13g2_fill_8 FILLER_53_248 ();
 sg13g2_fill_8 FILLER_53_256 ();
 sg13g2_fill_8 FILLER_53_264 ();
 sg13g2_fill_8 FILLER_53_272 ();
 sg13g2_fill_8 FILLER_53_280 ();
 sg13g2_fill_8 FILLER_53_288 ();
 sg13g2_fill_8 FILLER_53_296 ();
 sg13g2_fill_4 FILLER_53_304 ();
 sg13g2_fill_4 FILLER_53_334 ();
 sg13g2_fill_2 FILLER_53_338 ();
 sg13g2_fill_1 FILLER_53_340 ();
 sg13g2_fill_8 FILLER_53_397 ();
 sg13g2_fill_8 FILLER_53_405 ();
 sg13g2_fill_8 FILLER_53_413 ();
 sg13g2_fill_4 FILLER_53_421 ();
 sg13g2_fill_2 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_427 ();
 sg13g2_fill_4 FILLER_53_432 ();
 sg13g2_fill_1 FILLER_53_436 ();
 sg13g2_fill_8 FILLER_53_443 ();
 sg13g2_fill_8 FILLER_53_451 ();
 sg13g2_fill_8 FILLER_53_459 ();
 sg13g2_fill_8 FILLER_53_467 ();
 sg13g2_fill_8 FILLER_53_475 ();
 sg13g2_fill_4 FILLER_53_483 ();
 sg13g2_fill_1 FILLER_53_487 ();
 sg13g2_fill_8 FILLER_53_491 ();
 sg13g2_fill_8 FILLER_53_505 ();
 sg13g2_fill_4 FILLER_53_513 ();
 sg13g2_fill_2 FILLER_53_517 ();
 sg13g2_fill_8 FILLER_53_545 ();
 sg13g2_fill_4 FILLER_53_553 ();
 sg13g2_fill_2 FILLER_53_557 ();
 sg13g2_fill_8 FILLER_53_585 ();
 sg13g2_fill_8 FILLER_53_593 ();
 sg13g2_fill_8 FILLER_53_601 ();
 sg13g2_fill_8 FILLER_53_609 ();
 sg13g2_fill_8 FILLER_53_617 ();
 sg13g2_fill_8 FILLER_53_625 ();
 sg13g2_fill_8 FILLER_53_633 ();
 sg13g2_fill_8 FILLER_53_641 ();
 sg13g2_fill_8 FILLER_53_649 ();
 sg13g2_fill_8 FILLER_53_657 ();
 sg13g2_fill_8 FILLER_53_665 ();
 sg13g2_fill_8 FILLER_53_673 ();
 sg13g2_fill_8 FILLER_53_681 ();
 sg13g2_fill_8 FILLER_53_689 ();
 sg13g2_fill_8 FILLER_53_697 ();
 sg13g2_fill_8 FILLER_53_705 ();
 sg13g2_fill_8 FILLER_53_713 ();
 sg13g2_fill_8 FILLER_53_721 ();
 sg13g2_fill_8 FILLER_53_729 ();
 sg13g2_fill_8 FILLER_53_737 ();
 sg13g2_fill_8 FILLER_53_745 ();
 sg13g2_fill_8 FILLER_53_753 ();
 sg13g2_fill_8 FILLER_53_761 ();
 sg13g2_fill_8 FILLER_53_769 ();
 sg13g2_fill_8 FILLER_53_777 ();
 sg13g2_fill_8 FILLER_53_785 ();
 sg13g2_fill_8 FILLER_53_793 ();
 sg13g2_fill_8 FILLER_53_801 ();
 sg13g2_fill_8 FILLER_53_809 ();
 sg13g2_fill_8 FILLER_53_817 ();
 sg13g2_fill_8 FILLER_53_825 ();
 sg13g2_fill_8 FILLER_53_833 ();
 sg13g2_fill_8 FILLER_53_841 ();
 sg13g2_fill_8 FILLER_53_849 ();
 sg13g2_fill_8 FILLER_53_857 ();
 sg13g2_fill_8 FILLER_53_865 ();
 sg13g2_fill_8 FILLER_53_873 ();
 sg13g2_fill_8 FILLER_53_881 ();
 sg13g2_fill_8 FILLER_53_889 ();
 sg13g2_fill_8 FILLER_53_897 ();
 sg13g2_fill_8 FILLER_53_905 ();
 sg13g2_fill_8 FILLER_53_913 ();
 sg13g2_fill_8 FILLER_53_921 ();
 sg13g2_fill_8 FILLER_53_929 ();
 sg13g2_fill_8 FILLER_53_937 ();
 sg13g2_fill_8 FILLER_53_945 ();
 sg13g2_fill_8 FILLER_53_953 ();
 sg13g2_fill_8 FILLER_53_961 ();
 sg13g2_fill_8 FILLER_53_969 ();
 sg13g2_fill_8 FILLER_53_977 ();
 sg13g2_fill_8 FILLER_53_985 ();
 sg13g2_fill_8 FILLER_53_993 ();
 sg13g2_fill_8 FILLER_53_1001 ();
 sg13g2_fill_8 FILLER_53_1009 ();
 sg13g2_fill_8 FILLER_53_1017 ();
 sg13g2_fill_8 FILLER_53_1025 ();
 sg13g2_fill_8 FILLER_53_1033 ();
 sg13g2_fill_8 FILLER_53_1041 ();
 sg13g2_fill_8 FILLER_53_1049 ();
 sg13g2_fill_8 FILLER_53_1057 ();
 sg13g2_fill_8 FILLER_53_1065 ();
 sg13g2_fill_8 FILLER_53_1073 ();
 sg13g2_fill_8 FILLER_53_1081 ();
 sg13g2_fill_8 FILLER_53_1089 ();
 sg13g2_fill_8 FILLER_53_1097 ();
 sg13g2_fill_8 FILLER_53_1105 ();
 sg13g2_fill_8 FILLER_53_1113 ();
 sg13g2_fill_8 FILLER_53_1121 ();
 sg13g2_fill_8 FILLER_53_1129 ();
 sg13g2_fill_4 FILLER_53_1137 ();
 sg13g2_fill_2 FILLER_53_1141 ();
 sg13g2_fill_1 FILLER_53_1143 ();
 sg13g2_fill_8 FILLER_54_0 ();
 sg13g2_fill_8 FILLER_54_8 ();
 sg13g2_fill_8 FILLER_54_16 ();
 sg13g2_fill_8 FILLER_54_24 ();
 sg13g2_fill_8 FILLER_54_32 ();
 sg13g2_fill_8 FILLER_54_40 ();
 sg13g2_fill_8 FILLER_54_48 ();
 sg13g2_fill_8 FILLER_54_56 ();
 sg13g2_fill_8 FILLER_54_64 ();
 sg13g2_fill_8 FILLER_54_72 ();
 sg13g2_fill_8 FILLER_54_80 ();
 sg13g2_fill_8 FILLER_54_88 ();
 sg13g2_fill_8 FILLER_54_96 ();
 sg13g2_fill_8 FILLER_54_104 ();
 sg13g2_fill_8 FILLER_54_112 ();
 sg13g2_fill_8 FILLER_54_120 ();
 sg13g2_fill_8 FILLER_54_128 ();
 sg13g2_fill_8 FILLER_54_136 ();
 sg13g2_fill_8 FILLER_54_144 ();
 sg13g2_fill_8 FILLER_54_152 ();
 sg13g2_fill_8 FILLER_54_160 ();
 sg13g2_fill_8 FILLER_54_168 ();
 sg13g2_fill_8 FILLER_54_176 ();
 sg13g2_fill_8 FILLER_54_184 ();
 sg13g2_fill_8 FILLER_54_192 ();
 sg13g2_fill_8 FILLER_54_200 ();
 sg13g2_fill_8 FILLER_54_208 ();
 sg13g2_fill_8 FILLER_54_216 ();
 sg13g2_fill_8 FILLER_54_224 ();
 sg13g2_fill_8 FILLER_54_232 ();
 sg13g2_fill_8 FILLER_54_240 ();
 sg13g2_fill_8 FILLER_54_248 ();
 sg13g2_fill_8 FILLER_54_256 ();
 sg13g2_fill_8 FILLER_54_264 ();
 sg13g2_fill_8 FILLER_54_272 ();
 sg13g2_fill_8 FILLER_54_280 ();
 sg13g2_fill_8 FILLER_54_288 ();
 sg13g2_fill_8 FILLER_54_296 ();
 sg13g2_fill_8 FILLER_54_304 ();
 sg13g2_fill_8 FILLER_54_312 ();
 sg13g2_fill_8 FILLER_54_320 ();
 sg13g2_fill_8 FILLER_54_334 ();
 sg13g2_fill_8 FILLER_54_342 ();
 sg13g2_fill_8 FILLER_54_350 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_fill_1 FILLER_54_373 ();
 sg13g2_fill_1 FILLER_54_416 ();
 sg13g2_fill_2 FILLER_54_454 ();
 sg13g2_fill_8 FILLER_54_466 ();
 sg13g2_fill_8 FILLER_54_474 ();
 sg13g2_fill_1 FILLER_54_482 ();
 sg13g2_fill_8 FILLER_54_509 ();
 sg13g2_fill_8 FILLER_54_517 ();
 sg13g2_fill_8 FILLER_54_551 ();
 sg13g2_fill_1 FILLER_54_559 ();
 sg13g2_fill_1 FILLER_54_571 ();
 sg13g2_fill_2 FILLER_54_578 ();
 sg13g2_fill_8 FILLER_54_606 ();
 sg13g2_fill_8 FILLER_54_614 ();
 sg13g2_fill_8 FILLER_54_622 ();
 sg13g2_fill_8 FILLER_54_630 ();
 sg13g2_fill_8 FILLER_54_638 ();
 sg13g2_fill_8 FILLER_54_646 ();
 sg13g2_fill_8 FILLER_54_654 ();
 sg13g2_fill_8 FILLER_54_662 ();
 sg13g2_fill_8 FILLER_54_670 ();
 sg13g2_fill_8 FILLER_54_678 ();
 sg13g2_fill_8 FILLER_54_686 ();
 sg13g2_fill_8 FILLER_54_694 ();
 sg13g2_fill_8 FILLER_54_702 ();
 sg13g2_fill_8 FILLER_54_710 ();
 sg13g2_fill_8 FILLER_54_718 ();
 sg13g2_fill_8 FILLER_54_726 ();
 sg13g2_fill_8 FILLER_54_734 ();
 sg13g2_fill_8 FILLER_54_742 ();
 sg13g2_fill_8 FILLER_54_750 ();
 sg13g2_fill_8 FILLER_54_758 ();
 sg13g2_fill_8 FILLER_54_766 ();
 sg13g2_fill_8 FILLER_54_774 ();
 sg13g2_fill_8 FILLER_54_782 ();
 sg13g2_fill_8 FILLER_54_790 ();
 sg13g2_fill_8 FILLER_54_798 ();
 sg13g2_fill_8 FILLER_54_806 ();
 sg13g2_fill_8 FILLER_54_814 ();
 sg13g2_fill_8 FILLER_54_822 ();
 sg13g2_fill_8 FILLER_54_830 ();
 sg13g2_fill_8 FILLER_54_838 ();
 sg13g2_fill_8 FILLER_54_846 ();
 sg13g2_fill_8 FILLER_54_854 ();
 sg13g2_fill_8 FILLER_54_862 ();
 sg13g2_fill_8 FILLER_54_870 ();
 sg13g2_fill_8 FILLER_54_878 ();
 sg13g2_fill_8 FILLER_54_886 ();
 sg13g2_fill_8 FILLER_54_894 ();
 sg13g2_fill_8 FILLER_54_902 ();
 sg13g2_fill_8 FILLER_54_910 ();
 sg13g2_fill_8 FILLER_54_918 ();
 sg13g2_fill_8 FILLER_54_926 ();
 sg13g2_fill_8 FILLER_54_934 ();
 sg13g2_fill_8 FILLER_54_942 ();
 sg13g2_fill_8 FILLER_54_950 ();
 sg13g2_fill_8 FILLER_54_958 ();
 sg13g2_fill_8 FILLER_54_966 ();
 sg13g2_fill_8 FILLER_54_974 ();
 sg13g2_fill_8 FILLER_54_982 ();
 sg13g2_fill_8 FILLER_54_990 ();
 sg13g2_fill_8 FILLER_54_998 ();
 sg13g2_fill_8 FILLER_54_1006 ();
 sg13g2_fill_8 FILLER_54_1014 ();
 sg13g2_fill_8 FILLER_54_1022 ();
 sg13g2_fill_8 FILLER_54_1030 ();
 sg13g2_fill_8 FILLER_54_1038 ();
 sg13g2_fill_8 FILLER_54_1046 ();
 sg13g2_fill_8 FILLER_54_1054 ();
 sg13g2_fill_8 FILLER_54_1062 ();
 sg13g2_fill_8 FILLER_54_1070 ();
 sg13g2_fill_8 FILLER_54_1078 ();
 sg13g2_fill_8 FILLER_54_1086 ();
 sg13g2_fill_8 FILLER_54_1094 ();
 sg13g2_fill_8 FILLER_54_1102 ();
 sg13g2_fill_8 FILLER_54_1110 ();
 sg13g2_fill_8 FILLER_54_1118 ();
 sg13g2_fill_8 FILLER_54_1126 ();
 sg13g2_fill_8 FILLER_54_1134 ();
 sg13g2_fill_2 FILLER_54_1142 ();
 sg13g2_fill_8 FILLER_55_0 ();
 sg13g2_fill_8 FILLER_55_8 ();
 sg13g2_fill_8 FILLER_55_16 ();
 sg13g2_fill_8 FILLER_55_24 ();
 sg13g2_fill_8 FILLER_55_32 ();
 sg13g2_fill_8 FILLER_55_40 ();
 sg13g2_fill_8 FILLER_55_48 ();
 sg13g2_fill_8 FILLER_55_56 ();
 sg13g2_fill_8 FILLER_55_64 ();
 sg13g2_fill_8 FILLER_55_72 ();
 sg13g2_fill_8 FILLER_55_80 ();
 sg13g2_fill_8 FILLER_55_88 ();
 sg13g2_fill_8 FILLER_55_96 ();
 sg13g2_fill_8 FILLER_55_104 ();
 sg13g2_fill_8 FILLER_55_112 ();
 sg13g2_fill_8 FILLER_55_120 ();
 sg13g2_fill_8 FILLER_55_128 ();
 sg13g2_fill_8 FILLER_55_136 ();
 sg13g2_fill_8 FILLER_55_144 ();
 sg13g2_fill_8 FILLER_55_152 ();
 sg13g2_fill_8 FILLER_55_160 ();
 sg13g2_fill_8 FILLER_55_168 ();
 sg13g2_fill_8 FILLER_55_176 ();
 sg13g2_fill_8 FILLER_55_184 ();
 sg13g2_fill_8 FILLER_55_192 ();
 sg13g2_fill_8 FILLER_55_200 ();
 sg13g2_fill_8 FILLER_55_208 ();
 sg13g2_fill_8 FILLER_55_216 ();
 sg13g2_fill_8 FILLER_55_224 ();
 sg13g2_fill_8 FILLER_55_232 ();
 sg13g2_fill_8 FILLER_55_240 ();
 sg13g2_fill_8 FILLER_55_248 ();
 sg13g2_fill_8 FILLER_55_256 ();
 sg13g2_fill_8 FILLER_55_264 ();
 sg13g2_fill_8 FILLER_55_272 ();
 sg13g2_fill_8 FILLER_55_280 ();
 sg13g2_fill_8 FILLER_55_288 ();
 sg13g2_fill_8 FILLER_55_296 ();
 sg13g2_fill_4 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_308 ();
 sg13g2_fill_4 FILLER_55_341 ();
 sg13g2_fill_1 FILLER_55_345 ();
 sg13g2_fill_8 FILLER_55_372 ();
 sg13g2_fill_4 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_384 ();
 sg13g2_fill_2 FILLER_55_411 ();
 sg13g2_fill_1 FILLER_55_413 ();
 sg13g2_fill_4 FILLER_55_445 ();
 sg13g2_fill_2 FILLER_55_483 ();
 sg13g2_fill_1 FILLER_55_485 ();
 sg13g2_fill_1 FILLER_55_521 ();
 sg13g2_fill_1 FILLER_55_531 ();
 sg13g2_fill_8 FILLER_55_541 ();
 sg13g2_fill_4 FILLER_55_549 ();
 sg13g2_fill_1 FILLER_55_553 ();
 sg13g2_fill_8 FILLER_55_585 ();
 sg13g2_fill_8 FILLER_55_593 ();
 sg13g2_fill_8 FILLER_55_601 ();
 sg13g2_fill_8 FILLER_55_609 ();
 sg13g2_fill_8 FILLER_55_617 ();
 sg13g2_fill_8 FILLER_55_625 ();
 sg13g2_fill_8 FILLER_55_633 ();
 sg13g2_fill_8 FILLER_55_641 ();
 sg13g2_fill_8 FILLER_55_649 ();
 sg13g2_fill_8 FILLER_55_657 ();
 sg13g2_fill_8 FILLER_55_665 ();
 sg13g2_fill_8 FILLER_55_673 ();
 sg13g2_fill_8 FILLER_55_681 ();
 sg13g2_fill_8 FILLER_55_689 ();
 sg13g2_fill_8 FILLER_55_697 ();
 sg13g2_fill_8 FILLER_55_705 ();
 sg13g2_fill_8 FILLER_55_713 ();
 sg13g2_fill_8 FILLER_55_721 ();
 sg13g2_fill_8 FILLER_55_729 ();
 sg13g2_fill_8 FILLER_55_737 ();
 sg13g2_fill_8 FILLER_55_745 ();
 sg13g2_fill_8 FILLER_55_753 ();
 sg13g2_fill_8 FILLER_55_761 ();
 sg13g2_fill_8 FILLER_55_769 ();
 sg13g2_fill_8 FILLER_55_777 ();
 sg13g2_fill_8 FILLER_55_785 ();
 sg13g2_fill_8 FILLER_55_793 ();
 sg13g2_fill_8 FILLER_55_801 ();
 sg13g2_fill_8 FILLER_55_809 ();
 sg13g2_fill_8 FILLER_55_817 ();
 sg13g2_fill_8 FILLER_55_825 ();
 sg13g2_fill_8 FILLER_55_833 ();
 sg13g2_fill_8 FILLER_55_841 ();
 sg13g2_fill_8 FILLER_55_849 ();
 sg13g2_fill_8 FILLER_55_857 ();
 sg13g2_fill_8 FILLER_55_865 ();
 sg13g2_fill_8 FILLER_55_873 ();
 sg13g2_fill_8 FILLER_55_881 ();
 sg13g2_fill_8 FILLER_55_889 ();
 sg13g2_fill_8 FILLER_55_897 ();
 sg13g2_fill_8 FILLER_55_905 ();
 sg13g2_fill_8 FILLER_55_913 ();
 sg13g2_fill_8 FILLER_55_921 ();
 sg13g2_fill_8 FILLER_55_929 ();
 sg13g2_fill_8 FILLER_55_937 ();
 sg13g2_fill_8 FILLER_55_945 ();
 sg13g2_fill_8 FILLER_55_953 ();
 sg13g2_fill_8 FILLER_55_961 ();
 sg13g2_fill_8 FILLER_55_969 ();
 sg13g2_fill_8 FILLER_55_977 ();
 sg13g2_fill_8 FILLER_55_985 ();
 sg13g2_fill_8 FILLER_55_993 ();
 sg13g2_fill_8 FILLER_55_1001 ();
 sg13g2_fill_8 FILLER_55_1009 ();
 sg13g2_fill_8 FILLER_55_1017 ();
 sg13g2_fill_8 FILLER_55_1025 ();
 sg13g2_fill_8 FILLER_55_1033 ();
 sg13g2_fill_8 FILLER_55_1041 ();
 sg13g2_fill_8 FILLER_55_1049 ();
 sg13g2_fill_8 FILLER_55_1057 ();
 sg13g2_fill_8 FILLER_55_1065 ();
 sg13g2_fill_8 FILLER_55_1073 ();
 sg13g2_fill_8 FILLER_55_1081 ();
 sg13g2_fill_8 FILLER_55_1089 ();
 sg13g2_fill_8 FILLER_55_1097 ();
 sg13g2_fill_4 FILLER_55_1115 ();
 sg13g2_fill_2 FILLER_55_1119 ();
 sg13g2_fill_1 FILLER_55_1121 ();
 sg13g2_fill_8 FILLER_55_1130 ();
 sg13g2_fill_4 FILLER_55_1138 ();
 sg13g2_fill_2 FILLER_55_1142 ();
 sg13g2_fill_8 FILLER_56_0 ();
 sg13g2_fill_8 FILLER_56_8 ();
 sg13g2_fill_8 FILLER_56_16 ();
 sg13g2_fill_8 FILLER_56_24 ();
 sg13g2_fill_8 FILLER_56_32 ();
 sg13g2_fill_8 FILLER_56_40 ();
 sg13g2_fill_8 FILLER_56_48 ();
 sg13g2_fill_8 FILLER_56_56 ();
 sg13g2_fill_8 FILLER_56_64 ();
 sg13g2_fill_8 FILLER_56_72 ();
 sg13g2_fill_8 FILLER_56_80 ();
 sg13g2_fill_8 FILLER_56_88 ();
 sg13g2_fill_8 FILLER_56_96 ();
 sg13g2_fill_8 FILLER_56_104 ();
 sg13g2_fill_8 FILLER_56_112 ();
 sg13g2_fill_8 FILLER_56_120 ();
 sg13g2_fill_8 FILLER_56_128 ();
 sg13g2_fill_8 FILLER_56_136 ();
 sg13g2_fill_8 FILLER_56_144 ();
 sg13g2_fill_8 FILLER_56_152 ();
 sg13g2_fill_8 FILLER_56_160 ();
 sg13g2_fill_8 FILLER_56_168 ();
 sg13g2_fill_8 FILLER_56_176 ();
 sg13g2_fill_8 FILLER_56_184 ();
 sg13g2_fill_8 FILLER_56_192 ();
 sg13g2_fill_8 FILLER_56_200 ();
 sg13g2_fill_8 FILLER_56_208 ();
 sg13g2_fill_8 FILLER_56_216 ();
 sg13g2_fill_8 FILLER_56_224 ();
 sg13g2_fill_8 FILLER_56_232 ();
 sg13g2_fill_8 FILLER_56_240 ();
 sg13g2_fill_8 FILLER_56_248 ();
 sg13g2_fill_8 FILLER_56_256 ();
 sg13g2_fill_8 FILLER_56_264 ();
 sg13g2_fill_8 FILLER_56_272 ();
 sg13g2_fill_8 FILLER_56_280 ();
 sg13g2_fill_8 FILLER_56_288 ();
 sg13g2_fill_8 FILLER_56_296 ();
 sg13g2_fill_8 FILLER_56_304 ();
 sg13g2_fill_8 FILLER_56_312 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_8 FILLER_56_365 ();
 sg13g2_fill_8 FILLER_56_373 ();
 sg13g2_fill_8 FILLER_56_381 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_fill_4 FILLER_56_396 ();
 sg13g2_fill_2 FILLER_56_411 ();
 sg13g2_fill_1 FILLER_56_413 ();
 sg13g2_fill_8 FILLER_56_419 ();
 sg13g2_fill_1 FILLER_56_427 ();
 sg13g2_fill_8 FILLER_56_432 ();
 sg13g2_fill_4 FILLER_56_440 ();
 sg13g2_fill_1 FILLER_56_449 ();
 sg13g2_fill_8 FILLER_56_486 ();
 sg13g2_fill_4 FILLER_56_494 ();
 sg13g2_fill_1 FILLER_56_498 ();
 sg13g2_fill_2 FILLER_56_502 ();
 sg13g2_fill_2 FILLER_56_510 ();
 sg13g2_fill_8 FILLER_56_518 ();
 sg13g2_fill_4 FILLER_56_526 ();
 sg13g2_fill_1 FILLER_56_533 ();
 sg13g2_fill_8 FILLER_56_540 ();
 sg13g2_fill_8 FILLER_56_548 ();
 sg13g2_fill_1 FILLER_56_564 ();
 sg13g2_fill_8 FILLER_56_576 ();
 sg13g2_fill_8 FILLER_56_584 ();
 sg13g2_fill_8 FILLER_56_592 ();
 sg13g2_fill_8 FILLER_56_600 ();
 sg13g2_fill_8 FILLER_56_608 ();
 sg13g2_fill_8 FILLER_56_616 ();
 sg13g2_fill_8 FILLER_56_624 ();
 sg13g2_fill_8 FILLER_56_632 ();
 sg13g2_fill_8 FILLER_56_640 ();
 sg13g2_fill_8 FILLER_56_648 ();
 sg13g2_fill_8 FILLER_56_656 ();
 sg13g2_fill_8 FILLER_56_664 ();
 sg13g2_fill_8 FILLER_56_672 ();
 sg13g2_fill_8 FILLER_56_680 ();
 sg13g2_fill_8 FILLER_56_688 ();
 sg13g2_fill_8 FILLER_56_696 ();
 sg13g2_fill_8 FILLER_56_704 ();
 sg13g2_fill_8 FILLER_56_712 ();
 sg13g2_fill_8 FILLER_56_720 ();
 sg13g2_fill_8 FILLER_56_728 ();
 sg13g2_fill_8 FILLER_56_736 ();
 sg13g2_fill_8 FILLER_56_744 ();
 sg13g2_fill_8 FILLER_56_752 ();
 sg13g2_fill_8 FILLER_56_760 ();
 sg13g2_fill_8 FILLER_56_768 ();
 sg13g2_fill_8 FILLER_56_776 ();
 sg13g2_fill_8 FILLER_56_784 ();
 sg13g2_fill_8 FILLER_56_792 ();
 sg13g2_fill_8 FILLER_56_800 ();
 sg13g2_fill_8 FILLER_56_808 ();
 sg13g2_fill_8 FILLER_56_816 ();
 sg13g2_fill_8 FILLER_56_824 ();
 sg13g2_fill_8 FILLER_56_832 ();
 sg13g2_fill_8 FILLER_56_840 ();
 sg13g2_fill_8 FILLER_56_848 ();
 sg13g2_fill_8 FILLER_56_856 ();
 sg13g2_fill_8 FILLER_56_864 ();
 sg13g2_fill_8 FILLER_56_872 ();
 sg13g2_fill_8 FILLER_56_880 ();
 sg13g2_fill_8 FILLER_56_888 ();
 sg13g2_fill_8 FILLER_56_896 ();
 sg13g2_fill_8 FILLER_56_904 ();
 sg13g2_fill_8 FILLER_56_912 ();
 sg13g2_fill_8 FILLER_56_920 ();
 sg13g2_fill_8 FILLER_56_928 ();
 sg13g2_fill_4 FILLER_56_936 ();
 sg13g2_fill_8 FILLER_56_944 ();
 sg13g2_fill_8 FILLER_56_952 ();
 sg13g2_fill_8 FILLER_56_960 ();
 sg13g2_fill_8 FILLER_56_968 ();
 sg13g2_fill_4 FILLER_56_976 ();
 sg13g2_fill_1 FILLER_56_980 ();
 sg13g2_fill_8 FILLER_56_985 ();
 sg13g2_fill_4 FILLER_56_993 ();
 sg13g2_fill_1 FILLER_56_997 ();
 sg13g2_fill_4 FILLER_56_1008 ();
 sg13g2_fill_2 FILLER_56_1012 ();
 sg13g2_fill_1 FILLER_56_1014 ();
 sg13g2_fill_8 FILLER_56_1019 ();
 sg13g2_fill_8 FILLER_56_1027 ();
 sg13g2_fill_8 FILLER_56_1035 ();
 sg13g2_fill_8 FILLER_56_1043 ();
 sg13g2_fill_1 FILLER_56_1051 ();
 sg13g2_fill_2 FILLER_56_1062 ();
 sg13g2_fill_8 FILLER_57_0 ();
 sg13g2_fill_8 FILLER_57_8 ();
 sg13g2_fill_8 FILLER_57_16 ();
 sg13g2_fill_8 FILLER_57_24 ();
 sg13g2_fill_8 FILLER_57_32 ();
 sg13g2_fill_8 FILLER_57_40 ();
 sg13g2_fill_8 FILLER_57_48 ();
 sg13g2_fill_8 FILLER_57_56 ();
 sg13g2_fill_8 FILLER_57_64 ();
 sg13g2_fill_8 FILLER_57_72 ();
 sg13g2_fill_8 FILLER_57_80 ();
 sg13g2_fill_8 FILLER_57_88 ();
 sg13g2_fill_8 FILLER_57_96 ();
 sg13g2_fill_8 FILLER_57_104 ();
 sg13g2_fill_8 FILLER_57_112 ();
 sg13g2_fill_8 FILLER_57_120 ();
 sg13g2_fill_8 FILLER_57_128 ();
 sg13g2_fill_8 FILLER_57_136 ();
 sg13g2_fill_8 FILLER_57_144 ();
 sg13g2_fill_8 FILLER_57_152 ();
 sg13g2_fill_8 FILLER_57_160 ();
 sg13g2_fill_8 FILLER_57_168 ();
 sg13g2_fill_8 FILLER_57_176 ();
 sg13g2_fill_8 FILLER_57_184 ();
 sg13g2_fill_8 FILLER_57_192 ();
 sg13g2_fill_8 FILLER_57_200 ();
 sg13g2_fill_8 FILLER_57_208 ();
 sg13g2_fill_8 FILLER_57_216 ();
 sg13g2_fill_8 FILLER_57_224 ();
 sg13g2_fill_8 FILLER_57_232 ();
 sg13g2_fill_8 FILLER_57_240 ();
 sg13g2_fill_8 FILLER_57_248 ();
 sg13g2_fill_8 FILLER_57_256 ();
 sg13g2_fill_8 FILLER_57_264 ();
 sg13g2_fill_8 FILLER_57_272 ();
 sg13g2_fill_8 FILLER_57_280 ();
 sg13g2_fill_8 FILLER_57_288 ();
 sg13g2_fill_8 FILLER_57_296 ();
 sg13g2_fill_8 FILLER_57_304 ();
 sg13g2_fill_8 FILLER_57_312 ();
 sg13g2_fill_8 FILLER_57_320 ();
 sg13g2_fill_2 FILLER_57_332 ();
 sg13g2_fill_8 FILLER_57_340 ();
 sg13g2_fill_2 FILLER_57_348 ();
 sg13g2_fill_1 FILLER_57_350 ();
 sg13g2_fill_4 FILLER_57_355 ();
 sg13g2_fill_2 FILLER_57_359 ();
 sg13g2_fill_1 FILLER_57_361 ();
 sg13g2_fill_4 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_378 ();
 sg13g2_fill_8 FILLER_57_400 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_fill_8 FILLER_57_413 ();
 sg13g2_fill_4 FILLER_57_421 ();
 sg13g2_fill_2 FILLER_57_425 ();
 sg13g2_fill_1 FILLER_57_427 ();
 sg13g2_fill_1 FILLER_57_433 ();
 sg13g2_fill_8 FILLER_57_439 ();
 sg13g2_fill_8 FILLER_57_447 ();
 sg13g2_fill_8 FILLER_57_463 ();
 sg13g2_fill_8 FILLER_57_471 ();
 sg13g2_fill_8 FILLER_57_479 ();
 sg13g2_fill_8 FILLER_57_487 ();
 sg13g2_fill_4 FILLER_57_495 ();
 sg13g2_fill_8 FILLER_57_551 ();
 sg13g2_fill_8 FILLER_57_573 ();
 sg13g2_fill_8 FILLER_57_581 ();
 sg13g2_fill_2 FILLER_57_589 ();
 sg13g2_fill_1 FILLER_57_591 ();
 sg13g2_fill_8 FILLER_57_678 ();
 sg13g2_fill_8 FILLER_57_686 ();
 sg13g2_fill_8 FILLER_57_694 ();
 sg13g2_fill_8 FILLER_57_702 ();
 sg13g2_fill_8 FILLER_57_710 ();
 sg13g2_fill_8 FILLER_57_718 ();
 sg13g2_fill_8 FILLER_57_726 ();
 sg13g2_fill_8 FILLER_57_734 ();
 sg13g2_fill_8 FILLER_57_742 ();
 sg13g2_fill_8 FILLER_57_750 ();
 sg13g2_fill_8 FILLER_57_758 ();
 sg13g2_fill_8 FILLER_57_766 ();
 sg13g2_fill_8 FILLER_57_774 ();
 sg13g2_fill_8 FILLER_57_782 ();
 sg13g2_fill_8 FILLER_57_790 ();
 sg13g2_fill_8 FILLER_57_798 ();
 sg13g2_fill_8 FILLER_57_806 ();
 sg13g2_fill_8 FILLER_57_814 ();
 sg13g2_fill_8 FILLER_57_822 ();
 sg13g2_fill_8 FILLER_57_830 ();
 sg13g2_fill_8 FILLER_57_838 ();
 sg13g2_fill_8 FILLER_57_846 ();
 sg13g2_fill_8 FILLER_57_854 ();
 sg13g2_fill_8 FILLER_57_862 ();
 sg13g2_fill_8 FILLER_57_870 ();
 sg13g2_fill_8 FILLER_57_878 ();
 sg13g2_fill_8 FILLER_57_886 ();
 sg13g2_fill_8 FILLER_57_894 ();
 sg13g2_fill_8 FILLER_57_902 ();
 sg13g2_fill_8 FILLER_57_910 ();
 sg13g2_fill_8 FILLER_57_918 ();
 sg13g2_fill_4 FILLER_57_926 ();
 sg13g2_fill_2 FILLER_57_930 ();
 sg13g2_fill_1 FILLER_57_932 ();
 sg13g2_fill_8 FILLER_57_959 ();
 sg13g2_fill_4 FILLER_57_967 ();
 sg13g2_fill_2 FILLER_57_971 ();
 sg13g2_fill_1 FILLER_57_973 ();
 sg13g2_fill_4 FILLER_57_1000 ();
 sg13g2_fill_2 FILLER_57_1004 ();
 sg13g2_fill_1 FILLER_57_1006 ();
 sg13g2_fill_4 FILLER_57_1037 ();
 sg13g2_fill_1 FILLER_57_1041 ();
 sg13g2_fill_8 FILLER_57_1086 ();
 sg13g2_fill_8 FILLER_57_1094 ();
 sg13g2_fill_2 FILLER_57_1102 ();
 sg13g2_fill_8 FILLER_58_0 ();
 sg13g2_fill_8 FILLER_58_8 ();
 sg13g2_fill_8 FILLER_58_16 ();
 sg13g2_fill_8 FILLER_58_24 ();
 sg13g2_fill_4 FILLER_58_32 ();
 sg13g2_fill_1 FILLER_58_36 ();
 sg13g2_fill_8 FILLER_58_41 ();
 sg13g2_fill_8 FILLER_58_49 ();
 sg13g2_fill_8 FILLER_58_57 ();
 sg13g2_fill_8 FILLER_58_65 ();
 sg13g2_fill_8 FILLER_58_73 ();
 sg13g2_fill_8 FILLER_58_81 ();
 sg13g2_fill_8 FILLER_58_89 ();
 sg13g2_fill_8 FILLER_58_97 ();
 sg13g2_fill_8 FILLER_58_105 ();
 sg13g2_fill_8 FILLER_58_113 ();
 sg13g2_fill_8 FILLER_58_121 ();
 sg13g2_fill_8 FILLER_58_129 ();
 sg13g2_fill_8 FILLER_58_137 ();
 sg13g2_fill_8 FILLER_58_145 ();
 sg13g2_fill_8 FILLER_58_153 ();
 sg13g2_fill_8 FILLER_58_161 ();
 sg13g2_fill_8 FILLER_58_169 ();
 sg13g2_fill_8 FILLER_58_177 ();
 sg13g2_fill_8 FILLER_58_185 ();
 sg13g2_fill_8 FILLER_58_193 ();
 sg13g2_fill_8 FILLER_58_201 ();
 sg13g2_fill_8 FILLER_58_209 ();
 sg13g2_fill_8 FILLER_58_217 ();
 sg13g2_fill_8 FILLER_58_225 ();
 sg13g2_fill_8 FILLER_58_233 ();
 sg13g2_fill_8 FILLER_58_241 ();
 sg13g2_fill_8 FILLER_58_249 ();
 sg13g2_fill_8 FILLER_58_257 ();
 sg13g2_fill_8 FILLER_58_265 ();
 sg13g2_fill_8 FILLER_58_273 ();
 sg13g2_fill_8 FILLER_58_281 ();
 sg13g2_fill_8 FILLER_58_289 ();
 sg13g2_fill_8 FILLER_58_297 ();
 sg13g2_fill_8 FILLER_58_305 ();
 sg13g2_fill_8 FILLER_58_313 ();
 sg13g2_fill_2 FILLER_58_321 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_fill_8 FILLER_58_328 ();
 sg13g2_fill_4 FILLER_58_342 ();
 sg13g2_fill_2 FILLER_58_346 ();
 sg13g2_fill_1 FILLER_58_378 ();
 sg13g2_fill_8 FILLER_58_405 ();
 sg13g2_fill_4 FILLER_58_413 ();
 sg13g2_fill_4 FILLER_58_443 ();
 sg13g2_fill_1 FILLER_58_447 ();
 sg13g2_fill_8 FILLER_58_453 ();
 sg13g2_fill_4 FILLER_58_461 ();
 sg13g2_fill_1 FILLER_58_465 ();
 sg13g2_fill_4 FILLER_58_471 ();
 sg13g2_fill_2 FILLER_58_483 ();
 sg13g2_fill_8 FILLER_58_490 ();
 sg13g2_fill_8 FILLER_58_498 ();
 sg13g2_fill_1 FILLER_58_506 ();
 sg13g2_fill_8 FILLER_58_510 ();
 sg13g2_fill_4 FILLER_58_518 ();
 sg13g2_fill_2 FILLER_58_522 ();
 sg13g2_fill_4 FILLER_58_545 ();
 sg13g2_fill_1 FILLER_58_549 ();
 sg13g2_fill_4 FILLER_58_580 ();
 sg13g2_fill_8 FILLER_58_614 ();
 sg13g2_fill_8 FILLER_58_622 ();
 sg13g2_fill_4 FILLER_58_630 ();
 sg13g2_fill_2 FILLER_58_634 ();
 sg13g2_fill_8 FILLER_58_666 ();
 sg13g2_fill_4 FILLER_58_674 ();
 sg13g2_fill_8 FILLER_58_704 ();
 sg13g2_fill_8 FILLER_58_720 ();
 sg13g2_fill_8 FILLER_58_728 ();
 sg13g2_fill_8 FILLER_58_736 ();
 sg13g2_fill_8 FILLER_58_744 ();
 sg13g2_fill_8 FILLER_58_752 ();
 sg13g2_fill_8 FILLER_58_760 ();
 sg13g2_fill_8 FILLER_58_768 ();
 sg13g2_fill_8 FILLER_58_776 ();
 sg13g2_fill_8 FILLER_58_784 ();
 sg13g2_fill_8 FILLER_58_792 ();
 sg13g2_fill_8 FILLER_58_800 ();
 sg13g2_fill_8 FILLER_58_808 ();
 sg13g2_fill_8 FILLER_58_816 ();
 sg13g2_fill_8 FILLER_58_824 ();
 sg13g2_fill_8 FILLER_58_832 ();
 sg13g2_fill_8 FILLER_58_840 ();
 sg13g2_fill_8 FILLER_58_848 ();
 sg13g2_fill_8 FILLER_58_856 ();
 sg13g2_fill_8 FILLER_58_864 ();
 sg13g2_fill_8 FILLER_58_872 ();
 sg13g2_fill_8 FILLER_58_880 ();
 sg13g2_fill_8 FILLER_58_888 ();
 sg13g2_fill_8 FILLER_58_896 ();
 sg13g2_fill_8 FILLER_58_904 ();
 sg13g2_fill_2 FILLER_58_912 ();
 sg13g2_fill_8 FILLER_58_934 ();
 sg13g2_fill_8 FILLER_58_942 ();
 sg13g2_fill_8 FILLER_58_950 ();
 sg13g2_fill_1 FILLER_58_958 ();
 sg13g2_fill_8 FILLER_58_979 ();
 sg13g2_fill_8 FILLER_58_987 ();
 sg13g2_fill_2 FILLER_58_995 ();
 sg13g2_fill_1 FILLER_58_997 ();
 sg13g2_fill_2 FILLER_58_1008 ();
 sg13g2_fill_1 FILLER_58_1010 ();
 sg13g2_fill_4 FILLER_58_1037 ();
 sg13g2_fill_2 FILLER_58_1041 ();
 sg13g2_fill_1 FILLER_58_1043 ();
 sg13g2_fill_8 FILLER_58_1081 ();
 sg13g2_fill_8 FILLER_58_1089 ();
 sg13g2_fill_8 FILLER_58_1097 ();
 sg13g2_fill_8 FILLER_58_1115 ();
 sg13g2_fill_8 FILLER_58_1127 ();
 sg13g2_fill_8 FILLER_58_1135 ();
 sg13g2_fill_1 FILLER_58_1143 ();
 sg13g2_fill_8 FILLER_59_0 ();
 sg13g2_fill_8 FILLER_59_8 ();
 sg13g2_fill_2 FILLER_59_26 ();
 sg13g2_fill_1 FILLER_59_28 ();
 sg13g2_fill_8 FILLER_59_55 ();
 sg13g2_fill_8 FILLER_59_63 ();
 sg13g2_fill_8 FILLER_59_71 ();
 sg13g2_fill_8 FILLER_59_79 ();
 sg13g2_fill_8 FILLER_59_87 ();
 sg13g2_fill_8 FILLER_59_95 ();
 sg13g2_fill_8 FILLER_59_103 ();
 sg13g2_fill_8 FILLER_59_111 ();
 sg13g2_fill_8 FILLER_59_119 ();
 sg13g2_fill_8 FILLER_59_127 ();
 sg13g2_fill_8 FILLER_59_135 ();
 sg13g2_fill_8 FILLER_59_143 ();
 sg13g2_fill_8 FILLER_59_151 ();
 sg13g2_fill_8 FILLER_59_159 ();
 sg13g2_fill_8 FILLER_59_167 ();
 sg13g2_fill_8 FILLER_59_175 ();
 sg13g2_fill_8 FILLER_59_183 ();
 sg13g2_fill_8 FILLER_59_191 ();
 sg13g2_fill_1 FILLER_59_199 ();
 sg13g2_fill_8 FILLER_59_210 ();
 sg13g2_fill_4 FILLER_59_218 ();
 sg13g2_fill_8 FILLER_59_230 ();
 sg13g2_fill_8 FILLER_59_238 ();
 sg13g2_fill_8 FILLER_59_246 ();
 sg13g2_fill_8 FILLER_59_254 ();
 sg13g2_fill_8 FILLER_59_262 ();
 sg13g2_fill_8 FILLER_59_270 ();
 sg13g2_fill_8 FILLER_59_278 ();
 sg13g2_fill_8 FILLER_59_286 ();
 sg13g2_fill_8 FILLER_59_294 ();
 sg13g2_fill_8 FILLER_59_302 ();
 sg13g2_fill_4 FILLER_59_310 ();
 sg13g2_fill_2 FILLER_59_352 ();
 sg13g2_fill_8 FILLER_59_358 ();
 sg13g2_fill_8 FILLER_59_366 ();
 sg13g2_fill_8 FILLER_59_374 ();
 sg13g2_fill_2 FILLER_59_382 ();
 sg13g2_fill_4 FILLER_59_388 ();
 sg13g2_fill_2 FILLER_59_392 ();
 sg13g2_fill_8 FILLER_59_399 ();
 sg13g2_fill_8 FILLER_59_407 ();
 sg13g2_fill_4 FILLER_59_467 ();
 sg13g2_fill_8 FILLER_59_502 ();
 sg13g2_fill_8 FILLER_59_510 ();
 sg13g2_fill_2 FILLER_59_518 ();
 sg13g2_fill_1 FILLER_59_520 ();
 sg13g2_fill_8 FILLER_59_547 ();
 sg13g2_fill_2 FILLER_59_555 ();
 sg13g2_fill_1 FILLER_59_557 ();
 sg13g2_fill_8 FILLER_59_569 ();
 sg13g2_fill_8 FILLER_59_577 ();
 sg13g2_fill_4 FILLER_59_585 ();
 sg13g2_fill_2 FILLER_59_589 ();
 sg13g2_fill_2 FILLER_59_596 ();
 sg13g2_fill_8 FILLER_59_608 ();
 sg13g2_fill_4 FILLER_59_616 ();
 sg13g2_fill_2 FILLER_59_648 ();
 sg13g2_fill_1 FILLER_59_650 ();
 sg13g2_fill_8 FILLER_59_659 ();
 sg13g2_fill_4 FILLER_59_667 ();
 sg13g2_fill_2 FILLER_59_671 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_fill_8 FILLER_59_764 ();
 sg13g2_fill_8 FILLER_59_772 ();
 sg13g2_fill_8 FILLER_59_780 ();
 sg13g2_fill_8 FILLER_59_788 ();
 sg13g2_fill_8 FILLER_59_796 ();
 sg13g2_fill_8 FILLER_59_804 ();
 sg13g2_fill_8 FILLER_59_812 ();
 sg13g2_fill_8 FILLER_59_820 ();
 sg13g2_fill_8 FILLER_59_828 ();
 sg13g2_fill_8 FILLER_59_836 ();
 sg13g2_fill_8 FILLER_59_844 ();
 sg13g2_fill_8 FILLER_59_852 ();
 sg13g2_fill_8 FILLER_59_860 ();
 sg13g2_fill_8 FILLER_59_868 ();
 sg13g2_fill_8 FILLER_59_876 ();
 sg13g2_fill_8 FILLER_59_884 ();
 sg13g2_fill_2 FILLER_59_892 ();
 sg13g2_fill_1 FILLER_59_894 ();
 sg13g2_fill_2 FILLER_59_899 ();
 sg13g2_fill_2 FILLER_59_911 ();
 sg13g2_fill_8 FILLER_59_939 ();
 sg13g2_fill_8 FILLER_59_951 ();
 sg13g2_fill_4 FILLER_59_959 ();
 sg13g2_fill_1 FILLER_59_963 ();
 sg13g2_fill_8 FILLER_59_986 ();
 sg13g2_fill_4 FILLER_59_994 ();
 sg13g2_fill_2 FILLER_59_998 ();
 sg13g2_fill_8 FILLER_59_1024 ();
 sg13g2_fill_4 FILLER_59_1032 ();
 sg13g2_fill_2 FILLER_59_1036 ();
 sg13g2_fill_2 FILLER_59_1048 ();
 sg13g2_fill_1 FILLER_59_1050 ();
 sg13g2_fill_8 FILLER_59_1055 ();
 sg13g2_fill_8 FILLER_59_1063 ();
 sg13g2_fill_8 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1079 ();
 sg13g2_fill_1 FILLER_59_1081 ();
 sg13g2_fill_8 FILLER_59_1086 ();
 sg13g2_fill_2 FILLER_59_1094 ();
 sg13g2_fill_4 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_4 ();
 sg13g2_fill_8 FILLER_60_36 ();
 sg13g2_fill_8 FILLER_60_44 ();
 sg13g2_fill_8 FILLER_60_52 ();
 sg13g2_fill_8 FILLER_60_60 ();
 sg13g2_fill_8 FILLER_60_68 ();
 sg13g2_fill_8 FILLER_60_76 ();
 sg13g2_fill_8 FILLER_60_84 ();
 sg13g2_fill_8 FILLER_60_92 ();
 sg13g2_fill_8 FILLER_60_100 ();
 sg13g2_fill_8 FILLER_60_108 ();
 sg13g2_fill_8 FILLER_60_116 ();
 sg13g2_fill_8 FILLER_60_124 ();
 sg13g2_fill_1 FILLER_60_132 ();
 sg13g2_fill_8 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_151 ();
 sg13g2_fill_8 FILLER_60_157 ();
 sg13g2_fill_8 FILLER_60_165 ();
 sg13g2_fill_8 FILLER_60_173 ();
 sg13g2_fill_8 FILLER_60_181 ();
 sg13g2_fill_2 FILLER_60_189 ();
 sg13g2_fill_8 FILLER_60_237 ();
 sg13g2_fill_2 FILLER_60_255 ();
 sg13g2_fill_4 FILLER_60_261 ();
 sg13g2_fill_2 FILLER_60_265 ();
 sg13g2_fill_1 FILLER_60_267 ();
 sg13g2_fill_8 FILLER_60_278 ();
 sg13g2_fill_8 FILLER_60_290 ();
 sg13g2_fill_8 FILLER_60_298 ();
 sg13g2_fill_4 FILLER_60_306 ();
 sg13g2_fill_2 FILLER_60_310 ();
 sg13g2_fill_2 FILLER_60_342 ();
 sg13g2_fill_8 FILLER_60_376 ();
 sg13g2_fill_1 FILLER_60_384 ();
 sg13g2_fill_8 FILLER_60_389 ();
 sg13g2_fill_8 FILLER_60_397 ();
 sg13g2_fill_4 FILLER_60_405 ();
 sg13g2_fill_2 FILLER_60_449 ();
 sg13g2_fill_2 FILLER_60_463 ();
 sg13g2_fill_8 FILLER_60_502 ();
 sg13g2_fill_8 FILLER_60_510 ();
 sg13g2_fill_8 FILLER_60_518 ();
 sg13g2_fill_8 FILLER_60_526 ();
 sg13g2_fill_8 FILLER_60_534 ();
 sg13g2_fill_8 FILLER_60_542 ();
 sg13g2_fill_4 FILLER_60_550 ();
 sg13g2_fill_2 FILLER_60_554 ();
 sg13g2_fill_8 FILLER_60_560 ();
 sg13g2_fill_8 FILLER_60_568 ();
 sg13g2_fill_4 FILLER_60_576 ();
 sg13g2_fill_2 FILLER_60_580 ();
 sg13g2_fill_1 FILLER_60_582 ();
 sg13g2_fill_4 FILLER_60_590 ();
 sg13g2_fill_2 FILLER_60_594 ();
 sg13g2_fill_8 FILLER_60_600 ();
 sg13g2_fill_2 FILLER_60_608 ();
 sg13g2_fill_1 FILLER_60_620 ();
 sg13g2_fill_8 FILLER_60_635 ();
 sg13g2_fill_8 FILLER_60_643 ();
 sg13g2_fill_8 FILLER_60_683 ();
 sg13g2_fill_8 FILLER_60_691 ();
 sg13g2_fill_8 FILLER_60_699 ();
 sg13g2_fill_8 FILLER_60_707 ();
 sg13g2_fill_4 FILLER_60_715 ();
 sg13g2_fill_2 FILLER_60_719 ();
 sg13g2_fill_8 FILLER_60_726 ();
 sg13g2_fill_8 FILLER_60_734 ();
 sg13g2_fill_4 FILLER_60_742 ();
 sg13g2_fill_2 FILLER_60_746 ();
 sg13g2_fill_4 FILLER_60_778 ();
 sg13g2_fill_8 FILLER_60_808 ();
 sg13g2_fill_8 FILLER_60_816 ();
 sg13g2_fill_8 FILLER_60_824 ();
 sg13g2_fill_8 FILLER_60_832 ();
 sg13g2_fill_8 FILLER_60_840 ();
 sg13g2_fill_8 FILLER_60_848 ();
 sg13g2_fill_8 FILLER_60_856 ();
 sg13g2_fill_8 FILLER_60_864 ();
 sg13g2_fill_8 FILLER_60_872 ();
 sg13g2_fill_8 FILLER_60_880 ();
 sg13g2_fill_1 FILLER_60_888 ();
 sg13g2_fill_4 FILLER_60_915 ();
 sg13g2_fill_1 FILLER_60_919 ();
 sg13g2_fill_4 FILLER_60_924 ();
 sg13g2_fill_1 FILLER_60_928 ();
 sg13g2_fill_1 FILLER_60_939 ();
 sg13g2_fill_4 FILLER_60_966 ();
 sg13g2_fill_2 FILLER_60_970 ();
 sg13g2_fill_2 FILLER_60_998 ();
 sg13g2_fill_1 FILLER_60_1000 ();
 sg13g2_fill_4 FILLER_60_1011 ();
 sg13g2_fill_8 FILLER_60_1019 ();
 sg13g2_fill_4 FILLER_60_1027 ();
 sg13g2_fill_2 FILLER_60_1031 ();
 sg13g2_fill_1 FILLER_60_1073 ();
 sg13g2_fill_8 FILLER_60_1128 ();
 sg13g2_fill_8 FILLER_60_1136 ();
 sg13g2_fill_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_8 ();
 sg13g2_fill_4 FILLER_61_20 ();
 sg13g2_fill_2 FILLER_61_24 ();
 sg13g2_fill_4 FILLER_61_43 ();
 sg13g2_fill_2 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_49 ();
 sg13g2_fill_8 FILLER_61_54 ();
 sg13g2_fill_8 FILLER_61_62 ();
 sg13g2_fill_8 FILLER_61_70 ();
 sg13g2_fill_8 FILLER_61_78 ();
 sg13g2_fill_8 FILLER_61_86 ();
 sg13g2_fill_8 FILLER_61_94 ();
 sg13g2_fill_8 FILLER_61_102 ();
 sg13g2_fill_8 FILLER_61_110 ();
 sg13g2_fill_8 FILLER_61_118 ();
 sg13g2_fill_8 FILLER_61_126 ();
 sg13g2_fill_8 FILLER_61_174 ();
 sg13g2_fill_8 FILLER_61_182 ();
 sg13g2_fill_8 FILLER_61_190 ();
 sg13g2_fill_4 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_212 ();
 sg13g2_fill_1 FILLER_61_276 ();
 sg13g2_fill_8 FILLER_61_307 ();
 sg13g2_fill_4 FILLER_61_315 ();
 sg13g2_fill_1 FILLER_61_319 ();
 sg13g2_fill_1 FILLER_61_346 ();
 sg13g2_fill_8 FILLER_61_356 ();
 sg13g2_fill_8 FILLER_61_364 ();
 sg13g2_fill_4 FILLER_61_372 ();
 sg13g2_fill_2 FILLER_61_376 ();
 sg13g2_fill_8 FILLER_61_404 ();
 sg13g2_fill_4 FILLER_61_412 ();
 sg13g2_fill_8 FILLER_61_420 ();
 sg13g2_fill_8 FILLER_61_428 ();
 sg13g2_fill_8 FILLER_61_436 ();
 sg13g2_fill_4 FILLER_61_444 ();
 sg13g2_fill_2 FILLER_61_448 ();
 sg13g2_fill_2 FILLER_61_459 ();
 sg13g2_fill_1 FILLER_61_461 ();
 sg13g2_fill_8 FILLER_61_466 ();
 sg13g2_fill_8 FILLER_61_483 ();
 sg13g2_fill_8 FILLER_61_491 ();
 sg13g2_fill_2 FILLER_61_503 ();
 sg13g2_fill_1 FILLER_61_505 ();
 sg13g2_fill_4 FILLER_61_546 ();
 sg13g2_fill_1 FILLER_61_550 ();
 sg13g2_fill_8 FILLER_61_572 ();
 sg13g2_fill_1 FILLER_61_580 ();
 sg13g2_fill_4 FILLER_61_585 ();
 sg13g2_fill_1 FILLER_61_589 ();
 sg13g2_fill_4 FILLER_61_594 ();
 sg13g2_fill_1 FILLER_61_598 ();
 sg13g2_fill_2 FILLER_61_603 ();
 sg13g2_fill_1 FILLER_61_605 ();
 sg13g2_fill_2 FILLER_61_624 ();
 sg13g2_fill_4 FILLER_61_640 ();
 sg13g2_fill_2 FILLER_61_644 ();
 sg13g2_fill_8 FILLER_61_650 ();
 sg13g2_fill_4 FILLER_61_658 ();
 sg13g2_fill_2 FILLER_61_662 ();
 sg13g2_fill_1 FILLER_61_664 ();
 sg13g2_fill_4 FILLER_61_669 ();
 sg13g2_fill_8 FILLER_61_678 ();
 sg13g2_fill_8 FILLER_61_686 ();
 sg13g2_fill_8 FILLER_61_694 ();
 sg13g2_fill_8 FILLER_61_702 ();
 sg13g2_fill_8 FILLER_61_710 ();
 sg13g2_fill_4 FILLER_61_718 ();
 sg13g2_fill_2 FILLER_61_722 ();
 sg13g2_fill_1 FILLER_61_724 ();
 sg13g2_fill_1 FILLER_61_751 ();
 sg13g2_fill_8 FILLER_61_771 ();
 sg13g2_fill_2 FILLER_61_779 ();
 sg13g2_fill_4 FILLER_61_785 ();
 sg13g2_fill_2 FILLER_61_789 ();
 sg13g2_fill_8 FILLER_61_821 ();
 sg13g2_fill_8 FILLER_61_829 ();
 sg13g2_fill_8 FILLER_61_837 ();
 sg13g2_fill_1 FILLER_61_845 ();
 sg13g2_fill_8 FILLER_61_876 ();
 sg13g2_fill_2 FILLER_61_884 ();
 sg13g2_fill_1 FILLER_61_886 ();
 sg13g2_fill_8 FILLER_61_917 ();
 sg13g2_fill_4 FILLER_61_925 ();
 sg13g2_fill_1 FILLER_61_929 ();
 sg13g2_fill_8 FILLER_61_940 ();
 sg13g2_fill_8 FILLER_61_948 ();
 sg13g2_fill_8 FILLER_61_956 ();
 sg13g2_fill_8 FILLER_61_974 ();
 sg13g2_fill_4 FILLER_61_982 ();
 sg13g2_fill_2 FILLER_61_986 ();
 sg13g2_fill_4 FILLER_61_992 ();
 sg13g2_fill_1 FILLER_61_996 ();
 sg13g2_fill_2 FILLER_61_1033 ();
 sg13g2_fill_2 FILLER_61_1045 ();
 sg13g2_fill_8 FILLER_61_1051 ();
 sg13g2_fill_4 FILLER_61_1059 ();
 sg13g2_fill_2 FILLER_61_1063 ();
 sg13g2_fill_2 FILLER_61_1095 ();
 sg13g2_fill_1 FILLER_61_1097 ();
 sg13g2_fill_2 FILLER_61_1111 ();
 sg13g2_fill_1 FILLER_61_1113 ();
 sg13g2_fill_4 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_4 ();
 sg13g2_fill_8 FILLER_62_67 ();
 sg13g2_fill_8 FILLER_62_75 ();
 sg13g2_fill_8 FILLER_62_83 ();
 sg13g2_fill_8 FILLER_62_91 ();
 sg13g2_fill_8 FILLER_62_99 ();
 sg13g2_fill_8 FILLER_62_107 ();
 sg13g2_fill_8 FILLER_62_115 ();
 sg13g2_fill_8 FILLER_62_123 ();
 sg13g2_fill_8 FILLER_62_131 ();
 sg13g2_fill_2 FILLER_62_139 ();
 sg13g2_fill_2 FILLER_62_151 ();
 sg13g2_fill_4 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_187 ();
 sg13g2_fill_1 FILLER_62_199 ();
 sg13g2_fill_8 FILLER_62_210 ();
 sg13g2_fill_2 FILLER_62_218 ();
 sg13g2_fill_1 FILLER_62_220 ();
 sg13g2_fill_8 FILLER_62_225 ();
 sg13g2_fill_8 FILLER_62_233 ();
 sg13g2_fill_8 FILLER_62_241 ();
 sg13g2_fill_8 FILLER_62_249 ();
 sg13g2_fill_8 FILLER_62_257 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_fill_4 FILLER_62_322 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_8 FILLER_62_331 ();
 sg13g2_fill_2 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_341 ();
 sg13g2_fill_8 FILLER_62_368 ();
 sg13g2_fill_8 FILLER_62_376 ();
 sg13g2_fill_4 FILLER_62_411 ();
 sg13g2_fill_1 FILLER_62_415 ();
 sg13g2_fill_8 FILLER_62_442 ();
 sg13g2_fill_4 FILLER_62_450 ();
 sg13g2_fill_1 FILLER_62_468 ();
 sg13g2_fill_4 FILLER_62_474 ();
 sg13g2_fill_2 FILLER_62_478 ();
 sg13g2_fill_2 FILLER_62_492 ();
 sg13g2_fill_1 FILLER_62_494 ();
 sg13g2_fill_8 FILLER_62_514 ();
 sg13g2_fill_2 FILLER_62_522 ();
 sg13g2_fill_1 FILLER_62_524 ();
 sg13g2_fill_8 FILLER_62_542 ();
 sg13g2_fill_8 FILLER_62_550 ();
 sg13g2_fill_8 FILLER_62_558 ();
 sg13g2_fill_2 FILLER_62_566 ();
 sg13g2_fill_4 FILLER_62_573 ();
 sg13g2_fill_2 FILLER_62_577 ();
 sg13g2_fill_8 FILLER_62_584 ();
 sg13g2_fill_4 FILLER_62_618 ();
 sg13g2_fill_8 FILLER_62_626 ();
 sg13g2_fill_8 FILLER_62_634 ();
 sg13g2_fill_8 FILLER_62_642 ();
 sg13g2_fill_4 FILLER_62_650 ();
 sg13g2_fill_2 FILLER_62_658 ();
 sg13g2_fill_1 FILLER_62_660 ();
 sg13g2_fill_4 FILLER_62_714 ();
 sg13g2_fill_1 FILLER_62_718 ();
 sg13g2_fill_2 FILLER_62_728 ();
 sg13g2_fill_8 FILLER_62_749 ();
 sg13g2_fill_8 FILLER_62_761 ();
 sg13g2_fill_2 FILLER_62_769 ();
 sg13g2_fill_1 FILLER_62_776 ();
 sg13g2_fill_8 FILLER_62_796 ();
 sg13g2_fill_8 FILLER_62_804 ();
 sg13g2_fill_8 FILLER_62_812 ();
 sg13g2_fill_4 FILLER_62_820 ();
 sg13g2_fill_2 FILLER_62_824 ();
 sg13g2_fill_4 FILLER_62_856 ();
 sg13g2_fill_1 FILLER_62_860 ();
 sg13g2_fill_8 FILLER_62_865 ();
 sg13g2_fill_8 FILLER_62_873 ();
 sg13g2_fill_8 FILLER_62_881 ();
 sg13g2_fill_8 FILLER_62_889 ();
 sg13g2_fill_8 FILLER_62_897 ();
 sg13g2_fill_4 FILLER_62_915 ();
 sg13g2_fill_2 FILLER_62_919 ();
 sg13g2_fill_1 FILLER_62_925 ();
 sg13g2_fill_8 FILLER_62_936 ();
 sg13g2_fill_8 FILLER_62_948 ();
 sg13g2_fill_8 FILLER_62_956 ();
 sg13g2_fill_4 FILLER_62_964 ();
 sg13g2_fill_1 FILLER_62_968 ();
 sg13g2_fill_1 FILLER_62_979 ();
 sg13g2_fill_8 FILLER_62_1006 ();
 sg13g2_fill_8 FILLER_62_1014 ();
 sg13g2_fill_8 FILLER_62_1022 ();
 sg13g2_fill_2 FILLER_62_1070 ();
 sg13g2_fill_1 FILLER_62_1072 ();
 sg13g2_fill_8 FILLER_62_1090 ();
 sg13g2_fill_4 FILLER_62_1098 ();
 sg13g2_fill_1 FILLER_62_1102 ();
 sg13g2_fill_8 FILLER_62_1113 ();
 sg13g2_fill_2 FILLER_62_1121 ();
 sg13g2_fill_8 FILLER_62_1127 ();
 sg13g2_fill_8 FILLER_62_1135 ();
 sg13g2_fill_1 FILLER_62_1143 ();
 sg13g2_fill_8 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_22 ();
 sg13g2_fill_4 FILLER_63_63 ();
 sg13g2_fill_2 FILLER_63_67 ();
 sg13g2_fill_8 FILLER_63_73 ();
 sg13g2_fill_8 FILLER_63_81 ();
 sg13g2_fill_8 FILLER_63_89 ();
 sg13g2_fill_8 FILLER_63_97 ();
 sg13g2_fill_8 FILLER_63_105 ();
 sg13g2_fill_8 FILLER_63_113 ();
 sg13g2_fill_8 FILLER_63_121 ();
 sg13g2_fill_8 FILLER_63_129 ();
 sg13g2_fill_2 FILLER_63_137 ();
 sg13g2_fill_8 FILLER_63_149 ();
 sg13g2_fill_1 FILLER_63_157 ();
 sg13g2_fill_2 FILLER_63_172 ();
 sg13g2_fill_1 FILLER_63_174 ();
 sg13g2_fill_4 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_197 ();
 sg13g2_fill_4 FILLER_63_209 ();
 sg13g2_fill_8 FILLER_63_239 ();
 sg13g2_fill_1 FILLER_63_247 ();
 sg13g2_fill_8 FILLER_63_258 ();
 sg13g2_fill_1 FILLER_63_266 ();
 sg13g2_fill_8 FILLER_63_271 ();
 sg13g2_fill_8 FILLER_63_289 ();
 sg13g2_fill_2 FILLER_63_297 ();
 sg13g2_fill_1 FILLER_63_299 ();
 sg13g2_fill_8 FILLER_63_304 ();
 sg13g2_fill_8 FILLER_63_312 ();
 sg13g2_fill_8 FILLER_63_320 ();
 sg13g2_fill_8 FILLER_63_328 ();
 sg13g2_fill_8 FILLER_63_336 ();
 sg13g2_fill_8 FILLER_63_344 ();
 sg13g2_fill_8 FILLER_63_352 ();
 sg13g2_fill_8 FILLER_63_360 ();
 sg13g2_fill_4 FILLER_63_368 ();
 sg13g2_fill_2 FILLER_63_372 ();
 sg13g2_fill_1 FILLER_63_410 ();
 sg13g2_fill_1 FILLER_63_426 ();
 sg13g2_fill_4 FILLER_63_453 ();
 sg13g2_fill_1 FILLER_63_457 ();
 sg13g2_fill_2 FILLER_63_465 ();
 sg13g2_fill_1 FILLER_63_467 ();
 sg13g2_fill_2 FILLER_63_499 ();
 sg13g2_fill_1 FILLER_63_501 ();
 sg13g2_fill_2 FILLER_63_511 ();
 sg13g2_fill_1 FILLER_63_513 ();
 sg13g2_fill_4 FILLER_63_566 ();
 sg13g2_fill_2 FILLER_63_570 ();
 sg13g2_fill_1 FILLER_63_572 ();
 sg13g2_fill_4 FILLER_63_608 ();
 sg13g2_fill_1 FILLER_63_621 ();
 sg13g2_fill_8 FILLER_63_627 ();
 sg13g2_fill_4 FILLER_63_635 ();
 sg13g2_fill_1 FILLER_63_639 ();
 sg13g2_fill_4 FILLER_63_644 ();
 sg13g2_fill_4 FILLER_63_679 ();
 sg13g2_fill_2 FILLER_63_683 ();
 sg13g2_fill_2 FILLER_63_746 ();
 sg13g2_fill_1 FILLER_63_748 ();
 sg13g2_fill_1 FILLER_63_775 ();
 sg13g2_fill_4 FILLER_63_785 ();
 sg13g2_fill_2 FILLER_63_789 ();
 sg13g2_fill_8 FILLER_63_821 ();
 sg13g2_fill_8 FILLER_63_841 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_4 FILLER_63_893 ();
 sg13g2_fill_1 FILLER_63_912 ();
 sg13g2_fill_2 FILLER_63_990 ();
 sg13g2_fill_1 FILLER_63_992 ();
 sg13g2_fill_8 FILLER_63_997 ();
 sg13g2_fill_8 FILLER_63_1005 ();
 sg13g2_fill_8 FILLER_63_1013 ();
 sg13g2_fill_8 FILLER_63_1021 ();
 sg13g2_fill_8 FILLER_63_1029 ();
 sg13g2_fill_1 FILLER_63_1037 ();
 sg13g2_fill_8 FILLER_63_1046 ();
 sg13g2_fill_8 FILLER_63_1054 ();
 sg13g2_fill_1 FILLER_63_1062 ();
 sg13g2_fill_4 FILLER_63_1108 ();
 sg13g2_fill_2 FILLER_63_1112 ();
 sg13g2_fill_8 FILLER_64_0 ();
 sg13g2_fill_4 FILLER_64_18 ();
 sg13g2_fill_1 FILLER_64_22 ();
 sg13g2_fill_8 FILLER_64_31 ();
 sg13g2_fill_8 FILLER_64_39 ();
 sg13g2_fill_4 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_51 ();
 sg13g2_fill_8 FILLER_64_88 ();
 sg13g2_fill_8 FILLER_64_96 ();
 sg13g2_fill_4 FILLER_64_104 ();
 sg13g2_fill_2 FILLER_64_108 ();
 sg13g2_fill_4 FILLER_64_174 ();
 sg13g2_fill_2 FILLER_64_178 ();
 sg13g2_fill_8 FILLER_64_184 ();
 sg13g2_fill_8 FILLER_64_192 ();
 sg13g2_fill_8 FILLER_64_210 ();
 sg13g2_fill_2 FILLER_64_218 ();
 sg13g2_fill_8 FILLER_64_224 ();
 sg13g2_fill_8 FILLER_64_232 ();
 sg13g2_fill_1 FILLER_64_258 ();
 sg13g2_fill_4 FILLER_64_289 ();
 sg13g2_fill_8 FILLER_64_329 ();
 sg13g2_fill_8 FILLER_64_337 ();
 sg13g2_fill_8 FILLER_64_345 ();
 sg13g2_fill_8 FILLER_64_353 ();
 sg13g2_fill_8 FILLER_64_361 ();
 sg13g2_fill_4 FILLER_64_369 ();
 sg13g2_fill_2 FILLER_64_373 ();
 sg13g2_fill_1 FILLER_64_401 ();
 sg13g2_fill_4 FILLER_64_413 ();
 sg13g2_fill_2 FILLER_64_417 ();
 sg13g2_fill_8 FILLER_64_434 ();
 sg13g2_fill_8 FILLER_64_442 ();
 sg13g2_fill_4 FILLER_64_450 ();
 sg13g2_fill_1 FILLER_64_454 ();
 sg13g2_fill_8 FILLER_64_460 ();
 sg13g2_fill_8 FILLER_64_468 ();
 sg13g2_fill_4 FILLER_64_476 ();
 sg13g2_fill_2 FILLER_64_480 ();
 sg13g2_fill_2 FILLER_64_496 ();
 sg13g2_fill_4 FILLER_64_503 ();
 sg13g2_fill_2 FILLER_64_507 ();
 sg13g2_fill_1 FILLER_64_509 ();
 sg13g2_fill_2 FILLER_64_518 ();
 sg13g2_fill_1 FILLER_64_520 ();
 sg13g2_fill_4 FILLER_64_543 ();
 sg13g2_fill_2 FILLER_64_547 ();
 sg13g2_fill_8 FILLER_64_558 ();
 sg13g2_fill_4 FILLER_64_566 ();
 sg13g2_fill_2 FILLER_64_570 ();
 sg13g2_fill_1 FILLER_64_572 ();
 sg13g2_fill_1 FILLER_64_578 ();
 sg13g2_fill_4 FILLER_64_584 ();
 sg13g2_fill_2 FILLER_64_588 ();
 sg13g2_fill_1 FILLER_64_594 ();
 sg13g2_fill_2 FILLER_64_603 ();
 sg13g2_fill_1 FILLER_64_605 ();
 sg13g2_fill_4 FILLER_64_655 ();
 sg13g2_fill_2 FILLER_64_664 ();
 sg13g2_fill_4 FILLER_64_675 ();
 sg13g2_fill_8 FILLER_64_688 ();
 sg13g2_fill_4 FILLER_64_696 ();
 sg13g2_fill_1 FILLER_64_700 ();
 sg13g2_fill_4 FILLER_64_710 ();
 sg13g2_fill_1 FILLER_64_714 ();
 sg13g2_fill_2 FILLER_64_719 ();
 sg13g2_fill_2 FILLER_64_726 ();
 sg13g2_fill_1 FILLER_64_728 ();
 sg13g2_fill_8 FILLER_64_738 ();
 sg13g2_fill_8 FILLER_64_746 ();
 sg13g2_fill_8 FILLER_64_754 ();
 sg13g2_fill_8 FILLER_64_781 ();
 sg13g2_fill_8 FILLER_64_789 ();
 sg13g2_fill_1 FILLER_64_797 ();
 sg13g2_fill_8 FILLER_64_828 ();
 sg13g2_fill_2 FILLER_64_836 ();
 sg13g2_fill_1 FILLER_64_838 ();
 sg13g2_fill_1 FILLER_64_844 ();
 sg13g2_fill_2 FILLER_64_855 ();
 sg13g2_fill_1 FILLER_64_857 ();
 sg13g2_fill_8 FILLER_64_873 ();
 sg13g2_fill_8 FILLER_64_881 ();
 sg13g2_fill_8 FILLER_64_889 ();
 sg13g2_fill_8 FILLER_64_897 ();
 sg13g2_fill_4 FILLER_64_905 ();
 sg13g2_fill_2 FILLER_64_909 ();
 sg13g2_fill_1 FILLER_64_911 ();
 sg13g2_fill_4 FILLER_64_920 ();
 sg13g2_fill_1 FILLER_64_924 ();
 sg13g2_fill_8 FILLER_64_935 ();
 sg13g2_fill_4 FILLER_64_943 ();
 sg13g2_fill_2 FILLER_64_947 ();
 sg13g2_fill_8 FILLER_64_953 ();
 sg13g2_fill_4 FILLER_64_966 ();
 sg13g2_fill_2 FILLER_64_970 ();
 sg13g2_fill_4 FILLER_64_982 ();
 sg13g2_fill_2 FILLER_64_1012 ();
 sg13g2_fill_1 FILLER_64_1014 ();
 sg13g2_fill_8 FILLER_64_1035 ();
 sg13g2_fill_4 FILLER_64_1043 ();
 sg13g2_fill_8 FILLER_64_1057 ();
 sg13g2_fill_8 FILLER_64_1069 ();
 sg13g2_fill_8 FILLER_64_1077 ();
 sg13g2_fill_8 FILLER_64_1085 ();
 sg13g2_fill_8 FILLER_64_1093 ();
 sg13g2_fill_2 FILLER_64_1101 ();
 sg13g2_fill_1 FILLER_64_1103 ();
 sg13g2_fill_8 FILLER_64_1114 ();
 sg13g2_fill_1 FILLER_64_1122 ();
 sg13g2_fill_4 FILLER_64_1127 ();
 sg13g2_fill_8 FILLER_65_0 ();
 sg13g2_fill_8 FILLER_65_18 ();
 sg13g2_fill_8 FILLER_65_26 ();
 sg13g2_fill_8 FILLER_65_34 ();
 sg13g2_fill_8 FILLER_65_42 ();
 sg13g2_fill_8 FILLER_65_50 ();
 sg13g2_fill_8 FILLER_65_58 ();
 sg13g2_fill_8 FILLER_65_66 ();
 sg13g2_fill_8 FILLER_65_74 ();
 sg13g2_fill_8 FILLER_65_82 ();
 sg13g2_fill_8 FILLER_65_90 ();
 sg13g2_fill_8 FILLER_65_98 ();
 sg13g2_fill_8 FILLER_65_106 ();
 sg13g2_fill_8 FILLER_65_114 ();
 sg13g2_fill_2 FILLER_65_122 ();
 sg13g2_fill_1 FILLER_65_124 ();
 sg13g2_fill_4 FILLER_65_165 ();
 sg13g2_fill_2 FILLER_65_169 ();
 sg13g2_fill_8 FILLER_65_201 ();
 sg13g2_fill_2 FILLER_65_209 ();
 sg13g2_fill_1 FILLER_65_211 ();
 sg13g2_fill_4 FILLER_65_238 ();
 sg13g2_fill_1 FILLER_65_242 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_8 FILLER_65_258 ();
 sg13g2_fill_8 FILLER_65_266 ();
 sg13g2_fill_8 FILLER_65_274 ();
 sg13g2_fill_2 FILLER_65_282 ();
 sg13g2_fill_1 FILLER_65_284 ();
 sg13g2_fill_1 FILLER_65_305 ();
 sg13g2_fill_8 FILLER_65_332 ();
 sg13g2_fill_8 FILLER_65_340 ();
 sg13g2_fill_8 FILLER_65_348 ();
 sg13g2_fill_8 FILLER_65_356 ();
 sg13g2_fill_8 FILLER_65_364 ();
 sg13g2_fill_8 FILLER_65_372 ();
 sg13g2_fill_8 FILLER_65_380 ();
 sg13g2_fill_8 FILLER_65_388 ();
 sg13g2_fill_8 FILLER_65_396 ();
 sg13g2_fill_8 FILLER_65_404 ();
 sg13g2_fill_8 FILLER_65_412 ();
 sg13g2_fill_8 FILLER_65_420 ();
 sg13g2_fill_8 FILLER_65_428 ();
 sg13g2_fill_8 FILLER_65_470 ();
 sg13g2_fill_8 FILLER_65_478 ();
 sg13g2_fill_8 FILLER_65_486 ();
 sg13g2_fill_8 FILLER_65_494 ();
 sg13g2_fill_2 FILLER_65_502 ();
 sg13g2_fill_1 FILLER_65_504 ();
 sg13g2_fill_8 FILLER_65_510 ();
 sg13g2_fill_4 FILLER_65_518 ();
 sg13g2_fill_2 FILLER_65_522 ();
 sg13g2_fill_2 FILLER_65_528 ();
 sg13g2_fill_8 FILLER_65_534 ();
 sg13g2_fill_8 FILLER_65_542 ();
 sg13g2_fill_2 FILLER_65_550 ();
 sg13g2_fill_2 FILLER_65_557 ();
 sg13g2_fill_1 FILLER_65_613 ();
 sg13g2_fill_2 FILLER_65_628 ();
 sg13g2_fill_8 FILLER_65_635 ();
 sg13g2_fill_8 FILLER_65_643 ();
 sg13g2_fill_8 FILLER_65_651 ();
 sg13g2_fill_4 FILLER_65_672 ();
 sg13g2_fill_2 FILLER_65_676 ();
 sg13g2_fill_8 FILLER_65_682 ();
 sg13g2_fill_8 FILLER_65_690 ();
 sg13g2_fill_8 FILLER_65_698 ();
 sg13g2_fill_4 FILLER_65_706 ();
 sg13g2_fill_2 FILLER_65_710 ();
 sg13g2_fill_1 FILLER_65_712 ();
 sg13g2_fill_4 FILLER_65_721 ();
 sg13g2_fill_8 FILLER_65_735 ();
 sg13g2_fill_8 FILLER_65_743 ();
 sg13g2_fill_8 FILLER_65_751 ();
 sg13g2_fill_1 FILLER_65_759 ();
 sg13g2_fill_1 FILLER_65_768 ();
 sg13g2_fill_8 FILLER_65_781 ();
 sg13g2_fill_4 FILLER_65_789 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_799 ();
 sg13g2_fill_8 FILLER_65_808 ();
 sg13g2_fill_8 FILLER_65_816 ();
 sg13g2_fill_8 FILLER_65_824 ();
 sg13g2_fill_1 FILLER_65_845 ();
 sg13g2_fill_2 FILLER_65_876 ();
 sg13g2_fill_8 FILLER_65_914 ();
 sg13g2_fill_8 FILLER_65_922 ();
 sg13g2_fill_1 FILLER_65_930 ();
 sg13g2_fill_8 FILLER_65_967 ();
 sg13g2_fill_8 FILLER_65_975 ();
 sg13g2_fill_4 FILLER_65_983 ();
 sg13g2_fill_1 FILLER_65_987 ();
 sg13g2_fill_8 FILLER_65_998 ();
 sg13g2_fill_4 FILLER_65_1010 ();
 sg13g2_fill_2 FILLER_65_1014 ();
 sg13g2_fill_1 FILLER_65_1016 ();
 sg13g2_fill_8 FILLER_65_1087 ();
 sg13g2_fill_8 FILLER_65_1095 ();
 sg13g2_fill_1 FILLER_65_1103 ();
 sg13g2_fill_4 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_4 ();
 sg13g2_fill_2 FILLER_66_51 ();
 sg13g2_fill_8 FILLER_66_67 ();
 sg13g2_fill_1 FILLER_66_75 ();
 sg13g2_fill_8 FILLER_66_80 ();
 sg13g2_fill_8 FILLER_66_88 ();
 sg13g2_fill_8 FILLER_66_96 ();
 sg13g2_fill_8 FILLER_66_104 ();
 sg13g2_fill_8 FILLER_66_112 ();
 sg13g2_fill_4 FILLER_66_120 ();
 sg13g2_fill_4 FILLER_66_134 ();
 sg13g2_fill_2 FILLER_66_142 ();
 sg13g2_fill_4 FILLER_66_152 ();
 sg13g2_fill_2 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_158 ();
 sg13g2_fill_8 FILLER_66_183 ();
 sg13g2_fill_4 FILLER_66_191 ();
 sg13g2_fill_2 FILLER_66_195 ();
 sg13g2_fill_1 FILLER_66_197 ();
 sg13g2_fill_8 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_216 ();
 sg13g2_fill_8 FILLER_66_222 ();
 sg13g2_fill_4 FILLER_66_230 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_2 FILLER_66_281 ();
 sg13g2_fill_8 FILLER_66_293 ();
 sg13g2_fill_8 FILLER_66_301 ();
 sg13g2_fill_4 FILLER_66_309 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_fill_4 FILLER_66_322 ();
 sg13g2_fill_2 FILLER_66_326 ();
 sg13g2_fill_8 FILLER_66_347 ();
 sg13g2_fill_8 FILLER_66_355 ();
 sg13g2_fill_8 FILLER_66_363 ();
 sg13g2_fill_8 FILLER_66_371 ();
 sg13g2_fill_8 FILLER_66_379 ();
 sg13g2_fill_8 FILLER_66_387 ();
 sg13g2_fill_4 FILLER_66_395 ();
 sg13g2_fill_2 FILLER_66_399 ();
 sg13g2_fill_1 FILLER_66_401 ();
 sg13g2_fill_4 FILLER_66_412 ();
 sg13g2_fill_1 FILLER_66_416 ();
 sg13g2_fill_8 FILLER_66_435 ();
 sg13g2_fill_4 FILLER_66_443 ();
 sg13g2_fill_4 FILLER_66_465 ();
 sg13g2_fill_2 FILLER_66_469 ();
 sg13g2_fill_1 FILLER_66_471 ();
 sg13g2_fill_8 FILLER_66_492 ();
 sg13g2_fill_8 FILLER_66_500 ();
 sg13g2_fill_2 FILLER_66_508 ();
 sg13g2_fill_8 FILLER_66_534 ();
 sg13g2_fill_8 FILLER_66_542 ();
 sg13g2_fill_2 FILLER_66_550 ();
 sg13g2_fill_1 FILLER_66_552 ();
 sg13g2_fill_1 FILLER_66_557 ();
 sg13g2_fill_8 FILLER_66_563 ();
 sg13g2_fill_1 FILLER_66_571 ();
 sg13g2_fill_8 FILLER_66_576 ();
 sg13g2_fill_2 FILLER_66_584 ();
 sg13g2_fill_4 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_595 ();
 sg13g2_fill_1 FILLER_66_597 ();
 sg13g2_fill_2 FILLER_66_602 ();
 sg13g2_fill_8 FILLER_66_608 ();
 sg13g2_fill_8 FILLER_66_616 ();
 sg13g2_fill_8 FILLER_66_624 ();
 sg13g2_fill_8 FILLER_66_632 ();
 sg13g2_fill_8 FILLER_66_640 ();
 sg13g2_fill_8 FILLER_66_648 ();
 sg13g2_fill_4 FILLER_66_656 ();
 sg13g2_fill_1 FILLER_66_660 ();
 sg13g2_fill_8 FILLER_66_685 ();
 sg13g2_fill_2 FILLER_66_693 ();
 sg13g2_fill_1 FILLER_66_695 ();
 sg13g2_fill_4 FILLER_66_719 ();
 sg13g2_fill_2 FILLER_66_723 ();
 sg13g2_fill_1 FILLER_66_725 ();
 sg13g2_fill_2 FILLER_66_730 ();
 sg13g2_fill_8 FILLER_66_742 ();
 sg13g2_fill_4 FILLER_66_750 ();
 sg13g2_fill_2 FILLER_66_754 ();
 sg13g2_fill_2 FILLER_66_761 ();
 sg13g2_fill_1 FILLER_66_763 ();
 sg13g2_fill_4 FILLER_66_786 ();
 sg13g2_fill_1 FILLER_66_790 ();
 sg13g2_fill_8 FILLER_66_821 ();
 sg13g2_fill_2 FILLER_66_829 ();
 sg13g2_fill_1 FILLER_66_831 ();
 sg13g2_fill_8 FILLER_66_836 ();
 sg13g2_fill_8 FILLER_66_844 ();
 sg13g2_fill_2 FILLER_66_852 ();
 sg13g2_fill_8 FILLER_66_903 ();
 sg13g2_fill_8 FILLER_66_911 ();
 sg13g2_fill_4 FILLER_66_919 ();
 sg13g2_fill_2 FILLER_66_923 ();
 sg13g2_fill_1 FILLER_66_925 ();
 sg13g2_fill_4 FILLER_66_930 ();
 sg13g2_fill_2 FILLER_66_934 ();
 sg13g2_fill_8 FILLER_66_946 ();
 sg13g2_fill_4 FILLER_66_954 ();
 sg13g2_fill_2 FILLER_66_958 ();
 sg13g2_fill_4 FILLER_66_970 ();
 sg13g2_fill_2 FILLER_66_974 ();
 sg13g2_fill_1 FILLER_66_976 ();
 sg13g2_fill_4 FILLER_66_981 ();
 sg13g2_fill_1 FILLER_66_985 ();
 sg13g2_fill_2 FILLER_66_996 ();
 sg13g2_fill_1 FILLER_66_998 ();
 sg13g2_fill_4 FILLER_66_1029 ();
 sg13g2_fill_1 FILLER_66_1033 ();
 sg13g2_fill_8 FILLER_66_1081 ();
 sg13g2_fill_4 FILLER_66_1089 ();
 sg13g2_fill_1 FILLER_66_1093 ();
 sg13g2_fill_4 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_4 ();
 sg13g2_fill_8 FILLER_67_94 ();
 sg13g2_fill_8 FILLER_67_102 ();
 sg13g2_fill_8 FILLER_67_110 ();
 sg13g2_fill_2 FILLER_67_118 ();
 sg13g2_fill_8 FILLER_67_160 ();
 sg13g2_fill_1 FILLER_67_168 ();
 sg13g2_fill_4 FILLER_67_195 ();
 sg13g2_fill_1 FILLER_67_199 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_fill_8 FILLER_67_237 ();
 sg13g2_fill_8 FILLER_67_245 ();
 sg13g2_fill_8 FILLER_67_253 ();
 sg13g2_fill_8 FILLER_67_261 ();
 sg13g2_fill_8 FILLER_67_269 ();
 sg13g2_fill_4 FILLER_67_277 ();
 sg13g2_fill_2 FILLER_67_281 ();
 sg13g2_fill_8 FILLER_67_291 ();
 sg13g2_fill_8 FILLER_67_299 ();
 sg13g2_fill_8 FILLER_67_307 ();
 sg13g2_fill_8 FILLER_67_315 ();
 sg13g2_fill_4 FILLER_67_323 ();
 sg13g2_fill_1 FILLER_67_327 ();
 sg13g2_fill_4 FILLER_67_352 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_8 FILLER_67_392 ();
 sg13g2_fill_2 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_418 ();
 sg13g2_fill_1 FILLER_67_420 ();
 sg13g2_fill_4 FILLER_67_444 ();
 sg13g2_fill_1 FILLER_67_448 ();
 sg13g2_fill_1 FILLER_67_454 ();
 sg13g2_fill_1 FILLER_67_465 ();
 sg13g2_fill_2 FILLER_67_479 ();
 sg13g2_fill_1 FILLER_67_481 ();
 sg13g2_fill_8 FILLER_67_491 ();
 sg13g2_fill_2 FILLER_67_499 ();
 sg13g2_fill_1 FILLER_67_506 ();
 sg13g2_fill_4 FILLER_67_542 ();
 sg13g2_fill_8 FILLER_67_550 ();
 sg13g2_fill_4 FILLER_67_558 ();
 sg13g2_fill_2 FILLER_67_562 ();
 sg13g2_fill_1 FILLER_67_564 ();
 sg13g2_fill_2 FILLER_67_605 ();
 sg13g2_fill_4 FILLER_67_612 ();
 sg13g2_fill_2 FILLER_67_616 ();
 sg13g2_fill_2 FILLER_67_622 ();
 sg13g2_fill_4 FILLER_67_648 ();
 sg13g2_fill_1 FILLER_67_664 ();
 sg13g2_fill_1 FILLER_67_721 ();
 sg13g2_fill_1 FILLER_67_757 ();
 sg13g2_fill_2 FILLER_67_767 ();
 sg13g2_fill_1 FILLER_67_769 ();
 sg13g2_fill_4 FILLER_67_792 ();
 sg13g2_fill_2 FILLER_67_796 ();
 sg13g2_fill_2 FILLER_67_803 ();
 sg13g2_fill_1 FILLER_67_805 ();
 sg13g2_fill_8 FILLER_67_852 ();
 sg13g2_fill_2 FILLER_67_860 ();
 sg13g2_fill_4 FILLER_67_867 ();
 sg13g2_fill_2 FILLER_67_871 ();
 sg13g2_fill_2 FILLER_67_877 ();
 sg13g2_fill_4 FILLER_67_884 ();
 sg13g2_fill_8 FILLER_67_892 ();
 sg13g2_fill_8 FILLER_67_900 ();
 sg13g2_fill_4 FILLER_67_908 ();
 sg13g2_fill_8 FILLER_67_940 ();
 sg13g2_fill_8 FILLER_67_948 ();
 sg13g2_fill_2 FILLER_67_956 ();
 sg13g2_fill_1 FILLER_67_958 ();
 sg13g2_fill_8 FILLER_67_995 ();
 sg13g2_fill_8 FILLER_67_1003 ();
 sg13g2_fill_8 FILLER_67_1011 ();
 sg13g2_fill_8 FILLER_67_1019 ();
 sg13g2_fill_8 FILLER_67_1027 ();
 sg13g2_fill_8 FILLER_67_1035 ();
 sg13g2_fill_2 FILLER_67_1043 ();
 sg13g2_fill_1 FILLER_67_1055 ();
 sg13g2_fill_8 FILLER_67_1086 ();
 sg13g2_fill_8 FILLER_67_1094 ();
 sg13g2_fill_1 FILLER_67_1102 ();
 sg13g2_fill_8 FILLER_67_1113 ();
 sg13g2_fill_2 FILLER_67_1121 ();
 sg13g2_fill_4 FILLER_67_1127 ();
 sg13g2_fill_4 FILLER_68_36 ();
 sg13g2_fill_1 FILLER_68_40 ();
 sg13g2_fill_4 FILLER_68_51 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_fill_8 FILLER_68_74 ();
 sg13g2_fill_8 FILLER_68_82 ();
 sg13g2_fill_8 FILLER_68_90 ();
 sg13g2_fill_8 FILLER_68_98 ();
 sg13g2_fill_4 FILLER_68_106 ();
 sg13g2_fill_2 FILLER_68_110 ();
 sg13g2_fill_1 FILLER_68_112 ();
 sg13g2_fill_2 FILLER_68_117 ();
 sg13g2_fill_1 FILLER_68_119 ();
 sg13g2_fill_8 FILLER_68_133 ();
 sg13g2_fill_8 FILLER_68_141 ();
 sg13g2_fill_8 FILLER_68_149 ();
 sg13g2_fill_2 FILLER_68_157 ();
 sg13g2_fill_8 FILLER_68_169 ();
 sg13g2_fill_8 FILLER_68_177 ();
 sg13g2_fill_4 FILLER_68_185 ();
 sg13g2_fill_2 FILLER_68_202 ();
 sg13g2_fill_1 FILLER_68_214 ();
 sg13g2_fill_8 FILLER_68_232 ();
 sg13g2_fill_8 FILLER_68_240 ();
 sg13g2_fill_4 FILLER_68_258 ();
 sg13g2_fill_8 FILLER_68_302 ();
 sg13g2_fill_2 FILLER_68_310 ();
 sg13g2_fill_8 FILLER_68_316 ();
 sg13g2_fill_4 FILLER_68_324 ();
 sg13g2_fill_2 FILLER_68_328 ();
 sg13g2_fill_1 FILLER_68_330 ();
 sg13g2_fill_8 FILLER_68_340 ();
 sg13g2_fill_8 FILLER_68_348 ();
 sg13g2_fill_8 FILLER_68_356 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_fill_2 FILLER_68_408 ();
 sg13g2_fill_1 FILLER_68_427 ();
 sg13g2_fill_4 FILLER_68_493 ();
 sg13g2_fill_2 FILLER_68_497 ();
 sg13g2_fill_2 FILLER_68_509 ();
 sg13g2_fill_1 FILLER_68_511 ();
 sg13g2_fill_2 FILLER_68_543 ();
 sg13g2_fill_2 FILLER_68_550 ();
 sg13g2_fill_1 FILLER_68_552 ();
 sg13g2_fill_1 FILLER_68_558 ();
 sg13g2_fill_2 FILLER_68_569 ();
 sg13g2_fill_2 FILLER_68_584 ();
 sg13g2_fill_4 FILLER_68_590 ();
 sg13g2_fill_2 FILLER_68_618 ();
 sg13g2_fill_2 FILLER_68_630 ();
 sg13g2_fill_2 FILLER_68_637 ();
 sg13g2_fill_1 FILLER_68_639 ();
 sg13g2_fill_2 FILLER_68_670 ();
 sg13g2_fill_8 FILLER_68_681 ();
 sg13g2_fill_8 FILLER_68_689 ();
 sg13g2_fill_1 FILLER_68_697 ();
 sg13g2_fill_8 FILLER_68_712 ();
 sg13g2_fill_4 FILLER_68_720 ();
 sg13g2_fill_2 FILLER_68_724 ();
 sg13g2_fill_8 FILLER_68_742 ();
 sg13g2_fill_1 FILLER_68_750 ();
 sg13g2_fill_4 FILLER_68_756 ();
 sg13g2_fill_1 FILLER_68_760 ();
 sg13g2_fill_2 FILLER_68_769 ();
 sg13g2_fill_1 FILLER_68_771 ();
 sg13g2_fill_8 FILLER_68_785 ();
 sg13g2_fill_2 FILLER_68_793 ();
 sg13g2_fill_8 FILLER_68_805 ();
 sg13g2_fill_4 FILLER_68_813 ();
 sg13g2_fill_2 FILLER_68_817 ();
 sg13g2_fill_1 FILLER_68_819 ();
 sg13g2_fill_4 FILLER_68_824 ();
 sg13g2_fill_8 FILLER_68_838 ();
 sg13g2_fill_8 FILLER_68_846 ();
 sg13g2_fill_8 FILLER_68_854 ();
 sg13g2_fill_2 FILLER_68_871 ();
 sg13g2_fill_2 FILLER_68_878 ();
 sg13g2_fill_8 FILLER_68_888 ();
 sg13g2_fill_8 FILLER_68_896 ();
 sg13g2_fill_8 FILLER_68_904 ();
 sg13g2_fill_4 FILLER_68_912 ();
 sg13g2_fill_2 FILLER_68_916 ();
 sg13g2_fill_1 FILLER_68_918 ();
 sg13g2_fill_8 FILLER_68_968 ();
 sg13g2_fill_8 FILLER_68_976 ();
 sg13g2_fill_1 FILLER_68_1004 ();
 sg13g2_fill_8 FILLER_68_1009 ();
 sg13g2_fill_8 FILLER_68_1017 ();
 sg13g2_fill_2 FILLER_68_1025 ();
 sg13g2_fill_4 FILLER_68_1037 ();
 sg13g2_fill_4 FILLER_68_1045 ();
 sg13g2_fill_2 FILLER_68_1049 ();
 sg13g2_fill_1 FILLER_68_1051 ();
 sg13g2_fill_8 FILLER_68_1077 ();
 sg13g2_fill_4 FILLER_68_1099 ();
 sg13g2_fill_1 FILLER_68_1103 ();
 sg13g2_fill_8 FILLER_68_1124 ();
 sg13g2_fill_8 FILLER_68_1132 ();
 sg13g2_fill_4 FILLER_68_1140 ();
 sg13g2_fill_8 FILLER_69_0 ();
 sg13g2_fill_8 FILLER_69_8 ();
 sg13g2_fill_8 FILLER_69_16 ();
 sg13g2_fill_8 FILLER_69_24 ();
 sg13g2_fill_8 FILLER_69_32 ();
 sg13g2_fill_8 FILLER_69_40 ();
 sg13g2_fill_8 FILLER_69_48 ();
 sg13g2_fill_8 FILLER_69_56 ();
 sg13g2_fill_8 FILLER_69_64 ();
 sg13g2_fill_2 FILLER_69_72 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_8 FILLER_69_79 ();
 sg13g2_fill_8 FILLER_69_87 ();
 sg13g2_fill_1 FILLER_69_95 ();
 sg13g2_fill_8 FILLER_69_132 ();
 sg13g2_fill_8 FILLER_69_140 ();
 sg13g2_fill_8 FILLER_69_148 ();
 sg13g2_fill_1 FILLER_69_156 ();
 sg13g2_fill_4 FILLER_69_167 ();
 sg13g2_fill_2 FILLER_69_171 ();
 sg13g2_fill_8 FILLER_69_177 ();
 sg13g2_fill_1 FILLER_69_185 ();
 sg13g2_fill_2 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_193 ();
 sg13g2_fill_4 FILLER_69_202 ();
 sg13g2_fill_2 FILLER_69_216 ();
 sg13g2_fill_1 FILLER_69_302 ();
 sg13g2_fill_8 FILLER_69_338 ();
 sg13g2_fill_8 FILLER_69_372 ();
 sg13g2_fill_8 FILLER_69_380 ();
 sg13g2_fill_8 FILLER_69_388 ();
 sg13g2_fill_8 FILLER_69_396 ();
 sg13g2_fill_2 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_406 ();
 sg13g2_fill_2 FILLER_69_426 ();
 sg13g2_fill_1 FILLER_69_428 ();
 sg13g2_fill_1 FILLER_69_442 ();
 sg13g2_fill_2 FILLER_69_473 ();
 sg13g2_fill_2 FILLER_69_480 ();
 sg13g2_fill_8 FILLER_69_490 ();
 sg13g2_fill_8 FILLER_69_498 ();
 sg13g2_fill_4 FILLER_69_506 ();
 sg13g2_fill_2 FILLER_69_510 ();
 sg13g2_fill_2 FILLER_69_518 ();
 sg13g2_fill_2 FILLER_69_550 ();
 sg13g2_fill_1 FILLER_69_552 ();
 sg13g2_fill_8 FILLER_69_572 ();
 sg13g2_fill_8 FILLER_69_580 ();
 sg13g2_fill_4 FILLER_69_588 ();
 sg13g2_fill_2 FILLER_69_592 ();
 sg13g2_fill_4 FILLER_69_598 ();
 sg13g2_fill_1 FILLER_69_602 ();
 sg13g2_fill_8 FILLER_69_608 ();
 sg13g2_fill_8 FILLER_69_616 ();
 sg13g2_fill_8 FILLER_69_629 ();
 sg13g2_fill_4 FILLER_69_637 ();
 sg13g2_fill_4 FILLER_69_646 ();
 sg13g2_fill_2 FILLER_69_650 ();
 sg13g2_fill_8 FILLER_69_661 ();
 sg13g2_fill_1 FILLER_69_669 ();
 sg13g2_fill_8 FILLER_69_674 ();
 sg13g2_fill_4 FILLER_69_682 ();
 sg13g2_fill_2 FILLER_69_686 ();
 sg13g2_fill_2 FILLER_69_696 ();
 sg13g2_fill_1 FILLER_69_698 ();
 sg13g2_fill_8 FILLER_69_704 ();
 sg13g2_fill_8 FILLER_69_716 ();
 sg13g2_fill_8 FILLER_69_724 ();
 sg13g2_fill_4 FILLER_69_732 ();
 sg13g2_fill_1 FILLER_69_736 ();
 sg13g2_fill_8 FILLER_69_742 ();
 sg13g2_fill_8 FILLER_69_750 ();
 sg13g2_fill_4 FILLER_69_758 ();
 sg13g2_fill_2 FILLER_69_762 ();
 sg13g2_fill_8 FILLER_69_782 ();
 sg13g2_fill_4 FILLER_69_790 ();
 sg13g2_fill_2 FILLER_69_794 ();
 sg13g2_fill_1 FILLER_69_809 ();
 sg13g2_fill_8 FILLER_69_815 ();
 sg13g2_fill_8 FILLER_69_840 ();
 sg13g2_fill_8 FILLER_69_848 ();
 sg13g2_fill_2 FILLER_69_868 ();
 sg13g2_fill_1 FILLER_69_884 ();
 sg13g2_fill_1 FILLER_69_889 ();
 sg13g2_fill_2 FILLER_69_930 ();
 sg13g2_fill_1 FILLER_69_932 ();
 sg13g2_fill_4 FILLER_69_943 ();
 sg13g2_fill_2 FILLER_69_947 ();
 sg13g2_fill_1 FILLER_69_949 ();
 sg13g2_fill_4 FILLER_69_954 ();
 sg13g2_fill_2 FILLER_69_968 ();
 sg13g2_fill_4 FILLER_69_978 ();
 sg13g2_fill_4 FILLER_69_992 ();
 sg13g2_fill_1 FILLER_69_996 ();
 sg13g2_fill_8 FILLER_69_1063 ();
 sg13g2_fill_2 FILLER_69_1071 ();
 sg13g2_fill_8 FILLER_69_1134 ();
 sg13g2_fill_2 FILLER_69_1142 ();
 sg13g2_fill_8 FILLER_70_0 ();
 sg13g2_fill_8 FILLER_70_18 ();
 sg13g2_fill_8 FILLER_70_26 ();
 sg13g2_fill_4 FILLER_70_48 ();
 sg13g2_fill_1 FILLER_70_52 ();
 sg13g2_fill_4 FILLER_70_63 ();
 sg13g2_fill_4 FILLER_70_93 ();
 sg13g2_fill_2 FILLER_70_97 ();
 sg13g2_fill_2 FILLER_70_109 ();
 sg13g2_fill_4 FILLER_70_115 ();
 sg13g2_fill_2 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_121 ();
 sg13g2_fill_1 FILLER_70_126 ();
 sg13g2_fill_8 FILLER_70_132 ();
 sg13g2_fill_8 FILLER_70_140 ();
 sg13g2_fill_4 FILLER_70_148 ();
 sg13g2_fill_2 FILLER_70_152 ();
 sg13g2_fill_1 FILLER_70_154 ();
 sg13g2_fill_4 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_195 ();
 sg13g2_fill_8 FILLER_70_205 ();
 sg13g2_fill_8 FILLER_70_213 ();
 sg13g2_fill_2 FILLER_70_221 ();
 sg13g2_fill_1 FILLER_70_223 ();
 sg13g2_fill_8 FILLER_70_250 ();
 sg13g2_fill_2 FILLER_70_258 ();
 sg13g2_fill_1 FILLER_70_260 ();
 sg13g2_fill_4 FILLER_70_279 ();
 sg13g2_fill_4 FILLER_70_303 ();
 sg13g2_fill_2 FILLER_70_307 ();
 sg13g2_fill_1 FILLER_70_309 ();
 sg13g2_fill_8 FILLER_70_314 ();
 sg13g2_fill_8 FILLER_70_322 ();
 sg13g2_fill_8 FILLER_70_330 ();
 sg13g2_fill_8 FILLER_70_338 ();
 sg13g2_fill_4 FILLER_70_346 ();
 sg13g2_fill_2 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_352 ();
 sg13g2_fill_8 FILLER_70_367 ();
 sg13g2_fill_8 FILLER_70_375 ();
 sg13g2_fill_8 FILLER_70_383 ();
 sg13g2_fill_8 FILLER_70_391 ();
 sg13g2_fill_8 FILLER_70_399 ();
 sg13g2_fill_8 FILLER_70_407 ();
 sg13g2_fill_4 FILLER_70_415 ();
 sg13g2_fill_1 FILLER_70_419 ();
 sg13g2_fill_4 FILLER_70_439 ();
 sg13g2_fill_2 FILLER_70_443 ();
 sg13g2_fill_8 FILLER_70_461 ();
 sg13g2_fill_4 FILLER_70_469 ();
 sg13g2_fill_2 FILLER_70_473 ();
 sg13g2_fill_8 FILLER_70_480 ();
 sg13g2_fill_8 FILLER_70_488 ();
 sg13g2_fill_8 FILLER_70_496 ();
 sg13g2_fill_8 FILLER_70_504 ();
 sg13g2_fill_8 FILLER_70_512 ();
 sg13g2_fill_8 FILLER_70_528 ();
 sg13g2_fill_8 FILLER_70_574 ();
 sg13g2_fill_8 FILLER_70_582 ();
 sg13g2_fill_1 FILLER_70_590 ();
 sg13g2_fill_4 FILLER_70_617 ();
 sg13g2_fill_8 FILLER_70_626 ();
 sg13g2_fill_1 FILLER_70_634 ();
 sg13g2_fill_8 FILLER_70_640 ();
 sg13g2_fill_8 FILLER_70_648 ();
 sg13g2_fill_2 FILLER_70_656 ();
 sg13g2_fill_4 FILLER_70_672 ();
 sg13g2_fill_2 FILLER_70_676 ();
 sg13g2_fill_1 FILLER_70_678 ();
 sg13g2_fill_8 FILLER_70_719 ();
 sg13g2_fill_2 FILLER_70_727 ();
 sg13g2_fill_1 FILLER_70_729 ();
 sg13g2_fill_2 FILLER_70_735 ();
 sg13g2_fill_1 FILLER_70_737 ();
 sg13g2_fill_8 FILLER_70_743 ();
 sg13g2_fill_8 FILLER_70_755 ();
 sg13g2_fill_4 FILLER_70_763 ();
 sg13g2_fill_2 FILLER_70_767 ();
 sg13g2_fill_1 FILLER_70_769 ();
 sg13g2_fill_8 FILLER_70_774 ();
 sg13g2_fill_8 FILLER_70_782 ();
 sg13g2_fill_4 FILLER_70_790 ();
 sg13g2_fill_2 FILLER_70_794 ();
 sg13g2_fill_2 FILLER_70_823 ();
 sg13g2_fill_1 FILLER_70_825 ();
 sg13g2_fill_2 FILLER_70_838 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_fill_4 FILLER_70_850 ();
 sg13g2_fill_1 FILLER_70_854 ();
 sg13g2_fill_1 FILLER_70_869 ();
 sg13g2_fill_1 FILLER_70_879 ();
 sg13g2_fill_1 FILLER_70_906 ();
 sg13g2_fill_2 FILLER_70_1021 ();
 sg13g2_fill_8 FILLER_70_1047 ();
 sg13g2_fill_2 FILLER_70_1055 ();
 sg13g2_fill_2 FILLER_70_1072 ();
 sg13g2_fill_8 FILLER_70_1078 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_2 ();
 sg13g2_fill_2 FILLER_71_33 ();
 sg13g2_fill_1 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_72 ();
 sg13g2_fill_8 FILLER_71_78 ();
 sg13g2_fill_4 FILLER_71_106 ();
 sg13g2_fill_2 FILLER_71_110 ();
 sg13g2_fill_1 FILLER_71_112 ();
 sg13g2_fill_2 FILLER_71_143 ();
 sg13g2_fill_1 FILLER_71_145 ();
 sg13g2_fill_8 FILLER_71_180 ();
 sg13g2_fill_2 FILLER_71_188 ();
 sg13g2_fill_1 FILLER_71_190 ();
 sg13g2_fill_4 FILLER_71_195 ();
 sg13g2_fill_2 FILLER_71_199 ();
 sg13g2_fill_4 FILLER_71_206 ();
 sg13g2_fill_2 FILLER_71_210 ();
 sg13g2_fill_1 FILLER_71_212 ();
 sg13g2_fill_8 FILLER_71_237 ();
 sg13g2_fill_8 FILLER_71_245 ();
 sg13g2_fill_8 FILLER_71_253 ();
 sg13g2_fill_1 FILLER_71_261 ();
 sg13g2_fill_8 FILLER_71_266 ();
 sg13g2_fill_8 FILLER_71_274 ();
 sg13g2_fill_8 FILLER_71_282 ();
 sg13g2_fill_1 FILLER_71_290 ();
 sg13g2_fill_1 FILLER_71_301 ();
 sg13g2_fill_8 FILLER_71_328 ();
 sg13g2_fill_2 FILLER_71_336 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_fill_1 FILLER_71_409 ();
 sg13g2_fill_2 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_2 FILLER_71_442 ();
 sg13g2_fill_2 FILLER_71_448 ();
 sg13g2_fill_1 FILLER_71_450 ();
 sg13g2_fill_8 FILLER_71_481 ();
 sg13g2_fill_4 FILLER_71_489 ();
 sg13g2_fill_1 FILLER_71_493 ();
 sg13g2_fill_1 FILLER_71_505 ();
 sg13g2_fill_8 FILLER_71_511 ();
 sg13g2_fill_2 FILLER_71_519 ();
 sg13g2_fill_1 FILLER_71_521 ();
 sg13g2_fill_8 FILLER_71_526 ();
 sg13g2_fill_8 FILLER_71_534 ();
 sg13g2_fill_4 FILLER_71_542 ();
 sg13g2_fill_2 FILLER_71_546 ();
 sg13g2_fill_4 FILLER_71_579 ();
 sg13g2_fill_2 FILLER_71_583 ();
 sg13g2_fill_4 FILLER_71_590 ();
 sg13g2_fill_8 FILLER_71_598 ();
 sg13g2_fill_2 FILLER_71_606 ();
 sg13g2_fill_1 FILLER_71_608 ();
 sg13g2_fill_2 FILLER_71_618 ();
 sg13g2_fill_8 FILLER_71_637 ();
 sg13g2_fill_8 FILLER_71_645 ();
 sg13g2_fill_1 FILLER_71_662 ();
 sg13g2_fill_8 FILLER_71_676 ();
 sg13g2_fill_8 FILLER_71_684 ();
 sg13g2_fill_8 FILLER_71_707 ();
 sg13g2_fill_1 FILLER_71_719 ();
 sg13g2_fill_2 FILLER_71_750 ();
 sg13g2_fill_1 FILLER_71_752 ();
 sg13g2_fill_4 FILLER_71_761 ();
 sg13g2_fill_1 FILLER_71_765 ();
 sg13g2_fill_1 FILLER_71_770 ();
 sg13g2_fill_8 FILLER_71_797 ();
 sg13g2_fill_8 FILLER_71_805 ();
 sg13g2_fill_8 FILLER_71_813 ();
 sg13g2_fill_8 FILLER_71_847 ();
 sg13g2_fill_4 FILLER_71_855 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_8 FILLER_71_871 ();
 sg13g2_fill_4 FILLER_71_879 ();
 sg13g2_fill_1 FILLER_71_888 ();
 sg13g2_fill_8 FILLER_71_894 ();
 sg13g2_fill_8 FILLER_71_902 ();
 sg13g2_fill_8 FILLER_71_910 ();
 sg13g2_fill_4 FILLER_71_918 ();
 sg13g2_fill_2 FILLER_71_922 ();
 sg13g2_fill_4 FILLER_71_932 ();
 sg13g2_fill_8 FILLER_71_946 ();
 sg13g2_fill_8 FILLER_71_954 ();
 sg13g2_fill_8 FILLER_71_962 ();
 sg13g2_fill_8 FILLER_71_970 ();
 sg13g2_fill_4 FILLER_71_978 ();
 sg13g2_fill_1 FILLER_71_982 ();
 sg13g2_fill_8 FILLER_71_993 ();
 sg13g2_fill_1 FILLER_71_1001 ();
 sg13g2_fill_8 FILLER_71_1006 ();
 sg13g2_fill_8 FILLER_71_1014 ();
 sg13g2_fill_4 FILLER_71_1022 ();
 sg13g2_fill_2 FILLER_71_1026 ();
 sg13g2_fill_1 FILLER_71_1028 ();
 sg13g2_fill_8 FILLER_71_1059 ();
 sg13g2_fill_4 FILLER_71_1097 ();
 sg13g2_fill_2 FILLER_71_1101 ();
 sg13g2_fill_1 FILLER_71_1103 ();
 sg13g2_fill_8 FILLER_72_0 ();
 sg13g2_fill_8 FILLER_72_18 ();
 sg13g2_fill_4 FILLER_72_26 ();
 sg13g2_fill_1 FILLER_72_30 ();
 sg13g2_fill_4 FILLER_72_92 ();
 sg13g2_fill_8 FILLER_72_106 ();
 sg13g2_fill_8 FILLER_72_118 ();
 sg13g2_fill_8 FILLER_72_126 ();
 sg13g2_fill_1 FILLER_72_134 ();
 sg13g2_fill_8 FILLER_72_157 ();
 sg13g2_fill_2 FILLER_72_165 ();
 sg13g2_fill_8 FILLER_72_175 ();
 sg13g2_fill_8 FILLER_72_213 ();
 sg13g2_fill_8 FILLER_72_221 ();
 sg13g2_fill_8 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_241 ();
 sg13g2_fill_1 FILLER_72_283 ();
 sg13g2_fill_1 FILLER_72_292 ();
 sg13g2_fill_8 FILLER_72_297 ();
 sg13g2_fill_8 FILLER_72_305 ();
 sg13g2_fill_8 FILLER_72_313 ();
 sg13g2_fill_4 FILLER_72_321 ();
 sg13g2_fill_2 FILLER_72_325 ();
 sg13g2_fill_1 FILLER_72_327 ();
 sg13g2_fill_4 FILLER_72_338 ();
 sg13g2_fill_2 FILLER_72_358 ();
 sg13g2_fill_1 FILLER_72_377 ();
 sg13g2_fill_8 FILLER_72_404 ();
 sg13g2_fill_8 FILLER_72_412 ();
 sg13g2_fill_1 FILLER_72_420 ();
 sg13g2_fill_8 FILLER_72_425 ();
 sg13g2_fill_8 FILLER_72_433 ();
 sg13g2_fill_8 FILLER_72_441 ();
 sg13g2_fill_4 FILLER_72_449 ();
 sg13g2_fill_2 FILLER_72_453 ();
 sg13g2_fill_1 FILLER_72_459 ();
 sg13g2_fill_4 FILLER_72_495 ();
 sg13g2_fill_8 FILLER_72_517 ();
 sg13g2_fill_8 FILLER_72_525 ();
 sg13g2_fill_2 FILLER_72_533 ();
 sg13g2_fill_8 FILLER_72_540 ();
 sg13g2_fill_8 FILLER_72_548 ();
 sg13g2_fill_4 FILLER_72_556 ();
 sg13g2_fill_2 FILLER_72_560 ();
 sg13g2_fill_8 FILLER_72_570 ();
 sg13g2_fill_8 FILLER_72_578 ();
 sg13g2_fill_1 FILLER_72_586 ();
 sg13g2_fill_2 FILLER_72_613 ();
 sg13g2_fill_1 FILLER_72_615 ();
 sg13g2_fill_8 FILLER_72_646 ();
 sg13g2_fill_1 FILLER_72_654 ();
 sg13g2_fill_2 FILLER_72_665 ();
 sg13g2_fill_1 FILLER_72_667 ();
 sg13g2_fill_4 FILLER_72_681 ();
 sg13g2_fill_2 FILLER_72_685 ();
 sg13g2_fill_1 FILLER_72_687 ();
 sg13g2_fill_2 FILLER_72_693 ();
 sg13g2_fill_8 FILLER_72_719 ();
 sg13g2_fill_8 FILLER_72_727 ();
 sg13g2_fill_2 FILLER_72_735 ();
 sg13g2_fill_4 FILLER_72_741 ();
 sg13g2_fill_4 FILLER_72_754 ();
 sg13g2_fill_1 FILLER_72_758 ();
 sg13g2_fill_2 FILLER_72_764 ();
 sg13g2_fill_2 FILLER_72_774 ();
 sg13g2_fill_1 FILLER_72_776 ();
 sg13g2_fill_2 FILLER_72_800 ();
 sg13g2_fill_2 FILLER_72_836 ();
 sg13g2_fill_4 FILLER_72_843 ();
 sg13g2_fill_2 FILLER_72_847 ();
 sg13g2_fill_4 FILLER_72_859 ();
 sg13g2_fill_2 FILLER_72_863 ();
 sg13g2_fill_1 FILLER_72_865 ();
 sg13g2_fill_2 FILLER_72_871 ();
 sg13g2_fill_8 FILLER_72_882 ();
 sg13g2_fill_8 FILLER_72_890 ();
 sg13g2_fill_8 FILLER_72_898 ();
 sg13g2_fill_8 FILLER_72_906 ();
 sg13g2_fill_8 FILLER_72_914 ();
 sg13g2_fill_8 FILLER_72_922 ();
 sg13g2_fill_8 FILLER_72_930 ();
 sg13g2_fill_2 FILLER_72_938 ();
 sg13g2_fill_1 FILLER_72_940 ();
 sg13g2_fill_8 FILLER_72_946 ();
 sg13g2_fill_8 FILLER_72_954 ();
 sg13g2_fill_8 FILLER_72_962 ();
 sg13g2_fill_8 FILLER_72_970 ();
 sg13g2_fill_8 FILLER_72_978 ();
 sg13g2_fill_2 FILLER_72_986 ();
 sg13g2_fill_1 FILLER_72_988 ();
 sg13g2_fill_8 FILLER_72_999 ();
 sg13g2_fill_8 FILLER_72_1007 ();
 sg13g2_fill_8 FILLER_72_1015 ();
 sg13g2_fill_8 FILLER_72_1023 ();
 sg13g2_fill_4 FILLER_72_1031 ();
 sg13g2_fill_2 FILLER_72_1035 ();
 sg13g2_fill_8 FILLER_72_1042 ();
 sg13g2_fill_8 FILLER_72_1050 ();
 sg13g2_fill_4 FILLER_72_1058 ();
 sg13g2_fill_2 FILLER_72_1062 ();
 sg13g2_fill_1 FILLER_72_1064 ();
 sg13g2_fill_8 FILLER_72_1075 ();
 sg13g2_fill_8 FILLER_72_1083 ();
 sg13g2_fill_2 FILLER_72_1091 ();
 sg13g2_fill_8 FILLER_72_1118 ();
 sg13g2_fill_8 FILLER_72_1126 ();
 sg13g2_fill_8 FILLER_72_1134 ();
 sg13g2_fill_2 FILLER_72_1142 ();
 sg13g2_fill_2 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_2 ();
 sg13g2_fill_4 FILLER_73_13 ();
 sg13g2_fill_2 FILLER_73_17 ();
 sg13g2_fill_1 FILLER_73_19 ();
 sg13g2_fill_8 FILLER_73_24 ();
 sg13g2_fill_8 FILLER_73_32 ();
 sg13g2_fill_8 FILLER_73_74 ();
 sg13g2_fill_8 FILLER_73_82 ();
 sg13g2_fill_4 FILLER_73_90 ();
 sg13g2_fill_2 FILLER_73_104 ();
 sg13g2_fill_1 FILLER_73_106 ();
 sg13g2_fill_8 FILLER_73_133 ();
 sg13g2_fill_8 FILLER_73_151 ();
 sg13g2_fill_8 FILLER_73_159 ();
 sg13g2_fill_4 FILLER_73_167 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_fill_8 FILLER_73_197 ();
 sg13g2_fill_8 FILLER_73_209 ();
 sg13g2_fill_4 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_221 ();
 sg13g2_fill_8 FILLER_73_258 ();
 sg13g2_fill_4 FILLER_73_266 ();
 sg13g2_fill_2 FILLER_73_270 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_fill_2 FILLER_73_283 ();
 sg13g2_fill_8 FILLER_73_311 ();
 sg13g2_fill_4 FILLER_73_319 ();
 sg13g2_fill_1 FILLER_73_323 ();
 sg13g2_fill_4 FILLER_73_343 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_8 FILLER_73_382 ();
 sg13g2_fill_4 FILLER_73_399 ();
 sg13g2_fill_1 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_412 ();
 sg13g2_fill_1 FILLER_73_414 ();
 sg13g2_fill_8 FILLER_73_425 ();
 sg13g2_fill_4 FILLER_73_433 ();
 sg13g2_fill_8 FILLER_73_463 ();
 sg13g2_fill_8 FILLER_73_471 ();
 sg13g2_fill_8 FILLER_73_479 ();
 sg13g2_fill_4 FILLER_73_487 ();
 sg13g2_fill_1 FILLER_73_503 ();
 sg13g2_fill_4 FILLER_73_509 ();
 sg13g2_fill_1 FILLER_73_513 ();
 sg13g2_fill_2 FILLER_73_524 ();
 sg13g2_fill_2 FILLER_73_531 ();
 sg13g2_fill_1 FILLER_73_533 ();
 sg13g2_fill_8 FILLER_73_539 ();
 sg13g2_fill_8 FILLER_73_547 ();
 sg13g2_fill_1 FILLER_73_555 ();
 sg13g2_fill_4 FILLER_73_560 ();
 sg13g2_fill_1 FILLER_73_564 ();
 sg13g2_fill_4 FILLER_73_569 ();
 sg13g2_fill_2 FILLER_73_573 ();
 sg13g2_fill_2 FILLER_73_584 ();
 sg13g2_fill_1 FILLER_73_586 ();
 sg13g2_fill_4 FILLER_73_592 ();
 sg13g2_fill_1 FILLER_73_596 ();
 sg13g2_fill_8 FILLER_73_612 ();
 sg13g2_fill_2 FILLER_73_629 ();
 sg13g2_fill_8 FILLER_73_646 ();
 sg13g2_fill_8 FILLER_73_654 ();
 sg13g2_fill_4 FILLER_73_662 ();
 sg13g2_fill_2 FILLER_73_666 ();
 sg13g2_fill_4 FILLER_73_673 ();
 sg13g2_fill_1 FILLER_73_677 ();
 sg13g2_fill_1 FILLER_73_683 ();
 sg13g2_fill_4 FILLER_73_697 ();
 sg13g2_fill_2 FILLER_73_701 ();
 sg13g2_fill_1 FILLER_73_703 ();
 sg13g2_fill_2 FILLER_73_713 ();
 sg13g2_fill_1 FILLER_73_715 ();
 sg13g2_fill_8 FILLER_73_721 ();
 sg13g2_fill_1 FILLER_73_729 ();
 sg13g2_fill_8 FILLER_73_735 ();
 sg13g2_fill_2 FILLER_73_743 ();
 sg13g2_fill_8 FILLER_73_750 ();
 sg13g2_fill_8 FILLER_73_758 ();
 sg13g2_fill_2 FILLER_73_766 ();
 sg13g2_fill_4 FILLER_73_781 ();
 sg13g2_fill_2 FILLER_73_785 ();
 sg13g2_fill_2 FILLER_73_792 ();
 sg13g2_fill_1 FILLER_73_794 ();
 sg13g2_fill_8 FILLER_73_804 ();
 sg13g2_fill_8 FILLER_73_812 ();
 sg13g2_fill_8 FILLER_73_820 ();
 sg13g2_fill_8 FILLER_73_828 ();
 sg13g2_fill_8 FILLER_73_836 ();
 sg13g2_fill_8 FILLER_73_844 ();
 sg13g2_fill_8 FILLER_73_852 ();
 sg13g2_fill_4 FILLER_73_860 ();
 sg13g2_fill_1 FILLER_73_864 ();
 sg13g2_fill_8 FILLER_73_901 ();
 sg13g2_fill_4 FILLER_73_909 ();
 sg13g2_fill_2 FILLER_73_913 ();
 sg13g2_fill_1 FILLER_73_915 ();
 sg13g2_fill_4 FILLER_73_926 ();
 sg13g2_fill_2 FILLER_73_930 ();
 sg13g2_fill_8 FILLER_73_972 ();
 sg13g2_fill_4 FILLER_73_980 ();
 sg13g2_fill_2 FILLER_73_984 ();
 sg13g2_fill_1 FILLER_73_986 ();
 sg13g2_fill_4 FILLER_73_997 ();
 sg13g2_fill_4 FILLER_73_1027 ();
 sg13g2_fill_1 FILLER_73_1031 ();
 sg13g2_fill_8 FILLER_73_1046 ();
 sg13g2_fill_8 FILLER_73_1054 ();
 sg13g2_fill_4 FILLER_73_1062 ();
 sg13g2_fill_2 FILLER_73_1066 ();
 sg13g2_fill_1 FILLER_73_1068 ();
 sg13g2_fill_2 FILLER_73_1079 ();
 sg13g2_fill_1 FILLER_73_1081 ();
 sg13g2_fill_2 FILLER_73_1111 ();
 sg13g2_fill_1 FILLER_73_1113 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_2 ();
 sg13g2_fill_2 FILLER_74_39 ();
 sg13g2_fill_1 FILLER_74_41 ();
 sg13g2_fill_1 FILLER_74_50 ();
 sg13g2_fill_8 FILLER_74_87 ();
 sg13g2_fill_2 FILLER_74_95 ();
 sg13g2_fill_1 FILLER_74_97 ();
 sg13g2_fill_8 FILLER_74_116 ();
 sg13g2_fill_2 FILLER_74_124 ();
 sg13g2_fill_4 FILLER_74_142 ();
 sg13g2_fill_1 FILLER_74_146 ();
 sg13g2_fill_8 FILLER_74_151 ();
 sg13g2_fill_8 FILLER_74_159 ();
 sg13g2_fill_2 FILLER_74_167 ();
 sg13g2_fill_1 FILLER_74_169 ();
 sg13g2_fill_2 FILLER_74_183 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_fill_4 FILLER_74_233 ();
 sg13g2_fill_2 FILLER_74_237 ();
 sg13g2_fill_1 FILLER_74_239 ();
 sg13g2_fill_8 FILLER_74_258 ();
 sg13g2_fill_8 FILLER_74_266 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_8 FILLER_74_286 ();
 sg13g2_fill_8 FILLER_74_294 ();
 sg13g2_fill_4 FILLER_74_302 ();
 sg13g2_fill_8 FILLER_74_310 ();
 sg13g2_fill_4 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_322 ();
 sg13g2_fill_1 FILLER_74_324 ();
 sg13g2_fill_4 FILLER_74_339 ();
 sg13g2_fill_8 FILLER_74_373 ();
 sg13g2_fill_4 FILLER_74_381 ();
 sg13g2_fill_2 FILLER_74_385 ();
 sg13g2_fill_1 FILLER_74_387 ();
 sg13g2_fill_4 FILLER_74_414 ();
 sg13g2_fill_8 FILLER_74_433 ();
 sg13g2_fill_8 FILLER_74_441 ();
 sg13g2_fill_8 FILLER_74_449 ();
 sg13g2_fill_8 FILLER_74_457 ();
 sg13g2_fill_8 FILLER_74_465 ();
 sg13g2_fill_8 FILLER_74_473 ();
 sg13g2_fill_2 FILLER_74_481 ();
 sg13g2_fill_8 FILLER_74_497 ();
 sg13g2_fill_8 FILLER_74_505 ();
 sg13g2_fill_2 FILLER_74_513 ();
 sg13g2_fill_2 FILLER_74_533 ();
 sg13g2_fill_8 FILLER_74_567 ();
 sg13g2_fill_4 FILLER_74_580 ();
 sg13g2_fill_2 FILLER_74_584 ();
 sg13g2_fill_1 FILLER_74_586 ();
 sg13g2_fill_1 FILLER_74_591 ();
 sg13g2_fill_8 FILLER_74_600 ();
 sg13g2_fill_2 FILLER_74_608 ();
 sg13g2_fill_4 FILLER_74_614 ();
 sg13g2_fill_1 FILLER_74_618 ();
 sg13g2_fill_4 FILLER_74_624 ();
 sg13g2_fill_1 FILLER_74_628 ();
 sg13g2_fill_4 FILLER_74_638 ();
 sg13g2_fill_4 FILLER_74_646 ();
 sg13g2_fill_4 FILLER_74_654 ();
 sg13g2_fill_1 FILLER_74_658 ();
 sg13g2_fill_4 FILLER_74_664 ();
 sg13g2_fill_1 FILLER_74_704 ();
 sg13g2_fill_2 FILLER_74_740 ();
 sg13g2_fill_1 FILLER_74_742 ();
 sg13g2_fill_1 FILLER_74_782 ();
 sg13g2_fill_4 FILLER_74_788 ();
 sg13g2_fill_2 FILLER_74_792 ();
 sg13g2_fill_4 FILLER_74_799 ();
 sg13g2_fill_8 FILLER_74_833 ();
 sg13g2_fill_4 FILLER_74_851 ();
 sg13g2_fill_1 FILLER_74_855 ();
 sg13g2_fill_1 FILLER_74_860 ();
 sg13g2_fill_2 FILLER_74_876 ();
 sg13g2_fill_1 FILLER_74_914 ();
 sg13g2_fill_2 FILLER_74_925 ();
 sg13g2_fill_8 FILLER_74_953 ();
 sg13g2_fill_4 FILLER_74_987 ();
 sg13g2_fill_2 FILLER_74_991 ();
 sg13g2_fill_1 FILLER_74_993 ();
 sg13g2_fill_2 FILLER_74_1020 ();
 sg13g2_fill_1 FILLER_74_1022 ();
 sg13g2_fill_1 FILLER_74_1063 ();
 sg13g2_fill_4 FILLER_75_0 ();
 sg13g2_fill_4 FILLER_75_40 ();
 sg13g2_fill_1 FILLER_75_44 ();
 sg13g2_fill_4 FILLER_75_84 ();
 sg13g2_fill_1 FILLER_75_88 ();
 sg13g2_fill_2 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_171 ();
 sg13g2_fill_8 FILLER_75_190 ();
 sg13g2_fill_8 FILLER_75_198 ();
 sg13g2_fill_4 FILLER_75_206 ();
 sg13g2_fill_2 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_212 ();
 sg13g2_fill_8 FILLER_75_223 ();
 sg13g2_fill_4 FILLER_75_231 ();
 sg13g2_fill_4 FILLER_75_275 ();
 sg13g2_fill_1 FILLER_75_324 ();
 sg13g2_fill_8 FILLER_75_339 ();
 sg13g2_fill_8 FILLER_75_347 ();
 sg13g2_fill_4 FILLER_75_355 ();
 sg13g2_fill_2 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_fill_8 FILLER_75_366 ();
 sg13g2_fill_8 FILLER_75_374 ();
 sg13g2_fill_8 FILLER_75_382 ();
 sg13g2_fill_1 FILLER_75_390 ();
 sg13g2_fill_4 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_445 ();
 sg13g2_fill_8 FILLER_75_472 ();
 sg13g2_fill_2 FILLER_75_480 ();
 sg13g2_fill_8 FILLER_75_500 ();
 sg13g2_fill_8 FILLER_75_508 ();
 sg13g2_fill_4 FILLER_75_516 ();
 sg13g2_fill_1 FILLER_75_520 ();
 sg13g2_fill_4 FILLER_75_536 ();
 sg13g2_fill_1 FILLER_75_540 ();
 sg13g2_fill_2 FILLER_75_549 ();
 sg13g2_fill_1 FILLER_75_561 ();
 sg13g2_fill_2 FILLER_75_566 ();
 sg13g2_fill_8 FILLER_75_573 ();
 sg13g2_fill_1 FILLER_75_596 ();
 sg13g2_fill_2 FILLER_75_607 ();
 sg13g2_fill_1 FILLER_75_609 ();
 sg13g2_fill_4 FILLER_75_620 ();
 sg13g2_fill_1 FILLER_75_624 ();
 sg13g2_fill_4 FILLER_75_629 ();
 sg13g2_fill_2 FILLER_75_633 ();
 sg13g2_fill_1 FILLER_75_644 ();
 sg13g2_fill_1 FILLER_75_650 ();
 sg13g2_fill_8 FILLER_75_660 ();
 sg13g2_fill_8 FILLER_75_668 ();
 sg13g2_fill_8 FILLER_75_676 ();
 sg13g2_fill_8 FILLER_75_692 ();
 sg13g2_fill_8 FILLER_75_700 ();
 sg13g2_fill_2 FILLER_75_708 ();
 sg13g2_fill_1 FILLER_75_710 ();
 sg13g2_fill_4 FILLER_75_720 ();
 sg13g2_fill_1 FILLER_75_724 ();
 sg13g2_fill_1 FILLER_75_729 ();
 sg13g2_fill_4 FILLER_75_734 ();
 sg13g2_fill_2 FILLER_75_738 ();
 sg13g2_fill_1 FILLER_75_740 ();
 sg13g2_fill_4 FILLER_75_745 ();
 sg13g2_fill_1 FILLER_75_749 ();
 sg13g2_fill_2 FILLER_75_759 ();
 sg13g2_fill_4 FILLER_75_776 ();
 sg13g2_fill_4 FILLER_75_793 ();
 sg13g2_fill_8 FILLER_75_806 ();
 sg13g2_fill_8 FILLER_75_814 ();
 sg13g2_fill_8 FILLER_75_822 ();
 sg13g2_fill_4 FILLER_75_830 ();
 sg13g2_fill_1 FILLER_75_834 ();
 sg13g2_fill_8 FILLER_75_839 ();
 sg13g2_fill_2 FILLER_75_847 ();
 sg13g2_fill_8 FILLER_75_893 ();
 sg13g2_fill_8 FILLER_75_901 ();
 sg13g2_fill_8 FILLER_75_945 ();
 sg13g2_fill_4 FILLER_75_953 ();
 sg13g2_fill_2 FILLER_75_957 ();
 sg13g2_fill_1 FILLER_75_959 ();
 sg13g2_fill_8 FILLER_75_970 ();
 sg13g2_fill_4 FILLER_75_978 ();
 sg13g2_fill_2 FILLER_75_982 ();
 sg13g2_fill_1 FILLER_75_984 ();
 sg13g2_fill_4 FILLER_75_995 ();
 sg13g2_fill_4 FILLER_75_1017 ();
 sg13g2_fill_8 FILLER_75_1025 ();
 sg13g2_fill_4 FILLER_75_1033 ();
 sg13g2_fill_2 FILLER_75_1037 ();
 sg13g2_fill_8 FILLER_75_1087 ();
 sg13g2_fill_4 FILLER_75_1095 ();
 sg13g2_fill_2 FILLER_75_1099 ();
 sg13g2_fill_1 FILLER_75_1101 ();
 sg13g2_fill_8 FILLER_75_1130 ();
 sg13g2_fill_4 FILLER_75_1138 ();
 sg13g2_fill_2 FILLER_75_1142 ();
 sg13g2_fill_4 FILLER_76_13 ();
 sg13g2_fill_1 FILLER_76_17 ();
 sg13g2_fill_8 FILLER_76_32 ();
 sg13g2_fill_8 FILLER_76_40 ();
 sg13g2_fill_2 FILLER_76_48 ();
 sg13g2_fill_1 FILLER_76_50 ();
 sg13g2_fill_1 FILLER_76_111 ();
 sg13g2_fill_8 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_150 ();
 sg13g2_fill_8 FILLER_76_192 ();
 sg13g2_fill_4 FILLER_76_200 ();
 sg13g2_fill_1 FILLER_76_204 ();
 sg13g2_fill_4 FILLER_76_215 ();
 sg13g2_fill_2 FILLER_76_219 ();
 sg13g2_fill_1 FILLER_76_221 ();
 sg13g2_fill_8 FILLER_76_226 ();
 sg13g2_fill_8 FILLER_76_234 ();
 sg13g2_fill_2 FILLER_76_242 ();
 sg13g2_fill_1 FILLER_76_244 ();
 sg13g2_fill_8 FILLER_76_259 ();
 sg13g2_fill_8 FILLER_76_267 ();
 sg13g2_fill_1 FILLER_76_275 ();
 sg13g2_fill_8 FILLER_76_312 ();
 sg13g2_fill_4 FILLER_76_320 ();
 sg13g2_fill_2 FILLER_76_324 ();
 sg13g2_fill_8 FILLER_76_340 ();
 sg13g2_fill_8 FILLER_76_348 ();
 sg13g2_fill_8 FILLER_76_356 ();
 sg13g2_fill_2 FILLER_76_364 ();
 sg13g2_fill_1 FILLER_76_366 ();
 sg13g2_fill_4 FILLER_76_393 ();
 sg13g2_fill_2 FILLER_76_397 ();
 sg13g2_fill_2 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_418 ();
 sg13g2_fill_8 FILLER_76_431 ();
 sg13g2_fill_4 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_443 ();
 sg13g2_fill_1 FILLER_76_445 ();
 sg13g2_fill_8 FILLER_76_480 ();
 sg13g2_fill_8 FILLER_76_488 ();
 sg13g2_fill_1 FILLER_76_496 ();
 sg13g2_fill_1 FILLER_76_527 ();
 sg13g2_fill_2 FILLER_76_549 ();
 sg13g2_fill_1 FILLER_76_575 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_fill_1 FILLER_76_587 ();
 sg13g2_fill_4 FILLER_76_599 ();
 sg13g2_fill_2 FILLER_76_603 ();
 sg13g2_fill_1 FILLER_76_605 ();
 sg13g2_fill_1 FILLER_76_632 ();
 sg13g2_fill_1 FILLER_76_638 ();
 sg13g2_fill_2 FILLER_76_669 ();
 sg13g2_fill_1 FILLER_76_671 ();
 sg13g2_fill_1 FILLER_76_680 ();
 sg13g2_fill_1 FILLER_76_688 ();
 sg13g2_fill_1 FILLER_76_694 ();
 sg13g2_fill_8 FILLER_76_699 ();
 sg13g2_fill_4 FILLER_76_707 ();
 sg13g2_fill_2 FILLER_76_711 ();
 sg13g2_fill_1 FILLER_76_713 ();
 sg13g2_fill_2 FILLER_76_773 ();
 sg13g2_fill_4 FILLER_76_779 ();
 sg13g2_fill_2 FILLER_76_783 ();
 sg13g2_fill_1 FILLER_76_785 ();
 sg13g2_fill_4 FILLER_76_866 ();
 sg13g2_fill_2 FILLER_76_870 ();
 sg13g2_fill_2 FILLER_76_876 ();
 sg13g2_fill_1 FILLER_76_878 ();
 sg13g2_fill_2 FILLER_76_909 ();
 sg13g2_fill_8 FILLER_76_935 ();
 sg13g2_fill_8 FILLER_76_943 ();
 sg13g2_fill_8 FILLER_76_951 ();
 sg13g2_fill_1 FILLER_76_969 ();
 sg13g2_fill_8 FILLER_76_974 ();
 sg13g2_fill_4 FILLER_76_982 ();
 sg13g2_fill_2 FILLER_76_986 ();
 sg13g2_fill_4 FILLER_76_998 ();
 sg13g2_fill_1 FILLER_76_1012 ();
 sg13g2_fill_8 FILLER_76_1039 ();
 sg13g2_fill_2 FILLER_76_1047 ();
 sg13g2_fill_8 FILLER_76_1073 ();
 sg13g2_fill_8 FILLER_76_1081 ();
 sg13g2_fill_8 FILLER_76_1089 ();
 sg13g2_fill_4 FILLER_76_1097 ();
 sg13g2_fill_2 FILLER_76_1101 ();
 sg13g2_fill_1 FILLER_76_1103 ();
 sg13g2_fill_8 FILLER_76_1114 ();
 sg13g2_fill_8 FILLER_76_1122 ();
 sg13g2_fill_8 FILLER_76_1130 ();
 sg13g2_fill_4 FILLER_76_1138 ();
 sg13g2_fill_2 FILLER_76_1142 ();
 sg13g2_fill_8 FILLER_77_0 ();
 sg13g2_fill_8 FILLER_77_18 ();
 sg13g2_fill_2 FILLER_77_26 ();
 sg13g2_fill_1 FILLER_77_28 ();
 sg13g2_fill_8 FILLER_77_37 ();
 sg13g2_fill_8 FILLER_77_45 ();
 sg13g2_fill_8 FILLER_77_53 ();
 sg13g2_fill_8 FILLER_77_61 ();
 sg13g2_fill_8 FILLER_77_69 ();
 sg13g2_fill_8 FILLER_77_77 ();
 sg13g2_fill_8 FILLER_77_85 ();
 sg13g2_fill_8 FILLER_77_93 ();
 sg13g2_fill_8 FILLER_77_106 ();
 sg13g2_fill_8 FILLER_77_114 ();
 sg13g2_fill_2 FILLER_77_122 ();
 sg13g2_fill_8 FILLER_77_137 ();
 sg13g2_fill_4 FILLER_77_145 ();
 sg13g2_fill_2 FILLER_77_149 ();
 sg13g2_fill_1 FILLER_77_151 ();
 sg13g2_fill_8 FILLER_77_162 ();
 sg13g2_fill_2 FILLER_77_170 ();
 sg13g2_fill_4 FILLER_77_182 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_2 FILLER_77_192 ();
 sg13g2_fill_4 FILLER_77_240 ();
 sg13g2_fill_2 FILLER_77_244 ();
 sg13g2_fill_2 FILLER_77_264 ();
 sg13g2_fill_8 FILLER_77_286 ();
 sg13g2_fill_2 FILLER_77_294 ();
 sg13g2_fill_8 FILLER_77_300 ();
 sg13g2_fill_8 FILLER_77_308 ();
 sg13g2_fill_8 FILLER_77_316 ();
 sg13g2_fill_8 FILLER_77_324 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_334 ();
 sg13g2_fill_2 FILLER_77_370 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_fill_8 FILLER_77_399 ();
 sg13g2_fill_8 FILLER_77_407 ();
 sg13g2_fill_1 FILLER_77_415 ();
 sg13g2_fill_8 FILLER_77_421 ();
 sg13g2_fill_4 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_77_433 ();
 sg13g2_fill_2 FILLER_77_454 ();
 sg13g2_fill_1 FILLER_77_456 ();
 sg13g2_fill_1 FILLER_77_462 ();
 sg13g2_fill_8 FILLER_77_472 ();
 sg13g2_fill_8 FILLER_77_480 ();
 sg13g2_fill_2 FILLER_77_531 ();
 sg13g2_fill_1 FILLER_77_533 ();
 sg13g2_fill_8 FILLER_77_561 ();
 sg13g2_fill_2 FILLER_77_569 ();
 sg13g2_fill_1 FILLER_77_571 ();
 sg13g2_fill_1 FILLER_77_585 ();
 sg13g2_fill_2 FILLER_77_590 ();
 sg13g2_fill_1 FILLER_77_592 ();
 sg13g2_fill_1 FILLER_77_597 ();
 sg13g2_fill_8 FILLER_77_602 ();
 sg13g2_fill_4 FILLER_77_610 ();
 sg13g2_fill_2 FILLER_77_614 ();
 sg13g2_fill_1 FILLER_77_616 ();
 sg13g2_fill_8 FILLER_77_624 ();
 sg13g2_fill_2 FILLER_77_632 ();
 sg13g2_fill_1 FILLER_77_648 ();
 sg13g2_fill_4 FILLER_77_677 ();
 sg13g2_fill_2 FILLER_77_681 ();
 sg13g2_fill_4 FILLER_77_706 ();
 sg13g2_fill_4 FILLER_77_740 ();
 sg13g2_fill_2 FILLER_77_744 ();
 sg13g2_fill_1 FILLER_77_746 ();
 sg13g2_fill_4 FILLER_77_771 ();
 sg13g2_fill_2 FILLER_77_775 ();
 sg13g2_fill_2 FILLER_77_782 ();
 sg13g2_fill_8 FILLER_77_788 ();
 sg13g2_fill_2 FILLER_77_796 ();
 sg13g2_fill_1 FILLER_77_798 ();
 sg13g2_fill_8 FILLER_77_829 ();
 sg13g2_fill_4 FILLER_77_837 ();
 sg13g2_fill_8 FILLER_77_860 ();
 sg13g2_fill_8 FILLER_77_868 ();
 sg13g2_fill_8 FILLER_77_876 ();
 sg13g2_fill_8 FILLER_77_884 ();
 sg13g2_fill_8 FILLER_77_892 ();
 sg13g2_fill_8 FILLER_77_900 ();
 sg13g2_fill_4 FILLER_77_908 ();
 sg13g2_fill_1 FILLER_77_932 ();
 sg13g2_fill_4 FILLER_77_959 ();
 sg13g2_fill_8 FILLER_77_994 ();
 sg13g2_fill_1 FILLER_77_1002 ();
 sg13g2_fill_8 FILLER_77_1006 ();
 sg13g2_fill_8 FILLER_77_1014 ();
 sg13g2_fill_8 FILLER_77_1022 ();
 sg13g2_fill_8 FILLER_77_1030 ();
 sg13g2_fill_8 FILLER_77_1038 ();
 sg13g2_fill_4 FILLER_77_1046 ();
 sg13g2_fill_2 FILLER_77_1050 ();
 sg13g2_fill_1 FILLER_77_1052 ();
 sg13g2_fill_4 FILLER_77_1073 ();
 sg13g2_fill_1 FILLER_77_1077 ();
 sg13g2_fill_8 FILLER_77_1082 ();
 sg13g2_fill_2 FILLER_77_1090 ();
 sg13g2_fill_1 FILLER_77_1092 ();
 sg13g2_fill_1 FILLER_77_1113 ();
 sg13g2_fill_8 FILLER_78_0 ();
 sg13g2_fill_4 FILLER_78_44 ();
 sg13g2_fill_8 FILLER_78_67 ();
 sg13g2_fill_8 FILLER_78_75 ();
 sg13g2_fill_8 FILLER_78_83 ();
 sg13g2_fill_4 FILLER_78_91 ();
 sg13g2_fill_2 FILLER_78_95 ();
 sg13g2_fill_1 FILLER_78_97 ();
 sg13g2_fill_8 FILLER_78_108 ();
 sg13g2_fill_2 FILLER_78_116 ();
 sg13g2_fill_1 FILLER_78_118 ();
 sg13g2_fill_8 FILLER_78_123 ();
 sg13g2_fill_8 FILLER_78_131 ();
 sg13g2_fill_2 FILLER_78_139 ();
 sg13g2_fill_1 FILLER_78_151 ();
 sg13g2_fill_8 FILLER_78_156 ();
 sg13g2_fill_4 FILLER_78_164 ();
 sg13g2_fill_2 FILLER_78_168 ();
 sg13g2_fill_8 FILLER_78_206 ();
 sg13g2_fill_1 FILLER_78_214 ();
 sg13g2_fill_8 FILLER_78_241 ();
 sg13g2_fill_2 FILLER_78_249 ();
 sg13g2_fill_8 FILLER_78_277 ();
 sg13g2_fill_8 FILLER_78_285 ();
 sg13g2_fill_8 FILLER_78_293 ();
 sg13g2_fill_8 FILLER_78_301 ();
 sg13g2_fill_4 FILLER_78_309 ();
 sg13g2_fill_2 FILLER_78_313 ();
 sg13g2_fill_2 FILLER_78_353 ();
 sg13g2_fill_1 FILLER_78_355 ();
 sg13g2_fill_8 FILLER_78_364 ();
 sg13g2_fill_8 FILLER_78_395 ();
 sg13g2_fill_8 FILLER_78_403 ();
 sg13g2_fill_8 FILLER_78_411 ();
 sg13g2_fill_4 FILLER_78_419 ();
 sg13g2_fill_4 FILLER_78_462 ();
 sg13g2_fill_2 FILLER_78_466 ();
 sg13g2_fill_8 FILLER_78_498 ();
 sg13g2_fill_8 FILLER_78_506 ();
 sg13g2_fill_8 FILLER_78_514 ();
 sg13g2_fill_8 FILLER_78_522 ();
 sg13g2_fill_2 FILLER_78_530 ();
 sg13g2_fill_1 FILLER_78_532 ();
 sg13g2_fill_2 FILLER_78_563 ();
 sg13g2_fill_1 FILLER_78_565 ();
 sg13g2_fill_2 FILLER_78_583 ();
 sg13g2_fill_2 FILLER_78_590 ();
 sg13g2_fill_1 FILLER_78_592 ();
 sg13g2_fill_1 FILLER_78_598 ();
 sg13g2_fill_2 FILLER_78_604 ();
 sg13g2_fill_1 FILLER_78_606 ();
 sg13g2_fill_8 FILLER_78_611 ();
 sg13g2_fill_4 FILLER_78_624 ();
 sg13g2_fill_2 FILLER_78_628 ();
 sg13g2_fill_8 FILLER_78_634 ();
 sg13g2_fill_4 FILLER_78_642 ();
 sg13g2_fill_2 FILLER_78_646 ();
 sg13g2_fill_1 FILLER_78_648 ();
 sg13g2_fill_2 FILLER_78_654 ();
 sg13g2_fill_4 FILLER_78_669 ();
 sg13g2_fill_2 FILLER_78_673 ();
 sg13g2_fill_4 FILLER_78_710 ();
 sg13g2_fill_2 FILLER_78_714 ();
 sg13g2_fill_1 FILLER_78_716 ();
 sg13g2_fill_8 FILLER_78_727 ();
 sg13g2_fill_8 FILLER_78_735 ();
 sg13g2_fill_2 FILLER_78_743 ();
 sg13g2_fill_1 FILLER_78_745 ();
 sg13g2_fill_2 FILLER_78_772 ();
 sg13g2_fill_1 FILLER_78_774 ();
 sg13g2_fill_8 FILLER_78_801 ();
 sg13g2_fill_8 FILLER_78_809 ();
 sg13g2_fill_8 FILLER_78_817 ();
 sg13g2_fill_8 FILLER_78_825 ();
 sg13g2_fill_8 FILLER_78_833 ();
 sg13g2_fill_8 FILLER_78_841 ();
 sg13g2_fill_2 FILLER_78_849 ();
 sg13g2_fill_1 FILLER_78_851 ();
 sg13g2_fill_8 FILLER_78_878 ();
 sg13g2_fill_8 FILLER_78_886 ();
 sg13g2_fill_8 FILLER_78_894 ();
 sg13g2_fill_8 FILLER_78_902 ();
 sg13g2_fill_8 FILLER_78_910 ();
 sg13g2_fill_2 FILLER_78_918 ();
 sg13g2_fill_1 FILLER_78_920 ();
 sg13g2_fill_8 FILLER_78_951 ();
 sg13g2_fill_1 FILLER_78_959 ();
 sg13g2_fill_8 FILLER_78_978 ();
 sg13g2_fill_4 FILLER_78_996 ();
 sg13g2_fill_2 FILLER_78_1000 ();
 sg13g2_fill_1 FILLER_78_1002 ();
 sg13g2_fill_8 FILLER_78_1007 ();
 sg13g2_fill_2 FILLER_78_1015 ();
 sg13g2_fill_8 FILLER_78_1044 ();
 sg13g2_fill_4 FILLER_78_1062 ();
 sg13g2_fill_2 FILLER_78_1066 ();
 sg13g2_fill_1 FILLER_78_1068 ();
 sg13g2_fill_4 FILLER_78_1099 ();
 sg13g2_fill_1 FILLER_78_1143 ();
 sg13g2_fill_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_18 ();
 sg13g2_fill_8 FILLER_79_81 ();
 sg13g2_fill_8 FILLER_79_89 ();
 sg13g2_fill_2 FILLER_79_97 ();
 sg13g2_fill_2 FILLER_79_109 ();
 sg13g2_fill_4 FILLER_79_141 ();
 sg13g2_fill_8 FILLER_79_171 ();
 sg13g2_fill_8 FILLER_79_179 ();
 sg13g2_fill_8 FILLER_79_187 ();
 sg13g2_fill_8 FILLER_79_195 ();
 sg13g2_fill_2 FILLER_79_203 ();
 sg13g2_fill_1 FILLER_79_205 ();
 sg13g2_fill_4 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_220 ();
 sg13g2_fill_1 FILLER_79_222 ();
 sg13g2_fill_8 FILLER_79_227 ();
 sg13g2_fill_1 FILLER_79_235 ();
 sg13g2_fill_8 FILLER_79_271 ();
 sg13g2_fill_8 FILLER_79_279 ();
 sg13g2_fill_4 FILLER_79_287 ();
 sg13g2_fill_2 FILLER_79_291 ();
 sg13g2_fill_8 FILLER_79_319 ();
 sg13g2_fill_8 FILLER_79_327 ();
 sg13g2_fill_8 FILLER_79_335 ();
 sg13g2_fill_8 FILLER_79_343 ();
 sg13g2_fill_2 FILLER_79_351 ();
 sg13g2_fill_1 FILLER_79_353 ();
 sg13g2_fill_8 FILLER_79_358 ();
 sg13g2_fill_8 FILLER_79_366 ();
 sg13g2_fill_1 FILLER_79_374 ();
 sg13g2_fill_4 FILLER_79_378 ();
 sg13g2_fill_1 FILLER_79_382 ();
 sg13g2_fill_8 FILLER_79_393 ();
 sg13g2_fill_8 FILLER_79_401 ();
 sg13g2_fill_2 FILLER_79_409 ();
 sg13g2_fill_4 FILLER_79_415 ();
 sg13g2_fill_4 FILLER_79_435 ();
 sg13g2_fill_8 FILLER_79_455 ();
 sg13g2_fill_8 FILLER_79_463 ();
 sg13g2_fill_8 FILLER_79_471 ();
 sg13g2_fill_8 FILLER_79_479 ();
 sg13g2_fill_8 FILLER_79_487 ();
 sg13g2_fill_8 FILLER_79_495 ();
 sg13g2_fill_1 FILLER_79_503 ();
 sg13g2_fill_8 FILLER_79_542 ();
 sg13g2_fill_8 FILLER_79_550 ();
 sg13g2_fill_4 FILLER_79_558 ();
 sg13g2_fill_2 FILLER_79_562 ();
 sg13g2_fill_1 FILLER_79_564 ();
 sg13g2_fill_8 FILLER_79_625 ();
 sg13g2_fill_8 FILLER_79_633 ();
 sg13g2_fill_8 FILLER_79_641 ();
 sg13g2_fill_8 FILLER_79_649 ();
 sg13g2_fill_8 FILLER_79_657 ();
 sg13g2_fill_8 FILLER_79_665 ();
 sg13g2_fill_8 FILLER_79_673 ();
 sg13g2_fill_4 FILLER_79_681 ();
 sg13g2_fill_1 FILLER_79_685 ();
 sg13g2_fill_4 FILLER_79_691 ();
 sg13g2_fill_2 FILLER_79_695 ();
 sg13g2_fill_1 FILLER_79_697 ();
 sg13g2_fill_8 FILLER_79_702 ();
 sg13g2_fill_4 FILLER_79_710 ();
 sg13g2_fill_2 FILLER_79_714 ();
 sg13g2_fill_1 FILLER_79_721 ();
 sg13g2_fill_4 FILLER_79_726 ();
 sg13g2_fill_1 FILLER_79_730 ();
 sg13g2_fill_4 FILLER_79_736 ();
 sg13g2_fill_1 FILLER_79_744 ();
 sg13g2_fill_4 FILLER_79_749 ();
 sg13g2_fill_2 FILLER_79_757 ();
 sg13g2_fill_1 FILLER_79_759 ();
 sg13g2_fill_8 FILLER_79_790 ();
 sg13g2_fill_8 FILLER_79_798 ();
 sg13g2_fill_2 FILLER_79_806 ();
 sg13g2_fill_1 FILLER_79_808 ();
 sg13g2_fill_4 FILLER_79_819 ();
 sg13g2_fill_1 FILLER_79_823 ();
 sg13g2_fill_8 FILLER_79_829 ();
 sg13g2_fill_2 FILLER_79_837 ();
 sg13g2_fill_8 FILLER_79_843 ();
 sg13g2_fill_8 FILLER_79_851 ();
 sg13g2_fill_1 FILLER_79_859 ();
 sg13g2_fill_8 FILLER_79_886 ();
 sg13g2_fill_2 FILLER_79_894 ();
 sg13g2_fill_8 FILLER_79_922 ();
 sg13g2_fill_8 FILLER_79_930 ();
 sg13g2_fill_8 FILLER_79_938 ();
 sg13g2_fill_8 FILLER_79_946 ();
 sg13g2_fill_8 FILLER_79_958 ();
 sg13g2_fill_8 FILLER_79_966 ();
 sg13g2_fill_8 FILLER_79_974 ();
 sg13g2_fill_2 FILLER_79_982 ();
 sg13g2_fill_1 FILLER_79_984 ();
 sg13g2_fill_1 FILLER_79_995 ();
 sg13g2_fill_4 FILLER_79_1022 ();
 sg13g2_fill_2 FILLER_79_1026 ();
 sg13g2_fill_2 FILLER_79_1058 ();
 sg13g2_fill_1 FILLER_79_1060 ();
 sg13g2_fill_8 FILLER_79_1091 ();
 sg13g2_fill_8 FILLER_79_1099 ();
 sg13g2_fill_8 FILLER_79_1107 ();
 sg13g2_fill_4 FILLER_79_1115 ();
 sg13g2_fill_2 FILLER_79_1119 ();
 sg13g2_fill_1 FILLER_79_1121 ();
 sg13g2_fill_1 FILLER_79_1130 ();
 sg13g2_fill_8 FILLER_80_0 ();
 sg13g2_fill_8 FILLER_80_18 ();
 sg13g2_fill_8 FILLER_80_34 ();
 sg13g2_fill_8 FILLER_80_42 ();
 sg13g2_fill_8 FILLER_80_50 ();
 sg13g2_fill_8 FILLER_80_58 ();
 sg13g2_fill_8 FILLER_80_66 ();
 sg13g2_fill_8 FILLER_80_74 ();
 sg13g2_fill_8 FILLER_80_82 ();
 sg13g2_fill_8 FILLER_80_90 ();
 sg13g2_fill_8 FILLER_80_98 ();
 sg13g2_fill_8 FILLER_80_106 ();
 sg13g2_fill_8 FILLER_80_114 ();
 sg13g2_fill_1 FILLER_80_122 ();
 sg13g2_fill_4 FILLER_80_135 ();
 sg13g2_fill_1 FILLER_80_139 ();
 sg13g2_fill_1 FILLER_80_150 ();
 sg13g2_fill_8 FILLER_80_187 ();
 sg13g2_fill_8 FILLER_80_195 ();
 sg13g2_fill_8 FILLER_80_203 ();
 sg13g2_fill_8 FILLER_80_211 ();
 sg13g2_fill_8 FILLER_80_219 ();
 sg13g2_fill_8 FILLER_80_227 ();
 sg13g2_fill_8 FILLER_80_235 ();
 sg13g2_fill_4 FILLER_80_269 ();
 sg13g2_fill_2 FILLER_80_273 ();
 sg13g2_fill_1 FILLER_80_275 ();
 sg13g2_fill_4 FILLER_80_302 ();
 sg13g2_fill_8 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_332 ();
 sg13g2_fill_1 FILLER_80_334 ();
 sg13g2_fill_2 FILLER_80_345 ();
 sg13g2_fill_8 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_381 ();
 sg13g2_fill_1 FILLER_80_383 ();
 sg13g2_fill_4 FILLER_80_394 ();
 sg13g2_fill_4 FILLER_80_428 ();
 sg13g2_fill_8 FILLER_80_437 ();
 sg13g2_fill_8 FILLER_80_449 ();
 sg13g2_fill_1 FILLER_80_457 ();
 sg13g2_fill_1 FILLER_80_463 ();
 sg13g2_fill_8 FILLER_80_503 ();
 sg13g2_fill_8 FILLER_80_511 ();
 sg13g2_fill_8 FILLER_80_519 ();
 sg13g2_fill_8 FILLER_80_527 ();
 sg13g2_fill_8 FILLER_80_535 ();
 sg13g2_fill_8 FILLER_80_543 ();
 sg13g2_fill_8 FILLER_80_551 ();
 sg13g2_fill_8 FILLER_80_559 ();
 sg13g2_fill_8 FILLER_80_567 ();
 sg13g2_fill_8 FILLER_80_575 ();
 sg13g2_fill_2 FILLER_80_583 ();
 sg13g2_fill_1 FILLER_80_585 ();
 sg13g2_fill_8 FILLER_80_594 ();
 sg13g2_fill_8 FILLER_80_602 ();
 sg13g2_fill_4 FILLER_80_610 ();
 sg13g2_fill_2 FILLER_80_614 ();
 sg13g2_fill_1 FILLER_80_616 ();
 sg13g2_fill_2 FILLER_80_647 ();
 sg13g2_fill_8 FILLER_80_675 ();
 sg13g2_fill_4 FILLER_80_683 ();
 sg13g2_fill_1 FILLER_80_687 ();
 sg13g2_fill_8 FILLER_80_718 ();
 sg13g2_fill_4 FILLER_80_726 ();
 sg13g2_fill_1 FILLER_80_730 ();
 sg13g2_fill_8 FILLER_80_761 ();
 sg13g2_fill_8 FILLER_80_769 ();
 sg13g2_fill_8 FILLER_80_777 ();
 sg13g2_fill_8 FILLER_80_785 ();
 sg13g2_fill_8 FILLER_80_793 ();
 sg13g2_fill_2 FILLER_80_801 ();
 sg13g2_fill_2 FILLER_80_815 ();
 sg13g2_fill_8 FILLER_80_913 ();
 sg13g2_fill_8 FILLER_80_921 ();
 sg13g2_fill_4 FILLER_80_929 ();
 sg13g2_fill_8 FILLER_80_948 ();
 sg13g2_fill_2 FILLER_80_956 ();
 sg13g2_fill_8 FILLER_80_976 ();
 sg13g2_fill_4 FILLER_80_988 ();
 sg13g2_fill_4 FILLER_80_997 ();
 sg13g2_fill_1 FILLER_80_1001 ();
 sg13g2_fill_4 FILLER_80_1012 ();
 sg13g2_fill_1 FILLER_80_1016 ();
 sg13g2_fill_4 FILLER_80_1021 ();
 sg13g2_fill_2 FILLER_80_1025 ();
 sg13g2_fill_1 FILLER_80_1027 ();
 sg13g2_fill_8 FILLER_80_1046 ();
 sg13g2_fill_8 FILLER_80_1054 ();
 sg13g2_fill_8 FILLER_80_1062 ();
 sg13g2_fill_1 FILLER_80_1074 ();
 sg13g2_fill_2 FILLER_80_1085 ();
 sg13g2_fill_8 FILLER_80_1091 ();
 sg13g2_fill_4 FILLER_80_1099 ();
 sg13g2_fill_1 FILLER_80_1103 ();
 sg13g2_fill_8 FILLER_80_1114 ();
 sg13g2_fill_1 FILLER_80_1122 ();
 sg13g2_fill_8 FILLER_80_1127 ();
 sg13g2_fill_8 FILLER_80_1135 ();
 sg13g2_fill_1 FILLER_80_1143 ();
 sg13g2_fill_8 FILLER_81_0 ();
 sg13g2_fill_8 FILLER_81_8 ();
 sg13g2_fill_8 FILLER_81_16 ();
 sg13g2_fill_8 FILLER_81_24 ();
 sg13g2_fill_8 FILLER_81_32 ();
 sg13g2_fill_8 FILLER_81_40 ();
 sg13g2_fill_8 FILLER_81_48 ();
 sg13g2_fill_8 FILLER_81_56 ();
 sg13g2_fill_8 FILLER_81_64 ();
 sg13g2_fill_8 FILLER_81_72 ();
 sg13g2_fill_8 FILLER_81_80 ();
 sg13g2_fill_8 FILLER_81_88 ();
 sg13g2_fill_8 FILLER_81_96 ();
 sg13g2_fill_8 FILLER_81_104 ();
 sg13g2_fill_8 FILLER_81_112 ();
 sg13g2_fill_8 FILLER_81_120 ();
 sg13g2_fill_8 FILLER_81_128 ();
 sg13g2_fill_8 FILLER_81_136 ();
 sg13g2_fill_8 FILLER_81_144 ();
 sg13g2_fill_1 FILLER_81_152 ();
 sg13g2_fill_4 FILLER_81_163 ();
 sg13g2_fill_2 FILLER_81_167 ();
 sg13g2_fill_8 FILLER_81_173 ();
 sg13g2_fill_8 FILLER_81_181 ();
 sg13g2_fill_8 FILLER_81_189 ();
 sg13g2_fill_8 FILLER_81_197 ();
 sg13g2_fill_8 FILLER_81_205 ();
 sg13g2_fill_8 FILLER_81_213 ();
 sg13g2_fill_8 FILLER_81_221 ();
 sg13g2_fill_8 FILLER_81_229 ();
 sg13g2_fill_8 FILLER_81_237 ();
 sg13g2_fill_8 FILLER_81_245 ();
 sg13g2_fill_8 FILLER_81_253 ();
 sg13g2_fill_8 FILLER_81_287 ();
 sg13g2_fill_4 FILLER_81_295 ();
 sg13g2_fill_1 FILLER_81_325 ();
 sg13g2_fill_2 FILLER_81_348 ();
 sg13g2_fill_2 FILLER_81_355 ();
 sg13g2_fill_2 FILLER_81_362 ();
 sg13g2_fill_1 FILLER_81_369 ();
 sg13g2_fill_8 FILLER_81_382 ();
 sg13g2_fill_8 FILLER_81_431 ();
 sg13g2_fill_2 FILLER_81_439 ();
 sg13g2_fill_1 FILLER_81_446 ();
 sg13g2_fill_1 FILLER_81_472 ();
 sg13g2_fill_8 FILLER_81_519 ();
 sg13g2_fill_8 FILLER_81_527 ();
 sg13g2_fill_8 FILLER_81_535 ();
 sg13g2_fill_8 FILLER_81_543 ();
 sg13g2_fill_8 FILLER_81_551 ();
 sg13g2_fill_8 FILLER_81_559 ();
 sg13g2_fill_8 FILLER_81_567 ();
 sg13g2_fill_8 FILLER_81_575 ();
 sg13g2_fill_2 FILLER_81_583 ();
 sg13g2_fill_8 FILLER_81_589 ();
 sg13g2_fill_2 FILLER_81_597 ();
 sg13g2_fill_1 FILLER_81_599 ();
 sg13g2_fill_8 FILLER_81_630 ();
 sg13g2_fill_2 FILLER_81_638 ();
 sg13g2_fill_1 FILLER_81_640 ();
 sg13g2_fill_4 FILLER_81_679 ();
 sg13g2_fill_2 FILLER_81_683 ();
 sg13g2_fill_1 FILLER_81_685 ();
 sg13g2_fill_1 FILLER_81_716 ();
 sg13g2_fill_8 FILLER_81_747 ();
 sg13g2_fill_8 FILLER_81_755 ();
 sg13g2_fill_8 FILLER_81_763 ();
 sg13g2_fill_8 FILLER_81_771 ();
 sg13g2_fill_8 FILLER_81_779 ();
 sg13g2_fill_8 FILLER_81_787 ();
 sg13g2_fill_1 FILLER_81_795 ();
 sg13g2_fill_1 FILLER_81_827 ();
 sg13g2_fill_4 FILLER_81_841 ();
 sg13g2_fill_2 FILLER_81_845 ();
 sg13g2_fill_2 FILLER_81_851 ();
 sg13g2_fill_1 FILLER_81_853 ();
 sg13g2_fill_1 FILLER_81_875 ();
 sg13g2_fill_8 FILLER_81_920 ();
 sg13g2_fill_1 FILLER_81_964 ();
 sg13g2_fill_1 FILLER_81_975 ();
 sg13g2_fill_4 FILLER_81_1002 ();
 sg13g2_fill_2 FILLER_81_1006 ();
 sg13g2_fill_1 FILLER_81_1008 ();
 sg13g2_fill_2 FILLER_81_1035 ();
 sg13g2_fill_4 FILLER_81_1042 ();
 sg13g2_fill_8 FILLER_81_1056 ();
 sg13g2_fill_4 FILLER_81_1064 ();
 sg13g2_fill_1 FILLER_81_1068 ();
 sg13g2_fill_4 FILLER_81_1109 ();
 sg13g2_fill_1 FILLER_81_1113 ();
 sg13g2_fill_8 FILLER_82_0 ();
 sg13g2_fill_8 FILLER_82_8 ();
 sg13g2_fill_8 FILLER_82_16 ();
 sg13g2_fill_8 FILLER_82_24 ();
 sg13g2_fill_8 FILLER_82_32 ();
 sg13g2_fill_8 FILLER_82_40 ();
 sg13g2_fill_8 FILLER_82_48 ();
 sg13g2_fill_8 FILLER_82_56 ();
 sg13g2_fill_8 FILLER_82_64 ();
 sg13g2_fill_8 FILLER_82_72 ();
 sg13g2_fill_8 FILLER_82_80 ();
 sg13g2_fill_8 FILLER_82_88 ();
 sg13g2_fill_8 FILLER_82_96 ();
 sg13g2_fill_8 FILLER_82_104 ();
 sg13g2_fill_8 FILLER_82_112 ();
 sg13g2_fill_8 FILLER_82_120 ();
 sg13g2_fill_8 FILLER_82_128 ();
 sg13g2_fill_8 FILLER_82_136 ();
 sg13g2_fill_8 FILLER_82_144 ();
 sg13g2_fill_8 FILLER_82_152 ();
 sg13g2_fill_8 FILLER_82_160 ();
 sg13g2_fill_8 FILLER_82_168 ();
 sg13g2_fill_8 FILLER_82_176 ();
 sg13g2_fill_8 FILLER_82_184 ();
 sg13g2_fill_8 FILLER_82_192 ();
 sg13g2_fill_8 FILLER_82_200 ();
 sg13g2_fill_8 FILLER_82_208 ();
 sg13g2_fill_8 FILLER_82_216 ();
 sg13g2_fill_8 FILLER_82_224 ();
 sg13g2_fill_8 FILLER_82_232 ();
 sg13g2_fill_8 FILLER_82_240 ();
 sg13g2_fill_8 FILLER_82_248 ();
 sg13g2_fill_8 FILLER_82_256 ();
 sg13g2_fill_1 FILLER_82_264 ();
 sg13g2_fill_8 FILLER_82_302 ();
 sg13g2_fill_8 FILLER_82_310 ();
 sg13g2_fill_1 FILLER_82_318 ();
 sg13g2_fill_2 FILLER_82_324 ();
 sg13g2_fill_2 FILLER_82_356 ();
 sg13g2_fill_1 FILLER_82_358 ();
 sg13g2_fill_8 FILLER_82_388 ();
 sg13g2_fill_4 FILLER_82_396 ();
 sg13g2_fill_2 FILLER_82_400 ();
 sg13g2_fill_2 FILLER_82_407 ();
 sg13g2_fill_4 FILLER_82_435 ();
 sg13g2_fill_1 FILLER_82_439 ();
 sg13g2_fill_2 FILLER_82_447 ();
 sg13g2_fill_2 FILLER_82_459 ();
 sg13g2_fill_1 FILLER_82_461 ();
 sg13g2_fill_1 FILLER_82_467 ();
 sg13g2_fill_8 FILLER_82_471 ();
 sg13g2_fill_1 FILLER_82_479 ();
 sg13g2_fill_1 FILLER_82_485 ();
 sg13g2_fill_8 FILLER_82_516 ();
 sg13g2_fill_8 FILLER_82_524 ();
 sg13g2_fill_8 FILLER_82_532 ();
 sg13g2_fill_8 FILLER_82_540 ();
 sg13g2_fill_8 FILLER_82_548 ();
 sg13g2_fill_8 FILLER_82_556 ();
 sg13g2_fill_4 FILLER_82_564 ();
 sg13g2_fill_2 FILLER_82_568 ();
 sg13g2_fill_8 FILLER_82_600 ();
 sg13g2_fill_8 FILLER_82_608 ();
 sg13g2_fill_8 FILLER_82_616 ();
 sg13g2_fill_8 FILLER_82_624 ();
 sg13g2_fill_4 FILLER_82_632 ();
 sg13g2_fill_1 FILLER_82_636 ();
 sg13g2_fill_4 FILLER_82_642 ();
 sg13g2_fill_2 FILLER_82_646 ();
 sg13g2_fill_8 FILLER_82_683 ();
 sg13g2_fill_8 FILLER_82_691 ();
 sg13g2_fill_1 FILLER_82_699 ();
 sg13g2_fill_2 FILLER_82_708 ();
 sg13g2_fill_1 FILLER_82_710 ();
 sg13g2_fill_8 FILLER_82_732 ();
 sg13g2_fill_8 FILLER_82_740 ();
 sg13g2_fill_8 FILLER_82_748 ();
 sg13g2_fill_8 FILLER_82_756 ();
 sg13g2_fill_8 FILLER_82_764 ();
 sg13g2_fill_8 FILLER_82_772 ();
 sg13g2_fill_8 FILLER_82_780 ();
 sg13g2_fill_8 FILLER_82_788 ();
 sg13g2_fill_4 FILLER_82_796 ();
 sg13g2_fill_1 FILLER_82_800 ();
 sg13g2_fill_2 FILLER_82_813 ();
 sg13g2_fill_4 FILLER_82_838 ();
 sg13g2_fill_1 FILLER_82_842 ();
 sg13g2_fill_1 FILLER_82_877 ();
 sg13g2_fill_8 FILLER_82_887 ();
 sg13g2_fill_2 FILLER_82_895 ();
 sg13g2_fill_4 FILLER_82_927 ();
 sg13g2_fill_2 FILLER_82_931 ();
 sg13g2_fill_1 FILLER_82_933 ();
 sg13g2_fill_8 FILLER_82_952 ();
 sg13g2_fill_4 FILLER_82_996 ();
 sg13g2_fill_2 FILLER_82_1000 ();
 sg13g2_fill_8 FILLER_82_1012 ();
 sg13g2_fill_8 FILLER_82_1020 ();
 sg13g2_fill_8 FILLER_82_1028 ();
 sg13g2_fill_2 FILLER_82_1036 ();
 sg13g2_fill_8 FILLER_82_1078 ();
 sg13g2_fill_8 FILLER_82_1086 ();
 sg13g2_fill_8 FILLER_82_1094 ();
 sg13g2_fill_1 FILLER_82_1102 ();
 sg13g2_fill_8 FILLER_82_1130 ();
 sg13g2_fill_4 FILLER_82_1138 ();
 sg13g2_fill_2 FILLER_82_1142 ();
 sg13g2_fill_8 FILLER_83_0 ();
 sg13g2_fill_8 FILLER_83_8 ();
 sg13g2_fill_8 FILLER_83_16 ();
 sg13g2_fill_8 FILLER_83_24 ();
 sg13g2_fill_8 FILLER_83_32 ();
 sg13g2_fill_8 FILLER_83_40 ();
 sg13g2_fill_8 FILLER_83_48 ();
 sg13g2_fill_8 FILLER_83_56 ();
 sg13g2_fill_8 FILLER_83_64 ();
 sg13g2_fill_8 FILLER_83_72 ();
 sg13g2_fill_8 FILLER_83_80 ();
 sg13g2_fill_8 FILLER_83_88 ();
 sg13g2_fill_8 FILLER_83_96 ();
 sg13g2_fill_8 FILLER_83_104 ();
 sg13g2_fill_8 FILLER_83_112 ();
 sg13g2_fill_8 FILLER_83_120 ();
 sg13g2_fill_8 FILLER_83_128 ();
 sg13g2_fill_8 FILLER_83_136 ();
 sg13g2_fill_8 FILLER_83_144 ();
 sg13g2_fill_8 FILLER_83_152 ();
 sg13g2_fill_8 FILLER_83_160 ();
 sg13g2_fill_8 FILLER_83_168 ();
 sg13g2_fill_8 FILLER_83_176 ();
 sg13g2_fill_8 FILLER_83_184 ();
 sg13g2_fill_8 FILLER_83_192 ();
 sg13g2_fill_8 FILLER_83_200 ();
 sg13g2_fill_8 FILLER_83_208 ();
 sg13g2_fill_8 FILLER_83_216 ();
 sg13g2_fill_8 FILLER_83_224 ();
 sg13g2_fill_8 FILLER_83_232 ();
 sg13g2_fill_2 FILLER_83_240 ();
 sg13g2_fill_2 FILLER_83_260 ();
 sg13g2_fill_1 FILLER_83_262 ();
 sg13g2_fill_1 FILLER_83_279 ();
 sg13g2_fill_8 FILLER_83_293 ();
 sg13g2_fill_1 FILLER_83_318 ();
 sg13g2_fill_2 FILLER_83_344 ();
 sg13g2_fill_1 FILLER_83_346 ();
 sg13g2_fill_2 FILLER_83_355 ();
 sg13g2_fill_1 FILLER_83_357 ();
 sg13g2_fill_8 FILLER_83_395 ();
 sg13g2_fill_8 FILLER_83_403 ();
 sg13g2_fill_8 FILLER_83_411 ();
 sg13g2_fill_8 FILLER_83_419 ();
 sg13g2_fill_8 FILLER_83_427 ();
 sg13g2_fill_2 FILLER_83_470 ();
 sg13g2_fill_1 FILLER_83_472 ();
 sg13g2_fill_1 FILLER_83_495 ();
 sg13g2_fill_2 FILLER_83_505 ();
 sg13g2_fill_4 FILLER_83_512 ();
 sg13g2_fill_2 FILLER_83_516 ();
 sg13g2_fill_1 FILLER_83_518 ();
 sg13g2_fill_8 FILLER_83_522 ();
 sg13g2_fill_8 FILLER_83_530 ();
 sg13g2_fill_8 FILLER_83_538 ();
 sg13g2_fill_8 FILLER_83_546 ();
 sg13g2_fill_8 FILLER_83_554 ();
 sg13g2_fill_4 FILLER_83_562 ();
 sg13g2_fill_2 FILLER_83_566 ();
 sg13g2_fill_8 FILLER_83_588 ();
 sg13g2_fill_8 FILLER_83_596 ();
 sg13g2_fill_8 FILLER_83_604 ();
 sg13g2_fill_8 FILLER_83_612 ();
 sg13g2_fill_8 FILLER_83_620 ();
 sg13g2_fill_8 FILLER_83_628 ();
 sg13g2_fill_8 FILLER_83_636 ();
 sg13g2_fill_8 FILLER_83_644 ();
 sg13g2_fill_8 FILLER_83_652 ();
 sg13g2_fill_4 FILLER_83_660 ();
 sg13g2_fill_2 FILLER_83_664 ();
 sg13g2_fill_1 FILLER_83_666 ();
 sg13g2_fill_8 FILLER_83_671 ();
 sg13g2_fill_8 FILLER_83_679 ();
 sg13g2_fill_8 FILLER_83_687 ();
 sg13g2_fill_8 FILLER_83_695 ();
 sg13g2_fill_8 FILLER_83_703 ();
 sg13g2_fill_8 FILLER_83_711 ();
 sg13g2_fill_8 FILLER_83_719 ();
 sg13g2_fill_8 FILLER_83_727 ();
 sg13g2_fill_4 FILLER_83_735 ();
 sg13g2_fill_2 FILLER_83_739 ();
 sg13g2_fill_1 FILLER_83_741 ();
 sg13g2_fill_4 FILLER_83_773 ();
 sg13g2_fill_1 FILLER_83_777 ();
 sg13g2_fill_8 FILLER_83_800 ();
 sg13g2_fill_4 FILLER_83_808 ();
 sg13g2_fill_1 FILLER_83_812 ();
 sg13g2_fill_8 FILLER_83_843 ();
 sg13g2_fill_4 FILLER_83_856 ();
 sg13g2_fill_4 FILLER_83_868 ();
 sg13g2_fill_8 FILLER_83_880 ();
 sg13g2_fill_8 FILLER_83_888 ();
 sg13g2_fill_2 FILLER_83_896 ();
 sg13g2_fill_1 FILLER_83_898 ();
 sg13g2_fill_8 FILLER_83_908 ();
 sg13g2_fill_8 FILLER_83_923 ();
 sg13g2_fill_2 FILLER_83_931 ();
 sg13g2_fill_1 FILLER_83_933 ();
 sg13g2_fill_4 FILLER_83_944 ();
 sg13g2_fill_1 FILLER_83_948 ();
 sg13g2_fill_8 FILLER_83_953 ();
 sg13g2_fill_2 FILLER_83_961 ();
 sg13g2_fill_2 FILLER_83_973 ();
 sg13g2_fill_8 FILLER_83_983 ();
 sg13g2_fill_8 FILLER_83_991 ();
 sg13g2_fill_2 FILLER_83_999 ();
 sg13g2_fill_1 FILLER_83_1001 ();
 sg13g2_fill_8 FILLER_83_1012 ();
 sg13g2_fill_1 FILLER_83_1020 ();
 sg13g2_fill_8 FILLER_83_1025 ();
 sg13g2_fill_8 FILLER_83_1033 ();
 sg13g2_fill_4 FILLER_83_1041 ();
 sg13g2_fill_1 FILLER_83_1045 ();
 sg13g2_fill_1 FILLER_83_1054 ();
 sg13g2_fill_8 FILLER_83_1059 ();
 sg13g2_fill_8 FILLER_83_1067 ();
 sg13g2_fill_1 FILLER_83_1075 ();
 sg13g2_fill_8 FILLER_83_1089 ();
 sg13g2_fill_4 FILLER_83_1097 ();
 sg13g2_fill_2 FILLER_83_1101 ();
 sg13g2_fill_1 FILLER_83_1103 ();
 sg13g2_fill_8 FILLER_84_0 ();
 sg13g2_fill_8 FILLER_84_8 ();
 sg13g2_fill_8 FILLER_84_16 ();
 sg13g2_fill_8 FILLER_84_24 ();
 sg13g2_fill_8 FILLER_84_32 ();
 sg13g2_fill_8 FILLER_84_40 ();
 sg13g2_fill_8 FILLER_84_48 ();
 sg13g2_fill_8 FILLER_84_56 ();
 sg13g2_fill_8 FILLER_84_64 ();
 sg13g2_fill_8 FILLER_84_72 ();
 sg13g2_fill_8 FILLER_84_80 ();
 sg13g2_fill_8 FILLER_84_88 ();
 sg13g2_fill_8 FILLER_84_96 ();
 sg13g2_fill_8 FILLER_84_104 ();
 sg13g2_fill_8 FILLER_84_112 ();
 sg13g2_fill_8 FILLER_84_120 ();
 sg13g2_fill_8 FILLER_84_128 ();
 sg13g2_fill_8 FILLER_84_136 ();
 sg13g2_fill_8 FILLER_84_144 ();
 sg13g2_fill_8 FILLER_84_152 ();
 sg13g2_fill_8 FILLER_84_160 ();
 sg13g2_fill_8 FILLER_84_168 ();
 sg13g2_fill_8 FILLER_84_176 ();
 sg13g2_fill_8 FILLER_84_184 ();
 sg13g2_fill_8 FILLER_84_192 ();
 sg13g2_fill_8 FILLER_84_200 ();
 sg13g2_fill_8 FILLER_84_208 ();
 sg13g2_fill_8 FILLER_84_216 ();
 sg13g2_fill_8 FILLER_84_224 ();
 sg13g2_fill_8 FILLER_84_232 ();
 sg13g2_fill_8 FILLER_84_240 ();
 sg13g2_fill_8 FILLER_84_248 ();
 sg13g2_fill_8 FILLER_84_292 ();
 sg13g2_fill_8 FILLER_84_300 ();
 sg13g2_fill_8 FILLER_84_308 ();
 sg13g2_fill_2 FILLER_84_316 ();
 sg13g2_fill_8 FILLER_84_385 ();
 sg13g2_fill_4 FILLER_84_393 ();
 sg13g2_fill_2 FILLER_84_397 ();
 sg13g2_fill_1 FILLER_84_399 ();
 sg13g2_fill_8 FILLER_84_408 ();
 sg13g2_fill_8 FILLER_84_416 ();
 sg13g2_fill_4 FILLER_84_424 ();
 sg13g2_fill_2 FILLER_84_428 ();
 sg13g2_fill_1 FILLER_84_459 ();
 sg13g2_fill_2 FILLER_84_474 ();
 sg13g2_fill_2 FILLER_84_480 ();
 sg13g2_fill_2 FILLER_84_488 ();
 sg13g2_fill_1 FILLER_84_495 ();
 sg13g2_fill_8 FILLER_84_532 ();
 sg13g2_fill_8 FILLER_84_540 ();
 sg13g2_fill_8 FILLER_84_548 ();
 sg13g2_fill_8 FILLER_84_556 ();
 sg13g2_fill_8 FILLER_84_564 ();
 sg13g2_fill_8 FILLER_84_572 ();
 sg13g2_fill_8 FILLER_84_580 ();
 sg13g2_fill_8 FILLER_84_588 ();
 sg13g2_fill_8 FILLER_84_596 ();
 sg13g2_fill_8 FILLER_84_604 ();
 sg13g2_fill_8 FILLER_84_612 ();
 sg13g2_fill_8 FILLER_84_620 ();
 sg13g2_fill_8 FILLER_84_628 ();
 sg13g2_fill_8 FILLER_84_636 ();
 sg13g2_fill_8 FILLER_84_644 ();
 sg13g2_fill_8 FILLER_84_652 ();
 sg13g2_fill_8 FILLER_84_660 ();
 sg13g2_fill_8 FILLER_84_668 ();
 sg13g2_fill_8 FILLER_84_676 ();
 sg13g2_fill_8 FILLER_84_684 ();
 sg13g2_fill_8 FILLER_84_692 ();
 sg13g2_fill_8 FILLER_84_700 ();
 sg13g2_fill_8 FILLER_84_708 ();
 sg13g2_fill_8 FILLER_84_716 ();
 sg13g2_fill_8 FILLER_84_724 ();
 sg13g2_fill_8 FILLER_84_732 ();
 sg13g2_fill_8 FILLER_84_740 ();
 sg13g2_fill_2 FILLER_84_748 ();
 sg13g2_fill_4 FILLER_84_762 ();
 sg13g2_fill_2 FILLER_84_766 ();
 sg13g2_fill_1 FILLER_84_768 ();
 sg13g2_fill_2 FILLER_84_810 ();
 sg13g2_fill_1 FILLER_84_812 ();
 sg13g2_fill_8 FILLER_84_839 ();
 sg13g2_fill_8 FILLER_84_847 ();
 sg13g2_fill_4 FILLER_84_855 ();
 sg13g2_fill_4 FILLER_84_870 ();
 sg13g2_fill_8 FILLER_84_889 ();
 sg13g2_fill_1 FILLER_84_897 ();
 sg13g2_fill_8 FILLER_84_924 ();
 sg13g2_fill_8 FILLER_84_932 ();
 sg13g2_fill_1 FILLER_84_940 ();
 sg13g2_fill_8 FILLER_84_980 ();
 sg13g2_fill_8 FILLER_84_988 ();
 sg13g2_fill_4 FILLER_84_996 ();
 sg13g2_fill_1 FILLER_84_1000 ();
 sg13g2_fill_2 FILLER_84_1011 ();
 sg13g2_fill_8 FILLER_84_1039 ();
 sg13g2_fill_1 FILLER_84_1047 ();
 sg13g2_fill_1 FILLER_84_1058 ();
 sg13g2_fill_8 FILLER_84_1063 ();
 sg13g2_fill_8 FILLER_84_1071 ();
 sg13g2_fill_8 FILLER_84_1079 ();
 sg13g2_fill_8 FILLER_84_1087 ();
 sg13g2_fill_8 FILLER_84_1095 ();
 sg13g2_fill_1 FILLER_84_1103 ();
 sg13g2_fill_8 FILLER_84_1114 ();
 sg13g2_fill_1 FILLER_84_1122 ();
 sg13g2_fill_8 FILLER_84_1127 ();
 sg13g2_fill_8 FILLER_84_1135 ();
 sg13g2_fill_1 FILLER_84_1143 ();
 sg13g2_fill_8 FILLER_85_0 ();
 sg13g2_fill_8 FILLER_85_8 ();
 sg13g2_fill_8 FILLER_85_16 ();
 sg13g2_fill_8 FILLER_85_24 ();
 sg13g2_fill_8 FILLER_85_32 ();
 sg13g2_fill_8 FILLER_85_40 ();
 sg13g2_fill_8 FILLER_85_48 ();
 sg13g2_fill_8 FILLER_85_56 ();
 sg13g2_fill_8 FILLER_85_64 ();
 sg13g2_fill_8 FILLER_85_72 ();
 sg13g2_fill_8 FILLER_85_80 ();
 sg13g2_fill_8 FILLER_85_88 ();
 sg13g2_fill_8 FILLER_85_96 ();
 sg13g2_fill_8 FILLER_85_104 ();
 sg13g2_fill_8 FILLER_85_112 ();
 sg13g2_fill_8 FILLER_85_120 ();
 sg13g2_fill_8 FILLER_85_128 ();
 sg13g2_fill_8 FILLER_85_136 ();
 sg13g2_fill_8 FILLER_85_144 ();
 sg13g2_fill_8 FILLER_85_152 ();
 sg13g2_fill_8 FILLER_85_160 ();
 sg13g2_fill_8 FILLER_85_168 ();
 sg13g2_fill_8 FILLER_85_176 ();
 sg13g2_fill_8 FILLER_85_184 ();
 sg13g2_fill_8 FILLER_85_192 ();
 sg13g2_fill_8 FILLER_85_200 ();
 sg13g2_fill_8 FILLER_85_208 ();
 sg13g2_fill_8 FILLER_85_216 ();
 sg13g2_fill_8 FILLER_85_224 ();
 sg13g2_fill_8 FILLER_85_232 ();
 sg13g2_fill_8 FILLER_85_240 ();
 sg13g2_fill_8 FILLER_85_248 ();
 sg13g2_fill_8 FILLER_85_256 ();
 sg13g2_fill_8 FILLER_85_264 ();
 sg13g2_fill_4 FILLER_85_272 ();
 sg13g2_fill_1 FILLER_85_281 ();
 sg13g2_fill_4 FILLER_85_308 ();
 sg13g2_fill_1 FILLER_85_312 ();
 sg13g2_fill_2 FILLER_85_323 ();
 sg13g2_fill_2 FILLER_85_362 ();
 sg13g2_fill_1 FILLER_85_364 ();
 sg13g2_fill_8 FILLER_85_374 ();
 sg13g2_fill_4 FILLER_85_385 ();
 sg13g2_fill_2 FILLER_85_389 ();
 sg13g2_fill_8 FILLER_85_421 ();
 sg13g2_fill_4 FILLER_85_429 ();
 sg13g2_fill_2 FILLER_85_444 ();
 sg13g2_fill_8 FILLER_85_524 ();
 sg13g2_fill_8 FILLER_85_532 ();
 sg13g2_fill_8 FILLER_85_540 ();
 sg13g2_fill_2 FILLER_85_548 ();
 sg13g2_fill_1 FILLER_85_550 ();
 sg13g2_fill_8 FILLER_85_564 ();
 sg13g2_fill_8 FILLER_85_572 ();
 sg13g2_fill_8 FILLER_85_580 ();
 sg13g2_fill_8 FILLER_85_588 ();
 sg13g2_fill_8 FILLER_85_596 ();
 sg13g2_fill_8 FILLER_85_604 ();
 sg13g2_fill_8 FILLER_85_612 ();
 sg13g2_fill_8 FILLER_85_620 ();
 sg13g2_fill_8 FILLER_85_628 ();
 sg13g2_fill_8 FILLER_85_636 ();
 sg13g2_fill_8 FILLER_85_644 ();
 sg13g2_fill_8 FILLER_85_652 ();
 sg13g2_fill_8 FILLER_85_660 ();
 sg13g2_fill_8 FILLER_85_668 ();
 sg13g2_fill_8 FILLER_85_676 ();
 sg13g2_fill_8 FILLER_85_684 ();
 sg13g2_fill_8 FILLER_85_692 ();
 sg13g2_fill_8 FILLER_85_700 ();
 sg13g2_fill_8 FILLER_85_708 ();
 sg13g2_fill_8 FILLER_85_716 ();
 sg13g2_fill_4 FILLER_85_724 ();
 sg13g2_fill_1 FILLER_85_728 ();
 sg13g2_fill_4 FILLER_85_733 ();
 sg13g2_fill_2 FILLER_85_737 ();
 sg13g2_fill_1 FILLER_85_739 ();
 sg13g2_fill_4 FILLER_85_762 ();
 sg13g2_fill_2 FILLER_85_766 ();
 sg13g2_fill_1 FILLER_85_772 ();
 sg13g2_fill_8 FILLER_85_804 ();
 sg13g2_fill_4 FILLER_85_812 ();
 sg13g2_fill_2 FILLER_85_816 ();
 sg13g2_fill_8 FILLER_85_822 ();
 sg13g2_fill_8 FILLER_85_830 ();
 sg13g2_fill_8 FILLER_85_838 ();
 sg13g2_fill_8 FILLER_85_846 ();
 sg13g2_fill_8 FILLER_85_854 ();
 sg13g2_fill_1 FILLER_85_862 ();
 sg13g2_fill_4 FILLER_85_872 ();
 sg13g2_fill_8 FILLER_85_897 ();
 sg13g2_fill_4 FILLER_85_905 ();
 sg13g2_fill_1 FILLER_85_909 ();
 sg13g2_fill_8 FILLER_85_949 ();
 sg13g2_fill_2 FILLER_85_957 ();
 sg13g2_fill_1 FILLER_85_959 ();
 sg13g2_fill_2 FILLER_85_985 ();
 sg13g2_fill_8 FILLER_85_991 ();
 sg13g2_fill_2 FILLER_85_999 ();
 sg13g2_fill_1 FILLER_85_1001 ();
 sg13g2_fill_1 FILLER_85_1012 ();
 sg13g2_fill_2 FILLER_85_1039 ();
 sg13g2_fill_8 FILLER_85_1091 ();
 sg13g2_fill_4 FILLER_85_1099 ();
 sg13g2_fill_1 FILLER_85_1113 ();
 sg13g2_fill_8 FILLER_86_0 ();
 sg13g2_fill_8 FILLER_86_8 ();
 sg13g2_fill_8 FILLER_86_16 ();
 sg13g2_fill_8 FILLER_86_24 ();
 sg13g2_fill_8 FILLER_86_32 ();
 sg13g2_fill_8 FILLER_86_40 ();
 sg13g2_fill_8 FILLER_86_48 ();
 sg13g2_fill_8 FILLER_86_56 ();
 sg13g2_fill_8 FILLER_86_64 ();
 sg13g2_fill_8 FILLER_86_72 ();
 sg13g2_fill_8 FILLER_86_80 ();
 sg13g2_fill_8 FILLER_86_88 ();
 sg13g2_fill_8 FILLER_86_96 ();
 sg13g2_fill_8 FILLER_86_104 ();
 sg13g2_fill_8 FILLER_86_112 ();
 sg13g2_fill_8 FILLER_86_120 ();
 sg13g2_fill_8 FILLER_86_128 ();
 sg13g2_fill_8 FILLER_86_136 ();
 sg13g2_fill_8 FILLER_86_144 ();
 sg13g2_fill_8 FILLER_86_152 ();
 sg13g2_fill_8 FILLER_86_160 ();
 sg13g2_fill_8 FILLER_86_168 ();
 sg13g2_fill_8 FILLER_86_176 ();
 sg13g2_fill_8 FILLER_86_184 ();
 sg13g2_fill_8 FILLER_86_192 ();
 sg13g2_fill_8 FILLER_86_200 ();
 sg13g2_fill_8 FILLER_86_208 ();
 sg13g2_fill_8 FILLER_86_216 ();
 sg13g2_fill_8 FILLER_86_224 ();
 sg13g2_fill_8 FILLER_86_232 ();
 sg13g2_fill_8 FILLER_86_240 ();
 sg13g2_fill_8 FILLER_86_248 ();
 sg13g2_fill_8 FILLER_86_256 ();
 sg13g2_fill_8 FILLER_86_264 ();
 sg13g2_fill_8 FILLER_86_272 ();
 sg13g2_fill_2 FILLER_86_280 ();
 sg13g2_fill_1 FILLER_86_343 ();
 sg13g2_fill_8 FILLER_86_359 ();
 sg13g2_fill_1 FILLER_86_367 ();
 sg13g2_fill_4 FILLER_86_372 ();
 sg13g2_fill_2 FILLER_86_376 ();
 sg13g2_fill_1 FILLER_86_378 ();
 sg13g2_fill_8 FILLER_86_384 ();
 sg13g2_fill_4 FILLER_86_392 ();
 sg13g2_fill_2 FILLER_86_396 ();
 sg13g2_fill_1 FILLER_86_398 ();
 sg13g2_fill_4 FILLER_86_423 ();
 sg13g2_fill_1 FILLER_86_427 ();
 sg13g2_fill_8 FILLER_86_431 ();
 sg13g2_fill_4 FILLER_86_439 ();
 sg13g2_fill_2 FILLER_86_443 ();
 sg13g2_fill_1 FILLER_86_462 ();
 sg13g2_fill_1 FILLER_86_468 ();
 sg13g2_fill_1 FILLER_86_474 ();
 sg13g2_fill_4 FILLER_86_499 ();
 sg13g2_fill_1 FILLER_86_503 ();
 sg13g2_fill_8 FILLER_86_513 ();
 sg13g2_fill_8 FILLER_86_521 ();
 sg13g2_fill_8 FILLER_86_529 ();
 sg13g2_fill_8 FILLER_86_537 ();
 sg13g2_fill_8 FILLER_86_545 ();
 sg13g2_fill_8 FILLER_86_553 ();
 sg13g2_fill_8 FILLER_86_561 ();
 sg13g2_fill_8 FILLER_86_569 ();
 sg13g2_fill_8 FILLER_86_577 ();
 sg13g2_fill_8 FILLER_86_585 ();
 sg13g2_fill_8 FILLER_86_593 ();
 sg13g2_fill_8 FILLER_86_601 ();
 sg13g2_fill_8 FILLER_86_609 ();
 sg13g2_fill_8 FILLER_86_617 ();
 sg13g2_fill_8 FILLER_86_625 ();
 sg13g2_fill_8 FILLER_86_633 ();
 sg13g2_fill_8 FILLER_86_641 ();
 sg13g2_fill_8 FILLER_86_649 ();
 sg13g2_fill_8 FILLER_86_657 ();
 sg13g2_fill_8 FILLER_86_665 ();
 sg13g2_fill_8 FILLER_86_673 ();
 sg13g2_fill_8 FILLER_86_681 ();
 sg13g2_fill_8 FILLER_86_689 ();
 sg13g2_fill_8 FILLER_86_697 ();
 sg13g2_fill_8 FILLER_86_705 ();
 sg13g2_fill_2 FILLER_86_713 ();
 sg13g2_fill_2 FILLER_86_745 ();
 sg13g2_fill_1 FILLER_86_747 ();
 sg13g2_fill_2 FILLER_86_774 ();
 sg13g2_fill_1 FILLER_86_782 ();
 sg13g2_fill_4 FILLER_86_805 ();
 sg13g2_fill_2 FILLER_86_809 ();
 sg13g2_fill_1 FILLER_86_811 ();
 sg13g2_fill_4 FILLER_86_816 ();
 sg13g2_fill_2 FILLER_86_820 ();
 sg13g2_fill_4 FILLER_86_835 ();
 sg13g2_fill_1 FILLER_86_839 ();
 sg13g2_fill_8 FILLER_86_849 ();
 sg13g2_fill_1 FILLER_86_857 ();
 sg13g2_fill_8 FILLER_86_920 ();
 sg13g2_fill_8 FILLER_86_928 ();
 sg13g2_fill_8 FILLER_86_936 ();
 sg13g2_fill_8 FILLER_86_944 ();
 sg13g2_fill_8 FILLER_86_952 ();
 sg13g2_fill_4 FILLER_86_960 ();
 sg13g2_fill_1 FILLER_86_964 ();
 sg13g2_fill_4 FILLER_86_975 ();
 sg13g2_fill_4 FILLER_86_1015 ();
 sg13g2_fill_1 FILLER_86_1019 ();
 sg13g2_fill_8 FILLER_86_1024 ();
 sg13g2_fill_4 FILLER_86_1032 ();
 sg13g2_fill_2 FILLER_86_1036 ();
 sg13g2_fill_8 FILLER_86_1063 ();
 sg13g2_fill_4 FILLER_86_1071 ();
 sg13g2_fill_2 FILLER_86_1075 ();
 sg13g2_fill_4 FILLER_86_1117 ();
 sg13g2_fill_2 FILLER_86_1121 ();
 sg13g2_fill_8 FILLER_86_1127 ();
 sg13g2_fill_8 FILLER_86_1135 ();
 sg13g2_fill_1 FILLER_86_1143 ();
 sg13g2_fill_8 FILLER_87_0 ();
 sg13g2_fill_8 FILLER_87_8 ();
 sg13g2_fill_8 FILLER_87_16 ();
 sg13g2_fill_8 FILLER_87_24 ();
 sg13g2_fill_8 FILLER_87_32 ();
 sg13g2_fill_8 FILLER_87_40 ();
 sg13g2_fill_8 FILLER_87_48 ();
 sg13g2_fill_8 FILLER_87_56 ();
 sg13g2_fill_8 FILLER_87_64 ();
 sg13g2_fill_8 FILLER_87_72 ();
 sg13g2_fill_8 FILLER_87_80 ();
 sg13g2_fill_8 FILLER_87_88 ();
 sg13g2_fill_8 FILLER_87_96 ();
 sg13g2_fill_8 FILLER_87_104 ();
 sg13g2_fill_8 FILLER_87_112 ();
 sg13g2_fill_8 FILLER_87_120 ();
 sg13g2_fill_8 FILLER_87_128 ();
 sg13g2_fill_8 FILLER_87_136 ();
 sg13g2_fill_8 FILLER_87_144 ();
 sg13g2_fill_8 FILLER_87_152 ();
 sg13g2_fill_8 FILLER_87_160 ();
 sg13g2_fill_8 FILLER_87_168 ();
 sg13g2_fill_8 FILLER_87_176 ();
 sg13g2_fill_8 FILLER_87_184 ();
 sg13g2_fill_8 FILLER_87_192 ();
 sg13g2_fill_8 FILLER_87_200 ();
 sg13g2_fill_8 FILLER_87_208 ();
 sg13g2_fill_8 FILLER_87_216 ();
 sg13g2_fill_8 FILLER_87_224 ();
 sg13g2_fill_8 FILLER_87_232 ();
 sg13g2_fill_8 FILLER_87_240 ();
 sg13g2_fill_8 FILLER_87_248 ();
 sg13g2_fill_8 FILLER_87_256 ();
 sg13g2_fill_8 FILLER_87_264 ();
 sg13g2_fill_8 FILLER_87_272 ();
 sg13g2_fill_8 FILLER_87_280 ();
 sg13g2_fill_8 FILLER_87_288 ();
 sg13g2_fill_8 FILLER_87_296 ();
 sg13g2_fill_8 FILLER_87_304 ();
 sg13g2_fill_2 FILLER_87_312 ();
 sg13g2_fill_1 FILLER_87_314 ();
 sg13g2_fill_8 FILLER_87_345 ();
 sg13g2_fill_4 FILLER_87_371 ();
 sg13g2_fill_2 FILLER_87_375 ();
 sg13g2_fill_1 FILLER_87_377 ();
 sg13g2_fill_8 FILLER_87_382 ();
 sg13g2_fill_2 FILLER_87_390 ();
 sg13g2_fill_8 FILLER_87_432 ();
 sg13g2_fill_8 FILLER_87_440 ();
 sg13g2_fill_1 FILLER_87_448 ();
 sg13g2_fill_8 FILLER_87_456 ();
 sg13g2_fill_8 FILLER_87_464 ();
 sg13g2_fill_8 FILLER_87_480 ();
 sg13g2_fill_8 FILLER_87_488 ();
 sg13g2_fill_8 FILLER_87_496 ();
 sg13g2_fill_8 FILLER_87_504 ();
 sg13g2_fill_8 FILLER_87_512 ();
 sg13g2_fill_8 FILLER_87_520 ();
 sg13g2_fill_8 FILLER_87_528 ();
 sg13g2_fill_8 FILLER_87_536 ();
 sg13g2_fill_8 FILLER_87_544 ();
 sg13g2_fill_8 FILLER_87_552 ();
 sg13g2_fill_8 FILLER_87_560 ();
 sg13g2_fill_8 FILLER_87_568 ();
 sg13g2_fill_8 FILLER_87_576 ();
 sg13g2_fill_8 FILLER_87_584 ();
 sg13g2_fill_8 FILLER_87_592 ();
 sg13g2_fill_8 FILLER_87_600 ();
 sg13g2_fill_8 FILLER_87_608 ();
 sg13g2_fill_8 FILLER_87_616 ();
 sg13g2_fill_8 FILLER_87_624 ();
 sg13g2_fill_8 FILLER_87_632 ();
 sg13g2_fill_8 FILLER_87_640 ();
 sg13g2_fill_8 FILLER_87_648 ();
 sg13g2_fill_8 FILLER_87_656 ();
 sg13g2_fill_8 FILLER_87_664 ();
 sg13g2_fill_8 FILLER_87_672 ();
 sg13g2_fill_8 FILLER_87_680 ();
 sg13g2_fill_8 FILLER_87_688 ();
 sg13g2_fill_8 FILLER_87_696 ();
 sg13g2_fill_8 FILLER_87_704 ();
 sg13g2_fill_8 FILLER_87_712 ();
 sg13g2_fill_8 FILLER_87_720 ();
 sg13g2_fill_8 FILLER_87_728 ();
 sg13g2_fill_4 FILLER_87_736 ();
 sg13g2_fill_1 FILLER_87_740 ();
 sg13g2_fill_8 FILLER_87_796 ();
 sg13g2_fill_4 FILLER_87_804 ();
 sg13g2_fill_2 FILLER_87_808 ();
 sg13g2_fill_1 FILLER_87_810 ();
 sg13g2_fill_2 FILLER_87_852 ();
 sg13g2_fill_8 FILLER_87_897 ();
 sg13g2_fill_1 FILLER_87_905 ();
 sg13g2_fill_8 FILLER_87_932 ();
 sg13g2_fill_8 FILLER_87_940 ();
 sg13g2_fill_8 FILLER_87_948 ();
 sg13g2_fill_8 FILLER_87_956 ();
 sg13g2_fill_2 FILLER_87_964 ();
 sg13g2_fill_1 FILLER_87_966 ();
 sg13g2_fill_1 FILLER_87_977 ();
 sg13g2_fill_8 FILLER_87_1004 ();
 sg13g2_fill_8 FILLER_87_1012 ();
 sg13g2_fill_8 FILLER_87_1020 ();
 sg13g2_fill_8 FILLER_87_1028 ();
 sg13g2_fill_2 FILLER_87_1036 ();
 sg13g2_fill_8 FILLER_87_1063 ();
 sg13g2_fill_4 FILLER_87_1071 ();
 sg13g2_fill_4 FILLER_87_1089 ();
 sg13g2_fill_1 FILLER_87_1093 ();
 sg13g2_fill_8 FILLER_88_0 ();
 sg13g2_fill_8 FILLER_88_8 ();
 sg13g2_fill_8 FILLER_88_16 ();
 sg13g2_fill_8 FILLER_88_24 ();
 sg13g2_fill_8 FILLER_88_32 ();
 sg13g2_fill_8 FILLER_88_40 ();
 sg13g2_fill_8 FILLER_88_48 ();
 sg13g2_fill_8 FILLER_88_56 ();
 sg13g2_fill_8 FILLER_88_64 ();
 sg13g2_fill_8 FILLER_88_72 ();
 sg13g2_fill_8 FILLER_88_80 ();
 sg13g2_fill_8 FILLER_88_88 ();
 sg13g2_fill_8 FILLER_88_96 ();
 sg13g2_fill_8 FILLER_88_104 ();
 sg13g2_fill_8 FILLER_88_112 ();
 sg13g2_fill_8 FILLER_88_120 ();
 sg13g2_fill_8 FILLER_88_128 ();
 sg13g2_fill_8 FILLER_88_136 ();
 sg13g2_fill_8 FILLER_88_144 ();
 sg13g2_fill_8 FILLER_88_152 ();
 sg13g2_fill_8 FILLER_88_160 ();
 sg13g2_fill_8 FILLER_88_168 ();
 sg13g2_fill_8 FILLER_88_176 ();
 sg13g2_fill_8 FILLER_88_184 ();
 sg13g2_fill_8 FILLER_88_192 ();
 sg13g2_fill_8 FILLER_88_200 ();
 sg13g2_fill_8 FILLER_88_208 ();
 sg13g2_fill_8 FILLER_88_216 ();
 sg13g2_fill_8 FILLER_88_224 ();
 sg13g2_fill_8 FILLER_88_232 ();
 sg13g2_fill_8 FILLER_88_240 ();
 sg13g2_fill_8 FILLER_88_248 ();
 sg13g2_fill_8 FILLER_88_256 ();
 sg13g2_fill_8 FILLER_88_264 ();
 sg13g2_fill_8 FILLER_88_272 ();
 sg13g2_fill_8 FILLER_88_280 ();
 sg13g2_fill_8 FILLER_88_288 ();
 sg13g2_fill_8 FILLER_88_296 ();
 sg13g2_fill_8 FILLER_88_304 ();
 sg13g2_fill_8 FILLER_88_312 ();
 sg13g2_fill_8 FILLER_88_320 ();
 sg13g2_fill_8 FILLER_88_328 ();
 sg13g2_fill_8 FILLER_88_336 ();
 sg13g2_fill_4 FILLER_88_344 ();
 sg13g2_fill_8 FILLER_88_392 ();
 sg13g2_fill_8 FILLER_88_400 ();
 sg13g2_fill_4 FILLER_88_408 ();
 sg13g2_fill_8 FILLER_88_425 ();
 sg13g2_fill_8 FILLER_88_433 ();
 sg13g2_fill_4 FILLER_88_445 ();
 sg13g2_fill_1 FILLER_88_449 ();
 sg13g2_fill_8 FILLER_88_455 ();
 sg13g2_fill_8 FILLER_88_463 ();
 sg13g2_fill_8 FILLER_88_471 ();
 sg13g2_fill_8 FILLER_88_479 ();
 sg13g2_fill_8 FILLER_88_487 ();
 sg13g2_fill_8 FILLER_88_495 ();
 sg13g2_fill_8 FILLER_88_503 ();
 sg13g2_fill_8 FILLER_88_511 ();
 sg13g2_fill_8 FILLER_88_519 ();
 sg13g2_fill_8 FILLER_88_527 ();
 sg13g2_fill_8 FILLER_88_535 ();
 sg13g2_fill_8 FILLER_88_543 ();
 sg13g2_fill_8 FILLER_88_551 ();
 sg13g2_fill_8 FILLER_88_559 ();
 sg13g2_fill_8 FILLER_88_567 ();
 sg13g2_fill_8 FILLER_88_575 ();
 sg13g2_fill_8 FILLER_88_583 ();
 sg13g2_fill_8 FILLER_88_591 ();
 sg13g2_fill_8 FILLER_88_599 ();
 sg13g2_fill_8 FILLER_88_607 ();
 sg13g2_fill_8 FILLER_88_615 ();
 sg13g2_fill_8 FILLER_88_623 ();
 sg13g2_fill_8 FILLER_88_631 ();
 sg13g2_fill_8 FILLER_88_639 ();
 sg13g2_fill_8 FILLER_88_647 ();
 sg13g2_fill_8 FILLER_88_655 ();
 sg13g2_fill_8 FILLER_88_663 ();
 sg13g2_fill_8 FILLER_88_671 ();
 sg13g2_fill_8 FILLER_88_679 ();
 sg13g2_fill_8 FILLER_88_687 ();
 sg13g2_fill_8 FILLER_88_695 ();
 sg13g2_fill_8 FILLER_88_703 ();
 sg13g2_fill_8 FILLER_88_711 ();
 sg13g2_fill_4 FILLER_88_719 ();
 sg13g2_fill_2 FILLER_88_723 ();
 sg13g2_fill_8 FILLER_88_729 ();
 sg13g2_fill_8 FILLER_88_737 ();
 sg13g2_fill_2 FILLER_88_745 ();
 sg13g2_fill_1 FILLER_88_747 ();
 sg13g2_fill_4 FILLER_88_760 ();
 sg13g2_fill_2 FILLER_88_774 ();
 sg13g2_fill_8 FILLER_88_802 ();
 sg13g2_fill_2 FILLER_88_856 ();
 sg13g2_fill_1 FILLER_88_858 ();
 sg13g2_fill_4 FILLER_88_907 ();
 sg13g2_fill_8 FILLER_88_915 ();
 sg13g2_fill_1 FILLER_88_923 ();
 sg13g2_fill_8 FILLER_88_950 ();
 sg13g2_fill_8 FILLER_88_958 ();
 sg13g2_fill_8 FILLER_88_966 ();
 sg13g2_fill_8 FILLER_88_974 ();
 sg13g2_fill_4 FILLER_88_982 ();
 sg13g2_fill_8 FILLER_88_990 ();
 sg13g2_fill_8 FILLER_88_998 ();
 sg13g2_fill_8 FILLER_88_1006 ();
 sg13g2_fill_8 FILLER_88_1014 ();
 sg13g2_fill_8 FILLER_88_1022 ();
 sg13g2_fill_8 FILLER_88_1030 ();
 sg13g2_fill_8 FILLER_88_1038 ();
 sg13g2_fill_8 FILLER_88_1046 ();
 sg13g2_fill_8 FILLER_88_1054 ();
 sg13g2_fill_8 FILLER_88_1062 ();
 sg13g2_fill_8 FILLER_88_1070 ();
 sg13g2_fill_8 FILLER_88_1078 ();
 sg13g2_fill_8 FILLER_88_1086 ();
 sg13g2_fill_4 FILLER_88_1094 ();
 sg13g2_fill_8 FILLER_89_0 ();
 sg13g2_fill_8 FILLER_89_8 ();
 sg13g2_fill_8 FILLER_89_16 ();
 sg13g2_fill_8 FILLER_89_24 ();
 sg13g2_fill_8 FILLER_89_32 ();
 sg13g2_fill_8 FILLER_89_40 ();
 sg13g2_fill_8 FILLER_89_48 ();
 sg13g2_fill_8 FILLER_89_56 ();
 sg13g2_fill_8 FILLER_89_64 ();
 sg13g2_fill_8 FILLER_89_72 ();
 sg13g2_fill_8 FILLER_89_80 ();
 sg13g2_fill_8 FILLER_89_88 ();
 sg13g2_fill_8 FILLER_89_96 ();
 sg13g2_fill_8 FILLER_89_104 ();
 sg13g2_fill_8 FILLER_89_112 ();
 sg13g2_fill_8 FILLER_89_120 ();
 sg13g2_fill_8 FILLER_89_128 ();
 sg13g2_fill_8 FILLER_89_136 ();
 sg13g2_fill_8 FILLER_89_144 ();
 sg13g2_fill_8 FILLER_89_152 ();
 sg13g2_fill_8 FILLER_89_160 ();
 sg13g2_fill_8 FILLER_89_168 ();
 sg13g2_fill_8 FILLER_89_176 ();
 sg13g2_fill_8 FILLER_89_184 ();
 sg13g2_fill_8 FILLER_89_192 ();
 sg13g2_fill_8 FILLER_89_200 ();
 sg13g2_fill_8 FILLER_89_208 ();
 sg13g2_fill_8 FILLER_89_216 ();
 sg13g2_fill_8 FILLER_89_224 ();
 sg13g2_fill_8 FILLER_89_232 ();
 sg13g2_fill_8 FILLER_89_240 ();
 sg13g2_fill_8 FILLER_89_248 ();
 sg13g2_fill_8 FILLER_89_256 ();
 sg13g2_fill_8 FILLER_89_264 ();
 sg13g2_fill_8 FILLER_89_272 ();
 sg13g2_fill_8 FILLER_89_280 ();
 sg13g2_fill_8 FILLER_89_288 ();
 sg13g2_fill_8 FILLER_89_296 ();
 sg13g2_fill_8 FILLER_89_304 ();
 sg13g2_fill_8 FILLER_89_312 ();
 sg13g2_fill_4 FILLER_89_320 ();
 sg13g2_fill_1 FILLER_89_324 ();
 sg13g2_fill_8 FILLER_89_333 ();
 sg13g2_fill_8 FILLER_89_341 ();
 sg13g2_fill_4 FILLER_89_349 ();
 sg13g2_fill_1 FILLER_89_353 ();
 sg13g2_fill_4 FILLER_89_397 ();
 sg13g2_fill_2 FILLER_89_401 ();
 sg13g2_fill_1 FILLER_89_403 ();
 sg13g2_fill_8 FILLER_89_412 ();
 sg13g2_fill_8 FILLER_89_420 ();
 sg13g2_fill_4 FILLER_89_428 ();
 sg13g2_fill_1 FILLER_89_432 ();
 sg13g2_fill_2 FILLER_89_439 ();
 sg13g2_fill_8 FILLER_89_466 ();
 sg13g2_fill_8 FILLER_89_474 ();
 sg13g2_fill_8 FILLER_89_482 ();
 sg13g2_fill_8 FILLER_89_490 ();
 sg13g2_fill_8 FILLER_89_498 ();
 sg13g2_fill_8 FILLER_89_506 ();
 sg13g2_fill_8 FILLER_89_514 ();
 sg13g2_fill_8 FILLER_89_522 ();
 sg13g2_fill_8 FILLER_89_530 ();
 sg13g2_fill_8 FILLER_89_538 ();
 sg13g2_fill_8 FILLER_89_546 ();
 sg13g2_fill_8 FILLER_89_554 ();
 sg13g2_fill_8 FILLER_89_562 ();
 sg13g2_fill_8 FILLER_89_570 ();
 sg13g2_fill_8 FILLER_89_578 ();
 sg13g2_fill_8 FILLER_89_586 ();
 sg13g2_fill_8 FILLER_89_594 ();
 sg13g2_fill_8 FILLER_89_602 ();
 sg13g2_fill_8 FILLER_89_610 ();
 sg13g2_fill_8 FILLER_89_618 ();
 sg13g2_fill_8 FILLER_89_626 ();
 sg13g2_fill_8 FILLER_89_634 ();
 sg13g2_fill_8 FILLER_89_642 ();
 sg13g2_fill_8 FILLER_89_650 ();
 sg13g2_fill_8 FILLER_89_658 ();
 sg13g2_fill_8 FILLER_89_666 ();
 sg13g2_fill_8 FILLER_89_674 ();
 sg13g2_fill_8 FILLER_89_682 ();
 sg13g2_fill_4 FILLER_89_690 ();
 sg13g2_fill_2 FILLER_89_694 ();
 sg13g2_fill_1 FILLER_89_696 ();
 sg13g2_fill_8 FILLER_89_740 ();
 sg13g2_fill_8 FILLER_89_748 ();
 sg13g2_fill_8 FILLER_89_756 ();
 sg13g2_fill_1 FILLER_89_764 ();
 sg13g2_fill_8 FILLER_89_799 ();
 sg13g2_fill_8 FILLER_89_807 ();
 sg13g2_fill_8 FILLER_89_815 ();
 sg13g2_fill_1 FILLER_89_823 ();
 sg13g2_fill_8 FILLER_89_848 ();
 sg13g2_fill_4 FILLER_89_856 ();
 sg13g2_fill_2 FILLER_89_860 ();
 sg13g2_fill_2 FILLER_89_872 ();
 sg13g2_fill_8 FILLER_89_879 ();
 sg13g2_fill_8 FILLER_89_887 ();
 sg13g2_fill_8 FILLER_89_951 ();
 sg13g2_fill_8 FILLER_89_959 ();
 sg13g2_fill_8 FILLER_89_967 ();
 sg13g2_fill_8 FILLER_89_975 ();
 sg13g2_fill_8 FILLER_89_983 ();
 sg13g2_fill_8 FILLER_89_991 ();
 sg13g2_fill_8 FILLER_89_999 ();
 sg13g2_fill_8 FILLER_89_1007 ();
 sg13g2_fill_8 FILLER_89_1015 ();
 sg13g2_fill_8 FILLER_89_1023 ();
 sg13g2_fill_8 FILLER_89_1031 ();
 sg13g2_fill_8 FILLER_89_1039 ();
 sg13g2_fill_8 FILLER_89_1047 ();
 sg13g2_fill_8 FILLER_89_1055 ();
 sg13g2_fill_8 FILLER_89_1063 ();
 sg13g2_fill_8 FILLER_89_1071 ();
 sg13g2_fill_8 FILLER_89_1079 ();
 sg13g2_fill_8 FILLER_89_1087 ();
 sg13g2_fill_8 FILLER_89_1095 ();
 sg13g2_fill_1 FILLER_89_1103 ();
 sg13g2_fill_8 FILLER_89_1128 ();
 sg13g2_fill_8 FILLER_89_1136 ();
 sg13g2_fill_8 FILLER_90_0 ();
 sg13g2_fill_8 FILLER_90_8 ();
 sg13g2_fill_8 FILLER_90_16 ();
 sg13g2_fill_8 FILLER_90_24 ();
 sg13g2_fill_8 FILLER_90_32 ();
 sg13g2_fill_8 FILLER_90_40 ();
 sg13g2_fill_8 FILLER_90_48 ();
 sg13g2_fill_8 FILLER_90_56 ();
 sg13g2_fill_8 FILLER_90_64 ();
 sg13g2_fill_8 FILLER_90_72 ();
 sg13g2_fill_8 FILLER_90_80 ();
 sg13g2_fill_8 FILLER_90_88 ();
 sg13g2_fill_8 FILLER_90_96 ();
 sg13g2_fill_8 FILLER_90_104 ();
 sg13g2_fill_8 FILLER_90_112 ();
 sg13g2_fill_8 FILLER_90_120 ();
 sg13g2_fill_8 FILLER_90_128 ();
 sg13g2_fill_8 FILLER_90_136 ();
 sg13g2_fill_8 FILLER_90_144 ();
 sg13g2_fill_8 FILLER_90_152 ();
 sg13g2_fill_8 FILLER_90_160 ();
 sg13g2_fill_8 FILLER_90_168 ();
 sg13g2_fill_8 FILLER_90_176 ();
 sg13g2_fill_8 FILLER_90_184 ();
 sg13g2_fill_8 FILLER_90_192 ();
 sg13g2_fill_8 FILLER_90_200 ();
 sg13g2_fill_8 FILLER_90_208 ();
 sg13g2_fill_8 FILLER_90_216 ();
 sg13g2_fill_8 FILLER_90_224 ();
 sg13g2_fill_8 FILLER_90_232 ();
 sg13g2_fill_8 FILLER_90_240 ();
 sg13g2_fill_8 FILLER_90_248 ();
 sg13g2_fill_8 FILLER_90_256 ();
 sg13g2_fill_8 FILLER_90_264 ();
 sg13g2_fill_8 FILLER_90_272 ();
 sg13g2_fill_8 FILLER_90_280 ();
 sg13g2_fill_8 FILLER_90_288 ();
 sg13g2_fill_8 FILLER_90_296 ();
 sg13g2_fill_8 FILLER_90_304 ();
 sg13g2_fill_8 FILLER_90_312 ();
 sg13g2_fill_8 FILLER_90_320 ();
 sg13g2_fill_8 FILLER_90_328 ();
 sg13g2_fill_8 FILLER_90_336 ();
 sg13g2_fill_8 FILLER_90_344 ();
 sg13g2_fill_8 FILLER_90_352 ();
 sg13g2_fill_2 FILLER_90_360 ();
 sg13g2_fill_1 FILLER_90_362 ();
 sg13g2_fill_8 FILLER_90_387 ();
 sg13g2_fill_8 FILLER_90_395 ();
 sg13g2_fill_8 FILLER_90_403 ();
 sg13g2_fill_8 FILLER_90_476 ();
 sg13g2_fill_8 FILLER_90_484 ();
 sg13g2_fill_8 FILLER_90_492 ();
 sg13g2_fill_8 FILLER_90_500 ();
 sg13g2_fill_8 FILLER_90_508 ();
 sg13g2_fill_8 FILLER_90_516 ();
 sg13g2_fill_8 FILLER_90_524 ();
 sg13g2_fill_8 FILLER_90_532 ();
 sg13g2_fill_8 FILLER_90_540 ();
 sg13g2_fill_8 FILLER_90_548 ();
 sg13g2_fill_8 FILLER_90_556 ();
 sg13g2_fill_8 FILLER_90_564 ();
 sg13g2_fill_8 FILLER_90_572 ();
 sg13g2_fill_8 FILLER_90_580 ();
 sg13g2_fill_8 FILLER_90_588 ();
 sg13g2_fill_8 FILLER_90_596 ();
 sg13g2_fill_8 FILLER_90_604 ();
 sg13g2_fill_8 FILLER_90_612 ();
 sg13g2_fill_8 FILLER_90_620 ();
 sg13g2_fill_8 FILLER_90_628 ();
 sg13g2_fill_8 FILLER_90_636 ();
 sg13g2_fill_8 FILLER_90_644 ();
 sg13g2_fill_8 FILLER_90_652 ();
 sg13g2_fill_8 FILLER_90_660 ();
 sg13g2_fill_8 FILLER_90_668 ();
 sg13g2_fill_8 FILLER_90_676 ();
 sg13g2_fill_8 FILLER_90_684 ();
 sg13g2_fill_4 FILLER_90_692 ();
 sg13g2_fill_1 FILLER_90_696 ();
 sg13g2_fill_4 FILLER_90_746 ();
 sg13g2_fill_2 FILLER_90_780 ();
 sg13g2_fill_8 FILLER_90_792 ();
 sg13g2_fill_8 FILLER_90_800 ();
 sg13g2_fill_8 FILLER_90_808 ();
 sg13g2_fill_8 FILLER_90_816 ();
 sg13g2_fill_8 FILLER_90_824 ();
 sg13g2_fill_2 FILLER_90_832 ();
 sg13g2_fill_8 FILLER_90_838 ();
 sg13g2_fill_8 FILLER_90_846 ();
 sg13g2_fill_2 FILLER_90_854 ();
 sg13g2_fill_1 FILLER_90_856 ();
 sg13g2_fill_2 FILLER_90_860 ();
 sg13g2_fill_8 FILLER_90_872 ();
 sg13g2_fill_8 FILLER_90_880 ();
 sg13g2_fill_8 FILLER_90_888 ();
 sg13g2_fill_8 FILLER_90_896 ();
 sg13g2_fill_8 FILLER_90_904 ();
 sg13g2_fill_8 FILLER_90_912 ();
 sg13g2_fill_1 FILLER_90_920 ();
 sg13g2_fill_8 FILLER_90_935 ();
 sg13g2_fill_8 FILLER_90_943 ();
 sg13g2_fill_8 FILLER_90_951 ();
 sg13g2_fill_8 FILLER_90_959 ();
 sg13g2_fill_8 FILLER_90_980 ();
 sg13g2_fill_8 FILLER_90_988 ();
 sg13g2_fill_8 FILLER_90_996 ();
 sg13g2_fill_8 FILLER_90_1004 ();
 sg13g2_fill_8 FILLER_90_1012 ();
 sg13g2_fill_8 FILLER_90_1020 ();
 sg13g2_fill_8 FILLER_90_1028 ();
 sg13g2_fill_8 FILLER_90_1036 ();
 sg13g2_fill_8 FILLER_90_1044 ();
 sg13g2_fill_8 FILLER_90_1052 ();
 sg13g2_fill_8 FILLER_90_1060 ();
 sg13g2_fill_8 FILLER_90_1068 ();
 sg13g2_fill_8 FILLER_90_1076 ();
 sg13g2_fill_8 FILLER_90_1084 ();
 sg13g2_fill_8 FILLER_90_1092 ();
 sg13g2_fill_8 FILLER_90_1100 ();
 sg13g2_fill_8 FILLER_90_1108 ();
 sg13g2_fill_8 FILLER_90_1116 ();
 sg13g2_fill_8 FILLER_90_1124 ();
 sg13g2_fill_8 FILLER_90_1132 ();
 sg13g2_fill_4 FILLER_90_1140 ();
 sg13g2_fill_8 FILLER_91_0 ();
 sg13g2_fill_8 FILLER_91_8 ();
 sg13g2_fill_8 FILLER_91_16 ();
 sg13g2_fill_8 FILLER_91_24 ();
 sg13g2_fill_8 FILLER_91_32 ();
 sg13g2_fill_8 FILLER_91_40 ();
 sg13g2_fill_8 FILLER_91_48 ();
 sg13g2_fill_8 FILLER_91_56 ();
 sg13g2_fill_8 FILLER_91_64 ();
 sg13g2_fill_8 FILLER_91_72 ();
 sg13g2_fill_8 FILLER_91_80 ();
 sg13g2_fill_8 FILLER_91_88 ();
 sg13g2_fill_8 FILLER_91_96 ();
 sg13g2_fill_8 FILLER_91_104 ();
 sg13g2_fill_8 FILLER_91_112 ();
 sg13g2_fill_8 FILLER_91_120 ();
 sg13g2_fill_8 FILLER_91_128 ();
 sg13g2_fill_8 FILLER_91_136 ();
 sg13g2_fill_8 FILLER_91_144 ();
 sg13g2_fill_8 FILLER_91_152 ();
 sg13g2_fill_8 FILLER_91_160 ();
 sg13g2_fill_8 FILLER_91_168 ();
 sg13g2_fill_8 FILLER_91_176 ();
 sg13g2_fill_8 FILLER_91_184 ();
 sg13g2_fill_8 FILLER_91_192 ();
 sg13g2_fill_8 FILLER_91_200 ();
 sg13g2_fill_8 FILLER_91_208 ();
 sg13g2_fill_8 FILLER_91_216 ();
 sg13g2_fill_8 FILLER_91_224 ();
 sg13g2_fill_8 FILLER_91_232 ();
 sg13g2_fill_8 FILLER_91_240 ();
 sg13g2_fill_8 FILLER_91_248 ();
 sg13g2_fill_8 FILLER_91_256 ();
 sg13g2_fill_8 FILLER_91_264 ();
 sg13g2_fill_8 FILLER_91_272 ();
 sg13g2_fill_8 FILLER_91_280 ();
 sg13g2_fill_8 FILLER_91_288 ();
 sg13g2_fill_8 FILLER_91_296 ();
 sg13g2_fill_8 FILLER_91_304 ();
 sg13g2_fill_8 FILLER_91_312 ();
 sg13g2_fill_8 FILLER_91_320 ();
 sg13g2_fill_8 FILLER_91_328 ();
 sg13g2_fill_4 FILLER_91_336 ();
 sg13g2_fill_2 FILLER_91_349 ();
 sg13g2_fill_8 FILLER_91_361 ();
 sg13g2_fill_8 FILLER_91_369 ();
 sg13g2_fill_4 FILLER_91_377 ();
 sg13g2_fill_8 FILLER_91_398 ();
 sg13g2_fill_8 FILLER_91_406 ();
 sg13g2_fill_8 FILLER_91_414 ();
 sg13g2_fill_8 FILLER_91_422 ();
 sg13g2_fill_1 FILLER_91_430 ();
 sg13g2_fill_2 FILLER_91_451 ();
 sg13g2_fill_8 FILLER_91_467 ();
 sg13g2_fill_8 FILLER_91_475 ();
 sg13g2_fill_8 FILLER_91_483 ();
 sg13g2_fill_8 FILLER_91_491 ();
 sg13g2_fill_8 FILLER_91_499 ();
 sg13g2_fill_8 FILLER_91_507 ();
 sg13g2_fill_8 FILLER_91_515 ();
 sg13g2_fill_8 FILLER_91_523 ();
 sg13g2_fill_8 FILLER_91_531 ();
 sg13g2_fill_8 FILLER_91_539 ();
 sg13g2_fill_8 FILLER_91_547 ();
 sg13g2_fill_8 FILLER_91_555 ();
 sg13g2_fill_8 FILLER_91_563 ();
 sg13g2_fill_8 FILLER_91_571 ();
 sg13g2_fill_8 FILLER_91_579 ();
 sg13g2_fill_8 FILLER_91_587 ();
 sg13g2_fill_8 FILLER_91_595 ();
 sg13g2_fill_8 FILLER_91_603 ();
 sg13g2_fill_8 FILLER_91_611 ();
 sg13g2_fill_8 FILLER_91_619 ();
 sg13g2_fill_8 FILLER_91_627 ();
 sg13g2_fill_8 FILLER_91_635 ();
 sg13g2_fill_8 FILLER_91_643 ();
 sg13g2_fill_8 FILLER_91_651 ();
 sg13g2_fill_8 FILLER_91_659 ();
 sg13g2_fill_8 FILLER_91_667 ();
 sg13g2_fill_4 FILLER_91_675 ();
 sg13g2_fill_2 FILLER_91_679 ();
 sg13g2_fill_1 FILLER_91_681 ();
 sg13g2_fill_8 FILLER_91_690 ();
 sg13g2_fill_8 FILLER_91_698 ();
 sg13g2_fill_4 FILLER_91_706 ();
 sg13g2_fill_2 FILLER_91_710 ();
 sg13g2_fill_2 FILLER_91_744 ();
 sg13g2_fill_4 FILLER_91_780 ();
 sg13g2_fill_1 FILLER_91_784 ();
 sg13g2_fill_8 FILLER_91_810 ();
 sg13g2_fill_8 FILLER_91_818 ();
 sg13g2_fill_4 FILLER_91_826 ();
 sg13g2_fill_2 FILLER_91_830 ();
 sg13g2_fill_1 FILLER_91_832 ();
 sg13g2_fill_2 FILLER_91_869 ();
 sg13g2_fill_8 FILLER_91_901 ();
 sg13g2_fill_8 FILLER_91_909 ();
 sg13g2_fill_4 FILLER_91_917 ();
 sg13g2_fill_2 FILLER_91_921 ();
 sg13g2_fill_1 FILLER_91_923 ();
 sg13g2_fill_1 FILLER_91_930 ();
 sg13g2_fill_8 FILLER_91_946 ();
 sg13g2_fill_8 FILLER_91_954 ();
 sg13g2_fill_8 FILLER_91_962 ();
 sg13g2_fill_8 FILLER_91_970 ();
 sg13g2_fill_8 FILLER_91_978 ();
 sg13g2_fill_8 FILLER_91_986 ();
 sg13g2_fill_8 FILLER_91_994 ();
 sg13g2_fill_8 FILLER_91_1002 ();
 sg13g2_fill_8 FILLER_91_1010 ();
 sg13g2_fill_8 FILLER_91_1018 ();
 sg13g2_fill_8 FILLER_91_1026 ();
 sg13g2_fill_8 FILLER_91_1034 ();
 sg13g2_fill_8 FILLER_91_1042 ();
 sg13g2_fill_8 FILLER_91_1050 ();
 sg13g2_fill_8 FILLER_91_1058 ();
 sg13g2_fill_8 FILLER_91_1066 ();
 sg13g2_fill_8 FILLER_91_1074 ();
 sg13g2_fill_8 FILLER_91_1082 ();
 sg13g2_fill_8 FILLER_91_1090 ();
 sg13g2_fill_8 FILLER_91_1098 ();
 sg13g2_fill_8 FILLER_91_1106 ();
 sg13g2_fill_8 FILLER_91_1114 ();
 sg13g2_fill_8 FILLER_91_1122 ();
 sg13g2_fill_8 FILLER_91_1130 ();
 sg13g2_fill_4 FILLER_91_1138 ();
 sg13g2_fill_2 FILLER_91_1142 ();
 sg13g2_fill_8 FILLER_92_0 ();
 sg13g2_fill_8 FILLER_92_8 ();
 sg13g2_fill_8 FILLER_92_16 ();
 sg13g2_fill_8 FILLER_92_24 ();
 sg13g2_fill_8 FILLER_92_32 ();
 sg13g2_fill_8 FILLER_92_40 ();
 sg13g2_fill_8 FILLER_92_48 ();
 sg13g2_fill_8 FILLER_92_56 ();
 sg13g2_fill_8 FILLER_92_64 ();
 sg13g2_fill_8 FILLER_92_72 ();
 sg13g2_fill_8 FILLER_92_80 ();
 sg13g2_fill_8 FILLER_92_88 ();
 sg13g2_fill_8 FILLER_92_96 ();
 sg13g2_fill_8 FILLER_92_104 ();
 sg13g2_fill_8 FILLER_92_112 ();
 sg13g2_fill_8 FILLER_92_120 ();
 sg13g2_fill_8 FILLER_92_128 ();
 sg13g2_fill_8 FILLER_92_136 ();
 sg13g2_fill_8 FILLER_92_144 ();
 sg13g2_fill_8 FILLER_92_152 ();
 sg13g2_fill_8 FILLER_92_160 ();
 sg13g2_fill_8 FILLER_92_168 ();
 sg13g2_fill_8 FILLER_92_176 ();
 sg13g2_fill_8 FILLER_92_184 ();
 sg13g2_fill_8 FILLER_92_192 ();
 sg13g2_fill_8 FILLER_92_200 ();
 sg13g2_fill_8 FILLER_92_208 ();
 sg13g2_fill_8 FILLER_92_216 ();
 sg13g2_fill_8 FILLER_92_224 ();
 sg13g2_fill_8 FILLER_92_232 ();
 sg13g2_fill_8 FILLER_92_240 ();
 sg13g2_fill_8 FILLER_92_248 ();
 sg13g2_fill_8 FILLER_92_256 ();
 sg13g2_fill_4 FILLER_92_264 ();
 sg13g2_fill_1 FILLER_92_268 ();
 sg13g2_fill_8 FILLER_92_294 ();
 sg13g2_fill_8 FILLER_92_302 ();
 sg13g2_fill_8 FILLER_92_310 ();
 sg13g2_fill_8 FILLER_92_318 ();
 sg13g2_fill_1 FILLER_92_326 ();
 sg13g2_fill_4 FILLER_92_366 ();
 sg13g2_fill_4 FILLER_92_396 ();
 sg13g2_fill_1 FILLER_92_400 ();
 sg13g2_fill_8 FILLER_92_427 ();
 sg13g2_fill_1 FILLER_92_435 ();
 sg13g2_fill_2 FILLER_92_441 ();
 sg13g2_fill_1 FILLER_92_443 ();
 sg13g2_fill_8 FILLER_92_458 ();
 sg13g2_fill_8 FILLER_92_466 ();
 sg13g2_fill_8 FILLER_92_474 ();
 sg13g2_fill_8 FILLER_92_482 ();
 sg13g2_fill_8 FILLER_92_490 ();
 sg13g2_fill_8 FILLER_92_498 ();
 sg13g2_fill_8 FILLER_92_506 ();
 sg13g2_fill_8 FILLER_92_514 ();
 sg13g2_fill_8 FILLER_92_522 ();
 sg13g2_fill_8 FILLER_92_530 ();
 sg13g2_fill_8 FILLER_92_538 ();
 sg13g2_fill_8 FILLER_92_546 ();
 sg13g2_fill_8 FILLER_92_554 ();
 sg13g2_fill_8 FILLER_92_562 ();
 sg13g2_fill_8 FILLER_92_570 ();
 sg13g2_fill_8 FILLER_92_578 ();
 sg13g2_fill_8 FILLER_92_586 ();
 sg13g2_fill_8 FILLER_92_594 ();
 sg13g2_fill_8 FILLER_92_602 ();
 sg13g2_fill_8 FILLER_92_610 ();
 sg13g2_fill_8 FILLER_92_618 ();
 sg13g2_fill_8 FILLER_92_626 ();
 sg13g2_fill_8 FILLER_92_634 ();
 sg13g2_fill_8 FILLER_92_642 ();
 sg13g2_fill_8 FILLER_92_650 ();
 sg13g2_fill_8 FILLER_92_658 ();
 sg13g2_fill_8 FILLER_92_666 ();
 sg13g2_fill_8 FILLER_92_674 ();
 sg13g2_fill_8 FILLER_92_682 ();
 sg13g2_fill_8 FILLER_92_690 ();
 sg13g2_fill_8 FILLER_92_698 ();
 sg13g2_fill_8 FILLER_92_706 ();
 sg13g2_fill_2 FILLER_92_714 ();
 sg13g2_fill_1 FILLER_92_716 ();
 sg13g2_fill_1 FILLER_92_722 ();
 sg13g2_fill_2 FILLER_92_728 ();
 sg13g2_fill_1 FILLER_92_730 ();
 sg13g2_fill_8 FILLER_92_742 ();
 sg13g2_fill_8 FILLER_92_750 ();
 sg13g2_fill_8 FILLER_92_758 ();
 sg13g2_fill_8 FILLER_92_766 ();
 sg13g2_fill_4 FILLER_92_774 ();
 sg13g2_fill_1 FILLER_92_778 ();
 sg13g2_fill_2 FILLER_92_799 ();
 sg13g2_fill_1 FILLER_92_839 ();
 sg13g2_fill_4 FILLER_92_848 ();
 sg13g2_fill_8 FILLER_92_862 ();
 sg13g2_fill_1 FILLER_92_870 ();
 sg13g2_fill_4 FILLER_92_901 ();
 sg13g2_fill_1 FILLER_92_905 ();
 sg13g2_fill_8 FILLER_92_958 ();
 sg13g2_fill_8 FILLER_92_966 ();
 sg13g2_fill_8 FILLER_92_974 ();
 sg13g2_fill_8 FILLER_92_982 ();
 sg13g2_fill_8 FILLER_92_990 ();
 sg13g2_fill_8 FILLER_92_998 ();
 sg13g2_fill_8 FILLER_92_1006 ();
 sg13g2_fill_8 FILLER_92_1014 ();
 sg13g2_fill_8 FILLER_92_1022 ();
 sg13g2_fill_8 FILLER_92_1030 ();
 sg13g2_fill_8 FILLER_92_1038 ();
 sg13g2_fill_8 FILLER_92_1046 ();
 sg13g2_fill_8 FILLER_92_1054 ();
 sg13g2_fill_8 FILLER_92_1062 ();
 sg13g2_fill_8 FILLER_92_1070 ();
 sg13g2_fill_8 FILLER_92_1078 ();
 sg13g2_fill_8 FILLER_92_1086 ();
 sg13g2_fill_8 FILLER_92_1094 ();
 sg13g2_fill_8 FILLER_92_1102 ();
 sg13g2_fill_8 FILLER_92_1110 ();
 sg13g2_fill_8 FILLER_92_1118 ();
 sg13g2_fill_8 FILLER_92_1126 ();
 sg13g2_fill_8 FILLER_92_1134 ();
 sg13g2_fill_2 FILLER_92_1142 ();
 sg13g2_fill_8 FILLER_93_0 ();
 sg13g2_fill_8 FILLER_93_8 ();
 sg13g2_fill_8 FILLER_93_16 ();
 sg13g2_fill_8 FILLER_93_24 ();
 sg13g2_fill_8 FILLER_93_32 ();
 sg13g2_fill_8 FILLER_93_40 ();
 sg13g2_fill_8 FILLER_93_48 ();
 sg13g2_fill_8 FILLER_93_56 ();
 sg13g2_fill_8 FILLER_93_64 ();
 sg13g2_fill_8 FILLER_93_72 ();
 sg13g2_fill_8 FILLER_93_80 ();
 sg13g2_fill_8 FILLER_93_88 ();
 sg13g2_fill_8 FILLER_93_96 ();
 sg13g2_fill_8 FILLER_93_104 ();
 sg13g2_fill_8 FILLER_93_112 ();
 sg13g2_fill_8 FILLER_93_120 ();
 sg13g2_fill_8 FILLER_93_128 ();
 sg13g2_fill_8 FILLER_93_136 ();
 sg13g2_fill_8 FILLER_93_144 ();
 sg13g2_fill_8 FILLER_93_152 ();
 sg13g2_fill_8 FILLER_93_160 ();
 sg13g2_fill_8 FILLER_93_168 ();
 sg13g2_fill_8 FILLER_93_176 ();
 sg13g2_fill_8 FILLER_93_184 ();
 sg13g2_fill_8 FILLER_93_192 ();
 sg13g2_fill_8 FILLER_93_200 ();
 sg13g2_fill_8 FILLER_93_208 ();
 sg13g2_fill_8 FILLER_93_216 ();
 sg13g2_fill_8 FILLER_93_224 ();
 sg13g2_fill_8 FILLER_93_232 ();
 sg13g2_fill_8 FILLER_93_240 ();
 sg13g2_fill_8 FILLER_93_248 ();
 sg13g2_fill_8 FILLER_93_256 ();
 sg13g2_fill_8 FILLER_93_264 ();
 sg13g2_fill_8 FILLER_93_272 ();
 sg13g2_fill_8 FILLER_93_280 ();
 sg13g2_fill_8 FILLER_93_288 ();
 sg13g2_fill_8 FILLER_93_296 ();
 sg13g2_fill_8 FILLER_93_304 ();
 sg13g2_fill_8 FILLER_93_312 ();
 sg13g2_fill_4 FILLER_93_320 ();
 sg13g2_fill_2 FILLER_93_324 ();
 sg13g2_fill_8 FILLER_93_438 ();
 sg13g2_fill_8 FILLER_93_446 ();
 sg13g2_fill_8 FILLER_93_454 ();
 sg13g2_fill_8 FILLER_93_462 ();
 sg13g2_fill_8 FILLER_93_470 ();
 sg13g2_fill_8 FILLER_93_478 ();
 sg13g2_fill_8 FILLER_93_486 ();
 sg13g2_fill_8 FILLER_93_494 ();
 sg13g2_fill_8 FILLER_93_502 ();
 sg13g2_fill_8 FILLER_93_510 ();
 sg13g2_fill_8 FILLER_93_518 ();
 sg13g2_fill_8 FILLER_93_526 ();
 sg13g2_fill_8 FILLER_93_534 ();
 sg13g2_fill_8 FILLER_93_542 ();
 sg13g2_fill_8 FILLER_93_550 ();
 sg13g2_fill_8 FILLER_93_558 ();
 sg13g2_fill_8 FILLER_93_566 ();
 sg13g2_fill_8 FILLER_93_574 ();
 sg13g2_fill_8 FILLER_93_582 ();
 sg13g2_fill_8 FILLER_93_590 ();
 sg13g2_fill_8 FILLER_93_598 ();
 sg13g2_fill_8 FILLER_93_606 ();
 sg13g2_fill_8 FILLER_93_614 ();
 sg13g2_fill_8 FILLER_93_622 ();
 sg13g2_fill_8 FILLER_93_630 ();
 sg13g2_fill_8 FILLER_93_638 ();
 sg13g2_fill_8 FILLER_93_646 ();
 sg13g2_fill_8 FILLER_93_654 ();
 sg13g2_fill_8 FILLER_93_662 ();
 sg13g2_fill_8 FILLER_93_670 ();
 sg13g2_fill_8 FILLER_93_678 ();
 sg13g2_fill_8 FILLER_93_686 ();
 sg13g2_fill_8 FILLER_93_694 ();
 sg13g2_fill_8 FILLER_93_702 ();
 sg13g2_fill_8 FILLER_93_741 ();
 sg13g2_fill_1 FILLER_93_749 ();
 sg13g2_fill_8 FILLER_93_776 ();
 sg13g2_fill_4 FILLER_93_784 ();
 sg13g2_fill_2 FILLER_93_788 ();
 sg13g2_fill_1 FILLER_93_790 ();
 sg13g2_fill_8 FILLER_93_824 ();
 sg13g2_fill_8 FILLER_93_832 ();
 sg13g2_fill_8 FILLER_93_840 ();
 sg13g2_fill_8 FILLER_93_848 ();
 sg13g2_fill_8 FILLER_93_856 ();
 sg13g2_fill_1 FILLER_93_864 ();
 sg13g2_fill_8 FILLER_93_868 ();
 sg13g2_fill_4 FILLER_93_876 ();
 sg13g2_fill_8 FILLER_93_888 ();
 sg13g2_fill_8 FILLER_93_896 ();
 sg13g2_fill_8 FILLER_93_904 ();
 sg13g2_fill_8 FILLER_93_912 ();
 sg13g2_fill_2 FILLER_93_920 ();
 sg13g2_fill_1 FILLER_93_935 ();
 sg13g2_fill_8 FILLER_93_956 ();
 sg13g2_fill_8 FILLER_93_964 ();
 sg13g2_fill_8 FILLER_93_972 ();
 sg13g2_fill_8 FILLER_93_980 ();
 sg13g2_fill_8 FILLER_93_988 ();
 sg13g2_fill_8 FILLER_93_996 ();
 sg13g2_fill_8 FILLER_93_1004 ();
 sg13g2_fill_8 FILLER_93_1012 ();
 sg13g2_fill_8 FILLER_93_1020 ();
 sg13g2_fill_8 FILLER_93_1028 ();
 sg13g2_fill_8 FILLER_93_1036 ();
 sg13g2_fill_8 FILLER_93_1044 ();
 sg13g2_fill_8 FILLER_93_1052 ();
 sg13g2_fill_8 FILLER_93_1060 ();
 sg13g2_fill_8 FILLER_93_1068 ();
 sg13g2_fill_8 FILLER_93_1076 ();
 sg13g2_fill_8 FILLER_93_1084 ();
 sg13g2_fill_8 FILLER_93_1092 ();
 sg13g2_fill_8 FILLER_93_1100 ();
 sg13g2_fill_8 FILLER_93_1108 ();
 sg13g2_fill_8 FILLER_93_1116 ();
 sg13g2_fill_8 FILLER_93_1124 ();
 sg13g2_fill_8 FILLER_93_1132 ();
 sg13g2_fill_4 FILLER_93_1140 ();
 sg13g2_fill_8 FILLER_94_0 ();
 sg13g2_fill_8 FILLER_94_8 ();
 sg13g2_fill_8 FILLER_94_16 ();
 sg13g2_fill_8 FILLER_94_24 ();
 sg13g2_fill_8 FILLER_94_32 ();
 sg13g2_fill_8 FILLER_94_40 ();
 sg13g2_fill_8 FILLER_94_48 ();
 sg13g2_fill_8 FILLER_94_56 ();
 sg13g2_fill_8 FILLER_94_64 ();
 sg13g2_fill_8 FILLER_94_72 ();
 sg13g2_fill_8 FILLER_94_80 ();
 sg13g2_fill_8 FILLER_94_88 ();
 sg13g2_fill_8 FILLER_94_96 ();
 sg13g2_fill_8 FILLER_94_104 ();
 sg13g2_fill_8 FILLER_94_112 ();
 sg13g2_fill_8 FILLER_94_120 ();
 sg13g2_fill_8 FILLER_94_128 ();
 sg13g2_fill_8 FILLER_94_136 ();
 sg13g2_fill_8 FILLER_94_144 ();
 sg13g2_fill_8 FILLER_94_152 ();
 sg13g2_fill_8 FILLER_94_160 ();
 sg13g2_fill_8 FILLER_94_168 ();
 sg13g2_fill_8 FILLER_94_176 ();
 sg13g2_fill_8 FILLER_94_184 ();
 sg13g2_fill_8 FILLER_94_192 ();
 sg13g2_fill_8 FILLER_94_200 ();
 sg13g2_fill_8 FILLER_94_208 ();
 sg13g2_fill_8 FILLER_94_216 ();
 sg13g2_fill_8 FILLER_94_224 ();
 sg13g2_fill_8 FILLER_94_232 ();
 sg13g2_fill_8 FILLER_94_240 ();
 sg13g2_fill_8 FILLER_94_248 ();
 sg13g2_fill_8 FILLER_94_256 ();
 sg13g2_fill_8 FILLER_94_264 ();
 sg13g2_fill_8 FILLER_94_272 ();
 sg13g2_fill_8 FILLER_94_280 ();
 sg13g2_fill_4 FILLER_94_288 ();
 sg13g2_fill_2 FILLER_94_292 ();
 sg13g2_fill_1 FILLER_94_294 ();
 sg13g2_fill_8 FILLER_94_320 ();
 sg13g2_fill_4 FILLER_94_328 ();
 sg13g2_fill_2 FILLER_94_332 ();
 sg13g2_fill_1 FILLER_94_334 ();
 sg13g2_fill_2 FILLER_94_352 ();
 sg13g2_fill_2 FILLER_94_367 ();
 sg13g2_fill_8 FILLER_94_408 ();
 sg13g2_fill_8 FILLER_94_416 ();
 sg13g2_fill_8 FILLER_94_424 ();
 sg13g2_fill_8 FILLER_94_432 ();
 sg13g2_fill_8 FILLER_94_440 ();
 sg13g2_fill_8 FILLER_94_448 ();
 sg13g2_fill_8 FILLER_94_456 ();
 sg13g2_fill_8 FILLER_94_464 ();
 sg13g2_fill_8 FILLER_94_472 ();
 sg13g2_fill_8 FILLER_94_480 ();
 sg13g2_fill_8 FILLER_94_488 ();
 sg13g2_fill_8 FILLER_94_496 ();
 sg13g2_fill_8 FILLER_94_504 ();
 sg13g2_fill_8 FILLER_94_512 ();
 sg13g2_fill_8 FILLER_94_520 ();
 sg13g2_fill_8 FILLER_94_528 ();
 sg13g2_fill_8 FILLER_94_536 ();
 sg13g2_fill_8 FILLER_94_544 ();
 sg13g2_fill_8 FILLER_94_552 ();
 sg13g2_fill_8 FILLER_94_560 ();
 sg13g2_fill_8 FILLER_94_568 ();
 sg13g2_fill_8 FILLER_94_576 ();
 sg13g2_fill_8 FILLER_94_584 ();
 sg13g2_fill_8 FILLER_94_592 ();
 sg13g2_fill_8 FILLER_94_600 ();
 sg13g2_fill_8 FILLER_94_608 ();
 sg13g2_fill_8 FILLER_94_616 ();
 sg13g2_fill_8 FILLER_94_624 ();
 sg13g2_fill_8 FILLER_94_632 ();
 sg13g2_fill_8 FILLER_94_640 ();
 sg13g2_fill_8 FILLER_94_648 ();
 sg13g2_fill_8 FILLER_94_656 ();
 sg13g2_fill_8 FILLER_94_664 ();
 sg13g2_fill_8 FILLER_94_672 ();
 sg13g2_fill_8 FILLER_94_680 ();
 sg13g2_fill_8 FILLER_94_688 ();
 sg13g2_fill_8 FILLER_94_696 ();
 sg13g2_fill_4 FILLER_94_704 ();
 sg13g2_fill_2 FILLER_94_708 ();
 sg13g2_fill_8 FILLER_94_771 ();
 sg13g2_fill_8 FILLER_94_779 ();
 sg13g2_fill_8 FILLER_94_787 ();
 sg13g2_fill_8 FILLER_94_795 ();
 sg13g2_fill_8 FILLER_94_803 ();
 sg13g2_fill_8 FILLER_94_811 ();
 sg13g2_fill_2 FILLER_94_819 ();
 sg13g2_fill_4 FILLER_94_825 ();
 sg13g2_fill_2 FILLER_94_829 ();
 sg13g2_fill_4 FILLER_94_857 ();
 sg13g2_fill_1 FILLER_94_861 ();
 sg13g2_fill_8 FILLER_94_876 ();
 sg13g2_fill_8 FILLER_94_910 ();
 sg13g2_fill_8 FILLER_94_957 ();
 sg13g2_fill_8 FILLER_94_965 ();
 sg13g2_fill_8 FILLER_94_973 ();
 sg13g2_fill_8 FILLER_94_981 ();
 sg13g2_fill_8 FILLER_94_989 ();
 sg13g2_fill_8 FILLER_94_997 ();
 sg13g2_fill_8 FILLER_94_1005 ();
 sg13g2_fill_8 FILLER_94_1013 ();
 sg13g2_fill_8 FILLER_94_1021 ();
 sg13g2_fill_8 FILLER_94_1029 ();
 sg13g2_fill_8 FILLER_94_1037 ();
 sg13g2_fill_8 FILLER_94_1045 ();
 sg13g2_fill_8 FILLER_94_1053 ();
 sg13g2_fill_8 FILLER_94_1061 ();
 sg13g2_fill_8 FILLER_94_1069 ();
 sg13g2_fill_8 FILLER_94_1077 ();
 sg13g2_fill_8 FILLER_94_1085 ();
 sg13g2_fill_8 FILLER_94_1093 ();
 sg13g2_fill_8 FILLER_94_1101 ();
 sg13g2_fill_8 FILLER_94_1109 ();
 sg13g2_fill_8 FILLER_94_1117 ();
 sg13g2_fill_8 FILLER_94_1125 ();
 sg13g2_fill_8 FILLER_94_1133 ();
 sg13g2_fill_2 FILLER_94_1141 ();
 sg13g2_fill_1 FILLER_94_1143 ();
 sg13g2_fill_8 FILLER_95_0 ();
 sg13g2_fill_8 FILLER_95_8 ();
 sg13g2_fill_8 FILLER_95_16 ();
 sg13g2_fill_8 FILLER_95_24 ();
 sg13g2_fill_8 FILLER_95_32 ();
 sg13g2_fill_8 FILLER_95_40 ();
 sg13g2_fill_8 FILLER_95_48 ();
 sg13g2_fill_8 FILLER_95_56 ();
 sg13g2_fill_8 FILLER_95_64 ();
 sg13g2_fill_8 FILLER_95_72 ();
 sg13g2_fill_8 FILLER_95_80 ();
 sg13g2_fill_8 FILLER_95_88 ();
 sg13g2_fill_8 FILLER_95_96 ();
 sg13g2_fill_8 FILLER_95_104 ();
 sg13g2_fill_8 FILLER_95_112 ();
 sg13g2_fill_8 FILLER_95_120 ();
 sg13g2_fill_8 FILLER_95_128 ();
 sg13g2_fill_8 FILLER_95_136 ();
 sg13g2_fill_8 FILLER_95_144 ();
 sg13g2_fill_8 FILLER_95_152 ();
 sg13g2_fill_8 FILLER_95_160 ();
 sg13g2_fill_8 FILLER_95_168 ();
 sg13g2_fill_8 FILLER_95_176 ();
 sg13g2_fill_8 FILLER_95_184 ();
 sg13g2_fill_8 FILLER_95_192 ();
 sg13g2_fill_8 FILLER_95_200 ();
 sg13g2_fill_8 FILLER_95_208 ();
 sg13g2_fill_8 FILLER_95_216 ();
 sg13g2_fill_8 FILLER_95_224 ();
 sg13g2_fill_8 FILLER_95_232 ();
 sg13g2_fill_8 FILLER_95_240 ();
 sg13g2_fill_8 FILLER_95_248 ();
 sg13g2_fill_8 FILLER_95_256 ();
 sg13g2_fill_8 FILLER_95_264 ();
 sg13g2_fill_8 FILLER_95_272 ();
 sg13g2_fill_8 FILLER_95_280 ();
 sg13g2_fill_8 FILLER_95_288 ();
 sg13g2_fill_8 FILLER_95_296 ();
 sg13g2_fill_8 FILLER_95_304 ();
 sg13g2_fill_8 FILLER_95_312 ();
 sg13g2_fill_8 FILLER_95_320 ();
 sg13g2_fill_8 FILLER_95_328 ();
 sg13g2_fill_8 FILLER_95_336 ();
 sg13g2_fill_2 FILLER_95_349 ();
 sg13g2_fill_8 FILLER_95_356 ();
 sg13g2_fill_8 FILLER_95_364 ();
 sg13g2_fill_1 FILLER_95_372 ();
 sg13g2_fill_8 FILLER_95_378 ();
 sg13g2_fill_8 FILLER_95_386 ();
 sg13g2_fill_8 FILLER_95_394 ();
 sg13g2_fill_8 FILLER_95_402 ();
 sg13g2_fill_8 FILLER_95_410 ();
 sg13g2_fill_8 FILLER_95_418 ();
 sg13g2_fill_8 FILLER_95_426 ();
 sg13g2_fill_8 FILLER_95_434 ();
 sg13g2_fill_8 FILLER_95_442 ();
 sg13g2_fill_8 FILLER_95_450 ();
 sg13g2_fill_8 FILLER_95_458 ();
 sg13g2_fill_8 FILLER_95_466 ();
 sg13g2_fill_8 FILLER_95_474 ();
 sg13g2_fill_8 FILLER_95_482 ();
 sg13g2_fill_8 FILLER_95_490 ();
 sg13g2_fill_8 FILLER_95_498 ();
 sg13g2_fill_8 FILLER_95_506 ();
 sg13g2_fill_8 FILLER_95_514 ();
 sg13g2_fill_8 FILLER_95_522 ();
 sg13g2_fill_8 FILLER_95_530 ();
 sg13g2_fill_8 FILLER_95_538 ();
 sg13g2_fill_8 FILLER_95_546 ();
 sg13g2_fill_8 FILLER_95_554 ();
 sg13g2_fill_8 FILLER_95_562 ();
 sg13g2_fill_8 FILLER_95_570 ();
 sg13g2_fill_8 FILLER_95_578 ();
 sg13g2_fill_8 FILLER_95_586 ();
 sg13g2_fill_8 FILLER_95_594 ();
 sg13g2_fill_8 FILLER_95_602 ();
 sg13g2_fill_8 FILLER_95_610 ();
 sg13g2_fill_8 FILLER_95_618 ();
 sg13g2_fill_8 FILLER_95_626 ();
 sg13g2_fill_8 FILLER_95_634 ();
 sg13g2_fill_8 FILLER_95_642 ();
 sg13g2_fill_8 FILLER_95_650 ();
 sg13g2_fill_8 FILLER_95_658 ();
 sg13g2_fill_8 FILLER_95_666 ();
 sg13g2_fill_8 FILLER_95_674 ();
 sg13g2_fill_8 FILLER_95_682 ();
 sg13g2_fill_8 FILLER_95_690 ();
 sg13g2_fill_1 FILLER_95_698 ();
 sg13g2_fill_8 FILLER_95_725 ();
 sg13g2_fill_8 FILLER_95_733 ();
 sg13g2_fill_8 FILLER_95_741 ();
 sg13g2_fill_8 FILLER_95_749 ();
 sg13g2_fill_4 FILLER_95_757 ();
 sg13g2_fill_4 FILLER_95_766 ();
 sg13g2_fill_8 FILLER_95_780 ();
 sg13g2_fill_8 FILLER_95_788 ();
 sg13g2_fill_8 FILLER_95_806 ();
 sg13g2_fill_1 FILLER_95_814 ();
 sg13g2_fill_4 FILLER_95_845 ();
 sg13g2_fill_1 FILLER_95_849 ();
 sg13g2_fill_4 FILLER_95_894 ();
 sg13g2_fill_2 FILLER_95_898 ();
 sg13g2_fill_1 FILLER_95_900 ();
 sg13g2_fill_1 FILLER_95_906 ();
 sg13g2_fill_8 FILLER_95_911 ();
 sg13g2_fill_8 FILLER_95_919 ();
 sg13g2_fill_4 FILLER_95_927 ();
 sg13g2_fill_1 FILLER_95_931 ();
 sg13g2_fill_8 FILLER_95_949 ();
 sg13g2_fill_8 FILLER_95_957 ();
 sg13g2_fill_8 FILLER_95_965 ();
 sg13g2_fill_8 FILLER_95_973 ();
 sg13g2_fill_8 FILLER_95_981 ();
 sg13g2_fill_8 FILLER_95_989 ();
 sg13g2_fill_8 FILLER_95_997 ();
 sg13g2_fill_8 FILLER_95_1005 ();
 sg13g2_fill_8 FILLER_95_1013 ();
 sg13g2_fill_8 FILLER_95_1021 ();
 sg13g2_fill_8 FILLER_95_1029 ();
 sg13g2_fill_8 FILLER_95_1037 ();
 sg13g2_fill_8 FILLER_95_1045 ();
 sg13g2_fill_8 FILLER_95_1053 ();
 sg13g2_fill_8 FILLER_95_1061 ();
 sg13g2_fill_8 FILLER_95_1069 ();
 sg13g2_fill_8 FILLER_95_1077 ();
 sg13g2_fill_8 FILLER_95_1085 ();
 sg13g2_fill_8 FILLER_95_1093 ();
 sg13g2_fill_8 FILLER_95_1101 ();
 sg13g2_fill_8 FILLER_95_1109 ();
 sg13g2_fill_8 FILLER_95_1117 ();
 sg13g2_fill_8 FILLER_95_1125 ();
 sg13g2_fill_8 FILLER_95_1133 ();
 sg13g2_fill_2 FILLER_95_1141 ();
 sg13g2_fill_1 FILLER_95_1143 ();
 sg13g2_fill_8 FILLER_96_0 ();
 sg13g2_fill_8 FILLER_96_8 ();
 sg13g2_fill_8 FILLER_96_16 ();
 sg13g2_fill_8 FILLER_96_24 ();
 sg13g2_fill_8 FILLER_96_32 ();
 sg13g2_fill_8 FILLER_96_40 ();
 sg13g2_fill_8 FILLER_96_48 ();
 sg13g2_fill_8 FILLER_96_56 ();
 sg13g2_fill_8 FILLER_96_64 ();
 sg13g2_fill_8 FILLER_96_72 ();
 sg13g2_fill_8 FILLER_96_80 ();
 sg13g2_fill_8 FILLER_96_88 ();
 sg13g2_fill_8 FILLER_96_96 ();
 sg13g2_fill_8 FILLER_96_104 ();
 sg13g2_fill_8 FILLER_96_112 ();
 sg13g2_fill_8 FILLER_96_120 ();
 sg13g2_fill_8 FILLER_96_128 ();
 sg13g2_fill_8 FILLER_96_136 ();
 sg13g2_fill_8 FILLER_96_144 ();
 sg13g2_fill_8 FILLER_96_152 ();
 sg13g2_fill_8 FILLER_96_160 ();
 sg13g2_fill_8 FILLER_96_168 ();
 sg13g2_fill_8 FILLER_96_176 ();
 sg13g2_fill_8 FILLER_96_184 ();
 sg13g2_fill_8 FILLER_96_192 ();
 sg13g2_fill_8 FILLER_96_200 ();
 sg13g2_fill_8 FILLER_96_208 ();
 sg13g2_fill_8 FILLER_96_216 ();
 sg13g2_fill_8 FILLER_96_224 ();
 sg13g2_fill_8 FILLER_96_232 ();
 sg13g2_fill_8 FILLER_96_240 ();
 sg13g2_fill_8 FILLER_96_248 ();
 sg13g2_fill_8 FILLER_96_256 ();
 sg13g2_fill_8 FILLER_96_264 ();
 sg13g2_fill_8 FILLER_96_272 ();
 sg13g2_fill_8 FILLER_96_280 ();
 sg13g2_fill_8 FILLER_96_288 ();
 sg13g2_fill_8 FILLER_96_296 ();
 sg13g2_fill_8 FILLER_96_304 ();
 sg13g2_fill_8 FILLER_96_312 ();
 sg13g2_fill_8 FILLER_96_320 ();
 sg13g2_fill_8 FILLER_96_328 ();
 sg13g2_fill_8 FILLER_96_336 ();
 sg13g2_fill_8 FILLER_96_344 ();
 sg13g2_fill_8 FILLER_96_352 ();
 sg13g2_fill_8 FILLER_96_360 ();
 sg13g2_fill_8 FILLER_96_368 ();
 sg13g2_fill_8 FILLER_96_376 ();
 sg13g2_fill_8 FILLER_96_384 ();
 sg13g2_fill_8 FILLER_96_392 ();
 sg13g2_fill_8 FILLER_96_400 ();
 sg13g2_fill_8 FILLER_96_408 ();
 sg13g2_fill_8 FILLER_96_416 ();
 sg13g2_fill_8 FILLER_96_424 ();
 sg13g2_fill_8 FILLER_96_432 ();
 sg13g2_fill_8 FILLER_96_440 ();
 sg13g2_fill_8 FILLER_96_448 ();
 sg13g2_fill_8 FILLER_96_456 ();
 sg13g2_fill_8 FILLER_96_464 ();
 sg13g2_fill_8 FILLER_96_472 ();
 sg13g2_fill_8 FILLER_96_480 ();
 sg13g2_fill_8 FILLER_96_488 ();
 sg13g2_fill_8 FILLER_96_496 ();
 sg13g2_fill_8 FILLER_96_504 ();
 sg13g2_fill_8 FILLER_96_512 ();
 sg13g2_fill_8 FILLER_96_520 ();
 sg13g2_fill_8 FILLER_96_528 ();
 sg13g2_fill_8 FILLER_96_536 ();
 sg13g2_fill_8 FILLER_96_544 ();
 sg13g2_fill_8 FILLER_96_552 ();
 sg13g2_fill_8 FILLER_96_560 ();
 sg13g2_fill_8 FILLER_96_568 ();
 sg13g2_fill_8 FILLER_96_576 ();
 sg13g2_fill_8 FILLER_96_584 ();
 sg13g2_fill_8 FILLER_96_592 ();
 sg13g2_fill_8 FILLER_96_600 ();
 sg13g2_fill_8 FILLER_96_608 ();
 sg13g2_fill_8 FILLER_96_616 ();
 sg13g2_fill_8 FILLER_96_624 ();
 sg13g2_fill_8 FILLER_96_632 ();
 sg13g2_fill_8 FILLER_96_640 ();
 sg13g2_fill_8 FILLER_96_648 ();
 sg13g2_fill_8 FILLER_96_656 ();
 sg13g2_fill_8 FILLER_96_664 ();
 sg13g2_fill_8 FILLER_96_672 ();
 sg13g2_fill_4 FILLER_96_680 ();
 sg13g2_fill_8 FILLER_96_710 ();
 sg13g2_fill_8 FILLER_96_718 ();
 sg13g2_fill_8 FILLER_96_726 ();
 sg13g2_fill_8 FILLER_96_734 ();
 sg13g2_fill_8 FILLER_96_742 ();
 sg13g2_fill_4 FILLER_96_750 ();
 sg13g2_fill_2 FILLER_96_754 ();
 sg13g2_fill_1 FILLER_96_756 ();
 sg13g2_fill_2 FILLER_96_789 ();
 sg13g2_fill_1 FILLER_96_791 ();
 sg13g2_fill_8 FILLER_96_840 ();
 sg13g2_fill_4 FILLER_96_848 ();
 sg13g2_fill_2 FILLER_96_897 ();
 sg13g2_fill_1 FILLER_96_899 ();
 sg13g2_fill_2 FILLER_96_919 ();
 sg13g2_fill_8 FILLER_96_924 ();
 sg13g2_fill_8 FILLER_96_932 ();
 sg13g2_fill_8 FILLER_96_940 ();
 sg13g2_fill_8 FILLER_96_948 ();
 sg13g2_fill_8 FILLER_96_956 ();
 sg13g2_fill_8 FILLER_96_964 ();
 sg13g2_fill_8 FILLER_96_972 ();
 sg13g2_fill_8 FILLER_96_980 ();
 sg13g2_fill_8 FILLER_96_988 ();
 sg13g2_fill_8 FILLER_96_996 ();
 sg13g2_fill_8 FILLER_96_1004 ();
 sg13g2_fill_8 FILLER_96_1012 ();
 sg13g2_fill_8 FILLER_96_1020 ();
 sg13g2_fill_8 FILLER_96_1028 ();
 sg13g2_fill_8 FILLER_96_1036 ();
 sg13g2_fill_8 FILLER_96_1044 ();
 sg13g2_fill_8 FILLER_96_1052 ();
 sg13g2_fill_8 FILLER_96_1060 ();
 sg13g2_fill_8 FILLER_96_1068 ();
 sg13g2_fill_8 FILLER_96_1076 ();
 sg13g2_fill_8 FILLER_96_1084 ();
 sg13g2_fill_8 FILLER_96_1092 ();
 sg13g2_fill_8 FILLER_96_1100 ();
 sg13g2_fill_8 FILLER_96_1108 ();
 sg13g2_fill_8 FILLER_96_1116 ();
 sg13g2_fill_8 FILLER_96_1124 ();
 sg13g2_fill_8 FILLER_96_1132 ();
 sg13g2_fill_4 FILLER_96_1140 ();
 sg13g2_fill_8 FILLER_97_0 ();
 sg13g2_fill_8 FILLER_97_8 ();
 sg13g2_fill_8 FILLER_97_16 ();
 sg13g2_fill_8 FILLER_97_24 ();
 sg13g2_fill_8 FILLER_97_32 ();
 sg13g2_fill_8 FILLER_97_40 ();
 sg13g2_fill_8 FILLER_97_48 ();
 sg13g2_fill_8 FILLER_97_56 ();
 sg13g2_fill_8 FILLER_97_64 ();
 sg13g2_fill_8 FILLER_97_72 ();
 sg13g2_fill_8 FILLER_97_80 ();
 sg13g2_fill_8 FILLER_97_88 ();
 sg13g2_fill_8 FILLER_97_96 ();
 sg13g2_fill_8 FILLER_97_104 ();
 sg13g2_fill_8 FILLER_97_112 ();
 sg13g2_fill_8 FILLER_97_120 ();
 sg13g2_fill_8 FILLER_97_128 ();
 sg13g2_fill_8 FILLER_97_136 ();
 sg13g2_fill_8 FILLER_97_144 ();
 sg13g2_fill_8 FILLER_97_152 ();
 sg13g2_fill_8 FILLER_97_160 ();
 sg13g2_fill_8 FILLER_97_168 ();
 sg13g2_fill_8 FILLER_97_176 ();
 sg13g2_fill_8 FILLER_97_184 ();
 sg13g2_fill_8 FILLER_97_192 ();
 sg13g2_fill_8 FILLER_97_200 ();
 sg13g2_fill_8 FILLER_97_208 ();
 sg13g2_fill_8 FILLER_97_216 ();
 sg13g2_fill_8 FILLER_97_224 ();
 sg13g2_fill_8 FILLER_97_232 ();
 sg13g2_fill_8 FILLER_97_240 ();
 sg13g2_fill_8 FILLER_97_248 ();
 sg13g2_fill_8 FILLER_97_256 ();
 sg13g2_fill_8 FILLER_97_264 ();
 sg13g2_fill_8 FILLER_97_272 ();
 sg13g2_fill_8 FILLER_97_280 ();
 sg13g2_fill_8 FILLER_97_288 ();
 sg13g2_fill_8 FILLER_97_296 ();
 sg13g2_fill_8 FILLER_97_304 ();
 sg13g2_fill_8 FILLER_97_312 ();
 sg13g2_fill_8 FILLER_97_320 ();
 sg13g2_fill_8 FILLER_97_328 ();
 sg13g2_fill_8 FILLER_97_336 ();
 sg13g2_fill_8 FILLER_97_344 ();
 sg13g2_fill_8 FILLER_97_352 ();
 sg13g2_fill_8 FILLER_97_360 ();
 sg13g2_fill_8 FILLER_97_368 ();
 sg13g2_fill_8 FILLER_97_376 ();
 sg13g2_fill_8 FILLER_97_384 ();
 sg13g2_fill_8 FILLER_97_392 ();
 sg13g2_fill_8 FILLER_97_400 ();
 sg13g2_fill_8 FILLER_97_408 ();
 sg13g2_fill_8 FILLER_97_416 ();
 sg13g2_fill_8 FILLER_97_424 ();
 sg13g2_fill_8 FILLER_97_432 ();
 sg13g2_fill_8 FILLER_97_440 ();
 sg13g2_fill_8 FILLER_97_448 ();
 sg13g2_fill_8 FILLER_97_456 ();
 sg13g2_fill_8 FILLER_97_464 ();
 sg13g2_fill_8 FILLER_97_472 ();
 sg13g2_fill_8 FILLER_97_480 ();
 sg13g2_fill_8 FILLER_97_488 ();
 sg13g2_fill_8 FILLER_97_496 ();
 sg13g2_fill_8 FILLER_97_504 ();
 sg13g2_fill_8 FILLER_97_512 ();
 sg13g2_fill_8 FILLER_97_520 ();
 sg13g2_fill_8 FILLER_97_528 ();
 sg13g2_fill_8 FILLER_97_536 ();
 sg13g2_fill_8 FILLER_97_544 ();
 sg13g2_fill_8 FILLER_97_552 ();
 sg13g2_fill_8 FILLER_97_560 ();
 sg13g2_fill_8 FILLER_97_568 ();
 sg13g2_fill_8 FILLER_97_576 ();
 sg13g2_fill_8 FILLER_97_584 ();
 sg13g2_fill_8 FILLER_97_592 ();
 sg13g2_fill_8 FILLER_97_600 ();
 sg13g2_fill_8 FILLER_97_608 ();
 sg13g2_fill_8 FILLER_97_616 ();
 sg13g2_fill_8 FILLER_97_624 ();
 sg13g2_fill_8 FILLER_97_632 ();
 sg13g2_fill_8 FILLER_97_640 ();
 sg13g2_fill_8 FILLER_97_648 ();
 sg13g2_fill_8 FILLER_97_656 ();
 sg13g2_fill_8 FILLER_97_664 ();
 sg13g2_fill_8 FILLER_97_672 ();
 sg13g2_fill_8 FILLER_97_680 ();
 sg13g2_fill_8 FILLER_97_688 ();
 sg13g2_fill_8 FILLER_97_696 ();
 sg13g2_fill_8 FILLER_97_704 ();
 sg13g2_fill_8 FILLER_97_712 ();
 sg13g2_fill_8 FILLER_97_720 ();
 sg13g2_fill_8 FILLER_97_728 ();
 sg13g2_fill_2 FILLER_97_736 ();
 sg13g2_fill_1 FILLER_97_738 ();
 sg13g2_fill_2 FILLER_97_791 ();
 sg13g2_fill_1 FILLER_97_793 ();
 sg13g2_fill_8 FILLER_97_825 ();
 sg13g2_fill_8 FILLER_97_833 ();
 sg13g2_fill_2 FILLER_97_851 ();
 sg13g2_fill_2 FILLER_97_871 ();
 sg13g2_fill_8 FILLER_97_927 ();
 sg13g2_fill_8 FILLER_97_935 ();
 sg13g2_fill_8 FILLER_97_943 ();
 sg13g2_fill_8 FILLER_97_951 ();
 sg13g2_fill_8 FILLER_97_959 ();
 sg13g2_fill_8 FILLER_97_967 ();
 sg13g2_fill_8 FILLER_97_975 ();
 sg13g2_fill_8 FILLER_97_983 ();
 sg13g2_fill_8 FILLER_97_991 ();
 sg13g2_fill_8 FILLER_97_999 ();
 sg13g2_fill_8 FILLER_97_1007 ();
 sg13g2_fill_8 FILLER_97_1015 ();
 sg13g2_fill_8 FILLER_97_1023 ();
 sg13g2_fill_8 FILLER_97_1031 ();
 sg13g2_fill_8 FILLER_97_1039 ();
 sg13g2_fill_8 FILLER_97_1047 ();
 sg13g2_fill_8 FILLER_97_1055 ();
 sg13g2_fill_8 FILLER_97_1063 ();
 sg13g2_fill_8 FILLER_97_1071 ();
 sg13g2_fill_8 FILLER_97_1079 ();
 sg13g2_fill_8 FILLER_97_1087 ();
 sg13g2_fill_8 FILLER_97_1095 ();
 sg13g2_fill_8 FILLER_97_1103 ();
 sg13g2_fill_8 FILLER_97_1111 ();
 sg13g2_fill_8 FILLER_97_1119 ();
 sg13g2_fill_8 FILLER_97_1127 ();
 sg13g2_fill_8 FILLER_97_1135 ();
 sg13g2_fill_1 FILLER_97_1143 ();
 sg13g2_fill_8 FILLER_98_0 ();
 sg13g2_fill_8 FILLER_98_8 ();
 sg13g2_fill_8 FILLER_98_16 ();
 sg13g2_fill_8 FILLER_98_24 ();
 sg13g2_fill_8 FILLER_98_32 ();
 sg13g2_fill_8 FILLER_98_40 ();
 sg13g2_fill_8 FILLER_98_48 ();
 sg13g2_fill_8 FILLER_98_56 ();
 sg13g2_fill_8 FILLER_98_64 ();
 sg13g2_fill_8 FILLER_98_72 ();
 sg13g2_fill_8 FILLER_98_80 ();
 sg13g2_fill_8 FILLER_98_88 ();
 sg13g2_fill_8 FILLER_98_96 ();
 sg13g2_fill_8 FILLER_98_104 ();
 sg13g2_fill_8 FILLER_98_112 ();
 sg13g2_fill_8 FILLER_98_120 ();
 sg13g2_fill_8 FILLER_98_128 ();
 sg13g2_fill_8 FILLER_98_136 ();
 sg13g2_fill_8 FILLER_98_144 ();
 sg13g2_fill_8 FILLER_98_152 ();
 sg13g2_fill_8 FILLER_98_160 ();
 sg13g2_fill_8 FILLER_98_168 ();
 sg13g2_fill_8 FILLER_98_176 ();
 sg13g2_fill_8 FILLER_98_184 ();
 sg13g2_fill_8 FILLER_98_192 ();
 sg13g2_fill_8 FILLER_98_200 ();
 sg13g2_fill_8 FILLER_98_208 ();
 sg13g2_fill_8 FILLER_98_216 ();
 sg13g2_fill_8 FILLER_98_224 ();
 sg13g2_fill_8 FILLER_98_232 ();
 sg13g2_fill_8 FILLER_98_240 ();
 sg13g2_fill_8 FILLER_98_248 ();
 sg13g2_fill_8 FILLER_98_256 ();
 sg13g2_fill_8 FILLER_98_264 ();
 sg13g2_fill_8 FILLER_98_272 ();
 sg13g2_fill_8 FILLER_98_280 ();
 sg13g2_fill_8 FILLER_98_288 ();
 sg13g2_fill_8 FILLER_98_296 ();
 sg13g2_fill_8 FILLER_98_304 ();
 sg13g2_fill_8 FILLER_98_312 ();
 sg13g2_fill_8 FILLER_98_320 ();
 sg13g2_fill_8 FILLER_98_328 ();
 sg13g2_fill_8 FILLER_98_336 ();
 sg13g2_fill_8 FILLER_98_344 ();
 sg13g2_fill_8 FILLER_98_352 ();
 sg13g2_fill_8 FILLER_98_360 ();
 sg13g2_fill_8 FILLER_98_368 ();
 sg13g2_fill_8 FILLER_98_376 ();
 sg13g2_fill_8 FILLER_98_384 ();
 sg13g2_fill_8 FILLER_98_392 ();
 sg13g2_fill_8 FILLER_98_400 ();
 sg13g2_fill_8 FILLER_98_408 ();
 sg13g2_fill_8 FILLER_98_416 ();
 sg13g2_fill_8 FILLER_98_424 ();
 sg13g2_fill_8 FILLER_98_432 ();
 sg13g2_fill_8 FILLER_98_440 ();
 sg13g2_fill_8 FILLER_98_448 ();
 sg13g2_fill_8 FILLER_98_456 ();
 sg13g2_fill_8 FILLER_98_464 ();
 sg13g2_fill_8 FILLER_98_472 ();
 sg13g2_fill_8 FILLER_98_480 ();
 sg13g2_fill_8 FILLER_98_488 ();
 sg13g2_fill_8 FILLER_98_496 ();
 sg13g2_fill_8 FILLER_98_504 ();
 sg13g2_fill_8 FILLER_98_512 ();
 sg13g2_fill_8 FILLER_98_520 ();
 sg13g2_fill_8 FILLER_98_528 ();
 sg13g2_fill_8 FILLER_98_536 ();
 sg13g2_fill_8 FILLER_98_544 ();
 sg13g2_fill_8 FILLER_98_552 ();
 sg13g2_fill_8 FILLER_98_560 ();
 sg13g2_fill_8 FILLER_98_568 ();
 sg13g2_fill_8 FILLER_98_576 ();
 sg13g2_fill_8 FILLER_98_584 ();
 sg13g2_fill_8 FILLER_98_592 ();
 sg13g2_fill_8 FILLER_98_600 ();
 sg13g2_fill_8 FILLER_98_608 ();
 sg13g2_fill_8 FILLER_98_616 ();
 sg13g2_fill_8 FILLER_98_624 ();
 sg13g2_fill_8 FILLER_98_632 ();
 sg13g2_fill_8 FILLER_98_640 ();
 sg13g2_fill_8 FILLER_98_648 ();
 sg13g2_fill_8 FILLER_98_656 ();
 sg13g2_fill_8 FILLER_98_664 ();
 sg13g2_fill_8 FILLER_98_672 ();
 sg13g2_fill_8 FILLER_98_680 ();
 sg13g2_fill_8 FILLER_98_688 ();
 sg13g2_fill_8 FILLER_98_696 ();
 sg13g2_fill_8 FILLER_98_704 ();
 sg13g2_fill_8 FILLER_98_712 ();
 sg13g2_fill_8 FILLER_98_720 ();
 sg13g2_fill_8 FILLER_98_728 ();
 sg13g2_fill_4 FILLER_98_754 ();
 sg13g2_fill_2 FILLER_98_770 ();
 sg13g2_fill_8 FILLER_98_784 ();
 sg13g2_fill_2 FILLER_98_879 ();
 sg13g2_fill_1 FILLER_98_881 ();
 sg13g2_fill_8 FILLER_98_932 ();
 sg13g2_fill_8 FILLER_98_940 ();
 sg13g2_fill_8 FILLER_98_948 ();
 sg13g2_fill_8 FILLER_98_956 ();
 sg13g2_fill_8 FILLER_98_964 ();
 sg13g2_fill_8 FILLER_98_972 ();
 sg13g2_fill_8 FILLER_98_980 ();
 sg13g2_fill_8 FILLER_98_988 ();
 sg13g2_fill_8 FILLER_98_996 ();
 sg13g2_fill_8 FILLER_98_1004 ();
 sg13g2_fill_8 FILLER_98_1012 ();
 sg13g2_fill_8 FILLER_98_1020 ();
 sg13g2_fill_8 FILLER_98_1028 ();
 sg13g2_fill_8 FILLER_98_1036 ();
 sg13g2_fill_8 FILLER_98_1044 ();
 sg13g2_fill_8 FILLER_98_1052 ();
 sg13g2_fill_8 FILLER_98_1060 ();
 sg13g2_fill_8 FILLER_98_1068 ();
 sg13g2_fill_8 FILLER_98_1076 ();
 sg13g2_fill_8 FILLER_98_1084 ();
 sg13g2_fill_8 FILLER_98_1092 ();
 sg13g2_fill_8 FILLER_98_1100 ();
 sg13g2_fill_8 FILLER_98_1108 ();
 sg13g2_fill_8 FILLER_98_1116 ();
 sg13g2_fill_8 FILLER_98_1124 ();
 sg13g2_fill_8 FILLER_98_1132 ();
 sg13g2_fill_4 FILLER_98_1140 ();
 sg13g2_fill_8 FILLER_99_0 ();
 sg13g2_fill_8 FILLER_99_8 ();
 sg13g2_fill_8 FILLER_99_16 ();
 sg13g2_fill_8 FILLER_99_24 ();
 sg13g2_fill_8 FILLER_99_32 ();
 sg13g2_fill_8 FILLER_99_40 ();
 sg13g2_fill_8 FILLER_99_48 ();
 sg13g2_fill_8 FILLER_99_56 ();
 sg13g2_fill_8 FILLER_99_64 ();
 sg13g2_fill_8 FILLER_99_72 ();
 sg13g2_fill_8 FILLER_99_80 ();
 sg13g2_fill_8 FILLER_99_88 ();
 sg13g2_fill_8 FILLER_99_96 ();
 sg13g2_fill_8 FILLER_99_104 ();
 sg13g2_fill_8 FILLER_99_112 ();
 sg13g2_fill_8 FILLER_99_120 ();
 sg13g2_fill_8 FILLER_99_128 ();
 sg13g2_fill_8 FILLER_99_136 ();
 sg13g2_fill_8 FILLER_99_144 ();
 sg13g2_fill_8 FILLER_99_152 ();
 sg13g2_fill_8 FILLER_99_160 ();
 sg13g2_fill_8 FILLER_99_168 ();
 sg13g2_fill_8 FILLER_99_176 ();
 sg13g2_fill_8 FILLER_99_184 ();
 sg13g2_fill_8 FILLER_99_192 ();
 sg13g2_fill_8 FILLER_99_200 ();
 sg13g2_fill_8 FILLER_99_208 ();
 sg13g2_fill_8 FILLER_99_216 ();
 sg13g2_fill_8 FILLER_99_224 ();
 sg13g2_fill_8 FILLER_99_232 ();
 sg13g2_fill_8 FILLER_99_240 ();
 sg13g2_fill_8 FILLER_99_248 ();
 sg13g2_fill_8 FILLER_99_256 ();
 sg13g2_fill_8 FILLER_99_264 ();
 sg13g2_fill_8 FILLER_99_272 ();
 sg13g2_fill_8 FILLER_99_280 ();
 sg13g2_fill_8 FILLER_99_288 ();
 sg13g2_fill_8 FILLER_99_296 ();
 sg13g2_fill_8 FILLER_99_304 ();
 sg13g2_fill_8 FILLER_99_312 ();
 sg13g2_fill_8 FILLER_99_320 ();
 sg13g2_fill_8 FILLER_99_328 ();
 sg13g2_fill_8 FILLER_99_336 ();
 sg13g2_fill_8 FILLER_99_344 ();
 sg13g2_fill_8 FILLER_99_352 ();
 sg13g2_fill_8 FILLER_99_360 ();
 sg13g2_fill_8 FILLER_99_368 ();
 sg13g2_fill_8 FILLER_99_376 ();
 sg13g2_fill_8 FILLER_99_384 ();
 sg13g2_fill_8 FILLER_99_392 ();
 sg13g2_fill_8 FILLER_99_400 ();
 sg13g2_fill_8 FILLER_99_408 ();
 sg13g2_fill_8 FILLER_99_416 ();
 sg13g2_fill_8 FILLER_99_424 ();
 sg13g2_fill_8 FILLER_99_432 ();
 sg13g2_fill_8 FILLER_99_440 ();
 sg13g2_fill_8 FILLER_99_448 ();
 sg13g2_fill_8 FILLER_99_456 ();
 sg13g2_fill_8 FILLER_99_464 ();
 sg13g2_fill_8 FILLER_99_472 ();
 sg13g2_fill_8 FILLER_99_480 ();
 sg13g2_fill_8 FILLER_99_488 ();
 sg13g2_fill_8 FILLER_99_496 ();
 sg13g2_fill_8 FILLER_99_504 ();
 sg13g2_fill_8 FILLER_99_512 ();
 sg13g2_fill_8 FILLER_99_520 ();
 sg13g2_fill_8 FILLER_99_528 ();
 sg13g2_fill_8 FILLER_99_536 ();
 sg13g2_fill_8 FILLER_99_544 ();
 sg13g2_fill_8 FILLER_99_552 ();
 sg13g2_fill_8 FILLER_99_560 ();
 sg13g2_fill_8 FILLER_99_568 ();
 sg13g2_fill_8 FILLER_99_576 ();
 sg13g2_fill_8 FILLER_99_584 ();
 sg13g2_fill_8 FILLER_99_592 ();
 sg13g2_fill_8 FILLER_99_600 ();
 sg13g2_fill_8 FILLER_99_608 ();
 sg13g2_fill_8 FILLER_99_616 ();
 sg13g2_fill_8 FILLER_99_624 ();
 sg13g2_fill_8 FILLER_99_632 ();
 sg13g2_fill_8 FILLER_99_640 ();
 sg13g2_fill_8 FILLER_99_648 ();
 sg13g2_fill_8 FILLER_99_656 ();
 sg13g2_fill_8 FILLER_99_664 ();
 sg13g2_fill_8 FILLER_99_672 ();
 sg13g2_fill_8 FILLER_99_680 ();
 sg13g2_fill_8 FILLER_99_688 ();
 sg13g2_fill_8 FILLER_99_696 ();
 sg13g2_fill_8 FILLER_99_704 ();
 sg13g2_fill_8 FILLER_99_712 ();
 sg13g2_fill_8 FILLER_99_720 ();
 sg13g2_fill_8 FILLER_99_728 ();
 sg13g2_fill_8 FILLER_99_736 ();
 sg13g2_fill_8 FILLER_99_744 ();
 sg13g2_fill_8 FILLER_99_752 ();
 sg13g2_fill_8 FILLER_99_760 ();
 sg13g2_fill_1 FILLER_99_768 ();
 sg13g2_fill_8 FILLER_99_774 ();
 sg13g2_fill_8 FILLER_99_782 ();
 sg13g2_fill_8 FILLER_99_790 ();
 sg13g2_fill_8 FILLER_99_798 ();
 sg13g2_fill_8 FILLER_99_806 ();
 sg13g2_fill_2 FILLER_99_814 ();
 sg13g2_fill_8 FILLER_99_825 ();
 sg13g2_fill_8 FILLER_99_833 ();
 sg13g2_fill_4 FILLER_99_841 ();
 sg13g2_fill_1 FILLER_99_845 ();
 sg13g2_fill_1 FILLER_99_874 ();
 sg13g2_fill_1 FILLER_99_901 ();
 sg13g2_fill_8 FILLER_99_917 ();
 sg13g2_fill_8 FILLER_99_925 ();
 sg13g2_fill_8 FILLER_99_933 ();
 sg13g2_fill_8 FILLER_99_941 ();
 sg13g2_fill_8 FILLER_99_949 ();
 sg13g2_fill_8 FILLER_99_957 ();
 sg13g2_fill_8 FILLER_99_965 ();
 sg13g2_fill_8 FILLER_99_973 ();
 sg13g2_fill_8 FILLER_99_981 ();
 sg13g2_fill_8 FILLER_99_989 ();
 sg13g2_fill_8 FILLER_99_997 ();
 sg13g2_fill_8 FILLER_99_1005 ();
 sg13g2_fill_8 FILLER_99_1013 ();
 sg13g2_fill_8 FILLER_99_1021 ();
 sg13g2_fill_8 FILLER_99_1029 ();
 sg13g2_fill_8 FILLER_99_1037 ();
 sg13g2_fill_8 FILLER_99_1045 ();
 sg13g2_fill_8 FILLER_99_1053 ();
 sg13g2_fill_8 FILLER_99_1061 ();
 sg13g2_fill_8 FILLER_99_1069 ();
 sg13g2_fill_8 FILLER_99_1077 ();
 sg13g2_fill_8 FILLER_99_1085 ();
 sg13g2_fill_8 FILLER_99_1093 ();
 sg13g2_fill_8 FILLER_99_1101 ();
 sg13g2_fill_8 FILLER_99_1109 ();
 sg13g2_fill_8 FILLER_99_1117 ();
 sg13g2_fill_8 FILLER_99_1125 ();
 sg13g2_fill_8 FILLER_99_1133 ();
 sg13g2_fill_2 FILLER_99_1141 ();
 sg13g2_fill_1 FILLER_99_1143 ();
 sg13g2_fill_8 FILLER_100_0 ();
 sg13g2_fill_8 FILLER_100_8 ();
 sg13g2_fill_8 FILLER_100_16 ();
 sg13g2_fill_8 FILLER_100_24 ();
 sg13g2_fill_8 FILLER_100_32 ();
 sg13g2_fill_8 FILLER_100_40 ();
 sg13g2_fill_8 FILLER_100_48 ();
 sg13g2_fill_8 FILLER_100_56 ();
 sg13g2_fill_8 FILLER_100_64 ();
 sg13g2_fill_8 FILLER_100_72 ();
 sg13g2_fill_8 FILLER_100_80 ();
 sg13g2_fill_8 FILLER_100_88 ();
 sg13g2_fill_8 FILLER_100_96 ();
 sg13g2_fill_8 FILLER_100_104 ();
 sg13g2_fill_8 FILLER_100_112 ();
 sg13g2_fill_8 FILLER_100_120 ();
 sg13g2_fill_8 FILLER_100_128 ();
 sg13g2_fill_8 FILLER_100_136 ();
 sg13g2_fill_8 FILLER_100_144 ();
 sg13g2_fill_8 FILLER_100_152 ();
 sg13g2_fill_8 FILLER_100_160 ();
 sg13g2_fill_8 FILLER_100_168 ();
 sg13g2_fill_8 FILLER_100_176 ();
 sg13g2_fill_8 FILLER_100_184 ();
 sg13g2_fill_8 FILLER_100_192 ();
 sg13g2_fill_8 FILLER_100_200 ();
 sg13g2_fill_8 FILLER_100_208 ();
 sg13g2_fill_8 FILLER_100_216 ();
 sg13g2_fill_8 FILLER_100_224 ();
 sg13g2_fill_8 FILLER_100_232 ();
 sg13g2_fill_8 FILLER_100_240 ();
 sg13g2_fill_8 FILLER_100_248 ();
 sg13g2_fill_8 FILLER_100_256 ();
 sg13g2_fill_8 FILLER_100_264 ();
 sg13g2_fill_8 FILLER_100_272 ();
 sg13g2_fill_8 FILLER_100_280 ();
 sg13g2_fill_8 FILLER_100_288 ();
 sg13g2_fill_8 FILLER_100_296 ();
 sg13g2_fill_8 FILLER_100_304 ();
 sg13g2_fill_8 FILLER_100_312 ();
 sg13g2_fill_8 FILLER_100_320 ();
 sg13g2_fill_8 FILLER_100_328 ();
 sg13g2_fill_8 FILLER_100_336 ();
 sg13g2_fill_8 FILLER_100_344 ();
 sg13g2_fill_8 FILLER_100_352 ();
 sg13g2_fill_8 FILLER_100_360 ();
 sg13g2_fill_8 FILLER_100_368 ();
 sg13g2_fill_8 FILLER_100_376 ();
 sg13g2_fill_8 FILLER_100_384 ();
 sg13g2_fill_8 FILLER_100_392 ();
 sg13g2_fill_8 FILLER_100_400 ();
 sg13g2_fill_8 FILLER_100_408 ();
 sg13g2_fill_8 FILLER_100_416 ();
 sg13g2_fill_8 FILLER_100_424 ();
 sg13g2_fill_8 FILLER_100_432 ();
 sg13g2_fill_8 FILLER_100_440 ();
 sg13g2_fill_8 FILLER_100_448 ();
 sg13g2_fill_8 FILLER_100_456 ();
 sg13g2_fill_8 FILLER_100_464 ();
 sg13g2_fill_8 FILLER_100_472 ();
 sg13g2_fill_8 FILLER_100_480 ();
 sg13g2_fill_8 FILLER_100_488 ();
 sg13g2_fill_8 FILLER_100_496 ();
 sg13g2_fill_8 FILLER_100_504 ();
 sg13g2_fill_8 FILLER_100_512 ();
 sg13g2_fill_8 FILLER_100_520 ();
 sg13g2_fill_8 FILLER_100_528 ();
 sg13g2_fill_8 FILLER_100_536 ();
 sg13g2_fill_8 FILLER_100_544 ();
 sg13g2_fill_8 FILLER_100_552 ();
 sg13g2_fill_8 FILLER_100_560 ();
 sg13g2_fill_8 FILLER_100_568 ();
 sg13g2_fill_8 FILLER_100_576 ();
 sg13g2_fill_8 FILLER_100_584 ();
 sg13g2_fill_8 FILLER_100_592 ();
 sg13g2_fill_8 FILLER_100_600 ();
 sg13g2_fill_8 FILLER_100_608 ();
 sg13g2_fill_8 FILLER_100_616 ();
 sg13g2_fill_8 FILLER_100_624 ();
 sg13g2_fill_8 FILLER_100_632 ();
 sg13g2_fill_8 FILLER_100_640 ();
 sg13g2_fill_8 FILLER_100_648 ();
 sg13g2_fill_8 FILLER_100_656 ();
 sg13g2_fill_8 FILLER_100_664 ();
 sg13g2_fill_8 FILLER_100_672 ();
 sg13g2_fill_8 FILLER_100_680 ();
 sg13g2_fill_8 FILLER_100_688 ();
 sg13g2_fill_8 FILLER_100_696 ();
 sg13g2_fill_8 FILLER_100_704 ();
 sg13g2_fill_8 FILLER_100_712 ();
 sg13g2_fill_8 FILLER_100_720 ();
 sg13g2_fill_8 FILLER_100_728 ();
 sg13g2_fill_8 FILLER_100_736 ();
 sg13g2_fill_8 FILLER_100_744 ();
 sg13g2_fill_8 FILLER_100_752 ();
 sg13g2_fill_8 FILLER_100_760 ();
 sg13g2_fill_8 FILLER_100_768 ();
 sg13g2_fill_8 FILLER_100_776 ();
 sg13g2_fill_8 FILLER_100_784 ();
 sg13g2_fill_8 FILLER_100_792 ();
 sg13g2_fill_8 FILLER_100_800 ();
 sg13g2_fill_8 FILLER_100_808 ();
 sg13g2_fill_8 FILLER_100_816 ();
 sg13g2_fill_8 FILLER_100_824 ();
 sg13g2_fill_8 FILLER_100_832 ();
 sg13g2_fill_4 FILLER_100_840 ();
 sg13g2_fill_2 FILLER_100_844 ();
 sg13g2_fill_1 FILLER_100_846 ();
 sg13g2_fill_1 FILLER_100_851 ();
 sg13g2_fill_2 FILLER_100_856 ();
 sg13g2_fill_1 FILLER_100_858 ();
 sg13g2_fill_4 FILLER_100_864 ();
 sg13g2_fill_1 FILLER_100_868 ();
 sg13g2_fill_1 FILLER_100_899 ();
 sg13g2_fill_8 FILLER_100_907 ();
 sg13g2_fill_8 FILLER_100_915 ();
 sg13g2_fill_8 FILLER_100_923 ();
 sg13g2_fill_8 FILLER_100_931 ();
 sg13g2_fill_8 FILLER_100_939 ();
 sg13g2_fill_8 FILLER_100_947 ();
 sg13g2_fill_8 FILLER_100_955 ();
 sg13g2_fill_8 FILLER_100_963 ();
 sg13g2_fill_8 FILLER_100_971 ();
 sg13g2_fill_8 FILLER_100_979 ();
 sg13g2_fill_8 FILLER_100_987 ();
 sg13g2_fill_8 FILLER_100_995 ();
 sg13g2_fill_8 FILLER_100_1003 ();
 sg13g2_fill_8 FILLER_100_1011 ();
 sg13g2_fill_8 FILLER_100_1019 ();
 sg13g2_fill_8 FILLER_100_1027 ();
 sg13g2_fill_8 FILLER_100_1035 ();
 sg13g2_fill_8 FILLER_100_1043 ();
 sg13g2_fill_8 FILLER_100_1051 ();
 sg13g2_fill_8 FILLER_100_1059 ();
 sg13g2_fill_8 FILLER_100_1067 ();
 sg13g2_fill_8 FILLER_100_1075 ();
 sg13g2_fill_8 FILLER_100_1083 ();
 sg13g2_fill_8 FILLER_100_1091 ();
 sg13g2_fill_8 FILLER_100_1099 ();
 sg13g2_fill_8 FILLER_100_1107 ();
 sg13g2_fill_8 FILLER_100_1115 ();
 sg13g2_fill_8 FILLER_100_1123 ();
 sg13g2_fill_8 FILLER_100_1131 ();
 sg13g2_fill_4 FILLER_100_1139 ();
 sg13g2_fill_1 FILLER_100_1143 ();
 sg13g2_fill_8 FILLER_101_0 ();
 sg13g2_fill_8 FILLER_101_8 ();
 sg13g2_fill_8 FILLER_101_16 ();
 sg13g2_fill_8 FILLER_101_24 ();
 sg13g2_fill_8 FILLER_101_32 ();
 sg13g2_fill_8 FILLER_101_40 ();
 sg13g2_fill_8 FILLER_101_48 ();
 sg13g2_fill_8 FILLER_101_56 ();
 sg13g2_fill_8 FILLER_101_64 ();
 sg13g2_fill_8 FILLER_101_72 ();
 sg13g2_fill_8 FILLER_101_80 ();
 sg13g2_fill_8 FILLER_101_88 ();
 sg13g2_fill_8 FILLER_101_96 ();
 sg13g2_fill_8 FILLER_101_104 ();
 sg13g2_fill_8 FILLER_101_112 ();
 sg13g2_fill_8 FILLER_101_120 ();
 sg13g2_fill_8 FILLER_101_128 ();
 sg13g2_fill_8 FILLER_101_136 ();
 sg13g2_fill_8 FILLER_101_144 ();
 sg13g2_fill_8 FILLER_101_152 ();
 sg13g2_fill_8 FILLER_101_160 ();
 sg13g2_fill_8 FILLER_101_168 ();
 sg13g2_fill_8 FILLER_101_176 ();
 sg13g2_fill_8 FILLER_101_184 ();
 sg13g2_fill_8 FILLER_101_192 ();
 sg13g2_fill_8 FILLER_101_200 ();
 sg13g2_fill_8 FILLER_101_208 ();
 sg13g2_fill_8 FILLER_101_216 ();
 sg13g2_fill_8 FILLER_101_224 ();
 sg13g2_fill_8 FILLER_101_232 ();
 sg13g2_fill_8 FILLER_101_240 ();
 sg13g2_fill_8 FILLER_101_248 ();
 sg13g2_fill_8 FILLER_101_256 ();
 sg13g2_fill_8 FILLER_101_264 ();
 sg13g2_fill_8 FILLER_101_272 ();
 sg13g2_fill_8 FILLER_101_280 ();
 sg13g2_fill_8 FILLER_101_288 ();
 sg13g2_fill_8 FILLER_101_296 ();
 sg13g2_fill_8 FILLER_101_304 ();
 sg13g2_fill_8 FILLER_101_312 ();
 sg13g2_fill_8 FILLER_101_320 ();
 sg13g2_fill_8 FILLER_101_328 ();
 sg13g2_fill_8 FILLER_101_336 ();
 sg13g2_fill_8 FILLER_101_344 ();
 sg13g2_fill_8 FILLER_101_352 ();
 sg13g2_fill_8 FILLER_101_360 ();
 sg13g2_fill_8 FILLER_101_368 ();
 sg13g2_fill_8 FILLER_101_376 ();
 sg13g2_fill_8 FILLER_101_384 ();
 sg13g2_fill_8 FILLER_101_392 ();
 sg13g2_fill_8 FILLER_101_400 ();
 sg13g2_fill_8 FILLER_101_408 ();
 sg13g2_fill_8 FILLER_101_416 ();
 sg13g2_fill_8 FILLER_101_424 ();
 sg13g2_fill_8 FILLER_101_432 ();
 sg13g2_fill_8 FILLER_101_440 ();
 sg13g2_fill_8 FILLER_101_448 ();
 sg13g2_fill_8 FILLER_101_456 ();
 sg13g2_fill_8 FILLER_101_464 ();
 sg13g2_fill_8 FILLER_101_472 ();
 sg13g2_fill_8 FILLER_101_480 ();
 sg13g2_fill_8 FILLER_101_488 ();
 sg13g2_fill_8 FILLER_101_496 ();
 sg13g2_fill_8 FILLER_101_504 ();
 sg13g2_fill_8 FILLER_101_512 ();
 sg13g2_fill_8 FILLER_101_520 ();
 sg13g2_fill_8 FILLER_101_528 ();
 sg13g2_fill_8 FILLER_101_536 ();
 sg13g2_fill_8 FILLER_101_544 ();
 sg13g2_fill_8 FILLER_101_552 ();
 sg13g2_fill_8 FILLER_101_560 ();
 sg13g2_fill_8 FILLER_101_568 ();
 sg13g2_fill_8 FILLER_101_576 ();
 sg13g2_fill_8 FILLER_101_584 ();
 sg13g2_fill_8 FILLER_101_592 ();
 sg13g2_fill_8 FILLER_101_600 ();
 sg13g2_fill_8 FILLER_101_608 ();
 sg13g2_fill_8 FILLER_101_616 ();
 sg13g2_fill_8 FILLER_101_624 ();
 sg13g2_fill_8 FILLER_101_632 ();
 sg13g2_fill_8 FILLER_101_640 ();
 sg13g2_fill_8 FILLER_101_648 ();
 sg13g2_fill_8 FILLER_101_656 ();
 sg13g2_fill_8 FILLER_101_664 ();
 sg13g2_fill_8 FILLER_101_672 ();
 sg13g2_fill_8 FILLER_101_680 ();
 sg13g2_fill_8 FILLER_101_688 ();
 sg13g2_fill_8 FILLER_101_696 ();
 sg13g2_fill_8 FILLER_101_704 ();
 sg13g2_fill_8 FILLER_101_712 ();
 sg13g2_fill_8 FILLER_101_720 ();
 sg13g2_fill_8 FILLER_101_728 ();
 sg13g2_fill_8 FILLER_101_736 ();
 sg13g2_fill_8 FILLER_101_744 ();
 sg13g2_fill_8 FILLER_101_752 ();
 sg13g2_fill_8 FILLER_101_760 ();
 sg13g2_fill_8 FILLER_101_768 ();
 sg13g2_fill_8 FILLER_101_776 ();
 sg13g2_fill_8 FILLER_101_784 ();
 sg13g2_fill_8 FILLER_101_792 ();
 sg13g2_fill_8 FILLER_101_800 ();
 sg13g2_fill_8 FILLER_101_808 ();
 sg13g2_fill_8 FILLER_101_816 ();
 sg13g2_fill_8 FILLER_101_824 ();
 sg13g2_fill_8 FILLER_101_832 ();
 sg13g2_fill_8 FILLER_101_840 ();
 sg13g2_fill_8 FILLER_101_848 ();
 sg13g2_fill_8 FILLER_101_856 ();
 sg13g2_fill_4 FILLER_101_864 ();
 sg13g2_fill_2 FILLER_101_868 ();
 sg13g2_fill_2 FILLER_101_880 ();
 sg13g2_fill_1 FILLER_101_882 ();
 sg13g2_fill_8 FILLER_101_888 ();
 sg13g2_fill_8 FILLER_101_896 ();
 sg13g2_fill_8 FILLER_101_904 ();
 sg13g2_fill_8 FILLER_101_912 ();
 sg13g2_fill_8 FILLER_101_920 ();
 sg13g2_fill_8 FILLER_101_928 ();
 sg13g2_fill_8 FILLER_101_936 ();
 sg13g2_fill_8 FILLER_101_944 ();
 sg13g2_fill_8 FILLER_101_952 ();
 sg13g2_fill_8 FILLER_101_960 ();
 sg13g2_fill_8 FILLER_101_968 ();
 sg13g2_fill_8 FILLER_101_976 ();
 sg13g2_fill_8 FILLER_101_984 ();
 sg13g2_fill_8 FILLER_101_992 ();
 sg13g2_fill_8 FILLER_101_1000 ();
 sg13g2_fill_8 FILLER_101_1008 ();
 sg13g2_fill_8 FILLER_101_1016 ();
 sg13g2_fill_8 FILLER_101_1024 ();
 sg13g2_fill_8 FILLER_101_1032 ();
 sg13g2_fill_8 FILLER_101_1040 ();
 sg13g2_fill_8 FILLER_101_1048 ();
 sg13g2_fill_8 FILLER_101_1056 ();
 sg13g2_fill_8 FILLER_101_1064 ();
 sg13g2_fill_8 FILLER_101_1072 ();
 sg13g2_fill_8 FILLER_101_1080 ();
 sg13g2_fill_8 FILLER_101_1088 ();
 sg13g2_fill_8 FILLER_101_1096 ();
 sg13g2_fill_8 FILLER_101_1104 ();
 sg13g2_fill_8 FILLER_101_1112 ();
 sg13g2_fill_8 FILLER_101_1120 ();
 sg13g2_fill_8 FILLER_101_1128 ();
 sg13g2_fill_8 FILLER_101_1136 ();
 sg13g2_fill_8 FILLER_102_0 ();
 sg13g2_fill_8 FILLER_102_8 ();
 sg13g2_fill_8 FILLER_102_16 ();
 sg13g2_fill_8 FILLER_102_24 ();
 sg13g2_fill_8 FILLER_102_32 ();
 sg13g2_fill_8 FILLER_102_40 ();
 sg13g2_fill_8 FILLER_102_48 ();
 sg13g2_fill_8 FILLER_102_56 ();
 sg13g2_fill_8 FILLER_102_64 ();
 sg13g2_fill_8 FILLER_102_72 ();
 sg13g2_fill_8 FILLER_102_80 ();
 sg13g2_fill_8 FILLER_102_88 ();
 sg13g2_fill_8 FILLER_102_96 ();
 sg13g2_fill_8 FILLER_102_104 ();
 sg13g2_fill_8 FILLER_102_112 ();
 sg13g2_fill_8 FILLER_102_120 ();
 sg13g2_fill_8 FILLER_102_128 ();
 sg13g2_fill_8 FILLER_102_136 ();
 sg13g2_fill_8 FILLER_102_144 ();
 sg13g2_fill_8 FILLER_102_152 ();
 sg13g2_fill_8 FILLER_102_160 ();
 sg13g2_fill_8 FILLER_102_168 ();
 sg13g2_fill_8 FILLER_102_176 ();
 sg13g2_fill_8 FILLER_102_184 ();
 sg13g2_fill_8 FILLER_102_192 ();
 sg13g2_fill_8 FILLER_102_200 ();
 sg13g2_fill_8 FILLER_102_208 ();
 sg13g2_fill_8 FILLER_102_216 ();
 sg13g2_fill_8 FILLER_102_224 ();
 sg13g2_fill_8 FILLER_102_232 ();
 sg13g2_fill_8 FILLER_102_240 ();
 sg13g2_fill_8 FILLER_102_248 ();
 sg13g2_fill_8 FILLER_102_256 ();
 sg13g2_fill_8 FILLER_102_264 ();
 sg13g2_fill_8 FILLER_102_272 ();
 sg13g2_fill_8 FILLER_102_280 ();
 sg13g2_fill_8 FILLER_102_288 ();
 sg13g2_fill_8 FILLER_102_296 ();
 sg13g2_fill_8 FILLER_102_304 ();
 sg13g2_fill_8 FILLER_102_312 ();
 sg13g2_fill_8 FILLER_102_320 ();
 sg13g2_fill_8 FILLER_102_328 ();
 sg13g2_fill_8 FILLER_102_336 ();
 sg13g2_fill_8 FILLER_102_344 ();
 sg13g2_fill_8 FILLER_102_352 ();
 sg13g2_fill_8 FILLER_102_360 ();
 sg13g2_fill_8 FILLER_102_368 ();
 sg13g2_fill_8 FILLER_102_376 ();
 sg13g2_fill_8 FILLER_102_384 ();
 sg13g2_fill_8 FILLER_102_392 ();
 sg13g2_fill_8 FILLER_102_400 ();
 sg13g2_fill_8 FILLER_102_408 ();
 sg13g2_fill_8 FILLER_102_416 ();
 sg13g2_fill_8 FILLER_102_424 ();
 sg13g2_fill_8 FILLER_102_432 ();
 sg13g2_fill_8 FILLER_102_440 ();
 sg13g2_fill_8 FILLER_102_448 ();
 sg13g2_fill_8 FILLER_102_456 ();
 sg13g2_fill_8 FILLER_102_464 ();
 sg13g2_fill_8 FILLER_102_472 ();
 sg13g2_fill_8 FILLER_102_480 ();
 sg13g2_fill_8 FILLER_102_488 ();
 sg13g2_fill_8 FILLER_102_496 ();
 sg13g2_fill_8 FILLER_102_504 ();
 sg13g2_fill_8 FILLER_102_512 ();
 sg13g2_fill_8 FILLER_102_520 ();
 sg13g2_fill_8 FILLER_102_528 ();
 sg13g2_fill_8 FILLER_102_536 ();
 sg13g2_fill_8 FILLER_102_544 ();
 sg13g2_fill_8 FILLER_102_552 ();
 sg13g2_fill_8 FILLER_102_560 ();
 sg13g2_fill_8 FILLER_102_568 ();
 sg13g2_fill_8 FILLER_102_576 ();
 sg13g2_fill_8 FILLER_102_584 ();
 sg13g2_fill_8 FILLER_102_592 ();
 sg13g2_fill_8 FILLER_102_600 ();
 sg13g2_fill_8 FILLER_102_608 ();
 sg13g2_fill_8 FILLER_102_616 ();
 sg13g2_fill_8 FILLER_102_624 ();
 sg13g2_fill_8 FILLER_102_632 ();
 sg13g2_fill_8 FILLER_102_640 ();
 sg13g2_fill_8 FILLER_102_648 ();
 sg13g2_fill_8 FILLER_102_656 ();
 sg13g2_fill_8 FILLER_102_664 ();
 sg13g2_fill_8 FILLER_102_672 ();
 sg13g2_fill_8 FILLER_102_680 ();
 sg13g2_fill_8 FILLER_102_688 ();
 sg13g2_fill_8 FILLER_102_696 ();
 sg13g2_fill_8 FILLER_102_704 ();
 sg13g2_fill_8 FILLER_102_712 ();
 sg13g2_fill_8 FILLER_102_720 ();
 sg13g2_fill_8 FILLER_102_728 ();
 sg13g2_fill_8 FILLER_102_736 ();
 sg13g2_fill_8 FILLER_102_744 ();
 sg13g2_fill_8 FILLER_102_752 ();
 sg13g2_fill_8 FILLER_102_760 ();
 sg13g2_fill_8 FILLER_102_768 ();
 sg13g2_fill_8 FILLER_102_776 ();
 sg13g2_fill_8 FILLER_102_784 ();
 sg13g2_fill_8 FILLER_102_792 ();
 sg13g2_fill_8 FILLER_102_800 ();
 sg13g2_fill_8 FILLER_102_808 ();
 sg13g2_fill_8 FILLER_102_816 ();
 sg13g2_fill_8 FILLER_102_824 ();
 sg13g2_fill_8 FILLER_102_832 ();
 sg13g2_fill_8 FILLER_102_840 ();
 sg13g2_fill_8 FILLER_102_848 ();
 sg13g2_fill_8 FILLER_102_856 ();
 sg13g2_fill_8 FILLER_102_864 ();
 sg13g2_fill_8 FILLER_102_872 ();
 sg13g2_fill_8 FILLER_102_880 ();
 sg13g2_fill_8 FILLER_102_888 ();
 sg13g2_fill_8 FILLER_102_896 ();
 sg13g2_fill_8 FILLER_102_904 ();
 sg13g2_fill_8 FILLER_102_912 ();
 sg13g2_fill_8 FILLER_102_920 ();
 sg13g2_fill_8 FILLER_102_928 ();
 sg13g2_fill_8 FILLER_102_936 ();
 sg13g2_fill_8 FILLER_102_944 ();
 sg13g2_fill_8 FILLER_102_952 ();
 sg13g2_fill_8 FILLER_102_960 ();
 sg13g2_fill_8 FILLER_102_968 ();
 sg13g2_fill_8 FILLER_102_976 ();
 sg13g2_fill_8 FILLER_102_984 ();
 sg13g2_fill_8 FILLER_102_992 ();
 sg13g2_fill_8 FILLER_102_1000 ();
 sg13g2_fill_8 FILLER_102_1008 ();
 sg13g2_fill_8 FILLER_102_1016 ();
 sg13g2_fill_8 FILLER_102_1024 ();
 sg13g2_fill_8 FILLER_102_1032 ();
 sg13g2_fill_8 FILLER_102_1040 ();
 sg13g2_fill_8 FILLER_102_1048 ();
 sg13g2_fill_8 FILLER_102_1056 ();
 sg13g2_fill_8 FILLER_102_1064 ();
 sg13g2_fill_8 FILLER_102_1072 ();
 sg13g2_fill_8 FILLER_102_1080 ();
 sg13g2_fill_8 FILLER_102_1088 ();
 sg13g2_fill_8 FILLER_102_1096 ();
 sg13g2_fill_8 FILLER_102_1104 ();
 sg13g2_fill_8 FILLER_102_1112 ();
 sg13g2_fill_8 FILLER_102_1120 ();
 sg13g2_fill_8 FILLER_102_1128 ();
 sg13g2_fill_8 FILLER_102_1136 ();
 sg13g2_fill_8 FILLER_103_0 ();
 sg13g2_fill_8 FILLER_103_8 ();
 sg13g2_fill_8 FILLER_103_16 ();
 sg13g2_fill_8 FILLER_103_24 ();
 sg13g2_fill_8 FILLER_103_32 ();
 sg13g2_fill_8 FILLER_103_40 ();
 sg13g2_fill_8 FILLER_103_48 ();
 sg13g2_fill_8 FILLER_103_56 ();
 sg13g2_fill_8 FILLER_103_64 ();
 sg13g2_fill_8 FILLER_103_72 ();
 sg13g2_fill_8 FILLER_103_80 ();
 sg13g2_fill_8 FILLER_103_88 ();
 sg13g2_fill_8 FILLER_103_96 ();
 sg13g2_fill_8 FILLER_103_104 ();
 sg13g2_fill_8 FILLER_103_112 ();
 sg13g2_fill_8 FILLER_103_120 ();
 sg13g2_fill_8 FILLER_103_128 ();
 sg13g2_fill_8 FILLER_103_136 ();
 sg13g2_fill_8 FILLER_103_144 ();
 sg13g2_fill_8 FILLER_103_152 ();
 sg13g2_fill_8 FILLER_103_160 ();
 sg13g2_fill_8 FILLER_103_168 ();
 sg13g2_fill_8 FILLER_103_176 ();
 sg13g2_fill_8 FILLER_103_184 ();
 sg13g2_fill_8 FILLER_103_192 ();
 sg13g2_fill_8 FILLER_103_200 ();
 sg13g2_fill_8 FILLER_103_208 ();
 sg13g2_fill_8 FILLER_103_216 ();
 sg13g2_fill_8 FILLER_103_224 ();
 sg13g2_fill_8 FILLER_103_232 ();
 sg13g2_fill_8 FILLER_103_240 ();
 sg13g2_fill_8 FILLER_103_248 ();
 sg13g2_fill_8 FILLER_103_256 ();
 sg13g2_fill_8 FILLER_103_264 ();
 sg13g2_fill_8 FILLER_103_272 ();
 sg13g2_fill_8 FILLER_103_280 ();
 sg13g2_fill_8 FILLER_103_288 ();
 sg13g2_fill_8 FILLER_103_296 ();
 sg13g2_fill_8 FILLER_103_304 ();
 sg13g2_fill_8 FILLER_103_312 ();
 sg13g2_fill_8 FILLER_103_320 ();
 sg13g2_fill_8 FILLER_103_328 ();
 sg13g2_fill_8 FILLER_103_336 ();
 sg13g2_fill_8 FILLER_103_344 ();
 sg13g2_fill_8 FILLER_103_352 ();
 sg13g2_fill_8 FILLER_103_360 ();
 sg13g2_fill_8 FILLER_103_368 ();
 sg13g2_fill_8 FILLER_103_376 ();
 sg13g2_fill_8 FILLER_103_384 ();
 sg13g2_fill_8 FILLER_103_392 ();
 sg13g2_fill_8 FILLER_103_400 ();
 sg13g2_fill_8 FILLER_103_408 ();
 sg13g2_fill_8 FILLER_103_416 ();
 sg13g2_fill_8 FILLER_103_424 ();
 sg13g2_fill_8 FILLER_103_432 ();
 sg13g2_fill_8 FILLER_103_440 ();
 sg13g2_fill_8 FILLER_103_448 ();
 sg13g2_fill_8 FILLER_103_456 ();
 sg13g2_fill_8 FILLER_103_464 ();
 sg13g2_fill_8 FILLER_103_472 ();
 sg13g2_fill_8 FILLER_103_480 ();
 sg13g2_fill_8 FILLER_103_488 ();
 sg13g2_fill_8 FILLER_103_496 ();
 sg13g2_fill_8 FILLER_103_504 ();
 sg13g2_fill_8 FILLER_103_512 ();
 sg13g2_fill_8 FILLER_103_520 ();
 sg13g2_fill_8 FILLER_103_528 ();
 sg13g2_fill_8 FILLER_103_536 ();
 sg13g2_fill_8 FILLER_103_544 ();
 sg13g2_fill_8 FILLER_103_552 ();
 sg13g2_fill_8 FILLER_103_560 ();
 sg13g2_fill_8 FILLER_103_568 ();
 sg13g2_fill_8 FILLER_103_576 ();
 sg13g2_fill_8 FILLER_103_584 ();
 sg13g2_fill_8 FILLER_103_592 ();
 sg13g2_fill_8 FILLER_103_600 ();
 sg13g2_fill_8 FILLER_103_608 ();
 sg13g2_fill_8 FILLER_103_616 ();
 sg13g2_fill_8 FILLER_103_624 ();
 sg13g2_fill_8 FILLER_103_632 ();
 sg13g2_fill_8 FILLER_103_640 ();
 sg13g2_fill_8 FILLER_103_648 ();
 sg13g2_fill_8 FILLER_103_656 ();
 sg13g2_fill_8 FILLER_103_664 ();
 sg13g2_fill_8 FILLER_103_672 ();
 sg13g2_fill_8 FILLER_103_680 ();
 sg13g2_fill_8 FILLER_103_688 ();
 sg13g2_fill_8 FILLER_103_696 ();
 sg13g2_fill_8 FILLER_103_704 ();
 sg13g2_fill_8 FILLER_103_712 ();
 sg13g2_fill_8 FILLER_103_720 ();
 sg13g2_fill_8 FILLER_103_728 ();
 sg13g2_fill_8 FILLER_103_736 ();
 sg13g2_fill_8 FILLER_103_744 ();
 sg13g2_fill_8 FILLER_103_752 ();
 sg13g2_fill_8 FILLER_103_760 ();
 sg13g2_fill_8 FILLER_103_768 ();
 sg13g2_fill_8 FILLER_103_776 ();
 sg13g2_fill_8 FILLER_103_784 ();
 sg13g2_fill_8 FILLER_103_792 ();
 sg13g2_fill_8 FILLER_103_800 ();
 sg13g2_fill_8 FILLER_103_808 ();
 sg13g2_fill_8 FILLER_103_816 ();
 sg13g2_fill_8 FILLER_103_824 ();
 sg13g2_fill_8 FILLER_103_832 ();
 sg13g2_fill_8 FILLER_103_840 ();
 sg13g2_fill_8 FILLER_103_848 ();
 sg13g2_fill_8 FILLER_103_856 ();
 sg13g2_fill_8 FILLER_103_864 ();
 sg13g2_fill_8 FILLER_103_872 ();
 sg13g2_fill_8 FILLER_103_880 ();
 sg13g2_fill_8 FILLER_103_888 ();
 sg13g2_fill_8 FILLER_103_896 ();
 sg13g2_fill_8 FILLER_103_904 ();
 sg13g2_fill_8 FILLER_103_912 ();
 sg13g2_fill_8 FILLER_103_920 ();
 sg13g2_fill_8 FILLER_103_928 ();
 sg13g2_fill_8 FILLER_103_936 ();
 sg13g2_fill_8 FILLER_103_944 ();
 sg13g2_fill_8 FILLER_103_952 ();
 sg13g2_fill_8 FILLER_103_960 ();
 sg13g2_fill_8 FILLER_103_968 ();
 sg13g2_fill_8 FILLER_103_976 ();
 sg13g2_fill_8 FILLER_103_984 ();
 sg13g2_fill_8 FILLER_103_992 ();
 sg13g2_fill_8 FILLER_103_1000 ();
 sg13g2_fill_8 FILLER_103_1008 ();
 sg13g2_fill_8 FILLER_103_1016 ();
 sg13g2_fill_8 FILLER_103_1024 ();
 sg13g2_fill_8 FILLER_103_1032 ();
 sg13g2_fill_8 FILLER_103_1040 ();
 sg13g2_fill_8 FILLER_103_1048 ();
 sg13g2_fill_8 FILLER_103_1056 ();
 sg13g2_fill_8 FILLER_103_1064 ();
 sg13g2_fill_8 FILLER_103_1072 ();
 sg13g2_fill_8 FILLER_103_1080 ();
 sg13g2_fill_8 FILLER_103_1088 ();
 sg13g2_fill_8 FILLER_103_1096 ();
 sg13g2_fill_8 FILLER_103_1104 ();
 sg13g2_fill_8 FILLER_103_1112 ();
 sg13g2_fill_8 FILLER_103_1120 ();
 sg13g2_fill_8 FILLER_103_1128 ();
 sg13g2_fill_8 FILLER_103_1136 ();
 sg13g2_fill_8 FILLER_104_0 ();
 sg13g2_fill_8 FILLER_104_8 ();
 sg13g2_fill_8 FILLER_104_16 ();
 sg13g2_fill_8 FILLER_104_24 ();
 sg13g2_fill_8 FILLER_104_32 ();
 sg13g2_fill_8 FILLER_104_40 ();
 sg13g2_fill_8 FILLER_104_48 ();
 sg13g2_fill_8 FILLER_104_56 ();
 sg13g2_fill_8 FILLER_104_64 ();
 sg13g2_fill_8 FILLER_104_72 ();
 sg13g2_fill_8 FILLER_104_80 ();
 sg13g2_fill_8 FILLER_104_88 ();
 sg13g2_fill_8 FILLER_104_96 ();
 sg13g2_fill_8 FILLER_104_104 ();
 sg13g2_fill_8 FILLER_104_112 ();
 sg13g2_fill_8 FILLER_104_120 ();
 sg13g2_fill_8 FILLER_104_128 ();
 sg13g2_fill_8 FILLER_104_136 ();
 sg13g2_fill_8 FILLER_104_144 ();
 sg13g2_fill_8 FILLER_104_152 ();
 sg13g2_fill_8 FILLER_104_160 ();
 sg13g2_fill_8 FILLER_104_168 ();
 sg13g2_fill_8 FILLER_104_176 ();
 sg13g2_fill_8 FILLER_104_184 ();
 sg13g2_fill_8 FILLER_104_192 ();
 sg13g2_fill_8 FILLER_104_200 ();
 sg13g2_fill_8 FILLER_104_208 ();
 sg13g2_fill_8 FILLER_104_216 ();
 sg13g2_fill_8 FILLER_104_224 ();
 sg13g2_fill_8 FILLER_104_232 ();
 sg13g2_fill_8 FILLER_104_240 ();
 sg13g2_fill_8 FILLER_104_248 ();
 sg13g2_fill_8 FILLER_104_256 ();
 sg13g2_fill_8 FILLER_104_264 ();
 sg13g2_fill_8 FILLER_104_272 ();
 sg13g2_fill_8 FILLER_104_280 ();
 sg13g2_fill_8 FILLER_104_288 ();
 sg13g2_fill_8 FILLER_104_296 ();
 sg13g2_fill_8 FILLER_104_304 ();
 sg13g2_fill_8 FILLER_104_312 ();
 sg13g2_fill_8 FILLER_104_320 ();
 sg13g2_fill_8 FILLER_104_328 ();
 sg13g2_fill_8 FILLER_104_336 ();
 sg13g2_fill_8 FILLER_104_344 ();
 sg13g2_fill_8 FILLER_104_352 ();
 sg13g2_fill_8 FILLER_104_360 ();
 sg13g2_fill_8 FILLER_104_368 ();
 sg13g2_fill_8 FILLER_104_376 ();
 sg13g2_fill_8 FILLER_104_384 ();
 sg13g2_fill_8 FILLER_104_392 ();
 sg13g2_fill_8 FILLER_104_400 ();
 sg13g2_fill_8 FILLER_104_408 ();
 sg13g2_fill_8 FILLER_104_416 ();
 sg13g2_fill_8 FILLER_104_424 ();
 sg13g2_fill_8 FILLER_104_432 ();
 sg13g2_fill_8 FILLER_104_440 ();
 sg13g2_fill_8 FILLER_104_448 ();
 sg13g2_fill_8 FILLER_104_456 ();
 sg13g2_fill_8 FILLER_104_464 ();
 sg13g2_fill_8 FILLER_104_472 ();
 sg13g2_fill_8 FILLER_104_480 ();
 sg13g2_fill_8 FILLER_104_488 ();
 sg13g2_fill_8 FILLER_104_496 ();
 sg13g2_fill_8 FILLER_104_504 ();
 sg13g2_fill_8 FILLER_104_512 ();
 sg13g2_fill_8 FILLER_104_520 ();
 sg13g2_fill_8 FILLER_104_528 ();
 sg13g2_fill_8 FILLER_104_536 ();
 sg13g2_fill_8 FILLER_104_544 ();
 sg13g2_fill_8 FILLER_104_552 ();
 sg13g2_fill_8 FILLER_104_560 ();
 sg13g2_fill_8 FILLER_104_568 ();
 sg13g2_fill_8 FILLER_104_576 ();
 sg13g2_fill_8 FILLER_104_584 ();
 sg13g2_fill_8 FILLER_104_592 ();
 sg13g2_fill_8 FILLER_104_600 ();
 sg13g2_fill_8 FILLER_104_608 ();
 sg13g2_fill_8 FILLER_104_616 ();
 sg13g2_fill_8 FILLER_104_624 ();
 sg13g2_fill_8 FILLER_104_632 ();
 sg13g2_fill_8 FILLER_104_640 ();
 sg13g2_fill_8 FILLER_104_648 ();
 sg13g2_fill_8 FILLER_104_656 ();
 sg13g2_fill_8 FILLER_104_664 ();
 sg13g2_fill_8 FILLER_104_672 ();
 sg13g2_fill_8 FILLER_104_680 ();
 sg13g2_fill_8 FILLER_104_688 ();
 sg13g2_fill_8 FILLER_104_696 ();
 sg13g2_fill_8 FILLER_104_704 ();
 sg13g2_fill_8 FILLER_104_712 ();
 sg13g2_fill_8 FILLER_104_720 ();
 sg13g2_fill_8 FILLER_104_728 ();
 sg13g2_fill_8 FILLER_104_736 ();
 sg13g2_fill_8 FILLER_104_744 ();
 sg13g2_fill_8 FILLER_104_752 ();
 sg13g2_fill_8 FILLER_104_760 ();
 sg13g2_fill_8 FILLER_104_768 ();
 sg13g2_fill_8 FILLER_104_776 ();
 sg13g2_fill_8 FILLER_104_784 ();
 sg13g2_fill_8 FILLER_104_792 ();
 sg13g2_fill_8 FILLER_104_800 ();
 sg13g2_fill_8 FILLER_104_808 ();
 sg13g2_fill_8 FILLER_104_816 ();
 sg13g2_fill_8 FILLER_104_824 ();
 sg13g2_fill_8 FILLER_104_832 ();
 sg13g2_fill_8 FILLER_104_840 ();
 sg13g2_fill_8 FILLER_104_848 ();
 sg13g2_fill_8 FILLER_104_856 ();
 sg13g2_fill_8 FILLER_104_864 ();
 sg13g2_fill_8 FILLER_104_872 ();
 sg13g2_fill_8 FILLER_104_880 ();
 sg13g2_fill_8 FILLER_104_888 ();
 sg13g2_fill_8 FILLER_104_896 ();
 sg13g2_fill_8 FILLER_104_904 ();
 sg13g2_fill_8 FILLER_104_912 ();
 sg13g2_fill_8 FILLER_104_920 ();
 sg13g2_fill_8 FILLER_104_928 ();
 sg13g2_fill_8 FILLER_104_936 ();
 sg13g2_fill_8 FILLER_104_944 ();
 sg13g2_fill_8 FILLER_104_952 ();
 sg13g2_fill_8 FILLER_104_960 ();
 sg13g2_fill_8 FILLER_104_968 ();
 sg13g2_fill_8 FILLER_104_976 ();
 sg13g2_fill_8 FILLER_104_984 ();
 sg13g2_fill_8 FILLER_104_992 ();
 sg13g2_fill_8 FILLER_104_1000 ();
 sg13g2_fill_8 FILLER_104_1008 ();
 sg13g2_fill_8 FILLER_104_1016 ();
 sg13g2_fill_8 FILLER_104_1024 ();
 sg13g2_fill_8 FILLER_104_1032 ();
 sg13g2_fill_8 FILLER_104_1040 ();
 sg13g2_fill_8 FILLER_104_1048 ();
 sg13g2_fill_8 FILLER_104_1056 ();
 sg13g2_fill_8 FILLER_104_1064 ();
 sg13g2_fill_8 FILLER_104_1072 ();
 sg13g2_fill_8 FILLER_104_1080 ();
 sg13g2_fill_8 FILLER_104_1088 ();
 sg13g2_fill_8 FILLER_104_1096 ();
 sg13g2_fill_8 FILLER_104_1104 ();
 sg13g2_fill_8 FILLER_104_1112 ();
 sg13g2_fill_8 FILLER_104_1120 ();
 sg13g2_fill_8 FILLER_104_1128 ();
 sg13g2_fill_8 FILLER_104_1136 ();
 sg13g2_fill_8 FILLER_105_0 ();
 sg13g2_fill_8 FILLER_105_8 ();
 sg13g2_fill_8 FILLER_105_16 ();
 sg13g2_fill_8 FILLER_105_24 ();
 sg13g2_fill_8 FILLER_105_32 ();
 sg13g2_fill_8 FILLER_105_40 ();
 sg13g2_fill_8 FILLER_105_48 ();
 sg13g2_fill_8 FILLER_105_56 ();
 sg13g2_fill_8 FILLER_105_64 ();
 sg13g2_fill_8 FILLER_105_72 ();
 sg13g2_fill_8 FILLER_105_80 ();
 sg13g2_fill_8 FILLER_105_88 ();
 sg13g2_fill_8 FILLER_105_96 ();
 sg13g2_fill_8 FILLER_105_104 ();
 sg13g2_fill_8 FILLER_105_112 ();
 sg13g2_fill_8 FILLER_105_120 ();
 sg13g2_fill_8 FILLER_105_128 ();
 sg13g2_fill_8 FILLER_105_136 ();
 sg13g2_fill_8 FILLER_105_144 ();
 sg13g2_fill_8 FILLER_105_152 ();
 sg13g2_fill_8 FILLER_105_160 ();
 sg13g2_fill_8 FILLER_105_168 ();
 sg13g2_fill_8 FILLER_105_176 ();
 sg13g2_fill_8 FILLER_105_184 ();
 sg13g2_fill_8 FILLER_105_192 ();
 sg13g2_fill_8 FILLER_105_200 ();
 sg13g2_fill_8 FILLER_105_208 ();
 sg13g2_fill_8 FILLER_105_216 ();
 sg13g2_fill_8 FILLER_105_224 ();
 sg13g2_fill_8 FILLER_105_232 ();
 sg13g2_fill_8 FILLER_105_240 ();
 sg13g2_fill_8 FILLER_105_248 ();
 sg13g2_fill_8 FILLER_105_256 ();
 sg13g2_fill_8 FILLER_105_264 ();
 sg13g2_fill_8 FILLER_105_272 ();
 sg13g2_fill_8 FILLER_105_280 ();
 sg13g2_fill_8 FILLER_105_288 ();
 sg13g2_fill_8 FILLER_105_296 ();
 sg13g2_fill_8 FILLER_105_304 ();
 sg13g2_fill_8 FILLER_105_312 ();
 sg13g2_fill_8 FILLER_105_320 ();
 sg13g2_fill_8 FILLER_105_328 ();
 sg13g2_fill_8 FILLER_105_336 ();
 sg13g2_fill_8 FILLER_105_344 ();
 sg13g2_fill_8 FILLER_105_352 ();
 sg13g2_fill_8 FILLER_105_360 ();
 sg13g2_fill_8 FILLER_105_368 ();
 sg13g2_fill_8 FILLER_105_376 ();
 sg13g2_fill_8 FILLER_105_384 ();
 sg13g2_fill_8 FILLER_105_392 ();
 sg13g2_fill_8 FILLER_105_400 ();
 sg13g2_fill_8 FILLER_105_408 ();
 sg13g2_fill_8 FILLER_105_416 ();
 sg13g2_fill_8 FILLER_105_424 ();
 sg13g2_fill_8 FILLER_105_432 ();
 sg13g2_fill_8 FILLER_105_440 ();
 sg13g2_fill_8 FILLER_105_448 ();
 sg13g2_fill_8 FILLER_105_456 ();
 sg13g2_fill_8 FILLER_105_464 ();
 sg13g2_fill_8 FILLER_105_472 ();
 sg13g2_fill_8 FILLER_105_480 ();
 sg13g2_fill_8 FILLER_105_488 ();
 sg13g2_fill_8 FILLER_105_496 ();
 sg13g2_fill_8 FILLER_105_504 ();
 sg13g2_fill_8 FILLER_105_512 ();
 sg13g2_fill_8 FILLER_105_520 ();
 sg13g2_fill_8 FILLER_105_528 ();
 sg13g2_fill_8 FILLER_105_536 ();
 sg13g2_fill_8 FILLER_105_544 ();
 sg13g2_fill_8 FILLER_105_552 ();
 sg13g2_fill_8 FILLER_105_560 ();
 sg13g2_fill_8 FILLER_105_568 ();
 sg13g2_fill_8 FILLER_105_576 ();
 sg13g2_fill_8 FILLER_105_584 ();
 sg13g2_fill_8 FILLER_105_592 ();
 sg13g2_fill_8 FILLER_105_600 ();
 sg13g2_fill_8 FILLER_105_608 ();
 sg13g2_fill_8 FILLER_105_616 ();
 sg13g2_fill_8 FILLER_105_624 ();
 sg13g2_fill_8 FILLER_105_632 ();
 sg13g2_fill_8 FILLER_105_640 ();
 sg13g2_fill_8 FILLER_105_648 ();
 sg13g2_fill_8 FILLER_105_656 ();
 sg13g2_fill_8 FILLER_105_664 ();
 sg13g2_fill_8 FILLER_105_672 ();
 sg13g2_fill_8 FILLER_105_680 ();
 sg13g2_fill_8 FILLER_105_688 ();
 sg13g2_fill_8 FILLER_105_696 ();
 sg13g2_fill_8 FILLER_105_704 ();
 sg13g2_fill_8 FILLER_105_712 ();
 sg13g2_fill_8 FILLER_105_720 ();
 sg13g2_fill_8 FILLER_105_728 ();
 sg13g2_fill_8 FILLER_105_736 ();
 sg13g2_fill_8 FILLER_105_744 ();
 sg13g2_fill_8 FILLER_105_752 ();
 sg13g2_fill_8 FILLER_105_760 ();
 sg13g2_fill_8 FILLER_105_768 ();
 sg13g2_fill_8 FILLER_105_776 ();
 sg13g2_fill_8 FILLER_105_784 ();
 sg13g2_fill_8 FILLER_105_792 ();
 sg13g2_fill_8 FILLER_105_800 ();
 sg13g2_fill_8 FILLER_105_808 ();
 sg13g2_fill_8 FILLER_105_816 ();
 sg13g2_fill_8 FILLER_105_824 ();
 sg13g2_fill_8 FILLER_105_832 ();
 sg13g2_fill_8 FILLER_105_840 ();
 sg13g2_fill_8 FILLER_105_848 ();
 sg13g2_fill_8 FILLER_105_856 ();
 sg13g2_fill_8 FILLER_105_864 ();
 sg13g2_fill_8 FILLER_105_872 ();
 sg13g2_fill_8 FILLER_105_880 ();
 sg13g2_fill_8 FILLER_105_888 ();
 sg13g2_fill_8 FILLER_105_896 ();
 sg13g2_fill_8 FILLER_105_904 ();
 sg13g2_fill_8 FILLER_105_912 ();
 sg13g2_fill_8 FILLER_105_920 ();
 sg13g2_fill_8 FILLER_105_928 ();
 sg13g2_fill_8 FILLER_105_936 ();
 sg13g2_fill_8 FILLER_105_944 ();
 sg13g2_fill_8 FILLER_105_952 ();
 sg13g2_fill_8 FILLER_105_960 ();
 sg13g2_fill_8 FILLER_105_968 ();
 sg13g2_fill_8 FILLER_105_976 ();
 sg13g2_fill_8 FILLER_105_984 ();
 sg13g2_fill_8 FILLER_105_992 ();
 sg13g2_fill_8 FILLER_105_1000 ();
 sg13g2_fill_8 FILLER_105_1008 ();
 sg13g2_fill_8 FILLER_105_1016 ();
 sg13g2_fill_8 FILLER_105_1024 ();
 sg13g2_fill_8 FILLER_105_1032 ();
 sg13g2_fill_8 FILLER_105_1040 ();
 sg13g2_fill_8 FILLER_105_1048 ();
 sg13g2_fill_8 FILLER_105_1056 ();
 sg13g2_fill_8 FILLER_105_1064 ();
 sg13g2_fill_8 FILLER_105_1072 ();
 sg13g2_fill_8 FILLER_105_1080 ();
 sg13g2_fill_8 FILLER_105_1088 ();
 sg13g2_fill_8 FILLER_105_1096 ();
 sg13g2_fill_8 FILLER_105_1104 ();
 sg13g2_fill_8 FILLER_105_1112 ();
 sg13g2_fill_8 FILLER_105_1120 ();
 sg13g2_fill_8 FILLER_105_1128 ();
 sg13g2_fill_8 FILLER_105_1136 ();
 sg13g2_fill_8 FILLER_106_0 ();
 sg13g2_fill_8 FILLER_106_8 ();
 sg13g2_fill_8 FILLER_106_16 ();
 sg13g2_fill_8 FILLER_106_24 ();
 sg13g2_fill_8 FILLER_106_32 ();
 sg13g2_fill_8 FILLER_106_40 ();
 sg13g2_fill_8 FILLER_106_48 ();
 sg13g2_fill_8 FILLER_106_56 ();
 sg13g2_fill_8 FILLER_106_64 ();
 sg13g2_fill_8 FILLER_106_72 ();
 sg13g2_fill_8 FILLER_106_80 ();
 sg13g2_fill_8 FILLER_106_88 ();
 sg13g2_fill_8 FILLER_106_96 ();
 sg13g2_fill_8 FILLER_106_104 ();
 sg13g2_fill_8 FILLER_106_112 ();
 sg13g2_fill_8 FILLER_106_120 ();
 sg13g2_fill_8 FILLER_106_128 ();
 sg13g2_fill_8 FILLER_106_136 ();
 sg13g2_fill_8 FILLER_106_144 ();
 sg13g2_fill_8 FILLER_106_152 ();
 sg13g2_fill_8 FILLER_106_160 ();
 sg13g2_fill_8 FILLER_106_168 ();
 sg13g2_fill_8 FILLER_106_176 ();
 sg13g2_fill_8 FILLER_106_184 ();
 sg13g2_fill_8 FILLER_106_192 ();
 sg13g2_fill_8 FILLER_106_200 ();
 sg13g2_fill_8 FILLER_106_208 ();
 sg13g2_fill_8 FILLER_106_216 ();
 sg13g2_fill_8 FILLER_106_224 ();
 sg13g2_fill_8 FILLER_106_232 ();
 sg13g2_fill_8 FILLER_106_240 ();
 sg13g2_fill_8 FILLER_106_248 ();
 sg13g2_fill_8 FILLER_106_256 ();
 sg13g2_fill_8 FILLER_106_264 ();
 sg13g2_fill_8 FILLER_106_272 ();
 sg13g2_fill_8 FILLER_106_280 ();
 sg13g2_fill_8 FILLER_106_288 ();
 sg13g2_fill_8 FILLER_106_296 ();
 sg13g2_fill_8 FILLER_106_304 ();
 sg13g2_fill_8 FILLER_106_312 ();
 sg13g2_fill_8 FILLER_106_320 ();
 sg13g2_fill_8 FILLER_106_328 ();
 sg13g2_fill_8 FILLER_106_336 ();
 sg13g2_fill_8 FILLER_106_344 ();
 sg13g2_fill_8 FILLER_106_352 ();
 sg13g2_fill_8 FILLER_106_360 ();
 sg13g2_fill_8 FILLER_106_368 ();
 sg13g2_fill_8 FILLER_106_376 ();
 sg13g2_fill_8 FILLER_106_384 ();
 sg13g2_fill_8 FILLER_106_392 ();
 sg13g2_fill_8 FILLER_106_400 ();
 sg13g2_fill_8 FILLER_106_408 ();
 sg13g2_fill_8 FILLER_106_416 ();
 sg13g2_fill_8 FILLER_106_424 ();
 sg13g2_fill_8 FILLER_106_432 ();
 sg13g2_fill_8 FILLER_106_440 ();
 sg13g2_fill_8 FILLER_106_448 ();
 sg13g2_fill_8 FILLER_106_456 ();
 sg13g2_fill_8 FILLER_106_464 ();
 sg13g2_fill_8 FILLER_106_472 ();
 sg13g2_fill_8 FILLER_106_480 ();
 sg13g2_fill_8 FILLER_106_488 ();
 sg13g2_fill_8 FILLER_106_496 ();
 sg13g2_fill_8 FILLER_106_504 ();
 sg13g2_fill_8 FILLER_106_512 ();
 sg13g2_fill_8 FILLER_106_520 ();
 sg13g2_fill_8 FILLER_106_528 ();
 sg13g2_fill_8 FILLER_106_536 ();
 sg13g2_fill_8 FILLER_106_544 ();
 sg13g2_fill_8 FILLER_106_552 ();
 sg13g2_fill_8 FILLER_106_560 ();
 sg13g2_fill_8 FILLER_106_568 ();
 sg13g2_fill_8 FILLER_106_576 ();
 sg13g2_fill_8 FILLER_106_584 ();
 sg13g2_fill_8 FILLER_106_592 ();
 sg13g2_fill_8 FILLER_106_600 ();
 sg13g2_fill_8 FILLER_106_608 ();
 sg13g2_fill_8 FILLER_106_616 ();
 sg13g2_fill_8 FILLER_106_624 ();
 sg13g2_fill_8 FILLER_106_632 ();
 sg13g2_fill_8 FILLER_106_640 ();
 sg13g2_fill_8 FILLER_106_648 ();
 sg13g2_fill_8 FILLER_106_656 ();
 sg13g2_fill_8 FILLER_106_664 ();
 sg13g2_fill_8 FILLER_106_672 ();
 sg13g2_fill_8 FILLER_106_680 ();
 sg13g2_fill_8 FILLER_106_688 ();
 sg13g2_fill_8 FILLER_106_696 ();
 sg13g2_fill_8 FILLER_106_704 ();
 sg13g2_fill_8 FILLER_106_712 ();
 sg13g2_fill_8 FILLER_106_720 ();
 sg13g2_fill_8 FILLER_106_728 ();
 sg13g2_fill_8 FILLER_106_736 ();
 sg13g2_fill_8 FILLER_106_744 ();
 sg13g2_fill_8 FILLER_106_752 ();
 sg13g2_fill_8 FILLER_106_760 ();
 sg13g2_fill_8 FILLER_106_768 ();
 sg13g2_fill_8 FILLER_106_776 ();
 sg13g2_fill_8 FILLER_106_784 ();
 sg13g2_fill_8 FILLER_106_792 ();
 sg13g2_fill_8 FILLER_106_800 ();
 sg13g2_fill_8 FILLER_106_808 ();
 sg13g2_fill_8 FILLER_106_816 ();
 sg13g2_fill_8 FILLER_106_824 ();
 sg13g2_fill_8 FILLER_106_832 ();
 sg13g2_fill_8 FILLER_106_840 ();
 sg13g2_fill_8 FILLER_106_848 ();
 sg13g2_fill_8 FILLER_106_856 ();
 sg13g2_fill_8 FILLER_106_864 ();
 sg13g2_fill_8 FILLER_106_872 ();
 sg13g2_fill_8 FILLER_106_880 ();
 sg13g2_fill_8 FILLER_106_888 ();
 sg13g2_fill_8 FILLER_106_896 ();
 sg13g2_fill_8 FILLER_106_904 ();
 sg13g2_fill_8 FILLER_106_912 ();
 sg13g2_fill_8 FILLER_106_920 ();
 sg13g2_fill_8 FILLER_106_928 ();
 sg13g2_fill_8 FILLER_106_936 ();
 sg13g2_fill_8 FILLER_106_944 ();
 sg13g2_fill_8 FILLER_106_952 ();
 sg13g2_fill_8 FILLER_106_960 ();
 sg13g2_fill_8 FILLER_106_968 ();
 sg13g2_fill_8 FILLER_106_976 ();
 sg13g2_fill_8 FILLER_106_984 ();
 sg13g2_fill_8 FILLER_106_992 ();
 sg13g2_fill_8 FILLER_106_1000 ();
 sg13g2_fill_8 FILLER_106_1008 ();
 sg13g2_fill_8 FILLER_106_1016 ();
 sg13g2_fill_8 FILLER_106_1024 ();
 sg13g2_fill_8 FILLER_106_1032 ();
 sg13g2_fill_8 FILLER_106_1040 ();
 sg13g2_fill_8 FILLER_106_1048 ();
 sg13g2_fill_8 FILLER_106_1056 ();
 sg13g2_fill_8 FILLER_106_1064 ();
 sg13g2_fill_8 FILLER_106_1072 ();
 sg13g2_fill_8 FILLER_106_1080 ();
 sg13g2_fill_8 FILLER_106_1088 ();
 sg13g2_fill_8 FILLER_106_1096 ();
 sg13g2_fill_8 FILLER_106_1104 ();
 sg13g2_fill_8 FILLER_106_1112 ();
 sg13g2_fill_8 FILLER_106_1120 ();
 sg13g2_fill_8 FILLER_106_1128 ();
 sg13g2_fill_8 FILLER_106_1136 ();
 sg13g2_fill_8 FILLER_107_0 ();
 sg13g2_fill_8 FILLER_107_8 ();
 sg13g2_fill_8 FILLER_107_16 ();
 sg13g2_fill_8 FILLER_107_24 ();
 sg13g2_fill_8 FILLER_107_32 ();
 sg13g2_fill_8 FILLER_107_40 ();
 sg13g2_fill_8 FILLER_107_48 ();
 sg13g2_fill_8 FILLER_107_56 ();
 sg13g2_fill_8 FILLER_107_64 ();
 sg13g2_fill_8 FILLER_107_72 ();
 sg13g2_fill_8 FILLER_107_80 ();
 sg13g2_fill_8 FILLER_107_88 ();
 sg13g2_fill_8 FILLER_107_96 ();
 sg13g2_fill_8 FILLER_107_104 ();
 sg13g2_fill_8 FILLER_107_112 ();
 sg13g2_fill_8 FILLER_107_120 ();
 sg13g2_fill_8 FILLER_107_128 ();
 sg13g2_fill_8 FILLER_107_136 ();
 sg13g2_fill_8 FILLER_107_144 ();
 sg13g2_fill_8 FILLER_107_152 ();
 sg13g2_fill_8 FILLER_107_160 ();
 sg13g2_fill_8 FILLER_107_168 ();
 sg13g2_fill_8 FILLER_107_176 ();
 sg13g2_fill_8 FILLER_107_184 ();
 sg13g2_fill_8 FILLER_107_192 ();
 sg13g2_fill_8 FILLER_107_200 ();
 sg13g2_fill_8 FILLER_107_208 ();
 sg13g2_fill_8 FILLER_107_216 ();
 sg13g2_fill_8 FILLER_107_224 ();
 sg13g2_fill_8 FILLER_107_232 ();
 sg13g2_fill_8 FILLER_107_240 ();
 sg13g2_fill_8 FILLER_107_248 ();
 sg13g2_fill_8 FILLER_107_256 ();
 sg13g2_fill_8 FILLER_107_264 ();
 sg13g2_fill_8 FILLER_107_272 ();
 sg13g2_fill_8 FILLER_107_280 ();
 sg13g2_fill_8 FILLER_107_288 ();
 sg13g2_fill_8 FILLER_107_296 ();
 sg13g2_fill_8 FILLER_107_304 ();
 sg13g2_fill_8 FILLER_107_312 ();
 sg13g2_fill_8 FILLER_107_320 ();
 sg13g2_fill_8 FILLER_107_328 ();
 sg13g2_fill_8 FILLER_107_336 ();
 sg13g2_fill_8 FILLER_107_344 ();
 sg13g2_fill_8 FILLER_107_352 ();
 sg13g2_fill_8 FILLER_107_360 ();
 sg13g2_fill_8 FILLER_107_368 ();
 sg13g2_fill_8 FILLER_107_376 ();
 sg13g2_fill_8 FILLER_107_384 ();
 sg13g2_fill_8 FILLER_107_392 ();
 sg13g2_fill_8 FILLER_107_400 ();
 sg13g2_fill_8 FILLER_107_408 ();
 sg13g2_fill_8 FILLER_107_416 ();
 sg13g2_fill_8 FILLER_107_424 ();
 sg13g2_fill_8 FILLER_107_432 ();
 sg13g2_fill_8 FILLER_107_440 ();
 sg13g2_fill_8 FILLER_107_448 ();
 sg13g2_fill_8 FILLER_107_456 ();
 sg13g2_fill_8 FILLER_107_464 ();
 sg13g2_fill_8 FILLER_107_472 ();
 sg13g2_fill_8 FILLER_107_480 ();
 sg13g2_fill_8 FILLER_107_488 ();
 sg13g2_fill_8 FILLER_107_496 ();
 sg13g2_fill_8 FILLER_107_504 ();
 sg13g2_fill_8 FILLER_107_512 ();
 sg13g2_fill_8 FILLER_107_520 ();
 sg13g2_fill_8 FILLER_107_528 ();
 sg13g2_fill_8 FILLER_107_536 ();
 sg13g2_fill_8 FILLER_107_544 ();
 sg13g2_fill_8 FILLER_107_552 ();
 sg13g2_fill_8 FILLER_107_560 ();
 sg13g2_fill_8 FILLER_107_568 ();
 sg13g2_fill_8 FILLER_107_576 ();
 sg13g2_fill_8 FILLER_107_584 ();
 sg13g2_fill_8 FILLER_107_592 ();
 sg13g2_fill_8 FILLER_107_600 ();
 sg13g2_fill_8 FILLER_107_608 ();
 sg13g2_fill_8 FILLER_107_616 ();
 sg13g2_fill_8 FILLER_107_624 ();
 sg13g2_fill_8 FILLER_107_632 ();
 sg13g2_fill_8 FILLER_107_640 ();
 sg13g2_fill_8 FILLER_107_648 ();
 sg13g2_fill_8 FILLER_107_656 ();
 sg13g2_fill_8 FILLER_107_664 ();
 sg13g2_fill_8 FILLER_107_672 ();
 sg13g2_fill_8 FILLER_107_680 ();
 sg13g2_fill_8 FILLER_107_688 ();
 sg13g2_fill_8 FILLER_107_696 ();
 sg13g2_fill_8 FILLER_107_704 ();
 sg13g2_fill_8 FILLER_107_712 ();
 sg13g2_fill_8 FILLER_107_720 ();
 sg13g2_fill_8 FILLER_107_728 ();
 sg13g2_fill_8 FILLER_107_736 ();
 sg13g2_fill_8 FILLER_107_744 ();
 sg13g2_fill_8 FILLER_107_752 ();
 sg13g2_fill_8 FILLER_107_760 ();
 sg13g2_fill_8 FILLER_107_768 ();
 sg13g2_fill_8 FILLER_107_776 ();
 sg13g2_fill_8 FILLER_107_784 ();
 sg13g2_fill_8 FILLER_107_792 ();
 sg13g2_fill_8 FILLER_107_800 ();
 sg13g2_fill_8 FILLER_107_808 ();
 sg13g2_fill_8 FILLER_107_816 ();
 sg13g2_fill_8 FILLER_107_824 ();
 sg13g2_fill_8 FILLER_107_832 ();
 sg13g2_fill_8 FILLER_107_840 ();
 sg13g2_fill_8 FILLER_107_848 ();
 sg13g2_fill_8 FILLER_107_856 ();
 sg13g2_fill_8 FILLER_107_864 ();
 sg13g2_fill_8 FILLER_107_872 ();
 sg13g2_fill_8 FILLER_107_880 ();
 sg13g2_fill_8 FILLER_107_888 ();
 sg13g2_fill_8 FILLER_107_896 ();
 sg13g2_fill_8 FILLER_107_904 ();
 sg13g2_fill_8 FILLER_107_912 ();
 sg13g2_fill_8 FILLER_107_920 ();
 sg13g2_fill_8 FILLER_107_928 ();
 sg13g2_fill_8 FILLER_107_936 ();
 sg13g2_fill_8 FILLER_107_944 ();
 sg13g2_fill_8 FILLER_107_952 ();
 sg13g2_fill_8 FILLER_107_960 ();
 sg13g2_fill_8 FILLER_107_968 ();
 sg13g2_fill_8 FILLER_107_976 ();
 sg13g2_fill_8 FILLER_107_984 ();
 sg13g2_fill_8 FILLER_107_992 ();
 sg13g2_fill_8 FILLER_107_1000 ();
 sg13g2_fill_8 FILLER_107_1008 ();
 sg13g2_fill_8 FILLER_107_1016 ();
 sg13g2_fill_8 FILLER_107_1024 ();
 sg13g2_fill_8 FILLER_107_1032 ();
 sg13g2_fill_8 FILLER_107_1040 ();
 sg13g2_fill_8 FILLER_107_1048 ();
 sg13g2_fill_8 FILLER_107_1056 ();
 sg13g2_fill_8 FILLER_107_1064 ();
 sg13g2_fill_8 FILLER_107_1072 ();
 sg13g2_fill_8 FILLER_107_1080 ();
 sg13g2_fill_8 FILLER_107_1088 ();
 sg13g2_fill_8 FILLER_107_1096 ();
 sg13g2_fill_8 FILLER_107_1104 ();
 sg13g2_fill_8 FILLER_107_1112 ();
 sg13g2_fill_8 FILLER_107_1120 ();
 sg13g2_fill_8 FILLER_107_1128 ();
 sg13g2_fill_8 FILLER_107_1136 ();
 sg13g2_fill_8 FILLER_108_0 ();
 sg13g2_fill_8 FILLER_108_8 ();
 sg13g2_fill_8 FILLER_108_16 ();
 sg13g2_fill_8 FILLER_108_24 ();
 sg13g2_fill_8 FILLER_108_32 ();
 sg13g2_fill_8 FILLER_108_40 ();
 sg13g2_fill_8 FILLER_108_48 ();
 sg13g2_fill_8 FILLER_108_56 ();
 sg13g2_fill_8 FILLER_108_64 ();
 sg13g2_fill_8 FILLER_108_72 ();
 sg13g2_fill_8 FILLER_108_80 ();
 sg13g2_fill_8 FILLER_108_88 ();
 sg13g2_fill_8 FILLER_108_96 ();
 sg13g2_fill_8 FILLER_108_104 ();
 sg13g2_fill_8 FILLER_108_112 ();
 sg13g2_fill_8 FILLER_108_120 ();
 sg13g2_fill_8 FILLER_108_128 ();
 sg13g2_fill_8 FILLER_108_136 ();
 sg13g2_fill_8 FILLER_108_144 ();
 sg13g2_fill_8 FILLER_108_152 ();
 sg13g2_fill_8 FILLER_108_160 ();
 sg13g2_fill_8 FILLER_108_168 ();
 sg13g2_fill_8 FILLER_108_176 ();
 sg13g2_fill_8 FILLER_108_184 ();
 sg13g2_fill_8 FILLER_108_192 ();
 sg13g2_fill_8 FILLER_108_200 ();
 sg13g2_fill_8 FILLER_108_208 ();
 sg13g2_fill_8 FILLER_108_216 ();
 sg13g2_fill_8 FILLER_108_224 ();
 sg13g2_fill_8 FILLER_108_232 ();
 sg13g2_fill_8 FILLER_108_240 ();
 sg13g2_fill_8 FILLER_108_248 ();
 sg13g2_fill_8 FILLER_108_256 ();
 sg13g2_fill_8 FILLER_108_264 ();
 sg13g2_fill_8 FILLER_108_272 ();
 sg13g2_fill_8 FILLER_108_280 ();
 sg13g2_fill_8 FILLER_108_288 ();
 sg13g2_fill_8 FILLER_108_296 ();
 sg13g2_fill_8 FILLER_108_304 ();
 sg13g2_fill_8 FILLER_108_312 ();
 sg13g2_fill_8 FILLER_108_320 ();
 sg13g2_fill_8 FILLER_108_328 ();
 sg13g2_fill_8 FILLER_108_336 ();
 sg13g2_fill_8 FILLER_108_344 ();
 sg13g2_fill_8 FILLER_108_352 ();
 sg13g2_fill_8 FILLER_108_360 ();
 sg13g2_fill_8 FILLER_108_368 ();
 sg13g2_fill_8 FILLER_108_376 ();
 sg13g2_fill_8 FILLER_108_384 ();
 sg13g2_fill_8 FILLER_108_392 ();
 sg13g2_fill_8 FILLER_108_400 ();
 sg13g2_fill_8 FILLER_108_408 ();
 sg13g2_fill_8 FILLER_108_416 ();
 sg13g2_fill_8 FILLER_108_424 ();
 sg13g2_fill_8 FILLER_108_432 ();
 sg13g2_fill_8 FILLER_108_440 ();
 sg13g2_fill_8 FILLER_108_448 ();
 sg13g2_fill_8 FILLER_108_456 ();
 sg13g2_fill_8 FILLER_108_464 ();
 sg13g2_fill_8 FILLER_108_472 ();
 sg13g2_fill_8 FILLER_108_480 ();
 sg13g2_fill_8 FILLER_108_488 ();
 sg13g2_fill_8 FILLER_108_496 ();
 sg13g2_fill_8 FILLER_108_504 ();
 sg13g2_fill_8 FILLER_108_512 ();
 sg13g2_fill_8 FILLER_108_520 ();
 sg13g2_fill_8 FILLER_108_528 ();
 sg13g2_fill_8 FILLER_108_536 ();
 sg13g2_fill_8 FILLER_108_544 ();
 sg13g2_fill_8 FILLER_108_552 ();
 sg13g2_fill_8 FILLER_108_560 ();
 sg13g2_fill_8 FILLER_108_568 ();
 sg13g2_fill_8 FILLER_108_576 ();
 sg13g2_fill_8 FILLER_108_584 ();
 sg13g2_fill_8 FILLER_108_592 ();
 sg13g2_fill_8 FILLER_108_600 ();
 sg13g2_fill_8 FILLER_108_608 ();
 sg13g2_fill_8 FILLER_108_616 ();
 sg13g2_fill_8 FILLER_108_624 ();
 sg13g2_fill_8 FILLER_108_632 ();
 sg13g2_fill_8 FILLER_108_640 ();
 sg13g2_fill_8 FILLER_108_648 ();
 sg13g2_fill_8 FILLER_108_656 ();
 sg13g2_fill_8 FILLER_108_664 ();
 sg13g2_fill_8 FILLER_108_672 ();
 sg13g2_fill_8 FILLER_108_680 ();
 sg13g2_fill_8 FILLER_108_688 ();
 sg13g2_fill_8 FILLER_108_696 ();
 sg13g2_fill_8 FILLER_108_704 ();
 sg13g2_fill_8 FILLER_108_712 ();
 sg13g2_fill_8 FILLER_108_720 ();
 sg13g2_fill_8 FILLER_108_728 ();
 sg13g2_fill_8 FILLER_108_736 ();
 sg13g2_fill_8 FILLER_108_744 ();
 sg13g2_fill_8 FILLER_108_752 ();
 sg13g2_fill_8 FILLER_108_760 ();
 sg13g2_fill_8 FILLER_108_768 ();
 sg13g2_fill_8 FILLER_108_776 ();
 sg13g2_fill_8 FILLER_108_784 ();
 sg13g2_fill_8 FILLER_108_792 ();
 sg13g2_fill_8 FILLER_108_800 ();
 sg13g2_fill_8 FILLER_108_808 ();
 sg13g2_fill_8 FILLER_108_816 ();
 sg13g2_fill_8 FILLER_108_824 ();
 sg13g2_fill_8 FILLER_108_832 ();
 sg13g2_fill_8 FILLER_108_840 ();
 sg13g2_fill_8 FILLER_108_848 ();
 sg13g2_fill_8 FILLER_108_856 ();
 sg13g2_fill_8 FILLER_108_864 ();
 sg13g2_fill_8 FILLER_108_872 ();
 sg13g2_fill_8 FILLER_108_880 ();
 sg13g2_fill_8 FILLER_108_888 ();
 sg13g2_fill_8 FILLER_108_896 ();
 sg13g2_fill_8 FILLER_108_904 ();
 sg13g2_fill_8 FILLER_108_912 ();
 sg13g2_fill_8 FILLER_108_920 ();
 sg13g2_fill_8 FILLER_108_928 ();
 sg13g2_fill_8 FILLER_108_936 ();
 sg13g2_fill_8 FILLER_108_944 ();
 sg13g2_fill_8 FILLER_108_952 ();
 sg13g2_fill_8 FILLER_108_960 ();
 sg13g2_fill_8 FILLER_108_968 ();
 sg13g2_fill_8 FILLER_108_976 ();
 sg13g2_fill_8 FILLER_108_984 ();
 sg13g2_fill_8 FILLER_108_992 ();
 sg13g2_fill_8 FILLER_108_1000 ();
 sg13g2_fill_8 FILLER_108_1008 ();
 sg13g2_fill_8 FILLER_108_1016 ();
 sg13g2_fill_8 FILLER_108_1024 ();
 sg13g2_fill_8 FILLER_108_1032 ();
 sg13g2_fill_8 FILLER_108_1040 ();
 sg13g2_fill_8 FILLER_108_1048 ();
 sg13g2_fill_8 FILLER_108_1056 ();
 sg13g2_fill_8 FILLER_108_1064 ();
 sg13g2_fill_8 FILLER_108_1072 ();
 sg13g2_fill_8 FILLER_108_1080 ();
 sg13g2_fill_8 FILLER_108_1088 ();
 sg13g2_fill_8 FILLER_108_1096 ();
 sg13g2_fill_8 FILLER_108_1104 ();
 sg13g2_fill_8 FILLER_108_1112 ();
 sg13g2_fill_8 FILLER_108_1120 ();
 sg13g2_fill_8 FILLER_108_1128 ();
 sg13g2_fill_8 FILLER_108_1136 ();
 sg13g2_fill_8 FILLER_109_0 ();
 sg13g2_fill_8 FILLER_109_8 ();
 sg13g2_fill_8 FILLER_109_16 ();
 sg13g2_fill_8 FILLER_109_24 ();
 sg13g2_fill_8 FILLER_109_32 ();
 sg13g2_fill_8 FILLER_109_40 ();
 sg13g2_fill_8 FILLER_109_48 ();
 sg13g2_fill_8 FILLER_109_56 ();
 sg13g2_fill_8 FILLER_109_64 ();
 sg13g2_fill_8 FILLER_109_72 ();
 sg13g2_fill_8 FILLER_109_80 ();
 sg13g2_fill_8 FILLER_109_88 ();
 sg13g2_fill_8 FILLER_109_96 ();
 sg13g2_fill_8 FILLER_109_104 ();
 sg13g2_fill_8 FILLER_109_112 ();
 sg13g2_fill_8 FILLER_109_120 ();
 sg13g2_fill_8 FILLER_109_128 ();
 sg13g2_fill_8 FILLER_109_136 ();
 sg13g2_fill_8 FILLER_109_144 ();
 sg13g2_fill_8 FILLER_109_152 ();
 sg13g2_fill_8 FILLER_109_160 ();
 sg13g2_fill_8 FILLER_109_168 ();
 sg13g2_fill_8 FILLER_109_176 ();
 sg13g2_fill_8 FILLER_109_184 ();
 sg13g2_fill_8 FILLER_109_192 ();
 sg13g2_fill_8 FILLER_109_200 ();
 sg13g2_fill_8 FILLER_109_208 ();
 sg13g2_fill_8 FILLER_109_216 ();
 sg13g2_fill_8 FILLER_109_224 ();
 sg13g2_fill_8 FILLER_109_232 ();
 sg13g2_fill_8 FILLER_109_240 ();
 sg13g2_fill_8 FILLER_109_248 ();
 sg13g2_fill_8 FILLER_109_256 ();
 sg13g2_fill_8 FILLER_109_264 ();
 sg13g2_fill_8 FILLER_109_272 ();
 sg13g2_fill_8 FILLER_109_280 ();
 sg13g2_fill_8 FILLER_109_288 ();
 sg13g2_fill_8 FILLER_109_296 ();
 sg13g2_fill_8 FILLER_109_304 ();
 sg13g2_fill_8 FILLER_109_312 ();
 sg13g2_fill_8 FILLER_109_320 ();
 sg13g2_fill_8 FILLER_109_328 ();
 sg13g2_fill_8 FILLER_109_336 ();
 sg13g2_fill_8 FILLER_109_344 ();
 sg13g2_fill_8 FILLER_109_352 ();
 sg13g2_fill_8 FILLER_109_360 ();
 sg13g2_fill_8 FILLER_109_368 ();
 sg13g2_fill_8 FILLER_109_376 ();
 sg13g2_fill_8 FILLER_109_384 ();
 sg13g2_fill_8 FILLER_109_392 ();
 sg13g2_fill_8 FILLER_109_400 ();
 sg13g2_fill_8 FILLER_109_408 ();
 sg13g2_fill_8 FILLER_109_416 ();
 sg13g2_fill_8 FILLER_109_424 ();
 sg13g2_fill_8 FILLER_109_432 ();
 sg13g2_fill_8 FILLER_109_440 ();
 sg13g2_fill_8 FILLER_109_448 ();
 sg13g2_fill_8 FILLER_109_456 ();
 sg13g2_fill_8 FILLER_109_464 ();
 sg13g2_fill_8 FILLER_109_472 ();
 sg13g2_fill_8 FILLER_109_480 ();
 sg13g2_fill_8 FILLER_109_488 ();
 sg13g2_fill_8 FILLER_109_496 ();
 sg13g2_fill_8 FILLER_109_504 ();
 sg13g2_fill_8 FILLER_109_512 ();
 sg13g2_fill_8 FILLER_109_520 ();
 sg13g2_fill_8 FILLER_109_528 ();
 sg13g2_fill_8 FILLER_109_536 ();
 sg13g2_fill_8 FILLER_109_544 ();
 sg13g2_fill_8 FILLER_109_552 ();
 sg13g2_fill_8 FILLER_109_560 ();
 sg13g2_fill_8 FILLER_109_568 ();
 sg13g2_fill_8 FILLER_109_576 ();
 sg13g2_fill_8 FILLER_109_584 ();
 sg13g2_fill_8 FILLER_109_592 ();
 sg13g2_fill_8 FILLER_109_600 ();
 sg13g2_fill_8 FILLER_109_608 ();
 sg13g2_fill_8 FILLER_109_616 ();
 sg13g2_fill_8 FILLER_109_624 ();
 sg13g2_fill_8 FILLER_109_632 ();
 sg13g2_fill_8 FILLER_109_640 ();
 sg13g2_fill_8 FILLER_109_648 ();
 sg13g2_fill_8 FILLER_109_656 ();
 sg13g2_fill_8 FILLER_109_664 ();
 sg13g2_fill_8 FILLER_109_672 ();
 sg13g2_fill_8 FILLER_109_680 ();
 sg13g2_fill_8 FILLER_109_688 ();
 sg13g2_fill_8 FILLER_109_696 ();
 sg13g2_fill_8 FILLER_109_704 ();
 sg13g2_fill_8 FILLER_109_712 ();
 sg13g2_fill_8 FILLER_109_720 ();
 sg13g2_fill_8 FILLER_109_728 ();
 sg13g2_fill_8 FILLER_109_736 ();
 sg13g2_fill_8 FILLER_109_744 ();
 sg13g2_fill_8 FILLER_109_752 ();
 sg13g2_fill_8 FILLER_109_760 ();
 sg13g2_fill_8 FILLER_109_768 ();
 sg13g2_fill_8 FILLER_109_776 ();
 sg13g2_fill_8 FILLER_109_784 ();
 sg13g2_fill_8 FILLER_109_792 ();
 sg13g2_fill_8 FILLER_109_800 ();
 sg13g2_fill_8 FILLER_109_808 ();
 sg13g2_fill_8 FILLER_109_816 ();
 sg13g2_fill_8 FILLER_109_824 ();
 sg13g2_fill_8 FILLER_109_832 ();
 sg13g2_fill_8 FILLER_109_840 ();
 sg13g2_fill_8 FILLER_109_848 ();
 sg13g2_fill_8 FILLER_109_856 ();
 sg13g2_fill_8 FILLER_109_864 ();
 sg13g2_fill_8 FILLER_109_872 ();
 sg13g2_fill_8 FILLER_109_880 ();
 sg13g2_fill_8 FILLER_109_888 ();
 sg13g2_fill_8 FILLER_109_896 ();
 sg13g2_fill_8 FILLER_109_904 ();
 sg13g2_fill_8 FILLER_109_912 ();
 sg13g2_fill_8 FILLER_109_920 ();
 sg13g2_fill_8 FILLER_109_928 ();
 sg13g2_fill_8 FILLER_109_936 ();
 sg13g2_fill_8 FILLER_109_944 ();
 sg13g2_fill_8 FILLER_109_952 ();
 sg13g2_fill_8 FILLER_109_960 ();
 sg13g2_fill_8 FILLER_109_968 ();
 sg13g2_fill_8 FILLER_109_976 ();
 sg13g2_fill_8 FILLER_109_984 ();
 sg13g2_fill_8 FILLER_109_992 ();
 sg13g2_fill_8 FILLER_109_1000 ();
 sg13g2_fill_8 FILLER_109_1008 ();
 sg13g2_fill_8 FILLER_109_1016 ();
 sg13g2_fill_8 FILLER_109_1024 ();
 sg13g2_fill_8 FILLER_109_1032 ();
 sg13g2_fill_8 FILLER_109_1040 ();
 sg13g2_fill_8 FILLER_109_1048 ();
 sg13g2_fill_8 FILLER_109_1056 ();
 sg13g2_fill_8 FILLER_109_1064 ();
 sg13g2_fill_8 FILLER_109_1072 ();
 sg13g2_fill_8 FILLER_109_1080 ();
 sg13g2_fill_8 FILLER_109_1088 ();
 sg13g2_fill_8 FILLER_109_1096 ();
 sg13g2_fill_8 FILLER_109_1104 ();
 sg13g2_fill_8 FILLER_109_1112 ();
 sg13g2_fill_8 FILLER_109_1120 ();
 sg13g2_fill_8 FILLER_109_1128 ();
 sg13g2_fill_8 FILLER_109_1136 ();
 sg13g2_fill_8 FILLER_110_0 ();
 sg13g2_fill_8 FILLER_110_8 ();
 sg13g2_fill_8 FILLER_110_16 ();
 sg13g2_fill_8 FILLER_110_24 ();
 sg13g2_fill_8 FILLER_110_32 ();
 sg13g2_fill_8 FILLER_110_40 ();
 sg13g2_fill_8 FILLER_110_48 ();
 sg13g2_fill_8 FILLER_110_56 ();
 sg13g2_fill_8 FILLER_110_64 ();
 sg13g2_fill_8 FILLER_110_72 ();
 sg13g2_fill_8 FILLER_110_80 ();
 sg13g2_fill_8 FILLER_110_88 ();
 sg13g2_fill_8 FILLER_110_96 ();
 sg13g2_fill_8 FILLER_110_104 ();
 sg13g2_fill_8 FILLER_110_112 ();
 sg13g2_fill_8 FILLER_110_120 ();
 sg13g2_fill_8 FILLER_110_128 ();
 sg13g2_fill_8 FILLER_110_136 ();
 sg13g2_fill_8 FILLER_110_144 ();
 sg13g2_fill_8 FILLER_110_152 ();
 sg13g2_fill_8 FILLER_110_160 ();
 sg13g2_fill_8 FILLER_110_168 ();
 sg13g2_fill_8 FILLER_110_176 ();
 sg13g2_fill_8 FILLER_110_184 ();
 sg13g2_fill_8 FILLER_110_192 ();
 sg13g2_fill_8 FILLER_110_200 ();
 sg13g2_fill_8 FILLER_110_208 ();
 sg13g2_fill_8 FILLER_110_216 ();
 sg13g2_fill_8 FILLER_110_224 ();
 sg13g2_fill_8 FILLER_110_232 ();
 sg13g2_fill_8 FILLER_110_240 ();
 sg13g2_fill_8 FILLER_110_248 ();
 sg13g2_fill_8 FILLER_110_256 ();
 sg13g2_fill_8 FILLER_110_264 ();
 sg13g2_fill_8 FILLER_110_272 ();
 sg13g2_fill_8 FILLER_110_280 ();
 sg13g2_fill_8 FILLER_110_288 ();
 sg13g2_fill_8 FILLER_110_296 ();
 sg13g2_fill_8 FILLER_110_304 ();
 sg13g2_fill_8 FILLER_110_312 ();
 sg13g2_fill_8 FILLER_110_320 ();
 sg13g2_fill_8 FILLER_110_328 ();
 sg13g2_fill_8 FILLER_110_336 ();
 sg13g2_fill_8 FILLER_110_344 ();
 sg13g2_fill_8 FILLER_110_352 ();
 sg13g2_fill_8 FILLER_110_360 ();
 sg13g2_fill_8 FILLER_110_368 ();
 sg13g2_fill_8 FILLER_110_376 ();
 sg13g2_fill_8 FILLER_110_384 ();
 sg13g2_fill_8 FILLER_110_392 ();
 sg13g2_fill_8 FILLER_110_400 ();
 sg13g2_fill_8 FILLER_110_408 ();
 sg13g2_fill_8 FILLER_110_416 ();
 sg13g2_fill_8 FILLER_110_424 ();
 sg13g2_fill_8 FILLER_110_432 ();
 sg13g2_fill_8 FILLER_110_440 ();
 sg13g2_fill_8 FILLER_110_448 ();
 sg13g2_fill_8 FILLER_110_456 ();
 sg13g2_fill_8 FILLER_110_464 ();
 sg13g2_fill_8 FILLER_110_472 ();
 sg13g2_fill_8 FILLER_110_480 ();
 sg13g2_fill_8 FILLER_110_488 ();
 sg13g2_fill_8 FILLER_110_496 ();
 sg13g2_fill_8 FILLER_110_504 ();
 sg13g2_fill_8 FILLER_110_512 ();
 sg13g2_fill_8 FILLER_110_520 ();
 sg13g2_fill_8 FILLER_110_528 ();
 sg13g2_fill_8 FILLER_110_536 ();
 sg13g2_fill_8 FILLER_110_544 ();
 sg13g2_fill_8 FILLER_110_552 ();
 sg13g2_fill_8 FILLER_110_560 ();
 sg13g2_fill_8 FILLER_110_568 ();
 sg13g2_fill_8 FILLER_110_576 ();
 sg13g2_fill_8 FILLER_110_584 ();
 sg13g2_fill_8 FILLER_110_592 ();
 sg13g2_fill_8 FILLER_110_600 ();
 sg13g2_fill_8 FILLER_110_608 ();
 sg13g2_fill_8 FILLER_110_616 ();
 sg13g2_fill_8 FILLER_110_624 ();
 sg13g2_fill_8 FILLER_110_632 ();
 sg13g2_fill_8 FILLER_110_640 ();
 sg13g2_fill_8 FILLER_110_648 ();
 sg13g2_fill_8 FILLER_110_656 ();
 sg13g2_fill_8 FILLER_110_664 ();
 sg13g2_fill_8 FILLER_110_672 ();
 sg13g2_fill_8 FILLER_110_680 ();
 sg13g2_fill_8 FILLER_110_688 ();
 sg13g2_fill_8 FILLER_110_696 ();
 sg13g2_fill_8 FILLER_110_704 ();
 sg13g2_fill_8 FILLER_110_712 ();
 sg13g2_fill_8 FILLER_110_720 ();
 sg13g2_fill_8 FILLER_110_728 ();
 sg13g2_fill_8 FILLER_110_736 ();
 sg13g2_fill_8 FILLER_110_744 ();
 sg13g2_fill_8 FILLER_110_752 ();
 sg13g2_fill_8 FILLER_110_760 ();
 sg13g2_fill_8 FILLER_110_768 ();
 sg13g2_fill_8 FILLER_110_776 ();
 sg13g2_fill_8 FILLER_110_784 ();
 sg13g2_fill_8 FILLER_110_792 ();
 sg13g2_fill_8 FILLER_110_800 ();
 sg13g2_fill_8 FILLER_110_808 ();
 sg13g2_fill_8 FILLER_110_816 ();
 sg13g2_fill_8 FILLER_110_824 ();
 sg13g2_fill_8 FILLER_110_832 ();
 sg13g2_fill_8 FILLER_110_840 ();
 sg13g2_fill_8 FILLER_110_848 ();
 sg13g2_fill_8 FILLER_110_856 ();
 sg13g2_fill_8 FILLER_110_864 ();
 sg13g2_fill_8 FILLER_110_872 ();
 sg13g2_fill_8 FILLER_110_880 ();
 sg13g2_fill_8 FILLER_110_888 ();
 sg13g2_fill_8 FILLER_110_896 ();
 sg13g2_fill_8 FILLER_110_904 ();
 sg13g2_fill_8 FILLER_110_912 ();
 sg13g2_fill_8 FILLER_110_920 ();
 sg13g2_fill_8 FILLER_110_928 ();
 sg13g2_fill_8 FILLER_110_936 ();
 sg13g2_fill_8 FILLER_110_944 ();
 sg13g2_fill_8 FILLER_110_952 ();
 sg13g2_fill_8 FILLER_110_960 ();
 sg13g2_fill_8 FILLER_110_968 ();
 sg13g2_fill_8 FILLER_110_976 ();
 sg13g2_fill_8 FILLER_110_984 ();
 sg13g2_fill_8 FILLER_110_992 ();
 sg13g2_fill_8 FILLER_110_1000 ();
 sg13g2_fill_8 FILLER_110_1008 ();
 sg13g2_fill_8 FILLER_110_1016 ();
 sg13g2_fill_8 FILLER_110_1024 ();
 sg13g2_fill_8 FILLER_110_1032 ();
 sg13g2_fill_8 FILLER_110_1040 ();
 sg13g2_fill_8 FILLER_110_1048 ();
 sg13g2_fill_8 FILLER_110_1056 ();
 sg13g2_fill_8 FILLER_110_1064 ();
 sg13g2_fill_8 FILLER_110_1072 ();
 sg13g2_fill_8 FILLER_110_1080 ();
 sg13g2_fill_8 FILLER_110_1088 ();
 sg13g2_fill_8 FILLER_110_1096 ();
 sg13g2_fill_8 FILLER_110_1104 ();
 sg13g2_fill_8 FILLER_110_1112 ();
 sg13g2_fill_8 FILLER_110_1120 ();
 sg13g2_fill_8 FILLER_110_1128 ();
 sg13g2_fill_8 FILLER_110_1136 ();
 sg13g2_fill_8 FILLER_111_0 ();
 sg13g2_fill_8 FILLER_111_8 ();
 sg13g2_fill_8 FILLER_111_16 ();
 sg13g2_fill_8 FILLER_111_24 ();
 sg13g2_fill_8 FILLER_111_32 ();
 sg13g2_fill_8 FILLER_111_40 ();
 sg13g2_fill_8 FILLER_111_48 ();
 sg13g2_fill_8 FILLER_111_56 ();
 sg13g2_fill_8 FILLER_111_64 ();
 sg13g2_fill_8 FILLER_111_72 ();
 sg13g2_fill_8 FILLER_111_80 ();
 sg13g2_fill_8 FILLER_111_88 ();
 sg13g2_fill_8 FILLER_111_96 ();
 sg13g2_fill_8 FILLER_111_104 ();
 sg13g2_fill_8 FILLER_111_112 ();
 sg13g2_fill_8 FILLER_111_120 ();
 sg13g2_fill_8 FILLER_111_128 ();
 sg13g2_fill_8 FILLER_111_136 ();
 sg13g2_fill_8 FILLER_111_144 ();
 sg13g2_fill_8 FILLER_111_152 ();
 sg13g2_fill_8 FILLER_111_160 ();
 sg13g2_fill_8 FILLER_111_168 ();
 sg13g2_fill_8 FILLER_111_176 ();
 sg13g2_fill_8 FILLER_111_184 ();
 sg13g2_fill_8 FILLER_111_192 ();
 sg13g2_fill_8 FILLER_111_200 ();
 sg13g2_fill_8 FILLER_111_208 ();
 sg13g2_fill_8 FILLER_111_216 ();
 sg13g2_fill_8 FILLER_111_224 ();
 sg13g2_fill_8 FILLER_111_232 ();
 sg13g2_fill_8 FILLER_111_240 ();
 sg13g2_fill_8 FILLER_111_248 ();
 sg13g2_fill_8 FILLER_111_256 ();
 sg13g2_fill_8 FILLER_111_264 ();
 sg13g2_fill_8 FILLER_111_272 ();
 sg13g2_fill_8 FILLER_111_280 ();
 sg13g2_fill_8 FILLER_111_288 ();
 sg13g2_fill_8 FILLER_111_296 ();
 sg13g2_fill_8 FILLER_111_304 ();
 sg13g2_fill_8 FILLER_111_312 ();
 sg13g2_fill_8 FILLER_111_320 ();
 sg13g2_fill_8 FILLER_111_328 ();
 sg13g2_fill_8 FILLER_111_336 ();
 sg13g2_fill_8 FILLER_111_344 ();
 sg13g2_fill_8 FILLER_111_352 ();
 sg13g2_fill_8 FILLER_111_360 ();
 sg13g2_fill_8 FILLER_111_368 ();
 sg13g2_fill_8 FILLER_111_376 ();
 sg13g2_fill_8 FILLER_111_384 ();
 sg13g2_fill_8 FILLER_111_392 ();
 sg13g2_fill_8 FILLER_111_400 ();
 sg13g2_fill_8 FILLER_111_408 ();
 sg13g2_fill_8 FILLER_111_416 ();
 sg13g2_fill_8 FILLER_111_424 ();
 sg13g2_fill_8 FILLER_111_432 ();
 sg13g2_fill_8 FILLER_111_440 ();
 sg13g2_fill_8 FILLER_111_448 ();
 sg13g2_fill_8 FILLER_111_456 ();
 sg13g2_fill_8 FILLER_111_464 ();
 sg13g2_fill_8 FILLER_111_472 ();
 sg13g2_fill_8 FILLER_111_480 ();
 sg13g2_fill_8 FILLER_111_488 ();
 sg13g2_fill_8 FILLER_111_496 ();
 sg13g2_fill_8 FILLER_111_504 ();
 sg13g2_fill_8 FILLER_111_512 ();
 sg13g2_fill_8 FILLER_111_520 ();
 sg13g2_fill_8 FILLER_111_528 ();
 sg13g2_fill_8 FILLER_111_536 ();
 sg13g2_fill_8 FILLER_111_544 ();
 sg13g2_fill_8 FILLER_111_552 ();
 sg13g2_fill_8 FILLER_111_560 ();
 sg13g2_fill_8 FILLER_111_568 ();
 sg13g2_fill_8 FILLER_111_576 ();
 sg13g2_fill_8 FILLER_111_584 ();
 sg13g2_fill_8 FILLER_111_592 ();
 sg13g2_fill_8 FILLER_111_600 ();
 sg13g2_fill_8 FILLER_111_608 ();
 sg13g2_fill_8 FILLER_111_616 ();
 sg13g2_fill_8 FILLER_111_624 ();
 sg13g2_fill_8 FILLER_111_632 ();
 sg13g2_fill_8 FILLER_111_640 ();
 sg13g2_fill_8 FILLER_111_648 ();
 sg13g2_fill_8 FILLER_111_656 ();
 sg13g2_fill_8 FILLER_111_664 ();
 sg13g2_fill_8 FILLER_111_672 ();
 sg13g2_fill_8 FILLER_111_680 ();
 sg13g2_fill_8 FILLER_111_688 ();
 sg13g2_fill_8 FILLER_111_696 ();
 sg13g2_fill_8 FILLER_111_704 ();
 sg13g2_fill_8 FILLER_111_712 ();
 sg13g2_fill_8 FILLER_111_720 ();
 sg13g2_fill_8 FILLER_111_728 ();
 sg13g2_fill_8 FILLER_111_736 ();
 sg13g2_fill_8 FILLER_111_744 ();
 sg13g2_fill_8 FILLER_111_752 ();
 sg13g2_fill_8 FILLER_111_760 ();
 sg13g2_fill_8 FILLER_111_768 ();
 sg13g2_fill_8 FILLER_111_776 ();
 sg13g2_fill_8 FILLER_111_784 ();
 sg13g2_fill_8 FILLER_111_792 ();
 sg13g2_fill_8 FILLER_111_800 ();
 sg13g2_fill_8 FILLER_111_808 ();
 sg13g2_fill_8 FILLER_111_816 ();
 sg13g2_fill_8 FILLER_111_824 ();
 sg13g2_fill_8 FILLER_111_832 ();
 sg13g2_fill_8 FILLER_111_840 ();
 sg13g2_fill_8 FILLER_111_848 ();
 sg13g2_fill_8 FILLER_111_856 ();
 sg13g2_fill_8 FILLER_111_864 ();
 sg13g2_fill_8 FILLER_111_872 ();
 sg13g2_fill_8 FILLER_111_880 ();
 sg13g2_fill_8 FILLER_111_888 ();
 sg13g2_fill_8 FILLER_111_896 ();
 sg13g2_fill_8 FILLER_111_904 ();
 sg13g2_fill_8 FILLER_111_912 ();
 sg13g2_fill_8 FILLER_111_920 ();
 sg13g2_fill_8 FILLER_111_928 ();
 sg13g2_fill_8 FILLER_111_936 ();
 sg13g2_fill_8 FILLER_111_944 ();
 sg13g2_fill_8 FILLER_111_952 ();
 sg13g2_fill_8 FILLER_111_960 ();
 sg13g2_fill_8 FILLER_111_968 ();
 sg13g2_fill_8 FILLER_111_976 ();
 sg13g2_fill_8 FILLER_111_984 ();
 sg13g2_fill_8 FILLER_111_992 ();
 sg13g2_fill_8 FILLER_111_1000 ();
 sg13g2_fill_8 FILLER_111_1008 ();
 sg13g2_fill_8 FILLER_111_1016 ();
 sg13g2_fill_8 FILLER_111_1024 ();
 sg13g2_fill_8 FILLER_111_1032 ();
 sg13g2_fill_8 FILLER_111_1040 ();
 sg13g2_fill_8 FILLER_111_1048 ();
 sg13g2_fill_8 FILLER_111_1056 ();
 sg13g2_fill_8 FILLER_111_1064 ();
 sg13g2_fill_8 FILLER_111_1072 ();
 sg13g2_fill_8 FILLER_111_1080 ();
 sg13g2_fill_8 FILLER_111_1088 ();
 sg13g2_fill_8 FILLER_111_1096 ();
 sg13g2_fill_8 FILLER_111_1104 ();
 sg13g2_fill_8 FILLER_111_1112 ();
 sg13g2_fill_8 FILLER_111_1120 ();
 sg13g2_fill_8 FILLER_111_1128 ();
 sg13g2_fill_8 FILLER_111_1136 ();
 sg13g2_fill_8 FILLER_112_0 ();
 sg13g2_fill_8 FILLER_112_8 ();
 sg13g2_fill_8 FILLER_112_16 ();
 sg13g2_fill_8 FILLER_112_24 ();
 sg13g2_fill_8 FILLER_112_32 ();
 sg13g2_fill_8 FILLER_112_40 ();
 sg13g2_fill_8 FILLER_112_48 ();
 sg13g2_fill_8 FILLER_112_56 ();
 sg13g2_fill_8 FILLER_112_64 ();
 sg13g2_fill_8 FILLER_112_72 ();
 sg13g2_fill_8 FILLER_112_80 ();
 sg13g2_fill_8 FILLER_112_88 ();
 sg13g2_fill_8 FILLER_112_96 ();
 sg13g2_fill_8 FILLER_112_104 ();
 sg13g2_fill_8 FILLER_112_112 ();
 sg13g2_fill_8 FILLER_112_120 ();
 sg13g2_fill_8 FILLER_112_128 ();
 sg13g2_fill_8 FILLER_112_136 ();
 sg13g2_fill_8 FILLER_112_144 ();
 sg13g2_fill_8 FILLER_112_152 ();
 sg13g2_fill_8 FILLER_112_160 ();
 sg13g2_fill_8 FILLER_112_168 ();
 sg13g2_fill_8 FILLER_112_176 ();
 sg13g2_fill_8 FILLER_112_184 ();
 sg13g2_fill_8 FILLER_112_192 ();
 sg13g2_fill_8 FILLER_112_200 ();
 sg13g2_fill_8 FILLER_112_208 ();
 sg13g2_fill_8 FILLER_112_216 ();
 sg13g2_fill_8 FILLER_112_224 ();
 sg13g2_fill_8 FILLER_112_232 ();
 sg13g2_fill_8 FILLER_112_240 ();
 sg13g2_fill_8 FILLER_112_248 ();
 sg13g2_fill_8 FILLER_112_256 ();
 sg13g2_fill_8 FILLER_112_264 ();
 sg13g2_fill_8 FILLER_112_272 ();
 sg13g2_fill_8 FILLER_112_280 ();
 sg13g2_fill_8 FILLER_112_288 ();
 sg13g2_fill_8 FILLER_112_296 ();
 sg13g2_fill_8 FILLER_112_304 ();
 sg13g2_fill_8 FILLER_112_312 ();
 sg13g2_fill_8 FILLER_112_320 ();
 sg13g2_fill_8 FILLER_112_328 ();
 sg13g2_fill_8 FILLER_112_336 ();
 sg13g2_fill_8 FILLER_112_344 ();
 sg13g2_fill_8 FILLER_112_352 ();
 sg13g2_fill_8 FILLER_112_360 ();
 sg13g2_fill_8 FILLER_112_368 ();
 sg13g2_fill_8 FILLER_112_376 ();
 sg13g2_fill_8 FILLER_112_384 ();
 sg13g2_fill_8 FILLER_112_392 ();
 sg13g2_fill_8 FILLER_112_400 ();
 sg13g2_fill_8 FILLER_112_408 ();
 sg13g2_fill_8 FILLER_112_416 ();
 sg13g2_fill_8 FILLER_112_424 ();
 sg13g2_fill_8 FILLER_112_432 ();
 sg13g2_fill_8 FILLER_112_440 ();
 sg13g2_fill_8 FILLER_112_448 ();
 sg13g2_fill_8 FILLER_112_456 ();
 sg13g2_fill_8 FILLER_112_464 ();
 sg13g2_fill_8 FILLER_112_472 ();
 sg13g2_fill_8 FILLER_112_480 ();
 sg13g2_fill_8 FILLER_112_488 ();
 sg13g2_fill_8 FILLER_112_496 ();
 sg13g2_fill_8 FILLER_112_504 ();
 sg13g2_fill_8 FILLER_112_512 ();
 sg13g2_fill_8 FILLER_112_520 ();
 sg13g2_fill_8 FILLER_112_528 ();
 sg13g2_fill_8 FILLER_112_536 ();
 sg13g2_fill_8 FILLER_112_544 ();
 sg13g2_fill_8 FILLER_112_552 ();
 sg13g2_fill_8 FILLER_112_560 ();
 sg13g2_fill_8 FILLER_112_568 ();
 sg13g2_fill_8 FILLER_112_576 ();
 sg13g2_fill_8 FILLER_112_584 ();
 sg13g2_fill_8 FILLER_112_592 ();
 sg13g2_fill_8 FILLER_112_600 ();
 sg13g2_fill_8 FILLER_112_608 ();
 sg13g2_fill_8 FILLER_112_616 ();
 sg13g2_fill_8 FILLER_112_624 ();
 sg13g2_fill_8 FILLER_112_632 ();
 sg13g2_fill_8 FILLER_112_640 ();
 sg13g2_fill_8 FILLER_112_648 ();
 sg13g2_fill_8 FILLER_112_656 ();
 sg13g2_fill_8 FILLER_112_664 ();
 sg13g2_fill_8 FILLER_112_672 ();
 sg13g2_fill_8 FILLER_112_680 ();
 sg13g2_fill_8 FILLER_112_688 ();
 sg13g2_fill_8 FILLER_112_696 ();
 sg13g2_fill_8 FILLER_112_704 ();
 sg13g2_fill_8 FILLER_112_712 ();
 sg13g2_fill_8 FILLER_112_720 ();
 sg13g2_fill_8 FILLER_112_728 ();
 sg13g2_fill_8 FILLER_112_736 ();
 sg13g2_fill_8 FILLER_112_744 ();
 sg13g2_fill_8 FILLER_112_752 ();
 sg13g2_fill_8 FILLER_112_760 ();
 sg13g2_fill_8 FILLER_112_768 ();
 sg13g2_fill_8 FILLER_112_776 ();
 sg13g2_fill_8 FILLER_112_784 ();
 sg13g2_fill_8 FILLER_112_792 ();
 sg13g2_fill_8 FILLER_112_800 ();
 sg13g2_fill_8 FILLER_112_808 ();
 sg13g2_fill_8 FILLER_112_816 ();
 sg13g2_fill_8 FILLER_112_824 ();
 sg13g2_fill_8 FILLER_112_832 ();
 sg13g2_fill_8 FILLER_112_840 ();
 sg13g2_fill_8 FILLER_112_848 ();
 sg13g2_fill_8 FILLER_112_856 ();
 sg13g2_fill_8 FILLER_112_864 ();
 sg13g2_fill_8 FILLER_112_872 ();
 sg13g2_fill_8 FILLER_112_880 ();
 sg13g2_fill_8 FILLER_112_888 ();
 sg13g2_fill_8 FILLER_112_896 ();
 sg13g2_fill_8 FILLER_112_904 ();
 sg13g2_fill_8 FILLER_112_912 ();
 sg13g2_fill_8 FILLER_112_920 ();
 sg13g2_fill_8 FILLER_112_928 ();
 sg13g2_fill_8 FILLER_112_936 ();
 sg13g2_fill_8 FILLER_112_944 ();
 sg13g2_fill_8 FILLER_112_952 ();
 sg13g2_fill_8 FILLER_112_960 ();
 sg13g2_fill_8 FILLER_112_968 ();
 sg13g2_fill_8 FILLER_112_976 ();
 sg13g2_fill_8 FILLER_112_984 ();
 sg13g2_fill_8 FILLER_112_992 ();
 sg13g2_fill_8 FILLER_112_1000 ();
 sg13g2_fill_8 FILLER_112_1008 ();
 sg13g2_fill_8 FILLER_112_1016 ();
 sg13g2_fill_8 FILLER_112_1024 ();
 sg13g2_fill_8 FILLER_112_1032 ();
 sg13g2_fill_8 FILLER_112_1040 ();
 sg13g2_fill_8 FILLER_112_1048 ();
 sg13g2_fill_8 FILLER_112_1056 ();
 sg13g2_fill_8 FILLER_112_1064 ();
 sg13g2_fill_8 FILLER_112_1072 ();
 sg13g2_fill_8 FILLER_112_1080 ();
 sg13g2_fill_8 FILLER_112_1088 ();
 sg13g2_fill_8 FILLER_112_1096 ();
 sg13g2_fill_8 FILLER_112_1104 ();
 sg13g2_fill_8 FILLER_112_1112 ();
 sg13g2_fill_8 FILLER_112_1120 ();
 sg13g2_fill_8 FILLER_112_1128 ();
 sg13g2_fill_8 FILLER_112_1136 ();
 sg13g2_fill_8 FILLER_113_0 ();
 sg13g2_fill_8 FILLER_113_8 ();
 sg13g2_fill_8 FILLER_113_16 ();
 sg13g2_fill_8 FILLER_113_24 ();
 sg13g2_fill_8 FILLER_113_32 ();
 sg13g2_fill_8 FILLER_113_40 ();
 sg13g2_fill_8 FILLER_113_48 ();
 sg13g2_fill_8 FILLER_113_56 ();
 sg13g2_fill_8 FILLER_113_64 ();
 sg13g2_fill_8 FILLER_113_72 ();
 sg13g2_fill_8 FILLER_113_80 ();
 sg13g2_fill_8 FILLER_113_88 ();
 sg13g2_fill_8 FILLER_113_96 ();
 sg13g2_fill_8 FILLER_113_104 ();
 sg13g2_fill_8 FILLER_113_112 ();
 sg13g2_fill_8 FILLER_113_120 ();
 sg13g2_fill_8 FILLER_113_128 ();
 sg13g2_fill_8 FILLER_113_136 ();
 sg13g2_fill_8 FILLER_113_144 ();
 sg13g2_fill_8 FILLER_113_152 ();
 sg13g2_fill_8 FILLER_113_160 ();
 sg13g2_fill_8 FILLER_113_168 ();
 sg13g2_fill_8 FILLER_113_176 ();
 sg13g2_fill_8 FILLER_113_184 ();
 sg13g2_fill_8 FILLER_113_192 ();
 sg13g2_fill_8 FILLER_113_200 ();
 sg13g2_fill_8 FILLER_113_208 ();
 sg13g2_fill_8 FILLER_113_216 ();
 sg13g2_fill_8 FILLER_113_224 ();
 sg13g2_fill_8 FILLER_113_232 ();
 sg13g2_fill_8 FILLER_113_240 ();
 sg13g2_fill_8 FILLER_113_248 ();
 sg13g2_fill_8 FILLER_113_256 ();
 sg13g2_fill_8 FILLER_113_264 ();
 sg13g2_fill_8 FILLER_113_272 ();
 sg13g2_fill_8 FILLER_113_280 ();
 sg13g2_fill_8 FILLER_113_288 ();
 sg13g2_fill_8 FILLER_113_296 ();
 sg13g2_fill_8 FILLER_113_304 ();
 sg13g2_fill_8 FILLER_113_312 ();
 sg13g2_fill_8 FILLER_113_320 ();
 sg13g2_fill_8 FILLER_113_328 ();
 sg13g2_fill_8 FILLER_113_336 ();
 sg13g2_fill_8 FILLER_113_344 ();
 sg13g2_fill_8 FILLER_113_352 ();
 sg13g2_fill_8 FILLER_113_360 ();
 sg13g2_fill_8 FILLER_113_368 ();
 sg13g2_fill_8 FILLER_113_376 ();
 sg13g2_fill_8 FILLER_113_384 ();
 sg13g2_fill_8 FILLER_113_392 ();
 sg13g2_fill_8 FILLER_113_400 ();
 sg13g2_fill_8 FILLER_113_408 ();
 sg13g2_fill_8 FILLER_113_416 ();
 sg13g2_fill_8 FILLER_113_424 ();
 sg13g2_fill_8 FILLER_113_432 ();
 sg13g2_fill_8 FILLER_113_440 ();
 sg13g2_fill_8 FILLER_113_448 ();
 sg13g2_fill_8 FILLER_113_456 ();
 sg13g2_fill_8 FILLER_113_464 ();
 sg13g2_fill_8 FILLER_113_472 ();
 sg13g2_fill_8 FILLER_113_480 ();
 sg13g2_fill_8 FILLER_113_488 ();
 sg13g2_fill_8 FILLER_113_496 ();
 sg13g2_fill_8 FILLER_113_504 ();
 sg13g2_fill_8 FILLER_113_512 ();
 sg13g2_fill_8 FILLER_113_520 ();
 sg13g2_fill_8 FILLER_113_528 ();
 sg13g2_fill_8 FILLER_113_536 ();
 sg13g2_fill_8 FILLER_113_544 ();
 sg13g2_fill_8 FILLER_113_552 ();
 sg13g2_fill_8 FILLER_113_560 ();
 sg13g2_fill_8 FILLER_113_568 ();
 sg13g2_fill_8 FILLER_113_576 ();
 sg13g2_fill_8 FILLER_113_584 ();
 sg13g2_fill_8 FILLER_113_592 ();
 sg13g2_fill_8 FILLER_113_600 ();
 sg13g2_fill_8 FILLER_113_608 ();
 sg13g2_fill_8 FILLER_113_616 ();
 sg13g2_fill_8 FILLER_113_624 ();
 sg13g2_fill_8 FILLER_113_632 ();
 sg13g2_fill_8 FILLER_113_640 ();
 sg13g2_fill_8 FILLER_113_648 ();
 sg13g2_fill_8 FILLER_113_656 ();
 sg13g2_fill_8 FILLER_113_664 ();
 sg13g2_fill_8 FILLER_113_672 ();
 sg13g2_fill_8 FILLER_113_680 ();
 sg13g2_fill_8 FILLER_113_688 ();
 sg13g2_fill_8 FILLER_113_696 ();
 sg13g2_fill_8 FILLER_113_704 ();
 sg13g2_fill_8 FILLER_113_712 ();
 sg13g2_fill_8 FILLER_113_720 ();
 sg13g2_fill_8 FILLER_113_728 ();
 sg13g2_fill_8 FILLER_113_736 ();
 sg13g2_fill_8 FILLER_113_744 ();
 sg13g2_fill_8 FILLER_113_752 ();
 sg13g2_fill_8 FILLER_113_760 ();
 sg13g2_fill_8 FILLER_113_768 ();
 sg13g2_fill_8 FILLER_113_776 ();
 sg13g2_fill_8 FILLER_113_784 ();
 sg13g2_fill_8 FILLER_113_792 ();
 sg13g2_fill_8 FILLER_113_800 ();
 sg13g2_fill_8 FILLER_113_808 ();
 sg13g2_fill_8 FILLER_113_816 ();
 sg13g2_fill_8 FILLER_113_824 ();
 sg13g2_fill_8 FILLER_113_832 ();
 sg13g2_fill_8 FILLER_113_840 ();
 sg13g2_fill_8 FILLER_113_848 ();
 sg13g2_fill_8 FILLER_113_856 ();
 sg13g2_fill_8 FILLER_113_864 ();
 sg13g2_fill_8 FILLER_113_872 ();
 sg13g2_fill_8 FILLER_113_880 ();
 sg13g2_fill_8 FILLER_113_888 ();
 sg13g2_fill_8 FILLER_113_896 ();
 sg13g2_fill_8 FILLER_113_904 ();
 sg13g2_fill_8 FILLER_113_912 ();
 sg13g2_fill_8 FILLER_113_920 ();
 sg13g2_fill_8 FILLER_113_928 ();
 sg13g2_fill_8 FILLER_113_936 ();
 sg13g2_fill_8 FILLER_113_944 ();
 sg13g2_fill_8 FILLER_113_952 ();
 sg13g2_fill_8 FILLER_113_960 ();
 sg13g2_fill_8 FILLER_113_968 ();
 sg13g2_fill_8 FILLER_113_976 ();
 sg13g2_fill_8 FILLER_113_984 ();
 sg13g2_fill_8 FILLER_113_992 ();
 sg13g2_fill_8 FILLER_113_1000 ();
 sg13g2_fill_8 FILLER_113_1008 ();
 sg13g2_fill_8 FILLER_113_1016 ();
 sg13g2_fill_8 FILLER_113_1024 ();
 sg13g2_fill_8 FILLER_113_1032 ();
 sg13g2_fill_8 FILLER_113_1040 ();
 sg13g2_fill_8 FILLER_113_1048 ();
 sg13g2_fill_8 FILLER_113_1056 ();
 sg13g2_fill_8 FILLER_113_1064 ();
 sg13g2_fill_8 FILLER_113_1072 ();
 sg13g2_fill_8 FILLER_113_1080 ();
 sg13g2_fill_8 FILLER_113_1088 ();
 sg13g2_fill_8 FILLER_113_1096 ();
 sg13g2_fill_8 FILLER_113_1104 ();
 sg13g2_fill_8 FILLER_113_1112 ();
 sg13g2_fill_8 FILLER_113_1120 ();
 sg13g2_fill_8 FILLER_113_1128 ();
 sg13g2_fill_8 FILLER_113_1136 ();
 sg13g2_fill_8 FILLER_114_0 ();
 sg13g2_fill_8 FILLER_114_8 ();
 sg13g2_fill_8 FILLER_114_16 ();
 sg13g2_fill_8 FILLER_114_24 ();
 sg13g2_fill_8 FILLER_114_32 ();
 sg13g2_fill_8 FILLER_114_40 ();
 sg13g2_fill_8 FILLER_114_48 ();
 sg13g2_fill_8 FILLER_114_56 ();
 sg13g2_fill_8 FILLER_114_64 ();
 sg13g2_fill_8 FILLER_114_72 ();
 sg13g2_fill_8 FILLER_114_80 ();
 sg13g2_fill_8 FILLER_114_88 ();
 sg13g2_fill_8 FILLER_114_96 ();
 sg13g2_fill_8 FILLER_114_104 ();
 sg13g2_fill_8 FILLER_114_112 ();
 sg13g2_fill_8 FILLER_114_120 ();
 sg13g2_fill_8 FILLER_114_128 ();
 sg13g2_fill_8 FILLER_114_136 ();
 sg13g2_fill_8 FILLER_114_144 ();
 sg13g2_fill_8 FILLER_114_152 ();
 sg13g2_fill_8 FILLER_114_160 ();
 sg13g2_fill_8 FILLER_114_168 ();
 sg13g2_fill_8 FILLER_114_176 ();
 sg13g2_fill_8 FILLER_114_184 ();
 sg13g2_fill_8 FILLER_114_192 ();
 sg13g2_fill_8 FILLER_114_200 ();
 sg13g2_fill_8 FILLER_114_208 ();
 sg13g2_fill_8 FILLER_114_216 ();
 sg13g2_fill_8 FILLER_114_224 ();
 sg13g2_fill_8 FILLER_114_232 ();
 sg13g2_fill_8 FILLER_114_240 ();
 sg13g2_fill_8 FILLER_114_248 ();
 sg13g2_fill_8 FILLER_114_256 ();
 sg13g2_fill_8 FILLER_114_264 ();
 sg13g2_fill_8 FILLER_114_272 ();
 sg13g2_fill_8 FILLER_114_280 ();
 sg13g2_fill_8 FILLER_114_288 ();
 sg13g2_fill_8 FILLER_114_296 ();
 sg13g2_fill_8 FILLER_114_304 ();
 sg13g2_fill_8 FILLER_114_312 ();
 sg13g2_fill_8 FILLER_114_320 ();
 sg13g2_fill_8 FILLER_114_328 ();
 sg13g2_fill_8 FILLER_114_336 ();
 sg13g2_fill_8 FILLER_114_344 ();
 sg13g2_fill_8 FILLER_114_352 ();
 sg13g2_fill_8 FILLER_114_360 ();
 sg13g2_fill_8 FILLER_114_368 ();
 sg13g2_fill_8 FILLER_114_376 ();
 sg13g2_fill_8 FILLER_114_384 ();
 sg13g2_fill_8 FILLER_114_392 ();
 sg13g2_fill_8 FILLER_114_400 ();
 sg13g2_fill_8 FILLER_114_408 ();
 sg13g2_fill_8 FILLER_114_416 ();
 sg13g2_fill_8 FILLER_114_424 ();
 sg13g2_fill_8 FILLER_114_432 ();
 sg13g2_fill_8 FILLER_114_440 ();
 sg13g2_fill_8 FILLER_114_448 ();
 sg13g2_fill_8 FILLER_114_456 ();
 sg13g2_fill_8 FILLER_114_464 ();
 sg13g2_fill_8 FILLER_114_472 ();
 sg13g2_fill_8 FILLER_114_480 ();
 sg13g2_fill_8 FILLER_114_488 ();
 sg13g2_fill_8 FILLER_114_496 ();
 sg13g2_fill_8 FILLER_114_504 ();
 sg13g2_fill_8 FILLER_114_512 ();
 sg13g2_fill_8 FILLER_114_520 ();
 sg13g2_fill_8 FILLER_114_528 ();
 sg13g2_fill_8 FILLER_114_536 ();
 sg13g2_fill_8 FILLER_114_544 ();
 sg13g2_fill_8 FILLER_114_552 ();
 sg13g2_fill_8 FILLER_114_560 ();
 sg13g2_fill_8 FILLER_114_568 ();
 sg13g2_fill_8 FILLER_114_576 ();
 sg13g2_fill_8 FILLER_114_584 ();
 sg13g2_fill_8 FILLER_114_592 ();
 sg13g2_fill_8 FILLER_114_600 ();
 sg13g2_fill_8 FILLER_114_608 ();
 sg13g2_fill_8 FILLER_114_616 ();
 sg13g2_fill_8 FILLER_114_624 ();
 sg13g2_fill_8 FILLER_114_632 ();
 sg13g2_fill_8 FILLER_114_640 ();
 sg13g2_fill_8 FILLER_114_648 ();
 sg13g2_fill_8 FILLER_114_656 ();
 sg13g2_fill_8 FILLER_114_664 ();
 sg13g2_fill_8 FILLER_114_672 ();
 sg13g2_fill_8 FILLER_114_680 ();
 sg13g2_fill_8 FILLER_114_688 ();
 sg13g2_fill_8 FILLER_114_696 ();
 sg13g2_fill_8 FILLER_114_704 ();
 sg13g2_fill_8 FILLER_114_712 ();
 sg13g2_fill_8 FILLER_114_720 ();
 sg13g2_fill_8 FILLER_114_728 ();
 sg13g2_fill_8 FILLER_114_736 ();
 sg13g2_fill_8 FILLER_114_744 ();
 sg13g2_fill_8 FILLER_114_752 ();
 sg13g2_fill_8 FILLER_114_760 ();
 sg13g2_fill_8 FILLER_114_768 ();
 sg13g2_fill_8 FILLER_114_776 ();
 sg13g2_fill_8 FILLER_114_784 ();
 sg13g2_fill_8 FILLER_114_792 ();
 sg13g2_fill_8 FILLER_114_800 ();
 sg13g2_fill_8 FILLER_114_808 ();
 sg13g2_fill_8 FILLER_114_816 ();
 sg13g2_fill_8 FILLER_114_824 ();
 sg13g2_fill_8 FILLER_114_832 ();
 sg13g2_fill_8 FILLER_114_840 ();
 sg13g2_fill_8 FILLER_114_848 ();
 sg13g2_fill_8 FILLER_114_856 ();
 sg13g2_fill_8 FILLER_114_864 ();
 sg13g2_fill_8 FILLER_114_872 ();
 sg13g2_fill_8 FILLER_114_880 ();
 sg13g2_fill_8 FILLER_114_888 ();
 sg13g2_fill_8 FILLER_114_896 ();
 sg13g2_fill_8 FILLER_114_904 ();
 sg13g2_fill_8 FILLER_114_912 ();
 sg13g2_fill_8 FILLER_114_920 ();
 sg13g2_fill_8 FILLER_114_928 ();
 sg13g2_fill_8 FILLER_114_936 ();
 sg13g2_fill_8 FILLER_114_944 ();
 sg13g2_fill_8 FILLER_114_952 ();
 sg13g2_fill_8 FILLER_114_960 ();
 sg13g2_fill_8 FILLER_114_968 ();
 sg13g2_fill_8 FILLER_114_976 ();
 sg13g2_fill_8 FILLER_114_984 ();
 sg13g2_fill_8 FILLER_114_992 ();
 sg13g2_fill_8 FILLER_114_1000 ();
 sg13g2_fill_8 FILLER_114_1008 ();
 sg13g2_fill_8 FILLER_114_1016 ();
 sg13g2_fill_8 FILLER_114_1024 ();
 sg13g2_fill_8 FILLER_114_1032 ();
 sg13g2_fill_8 FILLER_114_1040 ();
 sg13g2_fill_8 FILLER_114_1048 ();
 sg13g2_fill_8 FILLER_114_1056 ();
 sg13g2_fill_8 FILLER_114_1064 ();
 sg13g2_fill_8 FILLER_114_1072 ();
 sg13g2_fill_8 FILLER_114_1080 ();
 sg13g2_fill_8 FILLER_114_1088 ();
 sg13g2_fill_8 FILLER_114_1096 ();
 sg13g2_fill_8 FILLER_114_1104 ();
 sg13g2_fill_8 FILLER_114_1112 ();
 sg13g2_fill_8 FILLER_114_1120 ();
 sg13g2_fill_8 FILLER_114_1128 ();
 sg13g2_fill_8 FILLER_114_1136 ();
 sg13g2_fill_8 FILLER_115_0 ();
 sg13g2_fill_8 FILLER_115_8 ();
 sg13g2_fill_8 FILLER_115_16 ();
 sg13g2_fill_8 FILLER_115_24 ();
 sg13g2_fill_8 FILLER_115_32 ();
 sg13g2_fill_8 FILLER_115_40 ();
 sg13g2_fill_8 FILLER_115_48 ();
 sg13g2_fill_8 FILLER_115_56 ();
 sg13g2_fill_8 FILLER_115_64 ();
 sg13g2_fill_8 FILLER_115_72 ();
 sg13g2_fill_8 FILLER_115_80 ();
 sg13g2_fill_8 FILLER_115_88 ();
 sg13g2_fill_8 FILLER_115_96 ();
 sg13g2_fill_8 FILLER_115_104 ();
 sg13g2_fill_8 FILLER_115_112 ();
 sg13g2_fill_8 FILLER_115_120 ();
 sg13g2_fill_8 FILLER_115_128 ();
 sg13g2_fill_8 FILLER_115_136 ();
 sg13g2_fill_8 FILLER_115_144 ();
 sg13g2_fill_8 FILLER_115_152 ();
 sg13g2_fill_8 FILLER_115_160 ();
 sg13g2_fill_8 FILLER_115_168 ();
 sg13g2_fill_8 FILLER_115_176 ();
 sg13g2_fill_8 FILLER_115_184 ();
 sg13g2_fill_8 FILLER_115_192 ();
 sg13g2_fill_8 FILLER_115_200 ();
 sg13g2_fill_8 FILLER_115_208 ();
 sg13g2_fill_8 FILLER_115_216 ();
 sg13g2_fill_8 FILLER_115_224 ();
 sg13g2_fill_8 FILLER_115_232 ();
 sg13g2_fill_8 FILLER_115_240 ();
 sg13g2_fill_8 FILLER_115_248 ();
 sg13g2_fill_8 FILLER_115_256 ();
 sg13g2_fill_8 FILLER_115_264 ();
 sg13g2_fill_8 FILLER_115_272 ();
 sg13g2_fill_8 FILLER_115_280 ();
 sg13g2_fill_8 FILLER_115_288 ();
 sg13g2_fill_8 FILLER_115_296 ();
 sg13g2_fill_8 FILLER_115_304 ();
 sg13g2_fill_8 FILLER_115_312 ();
 sg13g2_fill_8 FILLER_115_320 ();
 sg13g2_fill_8 FILLER_115_328 ();
 sg13g2_fill_8 FILLER_115_336 ();
 sg13g2_fill_8 FILLER_115_344 ();
 sg13g2_fill_8 FILLER_115_352 ();
 sg13g2_fill_8 FILLER_115_360 ();
 sg13g2_fill_8 FILLER_115_368 ();
 sg13g2_fill_8 FILLER_115_376 ();
 sg13g2_fill_8 FILLER_115_384 ();
 sg13g2_fill_8 FILLER_115_392 ();
 sg13g2_fill_8 FILLER_115_400 ();
 sg13g2_fill_8 FILLER_115_408 ();
 sg13g2_fill_8 FILLER_115_416 ();
 sg13g2_fill_8 FILLER_115_424 ();
 sg13g2_fill_8 FILLER_115_432 ();
 sg13g2_fill_8 FILLER_115_440 ();
 sg13g2_fill_8 FILLER_115_448 ();
 sg13g2_fill_8 FILLER_115_456 ();
 sg13g2_fill_8 FILLER_115_464 ();
 sg13g2_fill_8 FILLER_115_472 ();
 sg13g2_fill_8 FILLER_115_480 ();
 sg13g2_fill_8 FILLER_115_488 ();
 sg13g2_fill_8 FILLER_115_496 ();
 sg13g2_fill_8 FILLER_115_504 ();
 sg13g2_fill_8 FILLER_115_512 ();
 sg13g2_fill_8 FILLER_115_520 ();
 sg13g2_fill_8 FILLER_115_528 ();
 sg13g2_fill_8 FILLER_115_536 ();
 sg13g2_fill_8 FILLER_115_544 ();
 sg13g2_fill_8 FILLER_115_552 ();
 sg13g2_fill_8 FILLER_115_560 ();
 sg13g2_fill_8 FILLER_115_568 ();
 sg13g2_fill_8 FILLER_115_576 ();
 sg13g2_fill_8 FILLER_115_584 ();
 sg13g2_fill_8 FILLER_115_592 ();
 sg13g2_fill_8 FILLER_115_600 ();
 sg13g2_fill_8 FILLER_115_608 ();
 sg13g2_fill_8 FILLER_115_616 ();
 sg13g2_fill_8 FILLER_115_624 ();
 sg13g2_fill_8 FILLER_115_632 ();
 sg13g2_fill_8 FILLER_115_640 ();
 sg13g2_fill_8 FILLER_115_648 ();
 sg13g2_fill_8 FILLER_115_656 ();
 sg13g2_fill_8 FILLER_115_664 ();
 sg13g2_fill_8 FILLER_115_672 ();
 sg13g2_fill_8 FILLER_115_680 ();
 sg13g2_fill_8 FILLER_115_688 ();
 sg13g2_fill_8 FILLER_115_696 ();
 sg13g2_fill_8 FILLER_115_704 ();
 sg13g2_fill_8 FILLER_115_712 ();
 sg13g2_fill_8 FILLER_115_720 ();
 sg13g2_fill_8 FILLER_115_728 ();
 sg13g2_fill_8 FILLER_115_736 ();
 sg13g2_fill_8 FILLER_115_744 ();
 sg13g2_fill_8 FILLER_115_752 ();
 sg13g2_fill_8 FILLER_115_760 ();
 sg13g2_fill_8 FILLER_115_768 ();
 sg13g2_fill_8 FILLER_115_776 ();
 sg13g2_fill_8 FILLER_115_784 ();
 sg13g2_fill_8 FILLER_115_792 ();
 sg13g2_fill_8 FILLER_115_800 ();
 sg13g2_fill_8 FILLER_115_808 ();
 sg13g2_fill_8 FILLER_115_816 ();
 sg13g2_fill_8 FILLER_115_824 ();
 sg13g2_fill_8 FILLER_115_832 ();
 sg13g2_fill_8 FILLER_115_840 ();
 sg13g2_fill_8 FILLER_115_848 ();
 sg13g2_fill_8 FILLER_115_856 ();
 sg13g2_fill_8 FILLER_115_864 ();
 sg13g2_fill_8 FILLER_115_872 ();
 sg13g2_fill_8 FILLER_115_880 ();
 sg13g2_fill_8 FILLER_115_888 ();
 sg13g2_fill_8 FILLER_115_896 ();
 sg13g2_fill_8 FILLER_115_904 ();
 sg13g2_fill_8 FILLER_115_912 ();
 sg13g2_fill_8 FILLER_115_920 ();
 sg13g2_fill_8 FILLER_115_928 ();
 sg13g2_fill_8 FILLER_115_936 ();
 sg13g2_fill_8 FILLER_115_944 ();
 sg13g2_fill_8 FILLER_115_952 ();
 sg13g2_fill_8 FILLER_115_960 ();
 sg13g2_fill_8 FILLER_115_968 ();
 sg13g2_fill_8 FILLER_115_976 ();
 sg13g2_fill_8 FILLER_115_984 ();
 sg13g2_fill_8 FILLER_115_992 ();
 sg13g2_fill_8 FILLER_115_1000 ();
 sg13g2_fill_8 FILLER_115_1008 ();
 sg13g2_fill_8 FILLER_115_1016 ();
 sg13g2_fill_8 FILLER_115_1024 ();
 sg13g2_fill_8 FILLER_115_1032 ();
 sg13g2_fill_8 FILLER_115_1040 ();
 sg13g2_fill_8 FILLER_115_1048 ();
 sg13g2_fill_8 FILLER_115_1056 ();
 sg13g2_fill_8 FILLER_115_1064 ();
 sg13g2_fill_8 FILLER_115_1072 ();
 sg13g2_fill_8 FILLER_115_1080 ();
 sg13g2_fill_8 FILLER_115_1088 ();
 sg13g2_fill_8 FILLER_115_1096 ();
 sg13g2_fill_8 FILLER_115_1104 ();
 sg13g2_fill_8 FILLER_115_1112 ();
 sg13g2_fill_8 FILLER_115_1120 ();
 sg13g2_fill_8 FILLER_115_1128 ();
 sg13g2_fill_8 FILLER_115_1136 ();
 sg13g2_fill_8 FILLER_116_0 ();
 sg13g2_fill_8 FILLER_116_8 ();
 sg13g2_fill_8 FILLER_116_16 ();
 sg13g2_fill_8 FILLER_116_24 ();
 sg13g2_fill_8 FILLER_116_32 ();
 sg13g2_fill_8 FILLER_116_40 ();
 sg13g2_fill_8 FILLER_116_48 ();
 sg13g2_fill_8 FILLER_116_56 ();
 sg13g2_fill_8 FILLER_116_64 ();
 sg13g2_fill_8 FILLER_116_72 ();
 sg13g2_fill_8 FILLER_116_80 ();
 sg13g2_fill_8 FILLER_116_88 ();
 sg13g2_fill_8 FILLER_116_96 ();
 sg13g2_fill_8 FILLER_116_104 ();
 sg13g2_fill_8 FILLER_116_112 ();
 sg13g2_fill_8 FILLER_116_120 ();
 sg13g2_fill_8 FILLER_116_128 ();
 sg13g2_fill_8 FILLER_116_136 ();
 sg13g2_fill_8 FILLER_116_144 ();
 sg13g2_fill_8 FILLER_116_152 ();
 sg13g2_fill_8 FILLER_116_160 ();
 sg13g2_fill_8 FILLER_116_168 ();
 sg13g2_fill_8 FILLER_116_176 ();
 sg13g2_fill_8 FILLER_116_184 ();
 sg13g2_fill_8 FILLER_116_192 ();
 sg13g2_fill_8 FILLER_116_200 ();
 sg13g2_fill_8 FILLER_116_208 ();
 sg13g2_fill_8 FILLER_116_216 ();
 sg13g2_fill_8 FILLER_116_224 ();
 sg13g2_fill_8 FILLER_116_232 ();
 sg13g2_fill_8 FILLER_116_240 ();
 sg13g2_fill_8 FILLER_116_248 ();
 sg13g2_fill_8 FILLER_116_256 ();
 sg13g2_fill_8 FILLER_116_264 ();
 sg13g2_fill_8 FILLER_116_272 ();
 sg13g2_fill_8 FILLER_116_280 ();
 sg13g2_fill_8 FILLER_116_288 ();
 sg13g2_fill_8 FILLER_116_296 ();
 sg13g2_fill_8 FILLER_116_304 ();
 sg13g2_fill_8 FILLER_116_312 ();
 sg13g2_fill_8 FILLER_116_320 ();
 sg13g2_fill_8 FILLER_116_328 ();
 sg13g2_fill_8 FILLER_116_336 ();
 sg13g2_fill_8 FILLER_116_344 ();
 sg13g2_fill_8 FILLER_116_352 ();
 sg13g2_fill_8 FILLER_116_360 ();
 sg13g2_fill_8 FILLER_116_368 ();
 sg13g2_fill_8 FILLER_116_376 ();
 sg13g2_fill_8 FILLER_116_384 ();
 sg13g2_fill_8 FILLER_116_392 ();
 sg13g2_fill_8 FILLER_116_400 ();
 sg13g2_fill_8 FILLER_116_408 ();
 sg13g2_fill_8 FILLER_116_416 ();
 sg13g2_fill_8 FILLER_116_424 ();
 sg13g2_fill_8 FILLER_116_432 ();
 sg13g2_fill_8 FILLER_116_440 ();
 sg13g2_fill_8 FILLER_116_448 ();
 sg13g2_fill_8 FILLER_116_456 ();
 sg13g2_fill_8 FILLER_116_464 ();
 sg13g2_fill_8 FILLER_116_472 ();
 sg13g2_fill_8 FILLER_116_480 ();
 sg13g2_fill_8 FILLER_116_488 ();
 sg13g2_fill_8 FILLER_116_496 ();
 sg13g2_fill_8 FILLER_116_504 ();
 sg13g2_fill_8 FILLER_116_512 ();
 sg13g2_fill_8 FILLER_116_520 ();
 sg13g2_fill_8 FILLER_116_528 ();
 sg13g2_fill_8 FILLER_116_536 ();
 sg13g2_fill_8 FILLER_116_544 ();
 sg13g2_fill_8 FILLER_116_552 ();
 sg13g2_fill_8 FILLER_116_560 ();
 sg13g2_fill_8 FILLER_116_568 ();
 sg13g2_fill_8 FILLER_116_576 ();
 sg13g2_fill_8 FILLER_116_584 ();
 sg13g2_fill_8 FILLER_116_592 ();
 sg13g2_fill_8 FILLER_116_600 ();
 sg13g2_fill_8 FILLER_116_608 ();
 sg13g2_fill_8 FILLER_116_616 ();
 sg13g2_fill_8 FILLER_116_624 ();
 sg13g2_fill_8 FILLER_116_632 ();
 sg13g2_fill_8 FILLER_116_640 ();
 sg13g2_fill_8 FILLER_116_648 ();
 sg13g2_fill_8 FILLER_116_656 ();
 sg13g2_fill_8 FILLER_116_664 ();
 sg13g2_fill_8 FILLER_116_672 ();
 sg13g2_fill_8 FILLER_116_680 ();
 sg13g2_fill_8 FILLER_116_688 ();
 sg13g2_fill_8 FILLER_116_696 ();
 sg13g2_fill_8 FILLER_116_704 ();
 sg13g2_fill_8 FILLER_116_712 ();
 sg13g2_fill_8 FILLER_116_720 ();
 sg13g2_fill_8 FILLER_116_728 ();
 sg13g2_fill_8 FILLER_116_736 ();
 sg13g2_fill_8 FILLER_116_744 ();
 sg13g2_fill_8 FILLER_116_752 ();
 sg13g2_fill_8 FILLER_116_760 ();
 sg13g2_fill_8 FILLER_116_768 ();
 sg13g2_fill_8 FILLER_116_776 ();
 sg13g2_fill_8 FILLER_116_784 ();
 sg13g2_fill_8 FILLER_116_792 ();
 sg13g2_fill_8 FILLER_116_800 ();
 sg13g2_fill_8 FILLER_116_808 ();
 sg13g2_fill_8 FILLER_116_816 ();
 sg13g2_fill_8 FILLER_116_824 ();
 sg13g2_fill_8 FILLER_116_832 ();
 sg13g2_fill_8 FILLER_116_840 ();
 sg13g2_fill_8 FILLER_116_848 ();
 sg13g2_fill_8 FILLER_116_856 ();
 sg13g2_fill_8 FILLER_116_864 ();
 sg13g2_fill_8 FILLER_116_872 ();
 sg13g2_fill_8 FILLER_116_880 ();
 sg13g2_fill_8 FILLER_116_888 ();
 sg13g2_fill_8 FILLER_116_896 ();
 sg13g2_fill_8 FILLER_116_904 ();
 sg13g2_fill_8 FILLER_116_912 ();
 sg13g2_fill_8 FILLER_116_920 ();
 sg13g2_fill_8 FILLER_116_928 ();
 sg13g2_fill_8 FILLER_116_936 ();
 sg13g2_fill_8 FILLER_116_944 ();
 sg13g2_fill_8 FILLER_116_952 ();
 sg13g2_fill_8 FILLER_116_960 ();
 sg13g2_fill_8 FILLER_116_968 ();
 sg13g2_fill_8 FILLER_116_976 ();
 sg13g2_fill_8 FILLER_116_984 ();
 sg13g2_fill_8 FILLER_116_992 ();
 sg13g2_fill_8 FILLER_116_1000 ();
 sg13g2_fill_8 FILLER_116_1008 ();
 sg13g2_fill_8 FILLER_116_1016 ();
 sg13g2_fill_8 FILLER_116_1024 ();
 sg13g2_fill_8 FILLER_116_1032 ();
 sg13g2_fill_8 FILLER_116_1040 ();
 sg13g2_fill_8 FILLER_116_1048 ();
 sg13g2_fill_8 FILLER_116_1056 ();
 sg13g2_fill_8 FILLER_116_1064 ();
 sg13g2_fill_8 FILLER_116_1072 ();
 sg13g2_fill_8 FILLER_116_1080 ();
 sg13g2_fill_8 FILLER_116_1088 ();
 sg13g2_fill_8 FILLER_116_1096 ();
 sg13g2_fill_8 FILLER_116_1104 ();
 sg13g2_fill_8 FILLER_116_1112 ();
 sg13g2_fill_8 FILLER_116_1120 ();
 sg13g2_fill_8 FILLER_116_1128 ();
 sg13g2_fill_8 FILLER_116_1136 ();
 sg13g2_fill_8 FILLER_117_0 ();
 sg13g2_fill_8 FILLER_117_8 ();
 sg13g2_fill_8 FILLER_117_16 ();
 sg13g2_fill_8 FILLER_117_24 ();
 sg13g2_fill_8 FILLER_117_32 ();
 sg13g2_fill_8 FILLER_117_40 ();
 sg13g2_fill_8 FILLER_117_48 ();
 sg13g2_fill_8 FILLER_117_56 ();
 sg13g2_fill_8 FILLER_117_64 ();
 sg13g2_fill_8 FILLER_117_72 ();
 sg13g2_fill_8 FILLER_117_80 ();
 sg13g2_fill_8 FILLER_117_88 ();
 sg13g2_fill_8 FILLER_117_96 ();
 sg13g2_fill_8 FILLER_117_104 ();
 sg13g2_fill_8 FILLER_117_112 ();
 sg13g2_fill_8 FILLER_117_120 ();
 sg13g2_fill_8 FILLER_117_128 ();
 sg13g2_fill_8 FILLER_117_136 ();
 sg13g2_fill_8 FILLER_117_144 ();
 sg13g2_fill_8 FILLER_117_152 ();
 sg13g2_fill_8 FILLER_117_160 ();
 sg13g2_fill_8 FILLER_117_168 ();
 sg13g2_fill_8 FILLER_117_176 ();
 sg13g2_fill_8 FILLER_117_184 ();
 sg13g2_fill_8 FILLER_117_192 ();
 sg13g2_fill_8 FILLER_117_200 ();
 sg13g2_fill_8 FILLER_117_208 ();
 sg13g2_fill_8 FILLER_117_216 ();
 sg13g2_fill_8 FILLER_117_224 ();
 sg13g2_fill_8 FILLER_117_232 ();
 sg13g2_fill_8 FILLER_117_240 ();
 sg13g2_fill_8 FILLER_117_248 ();
 sg13g2_fill_8 FILLER_117_256 ();
 sg13g2_fill_8 FILLER_117_264 ();
 sg13g2_fill_8 FILLER_117_272 ();
 sg13g2_fill_8 FILLER_117_280 ();
 sg13g2_fill_8 FILLER_117_288 ();
 sg13g2_fill_8 FILLER_117_296 ();
 sg13g2_fill_8 FILLER_117_304 ();
 sg13g2_fill_8 FILLER_117_312 ();
 sg13g2_fill_8 FILLER_117_320 ();
 sg13g2_fill_8 FILLER_117_328 ();
 sg13g2_fill_8 FILLER_117_336 ();
 sg13g2_fill_8 FILLER_117_344 ();
 sg13g2_fill_8 FILLER_117_352 ();
 sg13g2_fill_8 FILLER_117_360 ();
 sg13g2_fill_8 FILLER_117_368 ();
 sg13g2_fill_8 FILLER_117_376 ();
 sg13g2_fill_8 FILLER_117_384 ();
 sg13g2_fill_8 FILLER_117_392 ();
 sg13g2_fill_8 FILLER_117_400 ();
 sg13g2_fill_8 FILLER_117_408 ();
 sg13g2_fill_8 FILLER_117_416 ();
 sg13g2_fill_8 FILLER_117_424 ();
 sg13g2_fill_8 FILLER_117_432 ();
 sg13g2_fill_8 FILLER_117_440 ();
 sg13g2_fill_8 FILLER_117_448 ();
 sg13g2_fill_8 FILLER_117_456 ();
 sg13g2_fill_8 FILLER_117_464 ();
 sg13g2_fill_8 FILLER_117_472 ();
 sg13g2_fill_8 FILLER_117_480 ();
 sg13g2_fill_8 FILLER_117_488 ();
 sg13g2_fill_8 FILLER_117_496 ();
 sg13g2_fill_8 FILLER_117_504 ();
 sg13g2_fill_8 FILLER_117_512 ();
 sg13g2_fill_8 FILLER_117_520 ();
 sg13g2_fill_8 FILLER_117_528 ();
 sg13g2_fill_8 FILLER_117_536 ();
 sg13g2_fill_8 FILLER_117_544 ();
 sg13g2_fill_8 FILLER_117_552 ();
 sg13g2_fill_8 FILLER_117_560 ();
 sg13g2_fill_8 FILLER_117_568 ();
 sg13g2_fill_8 FILLER_117_576 ();
 sg13g2_fill_8 FILLER_117_584 ();
 sg13g2_fill_8 FILLER_117_592 ();
 sg13g2_fill_8 FILLER_117_600 ();
 sg13g2_fill_8 FILLER_117_608 ();
 sg13g2_fill_8 FILLER_117_616 ();
 sg13g2_fill_8 FILLER_117_624 ();
 sg13g2_fill_8 FILLER_117_632 ();
 sg13g2_fill_8 FILLER_117_640 ();
 sg13g2_fill_8 FILLER_117_648 ();
 sg13g2_fill_8 FILLER_117_656 ();
 sg13g2_fill_8 FILLER_117_664 ();
 sg13g2_fill_8 FILLER_117_672 ();
 sg13g2_fill_8 FILLER_117_680 ();
 sg13g2_fill_8 FILLER_117_688 ();
 sg13g2_fill_8 FILLER_117_696 ();
 sg13g2_fill_8 FILLER_117_704 ();
 sg13g2_fill_8 FILLER_117_712 ();
 sg13g2_fill_8 FILLER_117_720 ();
 sg13g2_fill_8 FILLER_117_728 ();
 sg13g2_fill_8 FILLER_117_736 ();
 sg13g2_fill_8 FILLER_117_744 ();
 sg13g2_fill_8 FILLER_117_752 ();
 sg13g2_fill_8 FILLER_117_760 ();
 sg13g2_fill_8 FILLER_117_768 ();
 sg13g2_fill_8 FILLER_117_776 ();
 sg13g2_fill_8 FILLER_117_784 ();
 sg13g2_fill_8 FILLER_117_792 ();
 sg13g2_fill_8 FILLER_117_800 ();
 sg13g2_fill_8 FILLER_117_808 ();
 sg13g2_fill_8 FILLER_117_816 ();
 sg13g2_fill_8 FILLER_117_824 ();
 sg13g2_fill_8 FILLER_117_832 ();
 sg13g2_fill_8 FILLER_117_840 ();
 sg13g2_fill_8 FILLER_117_848 ();
 sg13g2_fill_8 FILLER_117_856 ();
 sg13g2_fill_8 FILLER_117_864 ();
 sg13g2_fill_8 FILLER_117_872 ();
 sg13g2_fill_8 FILLER_117_880 ();
 sg13g2_fill_8 FILLER_117_888 ();
 sg13g2_fill_8 FILLER_117_896 ();
 sg13g2_fill_8 FILLER_117_904 ();
 sg13g2_fill_8 FILLER_117_912 ();
 sg13g2_fill_8 FILLER_117_920 ();
 sg13g2_fill_8 FILLER_117_928 ();
 sg13g2_fill_8 FILLER_117_936 ();
 sg13g2_fill_8 FILLER_117_944 ();
 sg13g2_fill_8 FILLER_117_952 ();
 sg13g2_fill_8 FILLER_117_960 ();
 sg13g2_fill_8 FILLER_117_968 ();
 sg13g2_fill_8 FILLER_117_976 ();
 sg13g2_fill_8 FILLER_117_984 ();
 sg13g2_fill_8 FILLER_117_992 ();
 sg13g2_fill_8 FILLER_117_1000 ();
 sg13g2_fill_8 FILLER_117_1008 ();
 sg13g2_fill_8 FILLER_117_1016 ();
 sg13g2_fill_8 FILLER_117_1024 ();
 sg13g2_fill_8 FILLER_117_1032 ();
 sg13g2_fill_8 FILLER_117_1040 ();
 sg13g2_fill_8 FILLER_117_1048 ();
 sg13g2_fill_8 FILLER_117_1056 ();
 sg13g2_fill_8 FILLER_117_1064 ();
 sg13g2_fill_8 FILLER_117_1072 ();
 sg13g2_fill_8 FILLER_117_1080 ();
 sg13g2_fill_8 FILLER_117_1088 ();
 sg13g2_fill_8 FILLER_117_1096 ();
 sg13g2_fill_8 FILLER_117_1104 ();
 sg13g2_fill_8 FILLER_117_1112 ();
 sg13g2_fill_8 FILLER_117_1120 ();
 sg13g2_fill_8 FILLER_117_1128 ();
 sg13g2_fill_8 FILLER_117_1136 ();
 sg13g2_fill_8 FILLER_118_0 ();
 sg13g2_fill_8 FILLER_118_8 ();
 sg13g2_fill_8 FILLER_118_16 ();
 sg13g2_fill_8 FILLER_118_24 ();
 sg13g2_fill_8 FILLER_118_32 ();
 sg13g2_fill_8 FILLER_118_40 ();
 sg13g2_fill_8 FILLER_118_48 ();
 sg13g2_fill_8 FILLER_118_56 ();
 sg13g2_fill_8 FILLER_118_64 ();
 sg13g2_fill_8 FILLER_118_72 ();
 sg13g2_fill_8 FILLER_118_80 ();
 sg13g2_fill_8 FILLER_118_88 ();
 sg13g2_fill_8 FILLER_118_96 ();
 sg13g2_fill_8 FILLER_118_104 ();
 sg13g2_fill_8 FILLER_118_112 ();
 sg13g2_fill_8 FILLER_118_120 ();
 sg13g2_fill_8 FILLER_118_128 ();
 sg13g2_fill_8 FILLER_118_136 ();
 sg13g2_fill_8 FILLER_118_144 ();
 sg13g2_fill_8 FILLER_118_152 ();
 sg13g2_fill_8 FILLER_118_160 ();
 sg13g2_fill_8 FILLER_118_168 ();
 sg13g2_fill_8 FILLER_118_176 ();
 sg13g2_fill_8 FILLER_118_184 ();
 sg13g2_fill_8 FILLER_118_192 ();
 sg13g2_fill_8 FILLER_118_200 ();
 sg13g2_fill_8 FILLER_118_208 ();
 sg13g2_fill_8 FILLER_118_216 ();
 sg13g2_fill_8 FILLER_118_224 ();
 sg13g2_fill_8 FILLER_118_232 ();
 sg13g2_fill_8 FILLER_118_240 ();
 sg13g2_fill_8 FILLER_118_248 ();
 sg13g2_fill_8 FILLER_118_256 ();
 sg13g2_fill_8 FILLER_118_264 ();
 sg13g2_fill_8 FILLER_118_272 ();
 sg13g2_fill_8 FILLER_118_280 ();
 sg13g2_fill_8 FILLER_118_288 ();
 sg13g2_fill_8 FILLER_118_296 ();
 sg13g2_fill_8 FILLER_118_304 ();
 sg13g2_fill_8 FILLER_118_312 ();
 sg13g2_fill_8 FILLER_118_320 ();
 sg13g2_fill_8 FILLER_118_328 ();
 sg13g2_fill_8 FILLER_118_336 ();
 sg13g2_fill_8 FILLER_118_344 ();
 sg13g2_fill_8 FILLER_118_352 ();
 sg13g2_fill_8 FILLER_118_360 ();
 sg13g2_fill_8 FILLER_118_368 ();
 sg13g2_fill_8 FILLER_118_376 ();
 sg13g2_fill_8 FILLER_118_384 ();
 sg13g2_fill_8 FILLER_118_392 ();
 sg13g2_fill_8 FILLER_118_400 ();
 sg13g2_fill_8 FILLER_118_408 ();
 sg13g2_fill_8 FILLER_118_416 ();
 sg13g2_fill_8 FILLER_118_424 ();
 sg13g2_fill_8 FILLER_118_432 ();
 sg13g2_fill_8 FILLER_118_440 ();
 sg13g2_fill_8 FILLER_118_448 ();
 sg13g2_fill_8 FILLER_118_456 ();
 sg13g2_fill_8 FILLER_118_464 ();
 sg13g2_fill_8 FILLER_118_472 ();
 sg13g2_fill_8 FILLER_118_480 ();
 sg13g2_fill_8 FILLER_118_488 ();
 sg13g2_fill_8 FILLER_118_496 ();
 sg13g2_fill_8 FILLER_118_504 ();
 sg13g2_fill_8 FILLER_118_512 ();
 sg13g2_fill_8 FILLER_118_520 ();
 sg13g2_fill_8 FILLER_118_528 ();
 sg13g2_fill_8 FILLER_118_536 ();
 sg13g2_fill_8 FILLER_118_544 ();
 sg13g2_fill_8 FILLER_118_552 ();
 sg13g2_fill_8 FILLER_118_560 ();
 sg13g2_fill_8 FILLER_118_568 ();
 sg13g2_fill_8 FILLER_118_576 ();
 sg13g2_fill_8 FILLER_118_584 ();
 sg13g2_fill_8 FILLER_118_592 ();
 sg13g2_fill_8 FILLER_118_600 ();
 sg13g2_fill_8 FILLER_118_608 ();
 sg13g2_fill_8 FILLER_118_616 ();
 sg13g2_fill_8 FILLER_118_624 ();
 sg13g2_fill_8 FILLER_118_632 ();
 sg13g2_fill_8 FILLER_118_640 ();
 sg13g2_fill_8 FILLER_118_648 ();
 sg13g2_fill_8 FILLER_118_656 ();
 sg13g2_fill_8 FILLER_118_664 ();
 sg13g2_fill_8 FILLER_118_672 ();
 sg13g2_fill_8 FILLER_118_680 ();
 sg13g2_fill_8 FILLER_118_688 ();
 sg13g2_fill_8 FILLER_118_696 ();
 sg13g2_fill_8 FILLER_118_704 ();
 sg13g2_fill_8 FILLER_118_712 ();
 sg13g2_fill_8 FILLER_118_720 ();
 sg13g2_fill_8 FILLER_118_728 ();
 sg13g2_fill_8 FILLER_118_736 ();
 sg13g2_fill_8 FILLER_118_744 ();
 sg13g2_fill_8 FILLER_118_752 ();
 sg13g2_fill_8 FILLER_118_760 ();
 sg13g2_fill_8 FILLER_118_768 ();
 sg13g2_fill_8 FILLER_118_776 ();
 sg13g2_fill_8 FILLER_118_784 ();
 sg13g2_fill_8 FILLER_118_792 ();
 sg13g2_fill_8 FILLER_118_800 ();
 sg13g2_fill_8 FILLER_118_808 ();
 sg13g2_fill_8 FILLER_118_816 ();
 sg13g2_fill_8 FILLER_118_824 ();
 sg13g2_fill_8 FILLER_118_832 ();
 sg13g2_fill_8 FILLER_118_840 ();
 sg13g2_fill_8 FILLER_118_848 ();
 sg13g2_fill_8 FILLER_118_856 ();
 sg13g2_fill_8 FILLER_118_864 ();
 sg13g2_fill_8 FILLER_118_872 ();
 sg13g2_fill_8 FILLER_118_880 ();
 sg13g2_fill_8 FILLER_118_888 ();
 sg13g2_fill_8 FILLER_118_896 ();
 sg13g2_fill_8 FILLER_118_904 ();
 sg13g2_fill_8 FILLER_118_912 ();
 sg13g2_fill_8 FILLER_118_920 ();
 sg13g2_fill_8 FILLER_118_928 ();
 sg13g2_fill_8 FILLER_118_936 ();
 sg13g2_fill_8 FILLER_118_944 ();
 sg13g2_fill_8 FILLER_118_952 ();
 sg13g2_fill_8 FILLER_118_960 ();
 sg13g2_fill_8 FILLER_118_968 ();
 sg13g2_fill_8 FILLER_118_976 ();
 sg13g2_fill_8 FILLER_118_984 ();
 sg13g2_fill_8 FILLER_118_992 ();
 sg13g2_fill_8 FILLER_118_1000 ();
 sg13g2_fill_8 FILLER_118_1008 ();
 sg13g2_fill_8 FILLER_118_1016 ();
 sg13g2_fill_8 FILLER_118_1024 ();
 sg13g2_fill_8 FILLER_118_1032 ();
 sg13g2_fill_8 FILLER_118_1040 ();
 sg13g2_fill_8 FILLER_118_1048 ();
 sg13g2_fill_8 FILLER_118_1056 ();
 sg13g2_fill_8 FILLER_118_1064 ();
 sg13g2_fill_8 FILLER_118_1072 ();
 sg13g2_fill_8 FILLER_118_1080 ();
 sg13g2_fill_8 FILLER_118_1088 ();
 sg13g2_fill_8 FILLER_118_1096 ();
 sg13g2_fill_8 FILLER_118_1104 ();
 sg13g2_fill_8 FILLER_118_1112 ();
 sg13g2_fill_8 FILLER_118_1120 ();
 sg13g2_fill_8 FILLER_118_1128 ();
 sg13g2_fill_8 FILLER_118_1136 ();
 sg13g2_fill_8 FILLER_119_0 ();
 sg13g2_fill_8 FILLER_119_8 ();
 sg13g2_fill_8 FILLER_119_16 ();
 sg13g2_fill_8 FILLER_119_24 ();
 sg13g2_fill_8 FILLER_119_32 ();
 sg13g2_fill_8 FILLER_119_40 ();
 sg13g2_fill_8 FILLER_119_48 ();
 sg13g2_fill_8 FILLER_119_56 ();
 sg13g2_fill_8 FILLER_119_64 ();
 sg13g2_fill_8 FILLER_119_72 ();
 sg13g2_fill_8 FILLER_119_80 ();
 sg13g2_fill_8 FILLER_119_88 ();
 sg13g2_fill_8 FILLER_119_96 ();
 sg13g2_fill_8 FILLER_119_104 ();
 sg13g2_fill_8 FILLER_119_112 ();
 sg13g2_fill_8 FILLER_119_120 ();
 sg13g2_fill_8 FILLER_119_128 ();
 sg13g2_fill_8 FILLER_119_136 ();
 sg13g2_fill_8 FILLER_119_144 ();
 sg13g2_fill_8 FILLER_119_152 ();
 sg13g2_fill_8 FILLER_119_160 ();
 sg13g2_fill_8 FILLER_119_168 ();
 sg13g2_fill_8 FILLER_119_176 ();
 sg13g2_fill_8 FILLER_119_184 ();
 sg13g2_fill_8 FILLER_119_192 ();
 sg13g2_fill_8 FILLER_119_200 ();
 sg13g2_fill_8 FILLER_119_208 ();
 sg13g2_fill_8 FILLER_119_216 ();
 sg13g2_fill_8 FILLER_119_224 ();
 sg13g2_fill_8 FILLER_119_232 ();
 sg13g2_fill_8 FILLER_119_240 ();
 sg13g2_fill_8 FILLER_119_248 ();
 sg13g2_fill_8 FILLER_119_256 ();
 sg13g2_fill_8 FILLER_119_264 ();
 sg13g2_fill_8 FILLER_119_272 ();
 sg13g2_fill_8 FILLER_119_280 ();
 sg13g2_fill_8 FILLER_119_288 ();
 sg13g2_fill_8 FILLER_119_296 ();
 sg13g2_fill_8 FILLER_119_304 ();
 sg13g2_fill_8 FILLER_119_312 ();
 sg13g2_fill_8 FILLER_119_320 ();
 sg13g2_fill_8 FILLER_119_328 ();
 sg13g2_fill_8 FILLER_119_336 ();
 sg13g2_fill_8 FILLER_119_344 ();
 sg13g2_fill_8 FILLER_119_352 ();
 sg13g2_fill_8 FILLER_119_360 ();
 sg13g2_fill_8 FILLER_119_368 ();
 sg13g2_fill_8 FILLER_119_376 ();
 sg13g2_fill_8 FILLER_119_384 ();
 sg13g2_fill_8 FILLER_119_392 ();
 sg13g2_fill_8 FILLER_119_400 ();
 sg13g2_fill_8 FILLER_119_408 ();
 sg13g2_fill_8 FILLER_119_416 ();
 sg13g2_fill_8 FILLER_119_424 ();
 sg13g2_fill_8 FILLER_119_432 ();
 sg13g2_fill_8 FILLER_119_440 ();
 sg13g2_fill_8 FILLER_119_448 ();
 sg13g2_fill_8 FILLER_119_456 ();
 sg13g2_fill_8 FILLER_119_464 ();
 sg13g2_fill_8 FILLER_119_472 ();
 sg13g2_fill_8 FILLER_119_480 ();
 sg13g2_fill_8 FILLER_119_488 ();
 sg13g2_fill_8 FILLER_119_496 ();
 sg13g2_fill_8 FILLER_119_504 ();
 sg13g2_fill_8 FILLER_119_512 ();
 sg13g2_fill_8 FILLER_119_520 ();
 sg13g2_fill_8 FILLER_119_528 ();
 sg13g2_fill_8 FILLER_119_536 ();
 sg13g2_fill_8 FILLER_119_544 ();
 sg13g2_fill_8 FILLER_119_552 ();
 sg13g2_fill_8 FILLER_119_560 ();
 sg13g2_fill_8 FILLER_119_568 ();
 sg13g2_fill_8 FILLER_119_576 ();
 sg13g2_fill_8 FILLER_119_584 ();
 sg13g2_fill_8 FILLER_119_592 ();
 sg13g2_fill_8 FILLER_119_600 ();
 sg13g2_fill_8 FILLER_119_608 ();
 sg13g2_fill_8 FILLER_119_616 ();
 sg13g2_fill_8 FILLER_119_624 ();
 sg13g2_fill_8 FILLER_119_632 ();
 sg13g2_fill_8 FILLER_119_640 ();
 sg13g2_fill_8 FILLER_119_648 ();
 sg13g2_fill_8 FILLER_119_656 ();
 sg13g2_fill_8 FILLER_119_664 ();
 sg13g2_fill_8 FILLER_119_672 ();
 sg13g2_fill_8 FILLER_119_680 ();
 sg13g2_fill_8 FILLER_119_688 ();
 sg13g2_fill_8 FILLER_119_696 ();
 sg13g2_fill_8 FILLER_119_704 ();
 sg13g2_fill_8 FILLER_119_712 ();
 sg13g2_fill_8 FILLER_119_720 ();
 sg13g2_fill_8 FILLER_119_728 ();
 sg13g2_fill_8 FILLER_119_736 ();
 sg13g2_fill_8 FILLER_119_744 ();
 sg13g2_fill_8 FILLER_119_752 ();
 sg13g2_fill_8 FILLER_119_760 ();
 sg13g2_fill_8 FILLER_119_768 ();
 sg13g2_fill_8 FILLER_119_776 ();
 sg13g2_fill_8 FILLER_119_784 ();
 sg13g2_fill_8 FILLER_119_792 ();
 sg13g2_fill_8 FILLER_119_800 ();
 sg13g2_fill_8 FILLER_119_808 ();
 sg13g2_fill_8 FILLER_119_816 ();
 sg13g2_fill_8 FILLER_119_824 ();
 sg13g2_fill_8 FILLER_119_832 ();
 sg13g2_fill_8 FILLER_119_840 ();
 sg13g2_fill_8 FILLER_119_848 ();
 sg13g2_fill_8 FILLER_119_856 ();
 sg13g2_fill_8 FILLER_119_864 ();
 sg13g2_fill_8 FILLER_119_872 ();
 sg13g2_fill_8 FILLER_119_880 ();
 sg13g2_fill_8 FILLER_119_888 ();
 sg13g2_fill_8 FILLER_119_896 ();
 sg13g2_fill_8 FILLER_119_904 ();
 sg13g2_fill_8 FILLER_119_912 ();
 sg13g2_fill_8 FILLER_119_920 ();
 sg13g2_fill_8 FILLER_119_928 ();
 sg13g2_fill_8 FILLER_119_936 ();
 sg13g2_fill_8 FILLER_119_944 ();
 sg13g2_fill_8 FILLER_119_952 ();
 sg13g2_fill_8 FILLER_119_960 ();
 sg13g2_fill_8 FILLER_119_968 ();
 sg13g2_fill_8 FILLER_119_976 ();
 sg13g2_fill_8 FILLER_119_984 ();
 sg13g2_fill_8 FILLER_119_992 ();
 sg13g2_fill_8 FILLER_119_1000 ();
 sg13g2_fill_8 FILLER_119_1008 ();
 sg13g2_fill_8 FILLER_119_1016 ();
 sg13g2_fill_8 FILLER_119_1024 ();
 sg13g2_fill_8 FILLER_119_1032 ();
 sg13g2_fill_8 FILLER_119_1040 ();
 sg13g2_fill_8 FILLER_119_1048 ();
 sg13g2_fill_8 FILLER_119_1056 ();
 sg13g2_fill_8 FILLER_119_1064 ();
 sg13g2_fill_8 FILLER_119_1072 ();
 sg13g2_fill_8 FILLER_119_1080 ();
 sg13g2_fill_8 FILLER_119_1088 ();
 sg13g2_fill_8 FILLER_119_1096 ();
 sg13g2_fill_8 FILLER_119_1104 ();
 sg13g2_fill_8 FILLER_119_1112 ();
 sg13g2_fill_8 FILLER_119_1120 ();
 sg13g2_fill_8 FILLER_119_1128 ();
 sg13g2_fill_8 FILLER_119_1136 ();
 sg13g2_fill_8 FILLER_120_0 ();
 sg13g2_fill_8 FILLER_120_8 ();
 sg13g2_fill_8 FILLER_120_16 ();
 sg13g2_fill_8 FILLER_120_24 ();
 sg13g2_fill_8 FILLER_120_32 ();
 sg13g2_fill_8 FILLER_120_40 ();
 sg13g2_fill_8 FILLER_120_48 ();
 sg13g2_fill_8 FILLER_120_56 ();
 sg13g2_fill_8 FILLER_120_64 ();
 sg13g2_fill_8 FILLER_120_72 ();
 sg13g2_fill_8 FILLER_120_80 ();
 sg13g2_fill_8 FILLER_120_88 ();
 sg13g2_fill_8 FILLER_120_96 ();
 sg13g2_fill_8 FILLER_120_104 ();
 sg13g2_fill_8 FILLER_120_112 ();
 sg13g2_fill_8 FILLER_120_120 ();
 sg13g2_fill_8 FILLER_120_128 ();
 sg13g2_fill_8 FILLER_120_136 ();
 sg13g2_fill_8 FILLER_120_144 ();
 sg13g2_fill_8 FILLER_120_152 ();
 sg13g2_fill_8 FILLER_120_160 ();
 sg13g2_fill_8 FILLER_120_168 ();
 sg13g2_fill_8 FILLER_120_176 ();
 sg13g2_fill_8 FILLER_120_184 ();
 sg13g2_fill_8 FILLER_120_192 ();
 sg13g2_fill_8 FILLER_120_200 ();
 sg13g2_fill_8 FILLER_120_208 ();
 sg13g2_fill_8 FILLER_120_216 ();
 sg13g2_fill_8 FILLER_120_224 ();
 sg13g2_fill_8 FILLER_120_232 ();
 sg13g2_fill_8 FILLER_120_240 ();
 sg13g2_fill_8 FILLER_120_248 ();
 sg13g2_fill_8 FILLER_120_256 ();
 sg13g2_fill_8 FILLER_120_264 ();
 sg13g2_fill_8 FILLER_120_272 ();
 sg13g2_fill_8 FILLER_120_280 ();
 sg13g2_fill_8 FILLER_120_288 ();
 sg13g2_fill_8 FILLER_120_296 ();
 sg13g2_fill_8 FILLER_120_304 ();
 sg13g2_fill_8 FILLER_120_312 ();
 sg13g2_fill_8 FILLER_120_320 ();
 sg13g2_fill_8 FILLER_120_328 ();
 sg13g2_fill_8 FILLER_120_336 ();
 sg13g2_fill_8 FILLER_120_344 ();
 sg13g2_fill_8 FILLER_120_352 ();
 sg13g2_fill_8 FILLER_120_360 ();
 sg13g2_fill_8 FILLER_120_368 ();
 sg13g2_fill_8 FILLER_120_376 ();
 sg13g2_fill_8 FILLER_120_384 ();
 sg13g2_fill_8 FILLER_120_392 ();
 sg13g2_fill_8 FILLER_120_400 ();
 sg13g2_fill_8 FILLER_120_408 ();
 sg13g2_fill_8 FILLER_120_416 ();
 sg13g2_fill_8 FILLER_120_424 ();
 sg13g2_fill_8 FILLER_120_432 ();
 sg13g2_fill_8 FILLER_120_440 ();
 sg13g2_fill_8 FILLER_120_448 ();
 sg13g2_fill_8 FILLER_120_456 ();
 sg13g2_fill_8 FILLER_120_464 ();
 sg13g2_fill_8 FILLER_120_472 ();
 sg13g2_fill_8 FILLER_120_480 ();
 sg13g2_fill_8 FILLER_120_488 ();
 sg13g2_fill_8 FILLER_120_496 ();
 sg13g2_fill_8 FILLER_120_504 ();
 sg13g2_fill_8 FILLER_120_512 ();
 sg13g2_fill_8 FILLER_120_520 ();
 sg13g2_fill_8 FILLER_120_528 ();
 sg13g2_fill_8 FILLER_120_536 ();
 sg13g2_fill_8 FILLER_120_544 ();
 sg13g2_fill_8 FILLER_120_552 ();
 sg13g2_fill_8 FILLER_120_560 ();
 sg13g2_fill_8 FILLER_120_568 ();
 sg13g2_fill_8 FILLER_120_576 ();
 sg13g2_fill_8 FILLER_120_584 ();
 sg13g2_fill_8 FILLER_120_592 ();
 sg13g2_fill_8 FILLER_120_600 ();
 sg13g2_fill_8 FILLER_120_608 ();
 sg13g2_fill_8 FILLER_120_616 ();
 sg13g2_fill_8 FILLER_120_624 ();
 sg13g2_fill_8 FILLER_120_632 ();
 sg13g2_fill_8 FILLER_120_640 ();
 sg13g2_fill_8 FILLER_120_648 ();
 sg13g2_fill_8 FILLER_120_656 ();
 sg13g2_fill_8 FILLER_120_664 ();
 sg13g2_fill_8 FILLER_120_672 ();
 sg13g2_fill_8 FILLER_120_680 ();
 sg13g2_fill_8 FILLER_120_688 ();
 sg13g2_fill_8 FILLER_120_696 ();
 sg13g2_fill_8 FILLER_120_704 ();
 sg13g2_fill_8 FILLER_120_712 ();
 sg13g2_fill_8 FILLER_120_720 ();
 sg13g2_fill_8 FILLER_120_728 ();
 sg13g2_fill_8 FILLER_120_736 ();
 sg13g2_fill_8 FILLER_120_744 ();
 sg13g2_fill_8 FILLER_120_752 ();
 sg13g2_fill_8 FILLER_120_760 ();
 sg13g2_fill_8 FILLER_120_768 ();
 sg13g2_fill_8 FILLER_120_776 ();
 sg13g2_fill_8 FILLER_120_784 ();
 sg13g2_fill_8 FILLER_120_792 ();
 sg13g2_fill_8 FILLER_120_800 ();
 sg13g2_fill_8 FILLER_120_808 ();
 sg13g2_fill_8 FILLER_120_816 ();
 sg13g2_fill_8 FILLER_120_824 ();
 sg13g2_fill_8 FILLER_120_832 ();
 sg13g2_fill_8 FILLER_120_840 ();
 sg13g2_fill_8 FILLER_120_848 ();
 sg13g2_fill_8 FILLER_120_856 ();
 sg13g2_fill_8 FILLER_120_864 ();
 sg13g2_fill_8 FILLER_120_872 ();
 sg13g2_fill_8 FILLER_120_880 ();
 sg13g2_fill_8 FILLER_120_888 ();
 sg13g2_fill_8 FILLER_120_896 ();
 sg13g2_fill_8 FILLER_120_904 ();
 sg13g2_fill_8 FILLER_120_912 ();
 sg13g2_fill_8 FILLER_120_920 ();
 sg13g2_fill_8 FILLER_120_928 ();
 sg13g2_fill_8 FILLER_120_936 ();
 sg13g2_fill_8 FILLER_120_944 ();
 sg13g2_fill_8 FILLER_120_952 ();
 sg13g2_fill_8 FILLER_120_960 ();
 sg13g2_fill_8 FILLER_120_968 ();
 sg13g2_fill_8 FILLER_120_976 ();
 sg13g2_fill_8 FILLER_120_984 ();
 sg13g2_fill_8 FILLER_120_992 ();
 sg13g2_fill_8 FILLER_120_1000 ();
 sg13g2_fill_8 FILLER_120_1008 ();
 sg13g2_fill_8 FILLER_120_1016 ();
 sg13g2_fill_8 FILLER_120_1024 ();
 sg13g2_fill_8 FILLER_120_1032 ();
 sg13g2_fill_8 FILLER_120_1040 ();
 sg13g2_fill_8 FILLER_120_1048 ();
 sg13g2_fill_8 FILLER_120_1056 ();
 sg13g2_fill_8 FILLER_120_1064 ();
 sg13g2_fill_8 FILLER_120_1072 ();
 sg13g2_fill_8 FILLER_120_1080 ();
 sg13g2_fill_8 FILLER_120_1088 ();
 sg13g2_fill_8 FILLER_120_1096 ();
 sg13g2_fill_8 FILLER_120_1104 ();
 sg13g2_fill_8 FILLER_120_1112 ();
 sg13g2_fill_8 FILLER_120_1120 ();
 sg13g2_fill_8 FILLER_120_1128 ();
 sg13g2_fill_8 FILLER_120_1136 ();
 sg13g2_fill_8 FILLER_121_0 ();
 sg13g2_fill_8 FILLER_121_8 ();
 sg13g2_fill_8 FILLER_121_16 ();
 sg13g2_fill_8 FILLER_121_24 ();
 sg13g2_fill_8 FILLER_121_32 ();
 sg13g2_fill_8 FILLER_121_40 ();
 sg13g2_fill_8 FILLER_121_48 ();
 sg13g2_fill_8 FILLER_121_56 ();
 sg13g2_fill_8 FILLER_121_64 ();
 sg13g2_fill_8 FILLER_121_72 ();
 sg13g2_fill_8 FILLER_121_80 ();
 sg13g2_fill_8 FILLER_121_88 ();
 sg13g2_fill_8 FILLER_121_96 ();
 sg13g2_fill_8 FILLER_121_104 ();
 sg13g2_fill_8 FILLER_121_112 ();
 sg13g2_fill_8 FILLER_121_120 ();
 sg13g2_fill_8 FILLER_121_128 ();
 sg13g2_fill_8 FILLER_121_136 ();
 sg13g2_fill_8 FILLER_121_144 ();
 sg13g2_fill_8 FILLER_121_152 ();
 sg13g2_fill_8 FILLER_121_160 ();
 sg13g2_fill_8 FILLER_121_168 ();
 sg13g2_fill_8 FILLER_121_176 ();
 sg13g2_fill_8 FILLER_121_184 ();
 sg13g2_fill_8 FILLER_121_192 ();
 sg13g2_fill_8 FILLER_121_200 ();
 sg13g2_fill_8 FILLER_121_208 ();
 sg13g2_fill_8 FILLER_121_216 ();
 sg13g2_fill_8 FILLER_121_224 ();
 sg13g2_fill_8 FILLER_121_232 ();
 sg13g2_fill_8 FILLER_121_240 ();
 sg13g2_fill_8 FILLER_121_248 ();
 sg13g2_fill_8 FILLER_121_256 ();
 sg13g2_fill_8 FILLER_121_264 ();
 sg13g2_fill_8 FILLER_121_272 ();
 sg13g2_fill_8 FILLER_121_280 ();
 sg13g2_fill_8 FILLER_121_288 ();
 sg13g2_fill_8 FILLER_121_296 ();
 sg13g2_fill_8 FILLER_121_304 ();
 sg13g2_fill_8 FILLER_121_312 ();
 sg13g2_fill_8 FILLER_121_320 ();
 sg13g2_fill_8 FILLER_121_328 ();
 sg13g2_fill_8 FILLER_121_336 ();
 sg13g2_fill_8 FILLER_121_344 ();
 sg13g2_fill_8 FILLER_121_352 ();
 sg13g2_fill_8 FILLER_121_360 ();
 sg13g2_fill_8 FILLER_121_368 ();
 sg13g2_fill_8 FILLER_121_376 ();
 sg13g2_fill_8 FILLER_121_384 ();
 sg13g2_fill_8 FILLER_121_392 ();
 sg13g2_fill_8 FILLER_121_400 ();
 sg13g2_fill_8 FILLER_121_408 ();
 sg13g2_fill_8 FILLER_121_416 ();
 sg13g2_fill_8 FILLER_121_424 ();
 sg13g2_fill_8 FILLER_121_432 ();
 sg13g2_fill_8 FILLER_121_440 ();
 sg13g2_fill_8 FILLER_121_448 ();
 sg13g2_fill_8 FILLER_121_456 ();
 sg13g2_fill_8 FILLER_121_464 ();
 sg13g2_fill_8 FILLER_121_472 ();
 sg13g2_fill_8 FILLER_121_480 ();
 sg13g2_fill_8 FILLER_121_488 ();
 sg13g2_fill_8 FILLER_121_496 ();
 sg13g2_fill_8 FILLER_121_504 ();
 sg13g2_fill_8 FILLER_121_512 ();
 sg13g2_fill_8 FILLER_121_520 ();
 sg13g2_fill_8 FILLER_121_528 ();
 sg13g2_fill_8 FILLER_121_536 ();
 sg13g2_fill_8 FILLER_121_544 ();
 sg13g2_fill_8 FILLER_121_552 ();
 sg13g2_fill_8 FILLER_121_560 ();
 sg13g2_fill_8 FILLER_121_568 ();
 sg13g2_fill_8 FILLER_121_576 ();
 sg13g2_fill_8 FILLER_121_584 ();
 sg13g2_fill_8 FILLER_121_592 ();
 sg13g2_fill_8 FILLER_121_600 ();
 sg13g2_fill_8 FILLER_121_608 ();
 sg13g2_fill_8 FILLER_121_616 ();
 sg13g2_fill_8 FILLER_121_624 ();
 sg13g2_fill_8 FILLER_121_632 ();
 sg13g2_fill_8 FILLER_121_640 ();
 sg13g2_fill_8 FILLER_121_648 ();
 sg13g2_fill_8 FILLER_121_656 ();
 sg13g2_fill_8 FILLER_121_664 ();
 sg13g2_fill_8 FILLER_121_672 ();
 sg13g2_fill_8 FILLER_121_680 ();
 sg13g2_fill_8 FILLER_121_688 ();
 sg13g2_fill_8 FILLER_121_696 ();
 sg13g2_fill_8 FILLER_121_704 ();
 sg13g2_fill_8 FILLER_121_712 ();
 sg13g2_fill_8 FILLER_121_720 ();
 sg13g2_fill_8 FILLER_121_728 ();
 sg13g2_fill_8 FILLER_121_736 ();
 sg13g2_fill_8 FILLER_121_744 ();
 sg13g2_fill_8 FILLER_121_752 ();
 sg13g2_fill_8 FILLER_121_760 ();
 sg13g2_fill_8 FILLER_121_768 ();
 sg13g2_fill_8 FILLER_121_776 ();
 sg13g2_fill_8 FILLER_121_784 ();
 sg13g2_fill_8 FILLER_121_792 ();
 sg13g2_fill_8 FILLER_121_800 ();
 sg13g2_fill_8 FILLER_121_808 ();
 sg13g2_fill_8 FILLER_121_816 ();
 sg13g2_fill_8 FILLER_121_824 ();
 sg13g2_fill_8 FILLER_121_832 ();
 sg13g2_fill_8 FILLER_121_840 ();
 sg13g2_fill_8 FILLER_121_848 ();
 sg13g2_fill_8 FILLER_121_856 ();
 sg13g2_fill_8 FILLER_121_864 ();
 sg13g2_fill_8 FILLER_121_872 ();
 sg13g2_fill_8 FILLER_121_880 ();
 sg13g2_fill_8 FILLER_121_888 ();
 sg13g2_fill_8 FILLER_121_896 ();
 sg13g2_fill_8 FILLER_121_904 ();
 sg13g2_fill_8 FILLER_121_912 ();
 sg13g2_fill_8 FILLER_121_920 ();
 sg13g2_fill_8 FILLER_121_928 ();
 sg13g2_fill_8 FILLER_121_936 ();
 sg13g2_fill_8 FILLER_121_944 ();
 sg13g2_fill_8 FILLER_121_952 ();
 sg13g2_fill_8 FILLER_121_960 ();
 sg13g2_fill_8 FILLER_121_968 ();
 sg13g2_fill_8 FILLER_121_976 ();
 sg13g2_fill_8 FILLER_121_984 ();
 sg13g2_fill_8 FILLER_121_992 ();
 sg13g2_fill_8 FILLER_121_1000 ();
 sg13g2_fill_8 FILLER_121_1008 ();
 sg13g2_fill_8 FILLER_121_1016 ();
 sg13g2_fill_8 FILLER_121_1024 ();
 sg13g2_fill_8 FILLER_121_1032 ();
 sg13g2_fill_8 FILLER_121_1040 ();
 sg13g2_fill_8 FILLER_121_1048 ();
 sg13g2_fill_8 FILLER_121_1056 ();
 sg13g2_fill_8 FILLER_121_1064 ();
 sg13g2_fill_8 FILLER_121_1072 ();
 sg13g2_fill_8 FILLER_121_1080 ();
 sg13g2_fill_8 FILLER_121_1088 ();
 sg13g2_fill_8 FILLER_121_1096 ();
 sg13g2_fill_8 FILLER_121_1104 ();
 sg13g2_fill_8 FILLER_121_1112 ();
 sg13g2_fill_8 FILLER_121_1120 ();
 sg13g2_fill_8 FILLER_121_1128 ();
 sg13g2_fill_8 FILLER_121_1136 ();
 sg13g2_fill_8 FILLER_122_0 ();
 sg13g2_fill_8 FILLER_122_8 ();
 sg13g2_fill_8 FILLER_122_16 ();
 sg13g2_fill_8 FILLER_122_24 ();
 sg13g2_fill_8 FILLER_122_32 ();
 sg13g2_fill_8 FILLER_122_40 ();
 sg13g2_fill_8 FILLER_122_48 ();
 sg13g2_fill_8 FILLER_122_56 ();
 sg13g2_fill_8 FILLER_122_64 ();
 sg13g2_fill_8 FILLER_122_72 ();
 sg13g2_fill_8 FILLER_122_80 ();
 sg13g2_fill_8 FILLER_122_88 ();
 sg13g2_fill_8 FILLER_122_96 ();
 sg13g2_fill_8 FILLER_122_104 ();
 sg13g2_fill_8 FILLER_122_112 ();
 sg13g2_fill_8 FILLER_122_120 ();
 sg13g2_fill_8 FILLER_122_128 ();
 sg13g2_fill_8 FILLER_122_136 ();
 sg13g2_fill_8 FILLER_122_144 ();
 sg13g2_fill_8 FILLER_122_152 ();
 sg13g2_fill_8 FILLER_122_160 ();
 sg13g2_fill_8 FILLER_122_168 ();
 sg13g2_fill_8 FILLER_122_176 ();
 sg13g2_fill_8 FILLER_122_184 ();
 sg13g2_fill_8 FILLER_122_192 ();
 sg13g2_fill_8 FILLER_122_200 ();
 sg13g2_fill_8 FILLER_122_208 ();
 sg13g2_fill_8 FILLER_122_216 ();
 sg13g2_fill_8 FILLER_122_224 ();
 sg13g2_fill_8 FILLER_122_232 ();
 sg13g2_fill_8 FILLER_122_240 ();
 sg13g2_fill_8 FILLER_122_248 ();
 sg13g2_fill_8 FILLER_122_256 ();
 sg13g2_fill_8 FILLER_122_264 ();
 sg13g2_fill_8 FILLER_122_272 ();
 sg13g2_fill_8 FILLER_122_280 ();
 sg13g2_fill_8 FILLER_122_288 ();
 sg13g2_fill_8 FILLER_122_296 ();
 sg13g2_fill_8 FILLER_122_304 ();
 sg13g2_fill_8 FILLER_122_312 ();
 sg13g2_fill_8 FILLER_122_320 ();
 sg13g2_fill_8 FILLER_122_328 ();
 sg13g2_fill_8 FILLER_122_336 ();
 sg13g2_fill_8 FILLER_122_344 ();
 sg13g2_fill_8 FILLER_122_352 ();
 sg13g2_fill_8 FILLER_122_360 ();
 sg13g2_fill_8 FILLER_122_368 ();
 sg13g2_fill_8 FILLER_122_376 ();
 sg13g2_fill_8 FILLER_122_384 ();
 sg13g2_fill_8 FILLER_122_392 ();
 sg13g2_fill_8 FILLER_122_400 ();
 sg13g2_fill_8 FILLER_122_408 ();
 sg13g2_fill_8 FILLER_122_416 ();
 sg13g2_fill_8 FILLER_122_424 ();
 sg13g2_fill_8 FILLER_122_432 ();
 sg13g2_fill_8 FILLER_122_440 ();
 sg13g2_fill_8 FILLER_122_448 ();
 sg13g2_fill_8 FILLER_122_456 ();
 sg13g2_fill_8 FILLER_122_464 ();
 sg13g2_fill_8 FILLER_122_472 ();
 sg13g2_fill_8 FILLER_122_480 ();
 sg13g2_fill_8 FILLER_122_488 ();
 sg13g2_fill_8 FILLER_122_496 ();
 sg13g2_fill_8 FILLER_122_504 ();
 sg13g2_fill_8 FILLER_122_512 ();
 sg13g2_fill_8 FILLER_122_520 ();
 sg13g2_fill_8 FILLER_122_528 ();
 sg13g2_fill_8 FILLER_122_536 ();
 sg13g2_fill_8 FILLER_122_544 ();
 sg13g2_fill_8 FILLER_122_552 ();
 sg13g2_fill_8 FILLER_122_560 ();
 sg13g2_fill_8 FILLER_122_568 ();
 sg13g2_fill_8 FILLER_122_576 ();
 sg13g2_fill_8 FILLER_122_584 ();
 sg13g2_fill_8 FILLER_122_592 ();
 sg13g2_fill_8 FILLER_122_600 ();
 sg13g2_fill_8 FILLER_122_608 ();
 sg13g2_fill_8 FILLER_122_616 ();
 sg13g2_fill_8 FILLER_122_624 ();
 sg13g2_fill_8 FILLER_122_632 ();
 sg13g2_fill_8 FILLER_122_640 ();
 sg13g2_fill_8 FILLER_122_648 ();
 sg13g2_fill_8 FILLER_122_656 ();
 sg13g2_fill_8 FILLER_122_664 ();
 sg13g2_fill_8 FILLER_122_672 ();
 sg13g2_fill_8 FILLER_122_680 ();
 sg13g2_fill_8 FILLER_122_688 ();
 sg13g2_fill_8 FILLER_122_696 ();
 sg13g2_fill_8 FILLER_122_704 ();
 sg13g2_fill_8 FILLER_122_712 ();
 sg13g2_fill_8 FILLER_122_720 ();
 sg13g2_fill_8 FILLER_122_728 ();
 sg13g2_fill_8 FILLER_122_736 ();
 sg13g2_fill_8 FILLER_122_744 ();
 sg13g2_fill_8 FILLER_122_752 ();
 sg13g2_fill_8 FILLER_122_760 ();
 sg13g2_fill_8 FILLER_122_768 ();
 sg13g2_fill_8 FILLER_122_776 ();
 sg13g2_fill_8 FILLER_122_784 ();
 sg13g2_fill_8 FILLER_122_792 ();
 sg13g2_fill_8 FILLER_122_800 ();
 sg13g2_fill_8 FILLER_122_808 ();
 sg13g2_fill_8 FILLER_122_816 ();
 sg13g2_fill_8 FILLER_122_824 ();
 sg13g2_fill_8 FILLER_122_832 ();
 sg13g2_fill_8 FILLER_122_840 ();
 sg13g2_fill_8 FILLER_122_848 ();
 sg13g2_fill_8 FILLER_122_856 ();
 sg13g2_fill_8 FILLER_122_864 ();
 sg13g2_fill_8 FILLER_122_872 ();
 sg13g2_fill_8 FILLER_122_880 ();
 sg13g2_fill_8 FILLER_122_888 ();
 sg13g2_fill_8 FILLER_122_896 ();
 sg13g2_fill_8 FILLER_122_904 ();
 sg13g2_fill_8 FILLER_122_912 ();
 sg13g2_fill_8 FILLER_122_920 ();
 sg13g2_fill_8 FILLER_122_928 ();
 sg13g2_fill_8 FILLER_122_936 ();
 sg13g2_fill_8 FILLER_122_944 ();
 sg13g2_fill_8 FILLER_122_952 ();
 sg13g2_fill_8 FILLER_122_960 ();
 sg13g2_fill_8 FILLER_122_968 ();
 sg13g2_fill_8 FILLER_122_976 ();
 sg13g2_fill_8 FILLER_122_984 ();
 sg13g2_fill_8 FILLER_122_992 ();
 sg13g2_fill_8 FILLER_122_1000 ();
 sg13g2_fill_8 FILLER_122_1008 ();
 sg13g2_fill_8 FILLER_122_1016 ();
 sg13g2_fill_8 FILLER_122_1024 ();
 sg13g2_fill_8 FILLER_122_1032 ();
 sg13g2_fill_8 FILLER_122_1040 ();
 sg13g2_fill_8 FILLER_122_1048 ();
 sg13g2_fill_8 FILLER_122_1056 ();
 sg13g2_fill_8 FILLER_122_1064 ();
 sg13g2_fill_8 FILLER_122_1072 ();
 sg13g2_fill_8 FILLER_122_1080 ();
 sg13g2_fill_8 FILLER_122_1088 ();
 sg13g2_fill_8 FILLER_122_1096 ();
 sg13g2_fill_8 FILLER_122_1104 ();
 sg13g2_fill_8 FILLER_122_1112 ();
 sg13g2_fill_8 FILLER_122_1120 ();
 sg13g2_fill_8 FILLER_122_1128 ();
 sg13g2_fill_8 FILLER_122_1136 ();
 sg13g2_fill_8 FILLER_123_0 ();
 sg13g2_fill_8 FILLER_123_8 ();
 sg13g2_fill_8 FILLER_123_16 ();
 sg13g2_fill_8 FILLER_123_24 ();
 sg13g2_fill_8 FILLER_123_32 ();
 sg13g2_fill_8 FILLER_123_40 ();
 sg13g2_fill_8 FILLER_123_48 ();
 sg13g2_fill_8 FILLER_123_56 ();
 sg13g2_fill_8 FILLER_123_64 ();
 sg13g2_fill_8 FILLER_123_72 ();
 sg13g2_fill_8 FILLER_123_80 ();
 sg13g2_fill_8 FILLER_123_88 ();
 sg13g2_fill_8 FILLER_123_96 ();
 sg13g2_fill_8 FILLER_123_104 ();
 sg13g2_fill_8 FILLER_123_112 ();
 sg13g2_fill_8 FILLER_123_120 ();
 sg13g2_fill_8 FILLER_123_128 ();
 sg13g2_fill_8 FILLER_123_136 ();
 sg13g2_fill_8 FILLER_123_144 ();
 sg13g2_fill_8 FILLER_123_152 ();
 sg13g2_fill_8 FILLER_123_160 ();
 sg13g2_fill_8 FILLER_123_168 ();
 sg13g2_fill_8 FILLER_123_176 ();
 sg13g2_fill_8 FILLER_123_184 ();
 sg13g2_fill_8 FILLER_123_192 ();
 sg13g2_fill_8 FILLER_123_200 ();
 sg13g2_fill_8 FILLER_123_208 ();
 sg13g2_fill_8 FILLER_123_216 ();
 sg13g2_fill_8 FILLER_123_224 ();
 sg13g2_fill_8 FILLER_123_232 ();
 sg13g2_fill_8 FILLER_123_240 ();
 sg13g2_fill_8 FILLER_123_248 ();
 sg13g2_fill_8 FILLER_123_256 ();
 sg13g2_fill_8 FILLER_123_264 ();
 sg13g2_fill_8 FILLER_123_272 ();
 sg13g2_fill_8 FILLER_123_280 ();
 sg13g2_fill_8 FILLER_123_288 ();
 sg13g2_fill_8 FILLER_123_296 ();
 sg13g2_fill_8 FILLER_123_304 ();
 sg13g2_fill_8 FILLER_123_312 ();
 sg13g2_fill_8 FILLER_123_320 ();
 sg13g2_fill_8 FILLER_123_328 ();
 sg13g2_fill_8 FILLER_123_336 ();
 sg13g2_fill_8 FILLER_123_344 ();
 sg13g2_fill_8 FILLER_123_352 ();
 sg13g2_fill_8 FILLER_123_360 ();
 sg13g2_fill_8 FILLER_123_368 ();
 sg13g2_fill_8 FILLER_123_376 ();
 sg13g2_fill_8 FILLER_123_384 ();
 sg13g2_fill_8 FILLER_123_392 ();
 sg13g2_fill_8 FILLER_123_400 ();
 sg13g2_fill_8 FILLER_123_408 ();
 sg13g2_fill_8 FILLER_123_416 ();
 sg13g2_fill_8 FILLER_123_424 ();
 sg13g2_fill_8 FILLER_123_432 ();
 sg13g2_fill_8 FILLER_123_440 ();
 sg13g2_fill_8 FILLER_123_448 ();
 sg13g2_fill_8 FILLER_123_456 ();
 sg13g2_fill_8 FILLER_123_464 ();
 sg13g2_fill_8 FILLER_123_472 ();
 sg13g2_fill_8 FILLER_123_480 ();
 sg13g2_fill_8 FILLER_123_488 ();
 sg13g2_fill_8 FILLER_123_496 ();
 sg13g2_fill_8 FILLER_123_504 ();
 sg13g2_fill_8 FILLER_123_512 ();
 sg13g2_fill_8 FILLER_123_520 ();
 sg13g2_fill_8 FILLER_123_528 ();
 sg13g2_fill_8 FILLER_123_536 ();
 sg13g2_fill_8 FILLER_123_544 ();
 sg13g2_fill_8 FILLER_123_552 ();
 sg13g2_fill_8 FILLER_123_560 ();
 sg13g2_fill_8 FILLER_123_568 ();
 sg13g2_fill_8 FILLER_123_576 ();
 sg13g2_fill_8 FILLER_123_584 ();
 sg13g2_fill_8 FILLER_123_592 ();
 sg13g2_fill_8 FILLER_123_600 ();
 sg13g2_fill_8 FILLER_123_608 ();
 sg13g2_fill_8 FILLER_123_616 ();
 sg13g2_fill_8 FILLER_123_624 ();
 sg13g2_fill_8 FILLER_123_632 ();
 sg13g2_fill_8 FILLER_123_640 ();
 sg13g2_fill_8 FILLER_123_648 ();
 sg13g2_fill_8 FILLER_123_656 ();
 sg13g2_fill_8 FILLER_123_664 ();
 sg13g2_fill_8 FILLER_123_672 ();
 sg13g2_fill_8 FILLER_123_680 ();
 sg13g2_fill_8 FILLER_123_688 ();
 sg13g2_fill_8 FILLER_123_696 ();
 sg13g2_fill_8 FILLER_123_704 ();
 sg13g2_fill_8 FILLER_123_712 ();
 sg13g2_fill_8 FILLER_123_720 ();
 sg13g2_fill_8 FILLER_123_728 ();
 sg13g2_fill_8 FILLER_123_736 ();
 sg13g2_fill_8 FILLER_123_744 ();
 sg13g2_fill_8 FILLER_123_752 ();
 sg13g2_fill_8 FILLER_123_760 ();
 sg13g2_fill_8 FILLER_123_768 ();
 sg13g2_fill_8 FILLER_123_776 ();
 sg13g2_fill_8 FILLER_123_784 ();
 sg13g2_fill_8 FILLER_123_792 ();
 sg13g2_fill_8 FILLER_123_800 ();
 sg13g2_fill_8 FILLER_123_808 ();
 sg13g2_fill_8 FILLER_123_816 ();
 sg13g2_fill_8 FILLER_123_824 ();
 sg13g2_fill_8 FILLER_123_832 ();
 sg13g2_fill_8 FILLER_123_840 ();
 sg13g2_fill_8 FILLER_123_848 ();
 sg13g2_fill_8 FILLER_123_856 ();
 sg13g2_fill_8 FILLER_123_864 ();
 sg13g2_fill_8 FILLER_123_872 ();
 sg13g2_fill_8 FILLER_123_880 ();
 sg13g2_fill_8 FILLER_123_888 ();
 sg13g2_fill_8 FILLER_123_896 ();
 sg13g2_fill_8 FILLER_123_904 ();
 sg13g2_fill_8 FILLER_123_912 ();
 sg13g2_fill_8 FILLER_123_920 ();
 sg13g2_fill_8 FILLER_123_928 ();
 sg13g2_fill_8 FILLER_123_936 ();
 sg13g2_fill_8 FILLER_123_944 ();
 sg13g2_fill_8 FILLER_123_952 ();
 sg13g2_fill_8 FILLER_123_960 ();
 sg13g2_fill_8 FILLER_123_968 ();
 sg13g2_fill_8 FILLER_123_976 ();
 sg13g2_fill_8 FILLER_123_984 ();
 sg13g2_fill_8 FILLER_123_992 ();
 sg13g2_fill_8 FILLER_123_1000 ();
 sg13g2_fill_8 FILLER_123_1008 ();
 sg13g2_fill_8 FILLER_123_1016 ();
 sg13g2_fill_8 FILLER_123_1024 ();
 sg13g2_fill_8 FILLER_123_1032 ();
 sg13g2_fill_8 FILLER_123_1040 ();
 sg13g2_fill_8 FILLER_123_1048 ();
 sg13g2_fill_8 FILLER_123_1056 ();
 sg13g2_fill_8 FILLER_123_1064 ();
 sg13g2_fill_8 FILLER_123_1072 ();
 sg13g2_fill_8 FILLER_123_1080 ();
 sg13g2_fill_8 FILLER_123_1088 ();
 sg13g2_fill_8 FILLER_123_1096 ();
 sg13g2_fill_8 FILLER_123_1104 ();
 sg13g2_fill_8 FILLER_123_1112 ();
 sg13g2_fill_8 FILLER_123_1120 ();
 sg13g2_fill_8 FILLER_123_1128 ();
 sg13g2_fill_8 FILLER_123_1136 ();
 sg13g2_fill_8 FILLER_124_0 ();
 sg13g2_fill_8 FILLER_124_8 ();
 sg13g2_fill_8 FILLER_124_16 ();
 sg13g2_fill_8 FILLER_124_24 ();
 sg13g2_fill_8 FILLER_124_32 ();
 sg13g2_fill_8 FILLER_124_40 ();
 sg13g2_fill_8 FILLER_124_48 ();
 sg13g2_fill_8 FILLER_124_56 ();
 sg13g2_fill_8 FILLER_124_64 ();
 sg13g2_fill_8 FILLER_124_72 ();
 sg13g2_fill_8 FILLER_124_80 ();
 sg13g2_fill_8 FILLER_124_88 ();
 sg13g2_fill_8 FILLER_124_96 ();
 sg13g2_fill_8 FILLER_124_104 ();
 sg13g2_fill_8 FILLER_124_112 ();
 sg13g2_fill_8 FILLER_124_120 ();
 sg13g2_fill_8 FILLER_124_128 ();
 sg13g2_fill_8 FILLER_124_136 ();
 sg13g2_fill_8 FILLER_124_144 ();
 sg13g2_fill_8 FILLER_124_152 ();
 sg13g2_fill_8 FILLER_124_160 ();
 sg13g2_fill_8 FILLER_124_168 ();
 sg13g2_fill_8 FILLER_124_176 ();
 sg13g2_fill_8 FILLER_124_184 ();
 sg13g2_fill_8 FILLER_124_192 ();
 sg13g2_fill_8 FILLER_124_200 ();
 sg13g2_fill_8 FILLER_124_208 ();
 sg13g2_fill_8 FILLER_124_216 ();
 sg13g2_fill_8 FILLER_124_224 ();
 sg13g2_fill_8 FILLER_124_232 ();
 sg13g2_fill_8 FILLER_124_240 ();
 sg13g2_fill_8 FILLER_124_248 ();
 sg13g2_fill_8 FILLER_124_256 ();
 sg13g2_fill_8 FILLER_124_264 ();
 sg13g2_fill_8 FILLER_124_272 ();
 sg13g2_fill_8 FILLER_124_280 ();
 sg13g2_fill_8 FILLER_124_288 ();
 sg13g2_fill_8 FILLER_124_296 ();
 sg13g2_fill_8 FILLER_124_304 ();
 sg13g2_fill_8 FILLER_124_312 ();
 sg13g2_fill_8 FILLER_124_320 ();
 sg13g2_fill_8 FILLER_124_328 ();
 sg13g2_fill_8 FILLER_124_336 ();
 sg13g2_fill_8 FILLER_124_344 ();
 sg13g2_fill_8 FILLER_124_352 ();
 sg13g2_fill_8 FILLER_124_360 ();
 sg13g2_fill_8 FILLER_124_368 ();
 sg13g2_fill_8 FILLER_124_376 ();
 sg13g2_fill_8 FILLER_124_384 ();
 sg13g2_fill_8 FILLER_124_392 ();
 sg13g2_fill_8 FILLER_124_400 ();
 sg13g2_fill_8 FILLER_124_408 ();
 sg13g2_fill_8 FILLER_124_416 ();
 sg13g2_fill_8 FILLER_124_424 ();
 sg13g2_fill_8 FILLER_124_432 ();
 sg13g2_fill_8 FILLER_124_440 ();
 sg13g2_fill_8 FILLER_124_448 ();
 sg13g2_fill_8 FILLER_124_456 ();
 sg13g2_fill_8 FILLER_124_464 ();
 sg13g2_fill_8 FILLER_124_472 ();
 sg13g2_fill_8 FILLER_124_480 ();
 sg13g2_fill_8 FILLER_124_488 ();
 sg13g2_fill_8 FILLER_124_496 ();
 sg13g2_fill_8 FILLER_124_504 ();
 sg13g2_fill_8 FILLER_124_512 ();
 sg13g2_fill_8 FILLER_124_520 ();
 sg13g2_fill_8 FILLER_124_528 ();
 sg13g2_fill_8 FILLER_124_536 ();
 sg13g2_fill_8 FILLER_124_544 ();
 sg13g2_fill_8 FILLER_124_552 ();
 sg13g2_fill_8 FILLER_124_560 ();
 sg13g2_fill_8 FILLER_124_568 ();
 sg13g2_fill_8 FILLER_124_576 ();
 sg13g2_fill_8 FILLER_124_584 ();
 sg13g2_fill_8 FILLER_124_592 ();
 sg13g2_fill_8 FILLER_124_600 ();
 sg13g2_fill_8 FILLER_124_608 ();
 sg13g2_fill_8 FILLER_124_616 ();
 sg13g2_fill_8 FILLER_124_624 ();
 sg13g2_fill_8 FILLER_124_632 ();
 sg13g2_fill_8 FILLER_124_640 ();
 sg13g2_fill_8 FILLER_124_648 ();
 sg13g2_fill_8 FILLER_124_656 ();
 sg13g2_fill_8 FILLER_124_664 ();
 sg13g2_fill_8 FILLER_124_672 ();
 sg13g2_fill_8 FILLER_124_680 ();
 sg13g2_fill_8 FILLER_124_688 ();
 sg13g2_fill_8 FILLER_124_696 ();
 sg13g2_fill_8 FILLER_124_704 ();
 sg13g2_fill_8 FILLER_124_712 ();
 sg13g2_fill_8 FILLER_124_720 ();
 sg13g2_fill_8 FILLER_124_728 ();
 sg13g2_fill_8 FILLER_124_736 ();
 sg13g2_fill_8 FILLER_124_744 ();
 sg13g2_fill_8 FILLER_124_752 ();
 sg13g2_fill_8 FILLER_124_760 ();
 sg13g2_fill_8 FILLER_124_768 ();
 sg13g2_fill_8 FILLER_124_776 ();
 sg13g2_fill_8 FILLER_124_784 ();
 sg13g2_fill_8 FILLER_124_792 ();
 sg13g2_fill_8 FILLER_124_800 ();
 sg13g2_fill_8 FILLER_124_808 ();
 sg13g2_fill_8 FILLER_124_816 ();
 sg13g2_fill_8 FILLER_124_824 ();
 sg13g2_fill_8 FILLER_124_832 ();
 sg13g2_fill_8 FILLER_124_840 ();
 sg13g2_fill_8 FILLER_124_848 ();
 sg13g2_fill_8 FILLER_124_856 ();
 sg13g2_fill_8 FILLER_124_864 ();
 sg13g2_fill_8 FILLER_124_872 ();
 sg13g2_fill_8 FILLER_124_880 ();
 sg13g2_fill_8 FILLER_124_888 ();
 sg13g2_fill_8 FILLER_124_896 ();
 sg13g2_fill_8 FILLER_124_904 ();
 sg13g2_fill_8 FILLER_124_912 ();
 sg13g2_fill_8 FILLER_124_920 ();
 sg13g2_fill_8 FILLER_124_928 ();
 sg13g2_fill_8 FILLER_124_936 ();
 sg13g2_fill_8 FILLER_124_944 ();
 sg13g2_fill_8 FILLER_124_952 ();
 sg13g2_fill_8 FILLER_124_960 ();
 sg13g2_fill_8 FILLER_124_968 ();
 sg13g2_fill_8 FILLER_124_976 ();
 sg13g2_fill_8 FILLER_124_984 ();
 sg13g2_fill_8 FILLER_124_992 ();
 sg13g2_fill_8 FILLER_124_1000 ();
 sg13g2_fill_8 FILLER_124_1008 ();
 sg13g2_fill_8 FILLER_124_1016 ();
 sg13g2_fill_8 FILLER_124_1024 ();
 sg13g2_fill_8 FILLER_124_1032 ();
 sg13g2_fill_8 FILLER_124_1040 ();
 sg13g2_fill_8 FILLER_124_1048 ();
 sg13g2_fill_8 FILLER_124_1056 ();
 sg13g2_fill_8 FILLER_124_1064 ();
 sg13g2_fill_8 FILLER_124_1072 ();
 sg13g2_fill_8 FILLER_124_1080 ();
 sg13g2_fill_8 FILLER_124_1088 ();
 sg13g2_fill_8 FILLER_124_1096 ();
 sg13g2_fill_8 FILLER_124_1104 ();
 sg13g2_fill_8 FILLER_124_1112 ();
 sg13g2_fill_8 FILLER_124_1120 ();
 sg13g2_fill_8 FILLER_124_1128 ();
 sg13g2_fill_8 FILLER_124_1136 ();
 sg13g2_fill_8 FILLER_125_0 ();
 sg13g2_fill_8 FILLER_125_8 ();
 sg13g2_fill_8 FILLER_125_16 ();
 sg13g2_fill_8 FILLER_125_24 ();
 sg13g2_fill_8 FILLER_125_32 ();
 sg13g2_fill_8 FILLER_125_40 ();
 sg13g2_fill_8 FILLER_125_48 ();
 sg13g2_fill_8 FILLER_125_56 ();
 sg13g2_fill_8 FILLER_125_64 ();
 sg13g2_fill_8 FILLER_125_72 ();
 sg13g2_fill_8 FILLER_125_80 ();
 sg13g2_fill_8 FILLER_125_88 ();
 sg13g2_fill_8 FILLER_125_96 ();
 sg13g2_fill_8 FILLER_125_104 ();
 sg13g2_fill_8 FILLER_125_112 ();
 sg13g2_fill_8 FILLER_125_120 ();
 sg13g2_fill_8 FILLER_125_128 ();
 sg13g2_fill_8 FILLER_125_136 ();
 sg13g2_fill_8 FILLER_125_144 ();
 sg13g2_fill_8 FILLER_125_152 ();
 sg13g2_fill_8 FILLER_125_160 ();
 sg13g2_fill_8 FILLER_125_168 ();
 sg13g2_fill_8 FILLER_125_176 ();
 sg13g2_fill_8 FILLER_125_184 ();
 sg13g2_fill_8 FILLER_125_192 ();
 sg13g2_fill_8 FILLER_125_200 ();
 sg13g2_fill_8 FILLER_125_208 ();
 sg13g2_fill_8 FILLER_125_216 ();
 sg13g2_fill_8 FILLER_125_224 ();
 sg13g2_fill_8 FILLER_125_232 ();
 sg13g2_fill_8 FILLER_125_240 ();
 sg13g2_fill_8 FILLER_125_248 ();
 sg13g2_fill_8 FILLER_125_256 ();
 sg13g2_fill_8 FILLER_125_264 ();
 sg13g2_fill_8 FILLER_125_272 ();
 sg13g2_fill_8 FILLER_125_280 ();
 sg13g2_fill_8 FILLER_125_288 ();
 sg13g2_fill_8 FILLER_125_296 ();
 sg13g2_fill_8 FILLER_125_304 ();
 sg13g2_fill_8 FILLER_125_312 ();
 sg13g2_fill_8 FILLER_125_320 ();
 sg13g2_fill_8 FILLER_125_328 ();
 sg13g2_fill_8 FILLER_125_336 ();
 sg13g2_fill_8 FILLER_125_344 ();
 sg13g2_fill_8 FILLER_125_352 ();
 sg13g2_fill_8 FILLER_125_360 ();
 sg13g2_fill_8 FILLER_125_368 ();
 sg13g2_fill_8 FILLER_125_376 ();
 sg13g2_fill_8 FILLER_125_384 ();
 sg13g2_fill_8 FILLER_125_392 ();
 sg13g2_fill_8 FILLER_125_400 ();
 sg13g2_fill_8 FILLER_125_408 ();
 sg13g2_fill_8 FILLER_125_416 ();
 sg13g2_fill_8 FILLER_125_424 ();
 sg13g2_fill_8 FILLER_125_432 ();
 sg13g2_fill_8 FILLER_125_440 ();
 sg13g2_fill_8 FILLER_125_448 ();
 sg13g2_fill_8 FILLER_125_456 ();
 sg13g2_fill_8 FILLER_125_464 ();
 sg13g2_fill_8 FILLER_125_472 ();
 sg13g2_fill_8 FILLER_125_480 ();
 sg13g2_fill_8 FILLER_125_488 ();
 sg13g2_fill_8 FILLER_125_496 ();
 sg13g2_fill_8 FILLER_125_504 ();
 sg13g2_fill_8 FILLER_125_512 ();
 sg13g2_fill_8 FILLER_125_520 ();
 sg13g2_fill_8 FILLER_125_528 ();
 sg13g2_fill_8 FILLER_125_536 ();
 sg13g2_fill_8 FILLER_125_544 ();
 sg13g2_fill_8 FILLER_125_552 ();
 sg13g2_fill_8 FILLER_125_560 ();
 sg13g2_fill_8 FILLER_125_568 ();
 sg13g2_fill_8 FILLER_125_576 ();
 sg13g2_fill_8 FILLER_125_584 ();
 sg13g2_fill_8 FILLER_125_592 ();
 sg13g2_fill_8 FILLER_125_600 ();
 sg13g2_fill_8 FILLER_125_608 ();
 sg13g2_fill_8 FILLER_125_616 ();
 sg13g2_fill_8 FILLER_125_624 ();
 sg13g2_fill_8 FILLER_125_632 ();
 sg13g2_fill_8 FILLER_125_640 ();
 sg13g2_fill_8 FILLER_125_648 ();
 sg13g2_fill_8 FILLER_125_656 ();
 sg13g2_fill_8 FILLER_125_664 ();
 sg13g2_fill_8 FILLER_125_672 ();
 sg13g2_fill_8 FILLER_125_680 ();
 sg13g2_fill_8 FILLER_125_688 ();
 sg13g2_fill_8 FILLER_125_696 ();
 sg13g2_fill_8 FILLER_125_704 ();
 sg13g2_fill_8 FILLER_125_712 ();
 sg13g2_fill_8 FILLER_125_720 ();
 sg13g2_fill_8 FILLER_125_728 ();
 sg13g2_fill_8 FILLER_125_736 ();
 sg13g2_fill_8 FILLER_125_744 ();
 sg13g2_fill_8 FILLER_125_752 ();
 sg13g2_fill_8 FILLER_125_760 ();
 sg13g2_fill_8 FILLER_125_768 ();
 sg13g2_fill_8 FILLER_125_776 ();
 sg13g2_fill_8 FILLER_125_784 ();
 sg13g2_fill_8 FILLER_125_792 ();
 sg13g2_fill_8 FILLER_125_800 ();
 sg13g2_fill_8 FILLER_125_808 ();
 sg13g2_fill_8 FILLER_125_816 ();
 sg13g2_fill_8 FILLER_125_824 ();
 sg13g2_fill_8 FILLER_125_832 ();
 sg13g2_fill_8 FILLER_125_840 ();
 sg13g2_fill_8 FILLER_125_848 ();
 sg13g2_fill_8 FILLER_125_856 ();
 sg13g2_fill_8 FILLER_125_864 ();
 sg13g2_fill_8 FILLER_125_872 ();
 sg13g2_fill_8 FILLER_125_880 ();
 sg13g2_fill_8 FILLER_125_888 ();
 sg13g2_fill_8 FILLER_125_896 ();
 sg13g2_fill_8 FILLER_125_904 ();
 sg13g2_fill_8 FILLER_125_912 ();
 sg13g2_fill_8 FILLER_125_920 ();
 sg13g2_fill_8 FILLER_125_928 ();
 sg13g2_fill_8 FILLER_125_936 ();
 sg13g2_fill_8 FILLER_125_944 ();
 sg13g2_fill_8 FILLER_125_952 ();
 sg13g2_fill_8 FILLER_125_960 ();
 sg13g2_fill_8 FILLER_125_968 ();
 sg13g2_fill_8 FILLER_125_976 ();
 sg13g2_fill_8 FILLER_125_984 ();
 sg13g2_fill_8 FILLER_125_992 ();
 sg13g2_fill_8 FILLER_125_1000 ();
 sg13g2_fill_8 FILLER_125_1008 ();
 sg13g2_fill_8 FILLER_125_1016 ();
 sg13g2_fill_8 FILLER_125_1024 ();
 sg13g2_fill_8 FILLER_125_1032 ();
 sg13g2_fill_8 FILLER_125_1040 ();
 sg13g2_fill_8 FILLER_125_1048 ();
 sg13g2_fill_8 FILLER_125_1056 ();
 sg13g2_fill_8 FILLER_125_1064 ();
 sg13g2_fill_8 FILLER_125_1072 ();
 sg13g2_fill_8 FILLER_125_1080 ();
 sg13g2_fill_8 FILLER_125_1088 ();
 sg13g2_fill_8 FILLER_125_1096 ();
 sg13g2_fill_8 FILLER_125_1104 ();
 sg13g2_fill_8 FILLER_125_1112 ();
 sg13g2_fill_8 FILLER_125_1120 ();
 sg13g2_fill_8 FILLER_125_1128 ();
 sg13g2_fill_8 FILLER_125_1136 ();
 sg13g2_fill_8 FILLER_126_0 ();
 sg13g2_fill_8 FILLER_126_8 ();
 sg13g2_fill_8 FILLER_126_16 ();
 sg13g2_fill_8 FILLER_126_24 ();
 sg13g2_fill_8 FILLER_126_32 ();
 sg13g2_fill_8 FILLER_126_40 ();
 sg13g2_fill_8 FILLER_126_48 ();
 sg13g2_fill_8 FILLER_126_56 ();
 sg13g2_fill_8 FILLER_126_64 ();
 sg13g2_fill_8 FILLER_126_72 ();
 sg13g2_fill_8 FILLER_126_80 ();
 sg13g2_fill_8 FILLER_126_88 ();
 sg13g2_fill_8 FILLER_126_96 ();
 sg13g2_fill_8 FILLER_126_104 ();
 sg13g2_fill_8 FILLER_126_112 ();
 sg13g2_fill_8 FILLER_126_120 ();
 sg13g2_fill_8 FILLER_126_128 ();
 sg13g2_fill_8 FILLER_126_136 ();
 sg13g2_fill_8 FILLER_126_144 ();
 sg13g2_fill_8 FILLER_126_152 ();
 sg13g2_fill_8 FILLER_126_160 ();
 sg13g2_fill_8 FILLER_126_168 ();
 sg13g2_fill_8 FILLER_126_176 ();
 sg13g2_fill_8 FILLER_126_184 ();
 sg13g2_fill_8 FILLER_126_192 ();
 sg13g2_fill_8 FILLER_126_200 ();
 sg13g2_fill_8 FILLER_126_208 ();
 sg13g2_fill_8 FILLER_126_216 ();
 sg13g2_fill_8 FILLER_126_224 ();
 sg13g2_fill_8 FILLER_126_232 ();
 sg13g2_fill_8 FILLER_126_240 ();
 sg13g2_fill_8 FILLER_126_248 ();
 sg13g2_fill_8 FILLER_126_256 ();
 sg13g2_fill_8 FILLER_126_264 ();
 sg13g2_fill_8 FILLER_126_272 ();
 sg13g2_fill_8 FILLER_126_280 ();
 sg13g2_fill_8 FILLER_126_288 ();
 sg13g2_fill_8 FILLER_126_296 ();
 sg13g2_fill_8 FILLER_126_304 ();
 sg13g2_fill_8 FILLER_126_312 ();
 sg13g2_fill_8 FILLER_126_320 ();
 sg13g2_fill_8 FILLER_126_328 ();
 sg13g2_fill_8 FILLER_126_336 ();
 sg13g2_fill_8 FILLER_126_344 ();
 sg13g2_fill_8 FILLER_126_352 ();
 sg13g2_fill_8 FILLER_126_360 ();
 sg13g2_fill_8 FILLER_126_368 ();
 sg13g2_fill_8 FILLER_126_376 ();
 sg13g2_fill_8 FILLER_126_384 ();
 sg13g2_fill_8 FILLER_126_392 ();
 sg13g2_fill_8 FILLER_126_400 ();
 sg13g2_fill_8 FILLER_126_408 ();
 sg13g2_fill_8 FILLER_126_416 ();
 sg13g2_fill_8 FILLER_126_424 ();
 sg13g2_fill_8 FILLER_126_432 ();
 sg13g2_fill_8 FILLER_126_440 ();
 sg13g2_fill_8 FILLER_126_448 ();
 sg13g2_fill_8 FILLER_126_456 ();
 sg13g2_fill_8 FILLER_126_464 ();
 sg13g2_fill_8 FILLER_126_472 ();
 sg13g2_fill_8 FILLER_126_480 ();
 sg13g2_fill_8 FILLER_126_488 ();
 sg13g2_fill_8 FILLER_126_496 ();
 sg13g2_fill_8 FILLER_126_504 ();
 sg13g2_fill_8 FILLER_126_512 ();
 sg13g2_fill_8 FILLER_126_520 ();
 sg13g2_fill_8 FILLER_126_528 ();
 sg13g2_fill_8 FILLER_126_536 ();
 sg13g2_fill_8 FILLER_126_544 ();
 sg13g2_fill_8 FILLER_126_552 ();
 sg13g2_fill_8 FILLER_126_560 ();
 sg13g2_fill_8 FILLER_126_568 ();
 sg13g2_fill_8 FILLER_126_576 ();
 sg13g2_fill_8 FILLER_126_584 ();
 sg13g2_fill_8 FILLER_126_592 ();
 sg13g2_fill_8 FILLER_126_600 ();
 sg13g2_fill_8 FILLER_126_608 ();
 sg13g2_fill_8 FILLER_126_616 ();
 sg13g2_fill_8 FILLER_126_624 ();
 sg13g2_fill_8 FILLER_126_632 ();
 sg13g2_fill_8 FILLER_126_640 ();
 sg13g2_fill_8 FILLER_126_648 ();
 sg13g2_fill_8 FILLER_126_656 ();
 sg13g2_fill_8 FILLER_126_664 ();
 sg13g2_fill_8 FILLER_126_672 ();
 sg13g2_fill_8 FILLER_126_680 ();
 sg13g2_fill_8 FILLER_126_688 ();
 sg13g2_fill_8 FILLER_126_696 ();
 sg13g2_fill_8 FILLER_126_704 ();
 sg13g2_fill_8 FILLER_126_712 ();
 sg13g2_fill_8 FILLER_126_720 ();
 sg13g2_fill_8 FILLER_126_728 ();
 sg13g2_fill_8 FILLER_126_736 ();
 sg13g2_fill_8 FILLER_126_744 ();
 sg13g2_fill_8 FILLER_126_752 ();
 sg13g2_fill_8 FILLER_126_760 ();
 sg13g2_fill_8 FILLER_126_768 ();
 sg13g2_fill_8 FILLER_126_776 ();
 sg13g2_fill_8 FILLER_126_784 ();
 sg13g2_fill_8 FILLER_126_792 ();
 sg13g2_fill_8 FILLER_126_800 ();
 sg13g2_fill_8 FILLER_126_808 ();
 sg13g2_fill_8 FILLER_126_816 ();
 sg13g2_fill_8 FILLER_126_824 ();
 sg13g2_fill_8 FILLER_126_832 ();
 sg13g2_fill_8 FILLER_126_840 ();
 sg13g2_fill_8 FILLER_126_848 ();
 sg13g2_fill_8 FILLER_126_856 ();
 sg13g2_fill_8 FILLER_126_864 ();
 sg13g2_fill_8 FILLER_126_872 ();
 sg13g2_fill_8 FILLER_126_880 ();
 sg13g2_fill_8 FILLER_126_888 ();
 sg13g2_fill_8 FILLER_126_896 ();
 sg13g2_fill_8 FILLER_126_904 ();
 sg13g2_fill_8 FILLER_126_912 ();
 sg13g2_fill_8 FILLER_126_920 ();
 sg13g2_fill_8 FILLER_126_928 ();
 sg13g2_fill_8 FILLER_126_936 ();
 sg13g2_fill_8 FILLER_126_944 ();
 sg13g2_fill_8 FILLER_126_952 ();
 sg13g2_fill_8 FILLER_126_960 ();
 sg13g2_fill_8 FILLER_126_968 ();
 sg13g2_fill_8 FILLER_126_976 ();
 sg13g2_fill_8 FILLER_126_984 ();
 sg13g2_fill_8 FILLER_126_992 ();
 sg13g2_fill_8 FILLER_126_1000 ();
 sg13g2_fill_8 FILLER_126_1008 ();
 sg13g2_fill_8 FILLER_126_1016 ();
 sg13g2_fill_8 FILLER_126_1024 ();
 sg13g2_fill_8 FILLER_126_1032 ();
 sg13g2_fill_8 FILLER_126_1040 ();
 sg13g2_fill_8 FILLER_126_1048 ();
 sg13g2_fill_8 FILLER_126_1056 ();
 sg13g2_fill_8 FILLER_126_1064 ();
 sg13g2_fill_8 FILLER_126_1072 ();
 sg13g2_fill_8 FILLER_126_1080 ();
 sg13g2_fill_8 FILLER_126_1088 ();
 sg13g2_fill_8 FILLER_126_1096 ();
 sg13g2_fill_8 FILLER_126_1104 ();
 sg13g2_fill_8 FILLER_126_1112 ();
 sg13g2_fill_8 FILLER_126_1120 ();
 sg13g2_fill_8 FILLER_126_1128 ();
 sg13g2_fill_8 FILLER_126_1136 ();
 sg13g2_fill_8 FILLER_127_0 ();
 sg13g2_fill_8 FILLER_127_8 ();
 sg13g2_fill_8 FILLER_127_16 ();
 sg13g2_fill_8 FILLER_127_24 ();
 sg13g2_fill_8 FILLER_127_32 ();
 sg13g2_fill_8 FILLER_127_40 ();
 sg13g2_fill_8 FILLER_127_48 ();
 sg13g2_fill_8 FILLER_127_56 ();
 sg13g2_fill_8 FILLER_127_64 ();
 sg13g2_fill_8 FILLER_127_72 ();
 sg13g2_fill_8 FILLER_127_80 ();
 sg13g2_fill_8 FILLER_127_88 ();
 sg13g2_fill_8 FILLER_127_96 ();
 sg13g2_fill_8 FILLER_127_104 ();
 sg13g2_fill_8 FILLER_127_112 ();
 sg13g2_fill_8 FILLER_127_120 ();
 sg13g2_fill_8 FILLER_127_128 ();
 sg13g2_fill_8 FILLER_127_136 ();
 sg13g2_fill_8 FILLER_127_144 ();
 sg13g2_fill_8 FILLER_127_152 ();
 sg13g2_fill_8 FILLER_127_160 ();
 sg13g2_fill_8 FILLER_127_168 ();
 sg13g2_fill_8 FILLER_127_176 ();
 sg13g2_fill_8 FILLER_127_184 ();
 sg13g2_fill_8 FILLER_127_192 ();
 sg13g2_fill_8 FILLER_127_200 ();
 sg13g2_fill_8 FILLER_127_208 ();
 sg13g2_fill_8 FILLER_127_216 ();
 sg13g2_fill_8 FILLER_127_224 ();
 sg13g2_fill_8 FILLER_127_232 ();
 sg13g2_fill_8 FILLER_127_240 ();
 sg13g2_fill_8 FILLER_127_248 ();
 sg13g2_fill_8 FILLER_127_256 ();
 sg13g2_fill_8 FILLER_127_264 ();
 sg13g2_fill_8 FILLER_127_272 ();
 sg13g2_fill_8 FILLER_127_280 ();
 sg13g2_fill_8 FILLER_127_288 ();
 sg13g2_fill_8 FILLER_127_296 ();
 sg13g2_fill_8 FILLER_127_304 ();
 sg13g2_fill_8 FILLER_127_312 ();
 sg13g2_fill_8 FILLER_127_320 ();
 sg13g2_fill_8 FILLER_127_328 ();
 sg13g2_fill_8 FILLER_127_336 ();
 sg13g2_fill_8 FILLER_127_344 ();
 sg13g2_fill_8 FILLER_127_352 ();
 sg13g2_fill_8 FILLER_127_360 ();
 sg13g2_fill_8 FILLER_127_368 ();
 sg13g2_fill_8 FILLER_127_376 ();
 sg13g2_fill_8 FILLER_127_384 ();
 sg13g2_fill_8 FILLER_127_392 ();
 sg13g2_fill_8 FILLER_127_400 ();
 sg13g2_fill_8 FILLER_127_408 ();
 sg13g2_fill_8 FILLER_127_416 ();
 sg13g2_fill_8 FILLER_127_424 ();
 sg13g2_fill_8 FILLER_127_432 ();
 sg13g2_fill_8 FILLER_127_440 ();
 sg13g2_fill_8 FILLER_127_448 ();
 sg13g2_fill_8 FILLER_127_456 ();
 sg13g2_fill_8 FILLER_127_464 ();
 sg13g2_fill_8 FILLER_127_472 ();
 sg13g2_fill_8 FILLER_127_480 ();
 sg13g2_fill_8 FILLER_127_488 ();
 sg13g2_fill_8 FILLER_127_496 ();
 sg13g2_fill_8 FILLER_127_504 ();
 sg13g2_fill_8 FILLER_127_512 ();
 sg13g2_fill_8 FILLER_127_520 ();
 sg13g2_fill_8 FILLER_127_528 ();
 sg13g2_fill_8 FILLER_127_536 ();
 sg13g2_fill_8 FILLER_127_544 ();
 sg13g2_fill_8 FILLER_127_552 ();
 sg13g2_fill_8 FILLER_127_560 ();
 sg13g2_fill_8 FILLER_127_568 ();
 sg13g2_fill_8 FILLER_127_576 ();
 sg13g2_fill_8 FILLER_127_584 ();
 sg13g2_fill_8 FILLER_127_592 ();
 sg13g2_fill_8 FILLER_127_600 ();
 sg13g2_fill_8 FILLER_127_608 ();
 sg13g2_fill_8 FILLER_127_616 ();
 sg13g2_fill_8 FILLER_127_624 ();
 sg13g2_fill_8 FILLER_127_632 ();
 sg13g2_fill_8 FILLER_127_640 ();
 sg13g2_fill_8 FILLER_127_648 ();
 sg13g2_fill_8 FILLER_127_656 ();
 sg13g2_fill_8 FILLER_127_664 ();
 sg13g2_fill_8 FILLER_127_672 ();
 sg13g2_fill_8 FILLER_127_680 ();
 sg13g2_fill_8 FILLER_127_688 ();
 sg13g2_fill_8 FILLER_127_696 ();
 sg13g2_fill_8 FILLER_127_704 ();
 sg13g2_fill_8 FILLER_127_712 ();
 sg13g2_fill_8 FILLER_127_720 ();
 sg13g2_fill_8 FILLER_127_728 ();
 sg13g2_fill_8 FILLER_127_736 ();
 sg13g2_fill_8 FILLER_127_744 ();
 sg13g2_fill_8 FILLER_127_752 ();
 sg13g2_fill_8 FILLER_127_760 ();
 sg13g2_fill_8 FILLER_127_768 ();
 sg13g2_fill_8 FILLER_127_776 ();
 sg13g2_fill_8 FILLER_127_784 ();
 sg13g2_fill_8 FILLER_127_792 ();
 sg13g2_fill_8 FILLER_127_800 ();
 sg13g2_fill_8 FILLER_127_808 ();
 sg13g2_fill_8 FILLER_127_816 ();
 sg13g2_fill_8 FILLER_127_824 ();
 sg13g2_fill_8 FILLER_127_832 ();
 sg13g2_fill_8 FILLER_127_840 ();
 sg13g2_fill_8 FILLER_127_848 ();
 sg13g2_fill_8 FILLER_127_856 ();
 sg13g2_fill_8 FILLER_127_864 ();
 sg13g2_fill_8 FILLER_127_872 ();
 sg13g2_fill_8 FILLER_127_880 ();
 sg13g2_fill_8 FILLER_127_888 ();
 sg13g2_fill_8 FILLER_127_896 ();
 sg13g2_fill_8 FILLER_127_904 ();
 sg13g2_fill_8 FILLER_127_912 ();
 sg13g2_fill_8 FILLER_127_920 ();
 sg13g2_fill_8 FILLER_127_928 ();
 sg13g2_fill_8 FILLER_127_936 ();
 sg13g2_fill_8 FILLER_127_944 ();
 sg13g2_fill_8 FILLER_127_952 ();
 sg13g2_fill_8 FILLER_127_960 ();
 sg13g2_fill_8 FILLER_127_968 ();
 sg13g2_fill_8 FILLER_127_976 ();
 sg13g2_fill_8 FILLER_127_984 ();
 sg13g2_fill_8 FILLER_127_992 ();
 sg13g2_fill_8 FILLER_127_1000 ();
 sg13g2_fill_8 FILLER_127_1008 ();
 sg13g2_fill_8 FILLER_127_1016 ();
 sg13g2_fill_8 FILLER_127_1024 ();
 sg13g2_fill_8 FILLER_127_1032 ();
 sg13g2_fill_8 FILLER_127_1040 ();
 sg13g2_fill_8 FILLER_127_1048 ();
 sg13g2_fill_8 FILLER_127_1056 ();
 sg13g2_fill_8 FILLER_127_1064 ();
 sg13g2_fill_8 FILLER_127_1072 ();
 sg13g2_fill_8 FILLER_127_1080 ();
 sg13g2_fill_8 FILLER_127_1088 ();
 sg13g2_fill_8 FILLER_127_1096 ();
 sg13g2_fill_8 FILLER_127_1104 ();
 sg13g2_fill_8 FILLER_127_1112 ();
 sg13g2_fill_8 FILLER_127_1120 ();
 sg13g2_fill_8 FILLER_127_1128 ();
 sg13g2_fill_8 FILLER_127_1136 ();
 sg13g2_fill_8 FILLER_128_0 ();
 sg13g2_fill_8 FILLER_128_8 ();
 sg13g2_fill_8 FILLER_128_16 ();
 sg13g2_fill_8 FILLER_128_24 ();
 sg13g2_fill_8 FILLER_128_32 ();
 sg13g2_fill_8 FILLER_128_40 ();
 sg13g2_fill_8 FILLER_128_48 ();
 sg13g2_fill_8 FILLER_128_56 ();
 sg13g2_fill_8 FILLER_128_64 ();
 sg13g2_fill_8 FILLER_128_72 ();
 sg13g2_fill_8 FILLER_128_80 ();
 sg13g2_fill_8 FILLER_128_88 ();
 sg13g2_fill_8 FILLER_128_96 ();
 sg13g2_fill_8 FILLER_128_104 ();
 sg13g2_fill_8 FILLER_128_112 ();
 sg13g2_fill_8 FILLER_128_120 ();
 sg13g2_fill_8 FILLER_128_128 ();
 sg13g2_fill_8 FILLER_128_136 ();
 sg13g2_fill_8 FILLER_128_144 ();
 sg13g2_fill_8 FILLER_128_152 ();
 sg13g2_fill_8 FILLER_128_160 ();
 sg13g2_fill_8 FILLER_128_168 ();
 sg13g2_fill_8 FILLER_128_176 ();
 sg13g2_fill_8 FILLER_128_184 ();
 sg13g2_fill_8 FILLER_128_192 ();
 sg13g2_fill_8 FILLER_128_200 ();
 sg13g2_fill_8 FILLER_128_208 ();
 sg13g2_fill_8 FILLER_128_216 ();
 sg13g2_fill_8 FILLER_128_224 ();
 sg13g2_fill_8 FILLER_128_232 ();
 sg13g2_fill_8 FILLER_128_240 ();
 sg13g2_fill_8 FILLER_128_248 ();
 sg13g2_fill_8 FILLER_128_256 ();
 sg13g2_fill_8 FILLER_128_264 ();
 sg13g2_fill_8 FILLER_128_272 ();
 sg13g2_fill_8 FILLER_128_280 ();
 sg13g2_fill_8 FILLER_128_288 ();
 sg13g2_fill_8 FILLER_128_296 ();
 sg13g2_fill_8 FILLER_128_304 ();
 sg13g2_fill_8 FILLER_128_312 ();
 sg13g2_fill_8 FILLER_128_320 ();
 sg13g2_fill_8 FILLER_128_328 ();
 sg13g2_fill_8 FILLER_128_336 ();
 sg13g2_fill_8 FILLER_128_344 ();
 sg13g2_fill_8 FILLER_128_352 ();
 sg13g2_fill_8 FILLER_128_360 ();
 sg13g2_fill_8 FILLER_128_368 ();
 sg13g2_fill_8 FILLER_128_376 ();
 sg13g2_fill_8 FILLER_128_384 ();
 sg13g2_fill_8 FILLER_128_392 ();
 sg13g2_fill_8 FILLER_128_400 ();
 sg13g2_fill_8 FILLER_128_408 ();
 sg13g2_fill_8 FILLER_128_416 ();
 sg13g2_fill_8 FILLER_128_424 ();
 sg13g2_fill_8 FILLER_128_432 ();
 sg13g2_fill_8 FILLER_128_440 ();
 sg13g2_fill_8 FILLER_128_448 ();
 sg13g2_fill_8 FILLER_128_456 ();
 sg13g2_fill_8 FILLER_128_464 ();
 sg13g2_fill_8 FILLER_128_472 ();
 sg13g2_fill_8 FILLER_128_480 ();
 sg13g2_fill_8 FILLER_128_488 ();
 sg13g2_fill_8 FILLER_128_496 ();
 sg13g2_fill_8 FILLER_128_504 ();
 sg13g2_fill_8 FILLER_128_512 ();
 sg13g2_fill_8 FILLER_128_520 ();
 sg13g2_fill_8 FILLER_128_528 ();
 sg13g2_fill_8 FILLER_128_536 ();
 sg13g2_fill_8 FILLER_128_544 ();
 sg13g2_fill_8 FILLER_128_552 ();
 sg13g2_fill_8 FILLER_128_560 ();
 sg13g2_fill_8 FILLER_128_568 ();
 sg13g2_fill_8 FILLER_128_576 ();
 sg13g2_fill_8 FILLER_128_584 ();
 sg13g2_fill_8 FILLER_128_592 ();
 sg13g2_fill_8 FILLER_128_600 ();
 sg13g2_fill_8 FILLER_128_608 ();
 sg13g2_fill_8 FILLER_128_616 ();
 sg13g2_fill_8 FILLER_128_624 ();
 sg13g2_fill_8 FILLER_128_632 ();
 sg13g2_fill_8 FILLER_128_640 ();
 sg13g2_fill_8 FILLER_128_648 ();
 sg13g2_fill_8 FILLER_128_656 ();
 sg13g2_fill_8 FILLER_128_664 ();
 sg13g2_fill_8 FILLER_128_672 ();
 sg13g2_fill_8 FILLER_128_680 ();
 sg13g2_fill_8 FILLER_128_688 ();
 sg13g2_fill_8 FILLER_128_696 ();
 sg13g2_fill_8 FILLER_128_704 ();
 sg13g2_fill_8 FILLER_128_712 ();
 sg13g2_fill_8 FILLER_128_720 ();
 sg13g2_fill_8 FILLER_128_728 ();
 sg13g2_fill_8 FILLER_128_736 ();
 sg13g2_fill_8 FILLER_128_744 ();
 sg13g2_fill_8 FILLER_128_752 ();
 sg13g2_fill_8 FILLER_128_760 ();
 sg13g2_fill_8 FILLER_128_768 ();
 sg13g2_fill_8 FILLER_128_776 ();
 sg13g2_fill_8 FILLER_128_784 ();
 sg13g2_fill_8 FILLER_128_792 ();
 sg13g2_fill_8 FILLER_128_800 ();
 sg13g2_fill_8 FILLER_128_808 ();
 sg13g2_fill_8 FILLER_128_816 ();
 sg13g2_fill_8 FILLER_128_824 ();
 sg13g2_fill_8 FILLER_128_832 ();
 sg13g2_fill_8 FILLER_128_840 ();
 sg13g2_fill_8 FILLER_128_848 ();
 sg13g2_fill_8 FILLER_128_856 ();
 sg13g2_fill_8 FILLER_128_864 ();
 sg13g2_fill_8 FILLER_128_872 ();
 sg13g2_fill_8 FILLER_128_880 ();
 sg13g2_fill_8 FILLER_128_888 ();
 sg13g2_fill_8 FILLER_128_896 ();
 sg13g2_fill_8 FILLER_128_904 ();
 sg13g2_fill_8 FILLER_128_912 ();
 sg13g2_fill_8 FILLER_128_920 ();
 sg13g2_fill_8 FILLER_128_928 ();
 sg13g2_fill_8 FILLER_128_936 ();
 sg13g2_fill_8 FILLER_128_944 ();
 sg13g2_fill_8 FILLER_128_952 ();
 sg13g2_fill_8 FILLER_128_960 ();
 sg13g2_fill_8 FILLER_128_968 ();
 sg13g2_fill_8 FILLER_128_976 ();
 sg13g2_fill_8 FILLER_128_984 ();
 sg13g2_fill_8 FILLER_128_992 ();
 sg13g2_fill_8 FILLER_128_1000 ();
 sg13g2_fill_8 FILLER_128_1008 ();
 sg13g2_fill_8 FILLER_128_1016 ();
 sg13g2_fill_8 FILLER_128_1024 ();
 sg13g2_fill_8 FILLER_128_1032 ();
 sg13g2_fill_8 FILLER_128_1040 ();
 sg13g2_fill_8 FILLER_128_1048 ();
 sg13g2_fill_8 FILLER_128_1056 ();
 sg13g2_fill_8 FILLER_128_1064 ();
 sg13g2_fill_8 FILLER_128_1072 ();
 sg13g2_fill_8 FILLER_128_1080 ();
 sg13g2_fill_8 FILLER_128_1088 ();
 sg13g2_fill_8 FILLER_128_1096 ();
 sg13g2_fill_8 FILLER_128_1104 ();
 sg13g2_fill_8 FILLER_128_1112 ();
 sg13g2_fill_8 FILLER_128_1120 ();
 sg13g2_fill_8 FILLER_128_1128 ();
 sg13g2_fill_8 FILLER_128_1136 ();
 sg13g2_fill_8 FILLER_129_0 ();
 sg13g2_fill_8 FILLER_129_8 ();
 sg13g2_fill_8 FILLER_129_16 ();
 sg13g2_fill_8 FILLER_129_24 ();
 sg13g2_fill_8 FILLER_129_32 ();
 sg13g2_fill_8 FILLER_129_40 ();
 sg13g2_fill_8 FILLER_129_48 ();
 sg13g2_fill_8 FILLER_129_56 ();
 sg13g2_fill_8 FILLER_129_64 ();
 sg13g2_fill_8 FILLER_129_72 ();
 sg13g2_fill_8 FILLER_129_80 ();
 sg13g2_fill_8 FILLER_129_88 ();
 sg13g2_fill_8 FILLER_129_96 ();
 sg13g2_fill_8 FILLER_129_104 ();
 sg13g2_fill_8 FILLER_129_112 ();
 sg13g2_fill_8 FILLER_129_120 ();
 sg13g2_fill_8 FILLER_129_128 ();
 sg13g2_fill_8 FILLER_129_136 ();
 sg13g2_fill_8 FILLER_129_144 ();
 sg13g2_fill_8 FILLER_129_152 ();
 sg13g2_fill_8 FILLER_129_160 ();
 sg13g2_fill_8 FILLER_129_168 ();
 sg13g2_fill_8 FILLER_129_176 ();
 sg13g2_fill_8 FILLER_129_184 ();
 sg13g2_fill_8 FILLER_129_192 ();
 sg13g2_fill_8 FILLER_129_200 ();
 sg13g2_fill_8 FILLER_129_208 ();
 sg13g2_fill_8 FILLER_129_216 ();
 sg13g2_fill_8 FILLER_129_224 ();
 sg13g2_fill_8 FILLER_129_232 ();
 sg13g2_fill_8 FILLER_129_240 ();
 sg13g2_fill_8 FILLER_129_248 ();
 sg13g2_fill_8 FILLER_129_256 ();
 sg13g2_fill_8 FILLER_129_264 ();
 sg13g2_fill_8 FILLER_129_272 ();
 sg13g2_fill_8 FILLER_129_280 ();
 sg13g2_fill_8 FILLER_129_288 ();
 sg13g2_fill_8 FILLER_129_296 ();
 sg13g2_fill_8 FILLER_129_304 ();
 sg13g2_fill_8 FILLER_129_312 ();
 sg13g2_fill_8 FILLER_129_320 ();
 sg13g2_fill_8 FILLER_129_328 ();
 sg13g2_fill_8 FILLER_129_336 ();
 sg13g2_fill_8 FILLER_129_344 ();
 sg13g2_fill_8 FILLER_129_352 ();
 sg13g2_fill_8 FILLER_129_360 ();
 sg13g2_fill_8 FILLER_129_368 ();
 sg13g2_fill_8 FILLER_129_376 ();
 sg13g2_fill_8 FILLER_129_384 ();
 sg13g2_fill_8 FILLER_129_392 ();
 sg13g2_fill_8 FILLER_129_400 ();
 sg13g2_fill_8 FILLER_129_408 ();
 sg13g2_fill_8 FILLER_129_416 ();
 sg13g2_fill_8 FILLER_129_424 ();
 sg13g2_fill_8 FILLER_129_432 ();
 sg13g2_fill_8 FILLER_129_440 ();
 sg13g2_fill_8 FILLER_129_448 ();
 sg13g2_fill_8 FILLER_129_456 ();
 sg13g2_fill_8 FILLER_129_464 ();
 sg13g2_fill_8 FILLER_129_472 ();
 sg13g2_fill_8 FILLER_129_480 ();
 sg13g2_fill_8 FILLER_129_488 ();
 sg13g2_fill_8 FILLER_129_496 ();
 sg13g2_fill_8 FILLER_129_504 ();
 sg13g2_fill_8 FILLER_129_512 ();
 sg13g2_fill_8 FILLER_129_520 ();
 sg13g2_fill_8 FILLER_129_528 ();
 sg13g2_fill_8 FILLER_129_536 ();
 sg13g2_fill_8 FILLER_129_544 ();
 sg13g2_fill_8 FILLER_129_552 ();
 sg13g2_fill_8 FILLER_129_560 ();
 sg13g2_fill_8 FILLER_129_568 ();
 sg13g2_fill_8 FILLER_129_576 ();
 sg13g2_fill_8 FILLER_129_584 ();
 sg13g2_fill_8 FILLER_129_592 ();
 sg13g2_fill_8 FILLER_129_600 ();
 sg13g2_fill_8 FILLER_129_608 ();
 sg13g2_fill_8 FILLER_129_616 ();
 sg13g2_fill_8 FILLER_129_624 ();
 sg13g2_fill_8 FILLER_129_632 ();
 sg13g2_fill_8 FILLER_129_640 ();
 sg13g2_fill_8 FILLER_129_648 ();
 sg13g2_fill_8 FILLER_129_656 ();
 sg13g2_fill_8 FILLER_129_664 ();
 sg13g2_fill_8 FILLER_129_672 ();
 sg13g2_fill_8 FILLER_129_680 ();
 sg13g2_fill_8 FILLER_129_688 ();
 sg13g2_fill_8 FILLER_129_696 ();
 sg13g2_fill_8 FILLER_129_704 ();
 sg13g2_fill_8 FILLER_129_712 ();
 sg13g2_fill_8 FILLER_129_720 ();
 sg13g2_fill_8 FILLER_129_728 ();
 sg13g2_fill_8 FILLER_129_736 ();
 sg13g2_fill_8 FILLER_129_744 ();
 sg13g2_fill_8 FILLER_129_752 ();
 sg13g2_fill_8 FILLER_129_760 ();
 sg13g2_fill_8 FILLER_129_768 ();
 sg13g2_fill_8 FILLER_129_776 ();
 sg13g2_fill_8 FILLER_129_784 ();
 sg13g2_fill_8 FILLER_129_792 ();
 sg13g2_fill_8 FILLER_129_800 ();
 sg13g2_fill_8 FILLER_129_808 ();
 sg13g2_fill_8 FILLER_129_816 ();
 sg13g2_fill_8 FILLER_129_824 ();
 sg13g2_fill_8 FILLER_129_832 ();
 sg13g2_fill_8 FILLER_129_840 ();
 sg13g2_fill_8 FILLER_129_848 ();
 sg13g2_fill_8 FILLER_129_856 ();
 sg13g2_fill_8 FILLER_129_864 ();
 sg13g2_fill_8 FILLER_129_872 ();
 sg13g2_fill_8 FILLER_129_880 ();
 sg13g2_fill_8 FILLER_129_888 ();
 sg13g2_fill_8 FILLER_129_896 ();
 sg13g2_fill_8 FILLER_129_904 ();
 sg13g2_fill_8 FILLER_129_912 ();
 sg13g2_fill_8 FILLER_129_920 ();
 sg13g2_fill_8 FILLER_129_928 ();
 sg13g2_fill_8 FILLER_129_936 ();
 sg13g2_fill_8 FILLER_129_944 ();
 sg13g2_fill_8 FILLER_129_952 ();
 sg13g2_fill_8 FILLER_129_960 ();
 sg13g2_fill_8 FILLER_129_968 ();
 sg13g2_fill_8 FILLER_129_976 ();
 sg13g2_fill_8 FILLER_129_984 ();
 sg13g2_fill_8 FILLER_129_992 ();
 sg13g2_fill_8 FILLER_129_1000 ();
 sg13g2_fill_8 FILLER_129_1008 ();
 sg13g2_fill_8 FILLER_129_1016 ();
 sg13g2_fill_8 FILLER_129_1024 ();
 sg13g2_fill_8 FILLER_129_1032 ();
 sg13g2_fill_8 FILLER_129_1040 ();
 sg13g2_fill_8 FILLER_129_1048 ();
 sg13g2_fill_8 FILLER_129_1056 ();
 sg13g2_fill_8 FILLER_129_1064 ();
 sg13g2_fill_8 FILLER_129_1072 ();
 sg13g2_fill_8 FILLER_129_1080 ();
 sg13g2_fill_8 FILLER_129_1088 ();
 sg13g2_fill_8 FILLER_129_1096 ();
 sg13g2_fill_8 FILLER_129_1104 ();
 sg13g2_fill_8 FILLER_129_1112 ();
 sg13g2_fill_8 FILLER_129_1120 ();
 sg13g2_fill_8 FILLER_129_1128 ();
 sg13g2_fill_8 FILLER_129_1136 ();
 sg13g2_fill_8 FILLER_130_0 ();
 sg13g2_fill_8 FILLER_130_8 ();
 sg13g2_fill_8 FILLER_130_16 ();
 sg13g2_fill_8 FILLER_130_24 ();
 sg13g2_fill_8 FILLER_130_32 ();
 sg13g2_fill_8 FILLER_130_40 ();
 sg13g2_fill_8 FILLER_130_48 ();
 sg13g2_fill_8 FILLER_130_56 ();
 sg13g2_fill_8 FILLER_130_64 ();
 sg13g2_fill_8 FILLER_130_72 ();
 sg13g2_fill_8 FILLER_130_80 ();
 sg13g2_fill_8 FILLER_130_88 ();
 sg13g2_fill_8 FILLER_130_96 ();
 sg13g2_fill_8 FILLER_130_104 ();
 sg13g2_fill_8 FILLER_130_112 ();
 sg13g2_fill_8 FILLER_130_120 ();
 sg13g2_fill_8 FILLER_130_128 ();
 sg13g2_fill_8 FILLER_130_136 ();
 sg13g2_fill_8 FILLER_130_144 ();
 sg13g2_fill_8 FILLER_130_152 ();
 sg13g2_fill_8 FILLER_130_160 ();
 sg13g2_fill_8 FILLER_130_168 ();
 sg13g2_fill_8 FILLER_130_176 ();
 sg13g2_fill_8 FILLER_130_184 ();
 sg13g2_fill_8 FILLER_130_192 ();
 sg13g2_fill_8 FILLER_130_200 ();
 sg13g2_fill_8 FILLER_130_208 ();
 sg13g2_fill_8 FILLER_130_216 ();
 sg13g2_fill_8 FILLER_130_224 ();
 sg13g2_fill_8 FILLER_130_232 ();
 sg13g2_fill_8 FILLER_130_240 ();
 sg13g2_fill_8 FILLER_130_248 ();
 sg13g2_fill_8 FILLER_130_256 ();
 sg13g2_fill_8 FILLER_130_264 ();
 sg13g2_fill_8 FILLER_130_272 ();
 sg13g2_fill_8 FILLER_130_280 ();
 sg13g2_fill_8 FILLER_130_288 ();
 sg13g2_fill_8 FILLER_130_296 ();
 sg13g2_fill_8 FILLER_130_304 ();
 sg13g2_fill_8 FILLER_130_312 ();
 sg13g2_fill_8 FILLER_130_320 ();
 sg13g2_fill_8 FILLER_130_328 ();
 sg13g2_fill_8 FILLER_130_336 ();
 sg13g2_fill_8 FILLER_130_344 ();
 sg13g2_fill_8 FILLER_130_352 ();
 sg13g2_fill_8 FILLER_130_360 ();
 sg13g2_fill_8 FILLER_130_368 ();
 sg13g2_fill_8 FILLER_130_376 ();
 sg13g2_fill_8 FILLER_130_384 ();
 sg13g2_fill_8 FILLER_130_392 ();
 sg13g2_fill_8 FILLER_130_400 ();
 sg13g2_fill_8 FILLER_130_408 ();
 sg13g2_fill_8 FILLER_130_416 ();
 sg13g2_fill_8 FILLER_130_424 ();
 sg13g2_fill_8 FILLER_130_432 ();
 sg13g2_fill_8 FILLER_130_440 ();
 sg13g2_fill_8 FILLER_130_448 ();
 sg13g2_fill_8 FILLER_130_456 ();
 sg13g2_fill_8 FILLER_130_464 ();
 sg13g2_fill_8 FILLER_130_472 ();
 sg13g2_fill_8 FILLER_130_480 ();
 sg13g2_fill_8 FILLER_130_488 ();
 sg13g2_fill_8 FILLER_130_496 ();
 sg13g2_fill_8 FILLER_130_504 ();
 sg13g2_fill_8 FILLER_130_512 ();
 sg13g2_fill_8 FILLER_130_520 ();
 sg13g2_fill_8 FILLER_130_528 ();
 sg13g2_fill_8 FILLER_130_536 ();
 sg13g2_fill_8 FILLER_130_544 ();
 sg13g2_fill_8 FILLER_130_552 ();
 sg13g2_fill_8 FILLER_130_560 ();
 sg13g2_fill_8 FILLER_130_568 ();
 sg13g2_fill_8 FILLER_130_576 ();
 sg13g2_fill_8 FILLER_130_584 ();
 sg13g2_fill_8 FILLER_130_592 ();
 sg13g2_fill_8 FILLER_130_600 ();
 sg13g2_fill_8 FILLER_130_608 ();
 sg13g2_fill_8 FILLER_130_616 ();
 sg13g2_fill_8 FILLER_130_624 ();
 sg13g2_fill_8 FILLER_130_632 ();
 sg13g2_fill_8 FILLER_130_640 ();
 sg13g2_fill_8 FILLER_130_648 ();
 sg13g2_fill_8 FILLER_130_656 ();
 sg13g2_fill_8 FILLER_130_664 ();
 sg13g2_fill_8 FILLER_130_672 ();
 sg13g2_fill_8 FILLER_130_680 ();
 sg13g2_fill_8 FILLER_130_688 ();
 sg13g2_fill_8 FILLER_130_696 ();
 sg13g2_fill_8 FILLER_130_704 ();
 sg13g2_fill_8 FILLER_130_712 ();
 sg13g2_fill_8 FILLER_130_720 ();
 sg13g2_fill_8 FILLER_130_728 ();
 sg13g2_fill_8 FILLER_130_736 ();
 sg13g2_fill_8 FILLER_130_744 ();
 sg13g2_fill_8 FILLER_130_752 ();
 sg13g2_fill_8 FILLER_130_760 ();
 sg13g2_fill_8 FILLER_130_768 ();
 sg13g2_fill_8 FILLER_130_776 ();
 sg13g2_fill_8 FILLER_130_784 ();
 sg13g2_fill_8 FILLER_130_792 ();
 sg13g2_fill_8 FILLER_130_800 ();
 sg13g2_fill_8 FILLER_130_808 ();
 sg13g2_fill_8 FILLER_130_816 ();
 sg13g2_fill_8 FILLER_130_824 ();
 sg13g2_fill_8 FILLER_130_832 ();
 sg13g2_fill_8 FILLER_130_840 ();
 sg13g2_fill_8 FILLER_130_848 ();
 sg13g2_fill_8 FILLER_130_856 ();
 sg13g2_fill_8 FILLER_130_864 ();
 sg13g2_fill_8 FILLER_130_872 ();
 sg13g2_fill_8 FILLER_130_880 ();
 sg13g2_fill_8 FILLER_130_888 ();
 sg13g2_fill_8 FILLER_130_896 ();
 sg13g2_fill_8 FILLER_130_904 ();
 sg13g2_fill_8 FILLER_130_912 ();
 sg13g2_fill_8 FILLER_130_920 ();
 sg13g2_fill_8 FILLER_130_928 ();
 sg13g2_fill_8 FILLER_130_936 ();
 sg13g2_fill_8 FILLER_130_944 ();
 sg13g2_fill_8 FILLER_130_952 ();
 sg13g2_fill_8 FILLER_130_960 ();
 sg13g2_fill_8 FILLER_130_968 ();
 sg13g2_fill_8 FILLER_130_976 ();
 sg13g2_fill_8 FILLER_130_984 ();
 sg13g2_fill_8 FILLER_130_992 ();
 sg13g2_fill_8 FILLER_130_1000 ();
 sg13g2_fill_8 FILLER_130_1008 ();
 sg13g2_fill_8 FILLER_130_1016 ();
 sg13g2_fill_8 FILLER_130_1024 ();
 sg13g2_fill_8 FILLER_130_1032 ();
 sg13g2_fill_8 FILLER_130_1040 ();
 sg13g2_fill_8 FILLER_130_1048 ();
 sg13g2_fill_8 FILLER_130_1056 ();
 sg13g2_fill_8 FILLER_130_1064 ();
 sg13g2_fill_8 FILLER_130_1072 ();
 sg13g2_fill_8 FILLER_130_1080 ();
 sg13g2_fill_8 FILLER_130_1088 ();
 sg13g2_fill_8 FILLER_130_1096 ();
 sg13g2_fill_8 FILLER_130_1104 ();
 sg13g2_fill_8 FILLER_130_1112 ();
 sg13g2_fill_8 FILLER_130_1120 ();
 sg13g2_fill_8 FILLER_130_1128 ();
 sg13g2_fill_8 FILLER_130_1136 ();
 sg13g2_fill_8 FILLER_131_0 ();
 sg13g2_fill_8 FILLER_131_8 ();
 sg13g2_fill_8 FILLER_131_16 ();
 sg13g2_fill_8 FILLER_131_24 ();
 sg13g2_fill_8 FILLER_131_32 ();
 sg13g2_fill_8 FILLER_131_40 ();
 sg13g2_fill_8 FILLER_131_48 ();
 sg13g2_fill_8 FILLER_131_56 ();
 sg13g2_fill_8 FILLER_131_64 ();
 sg13g2_fill_8 FILLER_131_72 ();
 sg13g2_fill_8 FILLER_131_80 ();
 sg13g2_fill_8 FILLER_131_88 ();
 sg13g2_fill_8 FILLER_131_96 ();
 sg13g2_fill_8 FILLER_131_104 ();
 sg13g2_fill_8 FILLER_131_112 ();
 sg13g2_fill_8 FILLER_131_120 ();
 sg13g2_fill_8 FILLER_131_128 ();
 sg13g2_fill_8 FILLER_131_136 ();
 sg13g2_fill_8 FILLER_131_144 ();
 sg13g2_fill_8 FILLER_131_152 ();
 sg13g2_fill_8 FILLER_131_160 ();
 sg13g2_fill_8 FILLER_131_168 ();
 sg13g2_fill_8 FILLER_131_176 ();
 sg13g2_fill_8 FILLER_131_184 ();
 sg13g2_fill_8 FILLER_131_192 ();
 sg13g2_fill_8 FILLER_131_200 ();
 sg13g2_fill_8 FILLER_131_208 ();
 sg13g2_fill_8 FILLER_131_216 ();
 sg13g2_fill_8 FILLER_131_224 ();
 sg13g2_fill_8 FILLER_131_232 ();
 sg13g2_fill_8 FILLER_131_240 ();
 sg13g2_fill_8 FILLER_131_248 ();
 sg13g2_fill_8 FILLER_131_256 ();
 sg13g2_fill_8 FILLER_131_264 ();
 sg13g2_fill_8 FILLER_131_272 ();
 sg13g2_fill_8 FILLER_131_280 ();
 sg13g2_fill_8 FILLER_131_288 ();
 sg13g2_fill_8 FILLER_131_296 ();
 sg13g2_fill_8 FILLER_131_304 ();
 sg13g2_fill_8 FILLER_131_312 ();
 sg13g2_fill_8 FILLER_131_320 ();
 sg13g2_fill_8 FILLER_131_328 ();
 sg13g2_fill_8 FILLER_131_336 ();
 sg13g2_fill_8 FILLER_131_344 ();
 sg13g2_fill_8 FILLER_131_352 ();
 sg13g2_fill_8 FILLER_131_360 ();
 sg13g2_fill_8 FILLER_131_368 ();
 sg13g2_fill_8 FILLER_131_376 ();
 sg13g2_fill_8 FILLER_131_384 ();
 sg13g2_fill_8 FILLER_131_392 ();
 sg13g2_fill_8 FILLER_131_400 ();
 sg13g2_fill_8 FILLER_131_408 ();
 sg13g2_fill_8 FILLER_131_416 ();
 sg13g2_fill_8 FILLER_131_424 ();
 sg13g2_fill_8 FILLER_131_432 ();
 sg13g2_fill_8 FILLER_131_440 ();
 sg13g2_fill_8 FILLER_131_448 ();
 sg13g2_fill_8 FILLER_131_456 ();
 sg13g2_fill_8 FILLER_131_464 ();
 sg13g2_fill_8 FILLER_131_472 ();
 sg13g2_fill_8 FILLER_131_480 ();
 sg13g2_fill_8 FILLER_131_488 ();
 sg13g2_fill_8 FILLER_131_496 ();
 sg13g2_fill_8 FILLER_131_504 ();
 sg13g2_fill_8 FILLER_131_512 ();
 sg13g2_fill_8 FILLER_131_520 ();
 sg13g2_fill_8 FILLER_131_528 ();
 sg13g2_fill_8 FILLER_131_536 ();
 sg13g2_fill_8 FILLER_131_544 ();
 sg13g2_fill_8 FILLER_131_552 ();
 sg13g2_fill_8 FILLER_131_560 ();
 sg13g2_fill_8 FILLER_131_568 ();
 sg13g2_fill_8 FILLER_131_576 ();
 sg13g2_fill_8 FILLER_131_584 ();
 sg13g2_fill_8 FILLER_131_592 ();
 sg13g2_fill_8 FILLER_131_600 ();
 sg13g2_fill_8 FILLER_131_608 ();
 sg13g2_fill_8 FILLER_131_616 ();
 sg13g2_fill_8 FILLER_131_624 ();
 sg13g2_fill_8 FILLER_131_632 ();
 sg13g2_fill_8 FILLER_131_640 ();
 sg13g2_fill_8 FILLER_131_648 ();
 sg13g2_fill_8 FILLER_131_656 ();
 sg13g2_fill_8 FILLER_131_664 ();
 sg13g2_fill_8 FILLER_131_672 ();
 sg13g2_fill_8 FILLER_131_680 ();
 sg13g2_fill_8 FILLER_131_688 ();
 sg13g2_fill_8 FILLER_131_696 ();
 sg13g2_fill_8 FILLER_131_704 ();
 sg13g2_fill_8 FILLER_131_712 ();
 sg13g2_fill_8 FILLER_131_720 ();
 sg13g2_fill_8 FILLER_131_728 ();
 sg13g2_fill_8 FILLER_131_736 ();
 sg13g2_fill_8 FILLER_131_744 ();
 sg13g2_fill_8 FILLER_131_752 ();
 sg13g2_fill_8 FILLER_131_760 ();
 sg13g2_fill_8 FILLER_131_768 ();
 sg13g2_fill_8 FILLER_131_776 ();
 sg13g2_fill_8 FILLER_131_784 ();
 sg13g2_fill_8 FILLER_131_792 ();
 sg13g2_fill_8 FILLER_131_800 ();
 sg13g2_fill_8 FILLER_131_808 ();
 sg13g2_fill_8 FILLER_131_816 ();
 sg13g2_fill_8 FILLER_131_824 ();
 sg13g2_fill_8 FILLER_131_832 ();
 sg13g2_fill_8 FILLER_131_840 ();
 sg13g2_fill_8 FILLER_131_848 ();
 sg13g2_fill_8 FILLER_131_856 ();
 sg13g2_fill_8 FILLER_131_864 ();
 sg13g2_fill_8 FILLER_131_872 ();
 sg13g2_fill_8 FILLER_131_880 ();
 sg13g2_fill_8 FILLER_131_888 ();
 sg13g2_fill_8 FILLER_131_896 ();
 sg13g2_fill_8 FILLER_131_904 ();
 sg13g2_fill_8 FILLER_131_912 ();
 sg13g2_fill_8 FILLER_131_920 ();
 sg13g2_fill_8 FILLER_131_928 ();
 sg13g2_fill_8 FILLER_131_936 ();
 sg13g2_fill_8 FILLER_131_944 ();
 sg13g2_fill_8 FILLER_131_952 ();
 sg13g2_fill_8 FILLER_131_960 ();
 sg13g2_fill_8 FILLER_131_968 ();
 sg13g2_fill_8 FILLER_131_976 ();
 sg13g2_fill_8 FILLER_131_984 ();
 sg13g2_fill_8 FILLER_131_992 ();
 sg13g2_fill_8 FILLER_131_1000 ();
 sg13g2_fill_8 FILLER_131_1008 ();
 sg13g2_fill_8 FILLER_131_1016 ();
 sg13g2_fill_8 FILLER_131_1024 ();
 sg13g2_fill_8 FILLER_131_1032 ();
 sg13g2_fill_8 FILLER_131_1040 ();
 sg13g2_fill_8 FILLER_131_1048 ();
 sg13g2_fill_8 FILLER_131_1056 ();
 sg13g2_fill_8 FILLER_131_1064 ();
 sg13g2_fill_8 FILLER_131_1072 ();
 sg13g2_fill_8 FILLER_131_1080 ();
 sg13g2_fill_8 FILLER_131_1088 ();
 sg13g2_fill_8 FILLER_131_1096 ();
 sg13g2_fill_8 FILLER_131_1104 ();
 sg13g2_fill_8 FILLER_131_1112 ();
 sg13g2_fill_8 FILLER_131_1120 ();
 sg13g2_fill_8 FILLER_131_1128 ();
 sg13g2_fill_8 FILLER_131_1136 ();
 sg13g2_fill_8 FILLER_132_0 ();
 sg13g2_fill_8 FILLER_132_8 ();
 sg13g2_fill_8 FILLER_132_16 ();
 sg13g2_fill_8 FILLER_132_24 ();
 sg13g2_fill_8 FILLER_132_32 ();
 sg13g2_fill_8 FILLER_132_40 ();
 sg13g2_fill_8 FILLER_132_48 ();
 sg13g2_fill_8 FILLER_132_56 ();
 sg13g2_fill_8 FILLER_132_64 ();
 sg13g2_fill_8 FILLER_132_72 ();
 sg13g2_fill_8 FILLER_132_80 ();
 sg13g2_fill_8 FILLER_132_88 ();
 sg13g2_fill_8 FILLER_132_96 ();
 sg13g2_fill_8 FILLER_132_104 ();
 sg13g2_fill_8 FILLER_132_112 ();
 sg13g2_fill_8 FILLER_132_120 ();
 sg13g2_fill_8 FILLER_132_128 ();
 sg13g2_fill_8 FILLER_132_136 ();
 sg13g2_fill_8 FILLER_132_144 ();
 sg13g2_fill_8 FILLER_132_152 ();
 sg13g2_fill_8 FILLER_132_160 ();
 sg13g2_fill_8 FILLER_132_168 ();
 sg13g2_fill_8 FILLER_132_176 ();
 sg13g2_fill_8 FILLER_132_184 ();
 sg13g2_fill_8 FILLER_132_192 ();
 sg13g2_fill_8 FILLER_132_200 ();
 sg13g2_fill_8 FILLER_132_208 ();
 sg13g2_fill_8 FILLER_132_216 ();
 sg13g2_fill_8 FILLER_132_224 ();
 sg13g2_fill_8 FILLER_132_232 ();
 sg13g2_fill_8 FILLER_132_240 ();
 sg13g2_fill_8 FILLER_132_248 ();
 sg13g2_fill_8 FILLER_132_256 ();
 sg13g2_fill_8 FILLER_132_264 ();
 sg13g2_fill_8 FILLER_132_272 ();
 sg13g2_fill_8 FILLER_132_280 ();
 sg13g2_fill_8 FILLER_132_288 ();
 sg13g2_fill_8 FILLER_132_296 ();
 sg13g2_fill_8 FILLER_132_304 ();
 sg13g2_fill_8 FILLER_132_312 ();
 sg13g2_fill_8 FILLER_132_320 ();
 sg13g2_fill_8 FILLER_132_328 ();
 sg13g2_fill_8 FILLER_132_336 ();
 sg13g2_fill_8 FILLER_132_344 ();
 sg13g2_fill_8 FILLER_132_352 ();
 sg13g2_fill_8 FILLER_132_360 ();
 sg13g2_fill_8 FILLER_132_368 ();
 sg13g2_fill_8 FILLER_132_376 ();
 sg13g2_fill_8 FILLER_132_384 ();
 sg13g2_fill_8 FILLER_132_392 ();
 sg13g2_fill_8 FILLER_132_400 ();
 sg13g2_fill_8 FILLER_132_408 ();
 sg13g2_fill_8 FILLER_132_416 ();
 sg13g2_fill_8 FILLER_132_424 ();
 sg13g2_fill_8 FILLER_132_432 ();
 sg13g2_fill_8 FILLER_132_440 ();
 sg13g2_fill_8 FILLER_132_448 ();
 sg13g2_fill_8 FILLER_132_456 ();
 sg13g2_fill_8 FILLER_132_464 ();
 sg13g2_fill_8 FILLER_132_472 ();
 sg13g2_fill_8 FILLER_132_480 ();
 sg13g2_fill_8 FILLER_132_488 ();
 sg13g2_fill_8 FILLER_132_496 ();
 sg13g2_fill_8 FILLER_132_504 ();
 sg13g2_fill_8 FILLER_132_512 ();
 sg13g2_fill_8 FILLER_132_520 ();
 sg13g2_fill_8 FILLER_132_528 ();
 sg13g2_fill_8 FILLER_132_536 ();
 sg13g2_fill_8 FILLER_132_544 ();
 sg13g2_fill_8 FILLER_132_552 ();
 sg13g2_fill_8 FILLER_132_560 ();
 sg13g2_fill_8 FILLER_132_568 ();
 sg13g2_fill_8 FILLER_132_576 ();
 sg13g2_fill_8 FILLER_132_584 ();
 sg13g2_fill_8 FILLER_132_592 ();
 sg13g2_fill_8 FILLER_132_600 ();
 sg13g2_fill_8 FILLER_132_608 ();
 sg13g2_fill_8 FILLER_132_616 ();
 sg13g2_fill_8 FILLER_132_624 ();
 sg13g2_fill_8 FILLER_132_632 ();
 sg13g2_fill_8 FILLER_132_640 ();
 sg13g2_fill_8 FILLER_132_648 ();
 sg13g2_fill_8 FILLER_132_656 ();
 sg13g2_fill_8 FILLER_132_664 ();
 sg13g2_fill_8 FILLER_132_672 ();
 sg13g2_fill_8 FILLER_132_680 ();
 sg13g2_fill_8 FILLER_132_688 ();
 sg13g2_fill_8 FILLER_132_696 ();
 sg13g2_fill_8 FILLER_132_704 ();
 sg13g2_fill_8 FILLER_132_712 ();
 sg13g2_fill_8 FILLER_132_720 ();
 sg13g2_fill_8 FILLER_132_728 ();
 sg13g2_fill_8 FILLER_132_736 ();
 sg13g2_fill_8 FILLER_132_744 ();
 sg13g2_fill_8 FILLER_132_752 ();
 sg13g2_fill_8 FILLER_132_760 ();
 sg13g2_fill_8 FILLER_132_768 ();
 sg13g2_fill_8 FILLER_132_776 ();
 sg13g2_fill_8 FILLER_132_784 ();
 sg13g2_fill_8 FILLER_132_792 ();
 sg13g2_fill_8 FILLER_132_800 ();
 sg13g2_fill_8 FILLER_132_808 ();
 sg13g2_fill_8 FILLER_132_816 ();
 sg13g2_fill_8 FILLER_132_824 ();
 sg13g2_fill_8 FILLER_132_832 ();
 sg13g2_fill_8 FILLER_132_840 ();
 sg13g2_fill_8 FILLER_132_848 ();
 sg13g2_fill_8 FILLER_132_856 ();
 sg13g2_fill_8 FILLER_132_864 ();
 sg13g2_fill_8 FILLER_132_872 ();
 sg13g2_fill_8 FILLER_132_880 ();
 sg13g2_fill_8 FILLER_132_888 ();
 sg13g2_fill_8 FILLER_132_896 ();
 sg13g2_fill_8 FILLER_132_904 ();
 sg13g2_fill_8 FILLER_132_912 ();
 sg13g2_fill_8 FILLER_132_920 ();
 sg13g2_fill_8 FILLER_132_928 ();
 sg13g2_fill_8 FILLER_132_936 ();
 sg13g2_fill_8 FILLER_132_944 ();
 sg13g2_fill_8 FILLER_132_952 ();
 sg13g2_fill_8 FILLER_132_960 ();
 sg13g2_fill_8 FILLER_132_968 ();
 sg13g2_fill_8 FILLER_132_976 ();
 sg13g2_fill_8 FILLER_132_984 ();
 sg13g2_fill_8 FILLER_132_992 ();
 sg13g2_fill_8 FILLER_132_1000 ();
 sg13g2_fill_8 FILLER_132_1008 ();
 sg13g2_fill_8 FILLER_132_1016 ();
 sg13g2_fill_8 FILLER_132_1024 ();
 sg13g2_fill_8 FILLER_132_1032 ();
 sg13g2_fill_8 FILLER_132_1040 ();
 sg13g2_fill_8 FILLER_132_1048 ();
 sg13g2_fill_8 FILLER_132_1056 ();
 sg13g2_fill_8 FILLER_132_1064 ();
 sg13g2_fill_8 FILLER_132_1072 ();
 sg13g2_fill_8 FILLER_132_1080 ();
 sg13g2_fill_8 FILLER_132_1088 ();
 sg13g2_fill_8 FILLER_132_1096 ();
 sg13g2_fill_8 FILLER_132_1104 ();
 sg13g2_fill_8 FILLER_132_1112 ();
 sg13g2_fill_8 FILLER_132_1120 ();
 sg13g2_fill_8 FILLER_132_1128 ();
 sg13g2_fill_8 FILLER_132_1136 ();
 sg13g2_fill_8 FILLER_133_0 ();
 sg13g2_fill_8 FILLER_133_8 ();
 sg13g2_fill_8 FILLER_133_16 ();
 sg13g2_fill_8 FILLER_133_24 ();
 sg13g2_fill_8 FILLER_133_32 ();
 sg13g2_fill_8 FILLER_133_40 ();
 sg13g2_fill_8 FILLER_133_48 ();
 sg13g2_fill_8 FILLER_133_56 ();
 sg13g2_fill_8 FILLER_133_64 ();
 sg13g2_fill_8 FILLER_133_72 ();
 sg13g2_fill_8 FILLER_133_80 ();
 sg13g2_fill_8 FILLER_133_88 ();
 sg13g2_fill_8 FILLER_133_96 ();
 sg13g2_fill_8 FILLER_133_104 ();
 sg13g2_fill_8 FILLER_133_112 ();
 sg13g2_fill_8 FILLER_133_120 ();
 sg13g2_fill_8 FILLER_133_128 ();
 sg13g2_fill_8 FILLER_133_136 ();
 sg13g2_fill_8 FILLER_133_144 ();
 sg13g2_fill_8 FILLER_133_152 ();
 sg13g2_fill_8 FILLER_133_160 ();
 sg13g2_fill_8 FILLER_133_168 ();
 sg13g2_fill_8 FILLER_133_176 ();
 sg13g2_fill_8 FILLER_133_184 ();
 sg13g2_fill_8 FILLER_133_192 ();
 sg13g2_fill_8 FILLER_133_200 ();
 sg13g2_fill_8 FILLER_133_208 ();
 sg13g2_fill_8 FILLER_133_216 ();
 sg13g2_fill_8 FILLER_133_224 ();
 sg13g2_fill_8 FILLER_133_232 ();
 sg13g2_fill_8 FILLER_133_240 ();
 sg13g2_fill_8 FILLER_133_248 ();
 sg13g2_fill_8 FILLER_133_256 ();
 sg13g2_fill_8 FILLER_133_264 ();
 sg13g2_fill_8 FILLER_133_272 ();
 sg13g2_fill_8 FILLER_133_280 ();
 sg13g2_fill_8 FILLER_133_288 ();
 sg13g2_fill_8 FILLER_133_296 ();
 sg13g2_fill_8 FILLER_133_304 ();
 sg13g2_fill_8 FILLER_133_312 ();
 sg13g2_fill_8 FILLER_133_320 ();
 sg13g2_fill_8 FILLER_133_328 ();
 sg13g2_fill_8 FILLER_133_336 ();
 sg13g2_fill_8 FILLER_133_344 ();
 sg13g2_fill_8 FILLER_133_352 ();
 sg13g2_fill_8 FILLER_133_360 ();
 sg13g2_fill_8 FILLER_133_368 ();
 sg13g2_fill_8 FILLER_133_376 ();
 sg13g2_fill_8 FILLER_133_384 ();
 sg13g2_fill_8 FILLER_133_392 ();
 sg13g2_fill_8 FILLER_133_400 ();
 sg13g2_fill_8 FILLER_133_408 ();
 sg13g2_fill_8 FILLER_133_416 ();
 sg13g2_fill_8 FILLER_133_424 ();
 sg13g2_fill_8 FILLER_133_432 ();
 sg13g2_fill_8 FILLER_133_440 ();
 sg13g2_fill_8 FILLER_133_448 ();
 sg13g2_fill_8 FILLER_133_456 ();
 sg13g2_fill_8 FILLER_133_464 ();
 sg13g2_fill_8 FILLER_133_472 ();
 sg13g2_fill_8 FILLER_133_480 ();
 sg13g2_fill_8 FILLER_133_488 ();
 sg13g2_fill_8 FILLER_133_496 ();
 sg13g2_fill_8 FILLER_133_504 ();
 sg13g2_fill_8 FILLER_133_512 ();
 sg13g2_fill_8 FILLER_133_520 ();
 sg13g2_fill_8 FILLER_133_528 ();
 sg13g2_fill_8 FILLER_133_536 ();
 sg13g2_fill_8 FILLER_133_544 ();
 sg13g2_fill_8 FILLER_133_552 ();
 sg13g2_fill_8 FILLER_133_560 ();
 sg13g2_fill_8 FILLER_133_568 ();
 sg13g2_fill_8 FILLER_133_576 ();
 sg13g2_fill_8 FILLER_133_584 ();
 sg13g2_fill_8 FILLER_133_592 ();
 sg13g2_fill_8 FILLER_133_600 ();
 sg13g2_fill_8 FILLER_133_608 ();
 sg13g2_fill_8 FILLER_133_616 ();
 sg13g2_fill_8 FILLER_133_624 ();
 sg13g2_fill_8 FILLER_133_632 ();
 sg13g2_fill_8 FILLER_133_640 ();
 sg13g2_fill_8 FILLER_133_648 ();
 sg13g2_fill_8 FILLER_133_656 ();
 sg13g2_fill_8 FILLER_133_664 ();
 sg13g2_fill_8 FILLER_133_672 ();
 sg13g2_fill_8 FILLER_133_680 ();
 sg13g2_fill_8 FILLER_133_688 ();
 sg13g2_fill_8 FILLER_133_696 ();
 sg13g2_fill_8 FILLER_133_704 ();
 sg13g2_fill_8 FILLER_133_712 ();
 sg13g2_fill_8 FILLER_133_720 ();
 sg13g2_fill_8 FILLER_133_728 ();
 sg13g2_fill_8 FILLER_133_736 ();
 sg13g2_fill_8 FILLER_133_744 ();
 sg13g2_fill_8 FILLER_133_752 ();
 sg13g2_fill_8 FILLER_133_760 ();
 sg13g2_fill_8 FILLER_133_768 ();
 sg13g2_fill_8 FILLER_133_776 ();
 sg13g2_fill_8 FILLER_133_784 ();
 sg13g2_fill_8 FILLER_133_792 ();
 sg13g2_fill_8 FILLER_133_800 ();
 sg13g2_fill_8 FILLER_133_808 ();
 sg13g2_fill_8 FILLER_133_816 ();
 sg13g2_fill_8 FILLER_133_824 ();
 sg13g2_fill_8 FILLER_133_832 ();
 sg13g2_fill_8 FILLER_133_840 ();
 sg13g2_fill_8 FILLER_133_848 ();
 sg13g2_fill_8 FILLER_133_856 ();
 sg13g2_fill_8 FILLER_133_864 ();
 sg13g2_fill_8 FILLER_133_872 ();
 sg13g2_fill_8 FILLER_133_880 ();
 sg13g2_fill_8 FILLER_133_888 ();
 sg13g2_fill_8 FILLER_133_896 ();
 sg13g2_fill_8 FILLER_133_904 ();
 sg13g2_fill_8 FILLER_133_912 ();
 sg13g2_fill_8 FILLER_133_920 ();
 sg13g2_fill_8 FILLER_133_928 ();
 sg13g2_fill_8 FILLER_133_936 ();
 sg13g2_fill_8 FILLER_133_944 ();
 sg13g2_fill_8 FILLER_133_952 ();
 sg13g2_fill_8 FILLER_133_960 ();
 sg13g2_fill_8 FILLER_133_968 ();
 sg13g2_fill_8 FILLER_133_976 ();
 sg13g2_fill_8 FILLER_133_984 ();
 sg13g2_fill_8 FILLER_133_992 ();
 sg13g2_fill_8 FILLER_133_1000 ();
 sg13g2_fill_8 FILLER_133_1008 ();
 sg13g2_fill_8 FILLER_133_1016 ();
 sg13g2_fill_8 FILLER_133_1024 ();
 sg13g2_fill_8 FILLER_133_1032 ();
 sg13g2_fill_8 FILLER_133_1040 ();
 sg13g2_fill_8 FILLER_133_1048 ();
 sg13g2_fill_8 FILLER_133_1056 ();
 sg13g2_fill_8 FILLER_133_1064 ();
 sg13g2_fill_8 FILLER_133_1072 ();
 sg13g2_fill_8 FILLER_133_1080 ();
 sg13g2_fill_8 FILLER_133_1088 ();
 sg13g2_fill_8 FILLER_133_1096 ();
 sg13g2_fill_8 FILLER_133_1104 ();
 sg13g2_fill_8 FILLER_133_1112 ();
 sg13g2_fill_8 FILLER_133_1120 ();
 sg13g2_fill_8 FILLER_133_1128 ();
 sg13g2_fill_8 FILLER_133_1136 ();
 sg13g2_fill_8 FILLER_134_0 ();
 sg13g2_fill_8 FILLER_134_8 ();
 sg13g2_fill_8 FILLER_134_16 ();
 sg13g2_fill_8 FILLER_134_24 ();
 sg13g2_fill_8 FILLER_134_32 ();
 sg13g2_fill_8 FILLER_134_40 ();
 sg13g2_fill_8 FILLER_134_48 ();
 sg13g2_fill_8 FILLER_134_56 ();
 sg13g2_fill_8 FILLER_134_64 ();
 sg13g2_fill_8 FILLER_134_72 ();
 sg13g2_fill_8 FILLER_134_80 ();
 sg13g2_fill_8 FILLER_134_88 ();
 sg13g2_fill_8 FILLER_134_96 ();
 sg13g2_fill_8 FILLER_134_104 ();
 sg13g2_fill_8 FILLER_134_112 ();
 sg13g2_fill_8 FILLER_134_120 ();
 sg13g2_fill_8 FILLER_134_128 ();
 sg13g2_fill_8 FILLER_134_136 ();
 sg13g2_fill_8 FILLER_134_144 ();
 sg13g2_fill_8 FILLER_134_152 ();
 sg13g2_fill_8 FILLER_134_160 ();
 sg13g2_fill_8 FILLER_134_168 ();
 sg13g2_fill_8 FILLER_134_176 ();
 sg13g2_fill_8 FILLER_134_184 ();
 sg13g2_fill_8 FILLER_134_192 ();
 sg13g2_fill_8 FILLER_134_200 ();
 sg13g2_fill_8 FILLER_134_208 ();
 sg13g2_fill_8 FILLER_134_216 ();
 sg13g2_fill_8 FILLER_134_224 ();
 sg13g2_fill_8 FILLER_134_232 ();
 sg13g2_fill_8 FILLER_134_240 ();
 sg13g2_fill_8 FILLER_134_248 ();
 sg13g2_fill_8 FILLER_134_256 ();
 sg13g2_fill_8 FILLER_134_264 ();
 sg13g2_fill_8 FILLER_134_272 ();
 sg13g2_fill_8 FILLER_134_280 ();
 sg13g2_fill_8 FILLER_134_288 ();
 sg13g2_fill_8 FILLER_134_296 ();
 sg13g2_fill_8 FILLER_134_304 ();
 sg13g2_fill_8 FILLER_134_312 ();
 sg13g2_fill_8 FILLER_134_320 ();
 sg13g2_fill_8 FILLER_134_328 ();
 sg13g2_fill_8 FILLER_134_336 ();
 sg13g2_fill_8 FILLER_134_344 ();
 sg13g2_fill_8 FILLER_134_352 ();
 sg13g2_fill_8 FILLER_134_360 ();
 sg13g2_fill_8 FILLER_134_368 ();
 sg13g2_fill_8 FILLER_134_376 ();
 sg13g2_fill_8 FILLER_134_384 ();
 sg13g2_fill_8 FILLER_134_392 ();
 sg13g2_fill_8 FILLER_134_400 ();
 sg13g2_fill_8 FILLER_134_408 ();
 sg13g2_fill_8 FILLER_134_416 ();
 sg13g2_fill_8 FILLER_134_424 ();
 sg13g2_fill_8 FILLER_134_432 ();
 sg13g2_fill_8 FILLER_134_440 ();
 sg13g2_fill_8 FILLER_134_448 ();
 sg13g2_fill_8 FILLER_134_456 ();
 sg13g2_fill_8 FILLER_134_464 ();
 sg13g2_fill_8 FILLER_134_472 ();
 sg13g2_fill_8 FILLER_134_480 ();
 sg13g2_fill_8 FILLER_134_488 ();
 sg13g2_fill_8 FILLER_134_496 ();
 sg13g2_fill_8 FILLER_134_504 ();
 sg13g2_fill_8 FILLER_134_512 ();
 sg13g2_fill_8 FILLER_134_520 ();
 sg13g2_fill_8 FILLER_134_528 ();
 sg13g2_fill_8 FILLER_134_536 ();
 sg13g2_fill_8 FILLER_134_544 ();
 sg13g2_fill_8 FILLER_134_552 ();
 sg13g2_fill_8 FILLER_134_560 ();
 sg13g2_fill_8 FILLER_134_568 ();
 sg13g2_fill_8 FILLER_134_576 ();
 sg13g2_fill_8 FILLER_134_584 ();
 sg13g2_fill_8 FILLER_134_592 ();
 sg13g2_fill_8 FILLER_134_600 ();
 sg13g2_fill_8 FILLER_134_608 ();
 sg13g2_fill_8 FILLER_134_616 ();
 sg13g2_fill_8 FILLER_134_624 ();
 sg13g2_fill_8 FILLER_134_632 ();
 sg13g2_fill_8 FILLER_134_640 ();
 sg13g2_fill_8 FILLER_134_648 ();
 sg13g2_fill_8 FILLER_134_656 ();
 sg13g2_fill_8 FILLER_134_664 ();
 sg13g2_fill_8 FILLER_134_672 ();
 sg13g2_fill_8 FILLER_134_680 ();
 sg13g2_fill_8 FILLER_134_688 ();
 sg13g2_fill_8 FILLER_134_696 ();
 sg13g2_fill_8 FILLER_134_704 ();
 sg13g2_fill_8 FILLER_134_712 ();
 sg13g2_fill_8 FILLER_134_720 ();
 sg13g2_fill_8 FILLER_134_728 ();
 sg13g2_fill_8 FILLER_134_736 ();
 sg13g2_fill_8 FILLER_134_744 ();
 sg13g2_fill_8 FILLER_134_752 ();
 sg13g2_fill_8 FILLER_134_760 ();
 sg13g2_fill_8 FILLER_134_768 ();
 sg13g2_fill_8 FILLER_134_776 ();
 sg13g2_fill_8 FILLER_134_784 ();
 sg13g2_fill_8 FILLER_134_792 ();
 sg13g2_fill_8 FILLER_134_800 ();
 sg13g2_fill_8 FILLER_134_808 ();
 sg13g2_fill_8 FILLER_134_816 ();
 sg13g2_fill_8 FILLER_134_824 ();
 sg13g2_fill_8 FILLER_134_832 ();
 sg13g2_fill_8 FILLER_134_840 ();
 sg13g2_fill_8 FILLER_134_848 ();
 sg13g2_fill_8 FILLER_134_856 ();
 sg13g2_fill_8 FILLER_134_864 ();
 sg13g2_fill_8 FILLER_134_872 ();
 sg13g2_fill_8 FILLER_134_880 ();
 sg13g2_fill_8 FILLER_134_888 ();
 sg13g2_fill_8 FILLER_134_896 ();
 sg13g2_fill_8 FILLER_134_904 ();
 sg13g2_fill_8 FILLER_134_912 ();
 sg13g2_fill_8 FILLER_134_920 ();
 sg13g2_fill_8 FILLER_134_928 ();
 sg13g2_fill_8 FILLER_134_936 ();
 sg13g2_fill_8 FILLER_134_944 ();
 sg13g2_fill_8 FILLER_134_952 ();
 sg13g2_fill_8 FILLER_134_960 ();
 sg13g2_fill_8 FILLER_134_968 ();
 sg13g2_fill_8 FILLER_134_976 ();
 sg13g2_fill_8 FILLER_134_984 ();
 sg13g2_fill_8 FILLER_134_992 ();
 sg13g2_fill_8 FILLER_134_1000 ();
 sg13g2_fill_8 FILLER_134_1008 ();
 sg13g2_fill_8 FILLER_134_1016 ();
 sg13g2_fill_8 FILLER_134_1024 ();
 sg13g2_fill_8 FILLER_134_1032 ();
 sg13g2_fill_8 FILLER_134_1040 ();
 sg13g2_fill_8 FILLER_134_1048 ();
 sg13g2_fill_8 FILLER_134_1056 ();
 sg13g2_fill_8 FILLER_134_1064 ();
 sg13g2_fill_8 FILLER_134_1072 ();
 sg13g2_fill_8 FILLER_134_1080 ();
 sg13g2_fill_8 FILLER_134_1088 ();
 sg13g2_fill_8 FILLER_134_1096 ();
 sg13g2_fill_8 FILLER_134_1104 ();
 sg13g2_fill_8 FILLER_134_1112 ();
 sg13g2_fill_8 FILLER_134_1120 ();
 sg13g2_fill_8 FILLER_134_1128 ();
 sg13g2_fill_8 FILLER_134_1136 ();
 sg13g2_fill_8 FILLER_135_0 ();
 sg13g2_fill_8 FILLER_135_8 ();
 sg13g2_fill_8 FILLER_135_16 ();
 sg13g2_fill_8 FILLER_135_24 ();
 sg13g2_fill_8 FILLER_135_32 ();
 sg13g2_fill_8 FILLER_135_40 ();
 sg13g2_fill_8 FILLER_135_48 ();
 sg13g2_fill_8 FILLER_135_56 ();
 sg13g2_fill_8 FILLER_135_64 ();
 sg13g2_fill_8 FILLER_135_72 ();
 sg13g2_fill_8 FILLER_135_80 ();
 sg13g2_fill_8 FILLER_135_88 ();
 sg13g2_fill_8 FILLER_135_96 ();
 sg13g2_fill_8 FILLER_135_104 ();
 sg13g2_fill_8 FILLER_135_112 ();
 sg13g2_fill_8 FILLER_135_120 ();
 sg13g2_fill_8 FILLER_135_128 ();
 sg13g2_fill_8 FILLER_135_136 ();
 sg13g2_fill_8 FILLER_135_144 ();
 sg13g2_fill_8 FILLER_135_152 ();
 sg13g2_fill_8 FILLER_135_160 ();
 sg13g2_fill_8 FILLER_135_168 ();
 sg13g2_fill_8 FILLER_135_176 ();
 sg13g2_fill_8 FILLER_135_184 ();
 sg13g2_fill_8 FILLER_135_192 ();
 sg13g2_fill_8 FILLER_135_200 ();
 sg13g2_fill_8 FILLER_135_208 ();
 sg13g2_fill_8 FILLER_135_216 ();
 sg13g2_fill_8 FILLER_135_224 ();
 sg13g2_fill_8 FILLER_135_232 ();
 sg13g2_fill_8 FILLER_135_240 ();
 sg13g2_fill_8 FILLER_135_248 ();
 sg13g2_fill_8 FILLER_135_256 ();
 sg13g2_fill_8 FILLER_135_264 ();
 sg13g2_fill_8 FILLER_135_272 ();
 sg13g2_fill_8 FILLER_135_280 ();
 sg13g2_fill_8 FILLER_135_288 ();
 sg13g2_fill_8 FILLER_135_296 ();
 sg13g2_fill_8 FILLER_135_304 ();
 sg13g2_fill_8 FILLER_135_312 ();
 sg13g2_fill_8 FILLER_135_320 ();
 sg13g2_fill_8 FILLER_135_328 ();
 sg13g2_fill_8 FILLER_135_336 ();
 sg13g2_fill_8 FILLER_135_344 ();
 sg13g2_fill_8 FILLER_135_352 ();
 sg13g2_fill_8 FILLER_135_360 ();
 sg13g2_fill_8 FILLER_135_368 ();
 sg13g2_fill_8 FILLER_135_376 ();
 sg13g2_fill_8 FILLER_135_384 ();
 sg13g2_fill_8 FILLER_135_392 ();
 sg13g2_fill_8 FILLER_135_400 ();
 sg13g2_fill_8 FILLER_135_408 ();
 sg13g2_fill_8 FILLER_135_416 ();
 sg13g2_fill_8 FILLER_135_424 ();
 sg13g2_fill_8 FILLER_135_432 ();
 sg13g2_fill_8 FILLER_135_440 ();
 sg13g2_fill_8 FILLER_135_448 ();
 sg13g2_fill_8 FILLER_135_456 ();
 sg13g2_fill_8 FILLER_135_464 ();
 sg13g2_fill_8 FILLER_135_472 ();
 sg13g2_fill_8 FILLER_135_480 ();
 sg13g2_fill_8 FILLER_135_488 ();
 sg13g2_fill_8 FILLER_135_496 ();
 sg13g2_fill_8 FILLER_135_504 ();
 sg13g2_fill_8 FILLER_135_512 ();
 sg13g2_fill_8 FILLER_135_520 ();
 sg13g2_fill_8 FILLER_135_528 ();
 sg13g2_fill_8 FILLER_135_536 ();
 sg13g2_fill_8 FILLER_135_544 ();
 sg13g2_fill_8 FILLER_135_552 ();
 sg13g2_fill_8 FILLER_135_560 ();
 sg13g2_fill_8 FILLER_135_568 ();
 sg13g2_fill_8 FILLER_135_576 ();
 sg13g2_fill_8 FILLER_135_584 ();
 sg13g2_fill_8 FILLER_135_592 ();
 sg13g2_fill_8 FILLER_135_600 ();
 sg13g2_fill_8 FILLER_135_608 ();
 sg13g2_fill_8 FILLER_135_616 ();
 sg13g2_fill_8 FILLER_135_624 ();
 sg13g2_fill_8 FILLER_135_632 ();
 sg13g2_fill_8 FILLER_135_640 ();
 sg13g2_fill_8 FILLER_135_648 ();
 sg13g2_fill_8 FILLER_135_656 ();
 sg13g2_fill_8 FILLER_135_664 ();
 sg13g2_fill_8 FILLER_135_672 ();
 sg13g2_fill_8 FILLER_135_680 ();
 sg13g2_fill_8 FILLER_135_688 ();
 sg13g2_fill_8 FILLER_135_696 ();
 sg13g2_fill_8 FILLER_135_704 ();
 sg13g2_fill_8 FILLER_135_712 ();
 sg13g2_fill_8 FILLER_135_720 ();
 sg13g2_fill_8 FILLER_135_728 ();
 sg13g2_fill_8 FILLER_135_736 ();
 sg13g2_fill_8 FILLER_135_744 ();
 sg13g2_fill_8 FILLER_135_752 ();
 sg13g2_fill_8 FILLER_135_760 ();
 sg13g2_fill_8 FILLER_135_768 ();
 sg13g2_fill_8 FILLER_135_776 ();
 sg13g2_fill_8 FILLER_135_784 ();
 sg13g2_fill_8 FILLER_135_792 ();
 sg13g2_fill_8 FILLER_135_800 ();
 sg13g2_fill_8 FILLER_135_808 ();
 sg13g2_fill_8 FILLER_135_816 ();
 sg13g2_fill_8 FILLER_135_824 ();
 sg13g2_fill_8 FILLER_135_832 ();
 sg13g2_fill_8 FILLER_135_840 ();
 sg13g2_fill_8 FILLER_135_848 ();
 sg13g2_fill_8 FILLER_135_856 ();
 sg13g2_fill_8 FILLER_135_864 ();
 sg13g2_fill_8 FILLER_135_872 ();
 sg13g2_fill_8 FILLER_135_880 ();
 sg13g2_fill_8 FILLER_135_888 ();
 sg13g2_fill_8 FILLER_135_896 ();
 sg13g2_fill_8 FILLER_135_904 ();
 sg13g2_fill_8 FILLER_135_912 ();
 sg13g2_fill_8 FILLER_135_920 ();
 sg13g2_fill_8 FILLER_135_928 ();
 sg13g2_fill_8 FILLER_135_936 ();
 sg13g2_fill_8 FILLER_135_944 ();
 sg13g2_fill_8 FILLER_135_952 ();
 sg13g2_fill_8 FILLER_135_960 ();
 sg13g2_fill_8 FILLER_135_968 ();
 sg13g2_fill_8 FILLER_135_976 ();
 sg13g2_fill_8 FILLER_135_984 ();
 sg13g2_fill_8 FILLER_135_992 ();
 sg13g2_fill_8 FILLER_135_1000 ();
 sg13g2_fill_8 FILLER_135_1008 ();
 sg13g2_fill_8 FILLER_135_1016 ();
 sg13g2_fill_8 FILLER_135_1024 ();
 sg13g2_fill_8 FILLER_135_1032 ();
 sg13g2_fill_8 FILLER_135_1040 ();
 sg13g2_fill_8 FILLER_135_1048 ();
 sg13g2_fill_8 FILLER_135_1056 ();
 sg13g2_fill_8 FILLER_135_1064 ();
 sg13g2_fill_8 FILLER_135_1072 ();
 sg13g2_fill_8 FILLER_135_1080 ();
 sg13g2_fill_8 FILLER_135_1088 ();
 sg13g2_fill_8 FILLER_135_1096 ();
 sg13g2_fill_8 FILLER_135_1104 ();
 sg13g2_fill_8 FILLER_135_1112 ();
 sg13g2_fill_8 FILLER_135_1120 ();
 sg13g2_fill_8 FILLER_135_1128 ();
 sg13g2_fill_8 FILLER_135_1136 ();
 sg13g2_fill_8 FILLER_136_0 ();
 sg13g2_fill_8 FILLER_136_8 ();
 sg13g2_fill_8 FILLER_136_16 ();
 sg13g2_fill_8 FILLER_136_24 ();
 sg13g2_fill_8 FILLER_136_32 ();
 sg13g2_fill_8 FILLER_136_40 ();
 sg13g2_fill_8 FILLER_136_48 ();
 sg13g2_fill_8 FILLER_136_56 ();
 sg13g2_fill_8 FILLER_136_64 ();
 sg13g2_fill_8 FILLER_136_72 ();
 sg13g2_fill_8 FILLER_136_80 ();
 sg13g2_fill_8 FILLER_136_88 ();
 sg13g2_fill_8 FILLER_136_96 ();
 sg13g2_fill_8 FILLER_136_104 ();
 sg13g2_fill_8 FILLER_136_112 ();
 sg13g2_fill_8 FILLER_136_120 ();
 sg13g2_fill_8 FILLER_136_128 ();
 sg13g2_fill_8 FILLER_136_136 ();
 sg13g2_fill_8 FILLER_136_144 ();
 sg13g2_fill_8 FILLER_136_152 ();
 sg13g2_fill_8 FILLER_136_160 ();
 sg13g2_fill_8 FILLER_136_168 ();
 sg13g2_fill_8 FILLER_136_176 ();
 sg13g2_fill_8 FILLER_136_184 ();
 sg13g2_fill_8 FILLER_136_192 ();
 sg13g2_fill_8 FILLER_136_200 ();
 sg13g2_fill_8 FILLER_136_208 ();
 sg13g2_fill_8 FILLER_136_216 ();
 sg13g2_fill_8 FILLER_136_224 ();
 sg13g2_fill_8 FILLER_136_232 ();
 sg13g2_fill_8 FILLER_136_240 ();
 sg13g2_fill_8 FILLER_136_248 ();
 sg13g2_fill_8 FILLER_136_256 ();
 sg13g2_fill_8 FILLER_136_264 ();
 sg13g2_fill_8 FILLER_136_272 ();
 sg13g2_fill_8 FILLER_136_280 ();
 sg13g2_fill_8 FILLER_136_288 ();
 sg13g2_fill_8 FILLER_136_296 ();
 sg13g2_fill_8 FILLER_136_304 ();
 sg13g2_fill_8 FILLER_136_312 ();
 sg13g2_fill_8 FILLER_136_320 ();
 sg13g2_fill_8 FILLER_136_328 ();
 sg13g2_fill_8 FILLER_136_336 ();
 sg13g2_fill_8 FILLER_136_344 ();
 sg13g2_fill_8 FILLER_136_352 ();
 sg13g2_fill_8 FILLER_136_360 ();
 sg13g2_fill_8 FILLER_136_368 ();
 sg13g2_fill_8 FILLER_136_376 ();
 sg13g2_fill_8 FILLER_136_384 ();
 sg13g2_fill_8 FILLER_136_392 ();
 sg13g2_fill_8 FILLER_136_400 ();
 sg13g2_fill_8 FILLER_136_408 ();
 sg13g2_fill_8 FILLER_136_416 ();
 sg13g2_fill_8 FILLER_136_424 ();
 sg13g2_fill_8 FILLER_136_432 ();
 sg13g2_fill_8 FILLER_136_440 ();
 sg13g2_fill_8 FILLER_136_448 ();
 sg13g2_fill_8 FILLER_136_456 ();
 sg13g2_fill_8 FILLER_136_464 ();
 sg13g2_fill_8 FILLER_136_472 ();
 sg13g2_fill_8 FILLER_136_480 ();
 sg13g2_fill_8 FILLER_136_488 ();
 sg13g2_fill_8 FILLER_136_496 ();
 sg13g2_fill_8 FILLER_136_504 ();
 sg13g2_fill_8 FILLER_136_512 ();
 sg13g2_fill_8 FILLER_136_520 ();
 sg13g2_fill_8 FILLER_136_528 ();
 sg13g2_fill_8 FILLER_136_536 ();
 sg13g2_fill_8 FILLER_136_544 ();
 sg13g2_fill_8 FILLER_136_552 ();
 sg13g2_fill_8 FILLER_136_560 ();
 sg13g2_fill_8 FILLER_136_568 ();
 sg13g2_fill_8 FILLER_136_576 ();
 sg13g2_fill_8 FILLER_136_584 ();
 sg13g2_fill_8 FILLER_136_592 ();
 sg13g2_fill_8 FILLER_136_600 ();
 sg13g2_fill_8 FILLER_136_608 ();
 sg13g2_fill_8 FILLER_136_616 ();
 sg13g2_fill_8 FILLER_136_624 ();
 sg13g2_fill_8 FILLER_136_632 ();
 sg13g2_fill_8 FILLER_136_640 ();
 sg13g2_fill_8 FILLER_136_648 ();
 sg13g2_fill_8 FILLER_136_656 ();
 sg13g2_fill_8 FILLER_136_664 ();
 sg13g2_fill_8 FILLER_136_672 ();
 sg13g2_fill_8 FILLER_136_680 ();
 sg13g2_fill_8 FILLER_136_688 ();
 sg13g2_fill_8 FILLER_136_696 ();
 sg13g2_fill_8 FILLER_136_704 ();
 sg13g2_fill_8 FILLER_136_712 ();
 sg13g2_fill_8 FILLER_136_720 ();
 sg13g2_fill_8 FILLER_136_728 ();
 sg13g2_fill_8 FILLER_136_736 ();
 sg13g2_fill_8 FILLER_136_744 ();
 sg13g2_fill_8 FILLER_136_752 ();
 sg13g2_fill_8 FILLER_136_760 ();
 sg13g2_fill_8 FILLER_136_768 ();
 sg13g2_fill_8 FILLER_136_776 ();
 sg13g2_fill_8 FILLER_136_784 ();
 sg13g2_fill_8 FILLER_136_792 ();
 sg13g2_fill_8 FILLER_136_800 ();
 sg13g2_fill_8 FILLER_136_808 ();
 sg13g2_fill_8 FILLER_136_816 ();
 sg13g2_fill_8 FILLER_136_824 ();
 sg13g2_fill_8 FILLER_136_832 ();
 sg13g2_fill_8 FILLER_136_840 ();
 sg13g2_fill_8 FILLER_136_848 ();
 sg13g2_fill_8 FILLER_136_856 ();
 sg13g2_fill_8 FILLER_136_864 ();
 sg13g2_fill_8 FILLER_136_872 ();
 sg13g2_fill_8 FILLER_136_880 ();
 sg13g2_fill_8 FILLER_136_888 ();
 sg13g2_fill_8 FILLER_136_896 ();
 sg13g2_fill_8 FILLER_136_904 ();
 sg13g2_fill_8 FILLER_136_912 ();
 sg13g2_fill_8 FILLER_136_920 ();
 sg13g2_fill_8 FILLER_136_928 ();
 sg13g2_fill_8 FILLER_136_936 ();
 sg13g2_fill_8 FILLER_136_944 ();
 sg13g2_fill_8 FILLER_136_952 ();
 sg13g2_fill_8 FILLER_136_960 ();
 sg13g2_fill_8 FILLER_136_968 ();
 sg13g2_fill_8 FILLER_136_976 ();
 sg13g2_fill_8 FILLER_136_984 ();
 sg13g2_fill_8 FILLER_136_992 ();
 sg13g2_fill_8 FILLER_136_1000 ();
 sg13g2_fill_8 FILLER_136_1008 ();
 sg13g2_fill_8 FILLER_136_1016 ();
 sg13g2_fill_8 FILLER_136_1024 ();
 sg13g2_fill_8 FILLER_136_1032 ();
 sg13g2_fill_8 FILLER_136_1040 ();
 sg13g2_fill_8 FILLER_136_1048 ();
 sg13g2_fill_8 FILLER_136_1056 ();
 sg13g2_fill_8 FILLER_136_1064 ();
 sg13g2_fill_8 FILLER_136_1072 ();
 sg13g2_fill_8 FILLER_136_1080 ();
 sg13g2_fill_8 FILLER_136_1088 ();
 sg13g2_fill_8 FILLER_136_1096 ();
 sg13g2_fill_8 FILLER_136_1104 ();
 sg13g2_fill_8 FILLER_136_1112 ();
 sg13g2_fill_8 FILLER_136_1120 ();
 sg13g2_fill_8 FILLER_136_1128 ();
 sg13g2_fill_8 FILLER_136_1136 ();
 sg13g2_fill_8 FILLER_137_0 ();
 sg13g2_fill_8 FILLER_137_8 ();
 sg13g2_fill_8 FILLER_137_16 ();
 sg13g2_fill_8 FILLER_137_24 ();
 sg13g2_fill_8 FILLER_137_32 ();
 sg13g2_fill_8 FILLER_137_40 ();
 sg13g2_fill_8 FILLER_137_48 ();
 sg13g2_fill_8 FILLER_137_56 ();
 sg13g2_fill_8 FILLER_137_64 ();
 sg13g2_fill_8 FILLER_137_72 ();
 sg13g2_fill_8 FILLER_137_80 ();
 sg13g2_fill_8 FILLER_137_88 ();
 sg13g2_fill_8 FILLER_137_96 ();
 sg13g2_fill_8 FILLER_137_104 ();
 sg13g2_fill_8 FILLER_137_112 ();
 sg13g2_fill_8 FILLER_137_120 ();
 sg13g2_fill_8 FILLER_137_128 ();
 sg13g2_fill_8 FILLER_137_136 ();
 sg13g2_fill_8 FILLER_137_144 ();
 sg13g2_fill_8 FILLER_137_152 ();
 sg13g2_fill_8 FILLER_137_160 ();
 sg13g2_fill_8 FILLER_137_168 ();
 sg13g2_fill_8 FILLER_137_176 ();
 sg13g2_fill_8 FILLER_137_184 ();
 sg13g2_fill_8 FILLER_137_192 ();
 sg13g2_fill_8 FILLER_137_200 ();
 sg13g2_fill_8 FILLER_137_208 ();
 sg13g2_fill_8 FILLER_137_216 ();
 sg13g2_fill_8 FILLER_137_224 ();
 sg13g2_fill_8 FILLER_137_232 ();
 sg13g2_fill_8 FILLER_137_240 ();
 sg13g2_fill_8 FILLER_137_248 ();
 sg13g2_fill_8 FILLER_137_256 ();
 sg13g2_fill_8 FILLER_137_264 ();
 sg13g2_fill_8 FILLER_137_272 ();
 sg13g2_fill_8 FILLER_137_280 ();
 sg13g2_fill_8 FILLER_137_288 ();
 sg13g2_fill_8 FILLER_137_296 ();
 sg13g2_fill_8 FILLER_137_304 ();
 sg13g2_fill_8 FILLER_137_312 ();
 sg13g2_fill_8 FILLER_137_320 ();
 sg13g2_fill_8 FILLER_137_328 ();
 sg13g2_fill_8 FILLER_137_336 ();
 sg13g2_fill_8 FILLER_137_344 ();
 sg13g2_fill_8 FILLER_137_352 ();
 sg13g2_fill_8 FILLER_137_360 ();
 sg13g2_fill_8 FILLER_137_368 ();
 sg13g2_fill_8 FILLER_137_376 ();
 sg13g2_fill_8 FILLER_137_384 ();
 sg13g2_fill_8 FILLER_137_392 ();
 sg13g2_fill_8 FILLER_137_400 ();
 sg13g2_fill_8 FILLER_137_408 ();
 sg13g2_fill_8 FILLER_137_416 ();
 sg13g2_fill_8 FILLER_137_424 ();
 sg13g2_fill_8 FILLER_137_432 ();
 sg13g2_fill_8 FILLER_137_440 ();
 sg13g2_fill_8 FILLER_137_448 ();
 sg13g2_fill_8 FILLER_137_456 ();
 sg13g2_fill_8 FILLER_137_464 ();
 sg13g2_fill_8 FILLER_137_472 ();
 sg13g2_fill_8 FILLER_137_480 ();
 sg13g2_fill_8 FILLER_137_488 ();
 sg13g2_fill_8 FILLER_137_496 ();
 sg13g2_fill_8 FILLER_137_504 ();
 sg13g2_fill_8 FILLER_137_512 ();
 sg13g2_fill_8 FILLER_137_520 ();
 sg13g2_fill_8 FILLER_137_528 ();
 sg13g2_fill_8 FILLER_137_536 ();
 sg13g2_fill_8 FILLER_137_544 ();
 sg13g2_fill_8 FILLER_137_552 ();
 sg13g2_fill_8 FILLER_137_560 ();
 sg13g2_fill_8 FILLER_137_568 ();
 sg13g2_fill_8 FILLER_137_576 ();
 sg13g2_fill_8 FILLER_137_584 ();
 sg13g2_fill_8 FILLER_137_592 ();
 sg13g2_fill_8 FILLER_137_600 ();
 sg13g2_fill_8 FILLER_137_608 ();
 sg13g2_fill_8 FILLER_137_616 ();
 sg13g2_fill_8 FILLER_137_624 ();
 sg13g2_fill_8 FILLER_137_632 ();
 sg13g2_fill_8 FILLER_137_640 ();
 sg13g2_fill_8 FILLER_137_648 ();
 sg13g2_fill_8 FILLER_137_656 ();
 sg13g2_fill_8 FILLER_137_664 ();
 sg13g2_fill_8 FILLER_137_672 ();
 sg13g2_fill_8 FILLER_137_680 ();
 sg13g2_fill_8 FILLER_137_688 ();
 sg13g2_fill_8 FILLER_137_696 ();
 sg13g2_fill_8 FILLER_137_704 ();
 sg13g2_fill_8 FILLER_137_712 ();
 sg13g2_fill_8 FILLER_137_720 ();
 sg13g2_fill_8 FILLER_137_728 ();
 sg13g2_fill_8 FILLER_137_736 ();
 sg13g2_fill_8 FILLER_137_744 ();
 sg13g2_fill_8 FILLER_137_752 ();
 sg13g2_fill_8 FILLER_137_760 ();
 sg13g2_fill_8 FILLER_137_768 ();
 sg13g2_fill_8 FILLER_137_776 ();
 sg13g2_fill_8 FILLER_137_784 ();
 sg13g2_fill_8 FILLER_137_792 ();
 sg13g2_fill_8 FILLER_137_800 ();
 sg13g2_fill_8 FILLER_137_808 ();
 sg13g2_fill_8 FILLER_137_816 ();
 sg13g2_fill_8 FILLER_137_824 ();
 sg13g2_fill_8 FILLER_137_832 ();
 sg13g2_fill_8 FILLER_137_840 ();
 sg13g2_fill_8 FILLER_137_848 ();
 sg13g2_fill_8 FILLER_137_856 ();
 sg13g2_fill_8 FILLER_137_864 ();
 sg13g2_fill_8 FILLER_137_872 ();
 sg13g2_fill_8 FILLER_137_880 ();
 sg13g2_fill_8 FILLER_137_888 ();
 sg13g2_fill_8 FILLER_137_896 ();
 sg13g2_fill_8 FILLER_137_904 ();
 sg13g2_fill_8 FILLER_137_912 ();
 sg13g2_fill_8 FILLER_137_920 ();
 sg13g2_fill_8 FILLER_137_928 ();
 sg13g2_fill_8 FILLER_137_936 ();
 sg13g2_fill_8 FILLER_137_944 ();
 sg13g2_fill_8 FILLER_137_952 ();
 sg13g2_fill_8 FILLER_137_960 ();
 sg13g2_fill_8 FILLER_137_968 ();
 sg13g2_fill_8 FILLER_137_976 ();
 sg13g2_fill_8 FILLER_137_984 ();
 sg13g2_fill_8 FILLER_137_992 ();
 sg13g2_fill_8 FILLER_137_1000 ();
 sg13g2_fill_8 FILLER_137_1008 ();
 sg13g2_fill_8 FILLER_137_1016 ();
 sg13g2_fill_8 FILLER_137_1024 ();
 sg13g2_fill_8 FILLER_137_1032 ();
 sg13g2_fill_8 FILLER_137_1040 ();
 sg13g2_fill_8 FILLER_137_1048 ();
 sg13g2_fill_8 FILLER_137_1056 ();
 sg13g2_fill_8 FILLER_137_1064 ();
 sg13g2_fill_8 FILLER_137_1072 ();
 sg13g2_fill_8 FILLER_137_1080 ();
 sg13g2_fill_8 FILLER_137_1088 ();
 sg13g2_fill_8 FILLER_137_1096 ();
 sg13g2_fill_8 FILLER_137_1104 ();
 sg13g2_fill_8 FILLER_137_1112 ();
 sg13g2_fill_8 FILLER_137_1120 ();
 sg13g2_fill_8 FILLER_137_1128 ();
 sg13g2_fill_8 FILLER_137_1136 ();
 sg13g2_fill_8 FILLER_138_0 ();
 sg13g2_fill_8 FILLER_138_8 ();
 sg13g2_fill_8 FILLER_138_16 ();
 sg13g2_fill_8 FILLER_138_24 ();
 sg13g2_fill_8 FILLER_138_32 ();
 sg13g2_fill_8 FILLER_138_40 ();
 sg13g2_fill_8 FILLER_138_48 ();
 sg13g2_fill_8 FILLER_138_56 ();
 sg13g2_fill_8 FILLER_138_64 ();
 sg13g2_fill_8 FILLER_138_72 ();
 sg13g2_fill_8 FILLER_138_80 ();
 sg13g2_fill_8 FILLER_138_88 ();
 sg13g2_fill_8 FILLER_138_96 ();
 sg13g2_fill_8 FILLER_138_104 ();
 sg13g2_fill_8 FILLER_138_112 ();
 sg13g2_fill_8 FILLER_138_120 ();
 sg13g2_fill_8 FILLER_138_128 ();
 sg13g2_fill_8 FILLER_138_136 ();
 sg13g2_fill_8 FILLER_138_144 ();
 sg13g2_fill_8 FILLER_138_152 ();
 sg13g2_fill_8 FILLER_138_160 ();
 sg13g2_fill_8 FILLER_138_168 ();
 sg13g2_fill_8 FILLER_138_176 ();
 sg13g2_fill_8 FILLER_138_184 ();
 sg13g2_fill_8 FILLER_138_192 ();
 sg13g2_fill_8 FILLER_138_200 ();
 sg13g2_fill_8 FILLER_138_208 ();
 sg13g2_fill_8 FILLER_138_216 ();
 sg13g2_fill_8 FILLER_138_224 ();
 sg13g2_fill_8 FILLER_138_232 ();
 sg13g2_fill_8 FILLER_138_240 ();
 sg13g2_fill_8 FILLER_138_248 ();
 sg13g2_fill_8 FILLER_138_256 ();
 sg13g2_fill_8 FILLER_138_264 ();
 sg13g2_fill_8 FILLER_138_272 ();
 sg13g2_fill_8 FILLER_138_280 ();
 sg13g2_fill_8 FILLER_138_288 ();
 sg13g2_fill_8 FILLER_138_296 ();
 sg13g2_fill_8 FILLER_138_304 ();
 sg13g2_fill_8 FILLER_138_312 ();
 sg13g2_fill_8 FILLER_138_320 ();
 sg13g2_fill_8 FILLER_138_328 ();
 sg13g2_fill_8 FILLER_138_336 ();
 sg13g2_fill_8 FILLER_138_344 ();
 sg13g2_fill_8 FILLER_138_352 ();
 sg13g2_fill_8 FILLER_138_360 ();
 sg13g2_fill_8 FILLER_138_368 ();
 sg13g2_fill_8 FILLER_138_376 ();
 sg13g2_fill_8 FILLER_138_384 ();
 sg13g2_fill_8 FILLER_138_392 ();
 sg13g2_fill_8 FILLER_138_400 ();
 sg13g2_fill_8 FILLER_138_408 ();
 sg13g2_fill_8 FILLER_138_416 ();
 sg13g2_fill_8 FILLER_138_424 ();
 sg13g2_fill_8 FILLER_138_432 ();
 sg13g2_fill_8 FILLER_138_440 ();
 sg13g2_fill_8 FILLER_138_448 ();
 sg13g2_fill_8 FILLER_138_456 ();
 sg13g2_fill_8 FILLER_138_464 ();
 sg13g2_fill_8 FILLER_138_472 ();
 sg13g2_fill_8 FILLER_138_480 ();
 sg13g2_fill_8 FILLER_138_488 ();
 sg13g2_fill_8 FILLER_138_496 ();
 sg13g2_fill_8 FILLER_138_504 ();
 sg13g2_fill_8 FILLER_138_512 ();
 sg13g2_fill_8 FILLER_138_520 ();
 sg13g2_fill_8 FILLER_138_528 ();
 sg13g2_fill_8 FILLER_138_536 ();
 sg13g2_fill_8 FILLER_138_544 ();
 sg13g2_fill_8 FILLER_138_552 ();
 sg13g2_fill_8 FILLER_138_560 ();
 sg13g2_fill_8 FILLER_138_568 ();
 sg13g2_fill_8 FILLER_138_576 ();
 sg13g2_fill_8 FILLER_138_584 ();
 sg13g2_fill_8 FILLER_138_592 ();
 sg13g2_fill_8 FILLER_138_600 ();
 sg13g2_fill_8 FILLER_138_608 ();
 sg13g2_fill_8 FILLER_138_616 ();
 sg13g2_fill_8 FILLER_138_624 ();
 sg13g2_fill_8 FILLER_138_632 ();
 sg13g2_fill_8 FILLER_138_640 ();
 sg13g2_fill_8 FILLER_138_648 ();
 sg13g2_fill_8 FILLER_138_656 ();
 sg13g2_fill_8 FILLER_138_664 ();
 sg13g2_fill_8 FILLER_138_672 ();
 sg13g2_fill_8 FILLER_138_680 ();
 sg13g2_fill_8 FILLER_138_688 ();
 sg13g2_fill_8 FILLER_138_696 ();
 sg13g2_fill_8 FILLER_138_704 ();
 sg13g2_fill_8 FILLER_138_712 ();
 sg13g2_fill_8 FILLER_138_720 ();
 sg13g2_fill_8 FILLER_138_728 ();
 sg13g2_fill_8 FILLER_138_736 ();
 sg13g2_fill_8 FILLER_138_744 ();
 sg13g2_fill_8 FILLER_138_752 ();
 sg13g2_fill_8 FILLER_138_760 ();
 sg13g2_fill_8 FILLER_138_768 ();
 sg13g2_fill_8 FILLER_138_776 ();
 sg13g2_fill_8 FILLER_138_784 ();
 sg13g2_fill_8 FILLER_138_792 ();
 sg13g2_fill_8 FILLER_138_800 ();
 sg13g2_fill_8 FILLER_138_808 ();
 sg13g2_fill_8 FILLER_138_816 ();
 sg13g2_fill_8 FILLER_138_824 ();
 sg13g2_fill_8 FILLER_138_832 ();
 sg13g2_fill_8 FILLER_138_840 ();
 sg13g2_fill_8 FILLER_138_848 ();
 sg13g2_fill_8 FILLER_138_856 ();
 sg13g2_fill_8 FILLER_138_864 ();
 sg13g2_fill_8 FILLER_138_872 ();
 sg13g2_fill_8 FILLER_138_880 ();
 sg13g2_fill_8 FILLER_138_888 ();
 sg13g2_fill_8 FILLER_138_896 ();
 sg13g2_fill_8 FILLER_138_904 ();
 sg13g2_fill_8 FILLER_138_912 ();
 sg13g2_fill_8 FILLER_138_920 ();
 sg13g2_fill_8 FILLER_138_928 ();
 sg13g2_fill_8 FILLER_138_936 ();
 sg13g2_fill_8 FILLER_138_944 ();
 sg13g2_fill_8 FILLER_138_952 ();
 sg13g2_fill_8 FILLER_138_960 ();
 sg13g2_fill_8 FILLER_138_968 ();
 sg13g2_fill_8 FILLER_138_976 ();
 sg13g2_fill_8 FILLER_138_984 ();
 sg13g2_fill_8 FILLER_138_992 ();
 sg13g2_fill_8 FILLER_138_1000 ();
 sg13g2_fill_8 FILLER_138_1008 ();
 sg13g2_fill_8 FILLER_138_1016 ();
 sg13g2_fill_8 FILLER_138_1024 ();
 sg13g2_fill_8 FILLER_138_1032 ();
 sg13g2_fill_8 FILLER_138_1040 ();
 sg13g2_fill_8 FILLER_138_1048 ();
 sg13g2_fill_8 FILLER_138_1056 ();
 sg13g2_fill_8 FILLER_138_1064 ();
 sg13g2_fill_8 FILLER_138_1072 ();
 sg13g2_fill_8 FILLER_138_1080 ();
 sg13g2_fill_8 FILLER_138_1088 ();
 sg13g2_fill_8 FILLER_138_1096 ();
 sg13g2_fill_8 FILLER_138_1104 ();
 sg13g2_fill_8 FILLER_138_1112 ();
 sg13g2_fill_8 FILLER_138_1120 ();
 sg13g2_fill_8 FILLER_138_1128 ();
 sg13g2_fill_8 FILLER_138_1136 ();
 sg13g2_fill_8 FILLER_139_0 ();
 sg13g2_fill_8 FILLER_139_8 ();
 sg13g2_fill_8 FILLER_139_16 ();
 sg13g2_fill_8 FILLER_139_24 ();
 sg13g2_fill_8 FILLER_139_32 ();
 sg13g2_fill_8 FILLER_139_40 ();
 sg13g2_fill_8 FILLER_139_48 ();
 sg13g2_fill_8 FILLER_139_56 ();
 sg13g2_fill_8 FILLER_139_64 ();
 sg13g2_fill_8 FILLER_139_72 ();
 sg13g2_fill_8 FILLER_139_80 ();
 sg13g2_fill_8 FILLER_139_88 ();
 sg13g2_fill_8 FILLER_139_96 ();
 sg13g2_fill_8 FILLER_139_104 ();
 sg13g2_fill_8 FILLER_139_112 ();
 sg13g2_fill_8 FILLER_139_120 ();
 sg13g2_fill_8 FILLER_139_128 ();
 sg13g2_fill_8 FILLER_139_136 ();
 sg13g2_fill_8 FILLER_139_144 ();
 sg13g2_fill_8 FILLER_139_152 ();
 sg13g2_fill_8 FILLER_139_160 ();
 sg13g2_fill_8 FILLER_139_168 ();
 sg13g2_fill_8 FILLER_139_176 ();
 sg13g2_fill_8 FILLER_139_184 ();
 sg13g2_fill_8 FILLER_139_192 ();
 sg13g2_fill_8 FILLER_139_200 ();
 sg13g2_fill_8 FILLER_139_208 ();
 sg13g2_fill_8 FILLER_139_216 ();
 sg13g2_fill_8 FILLER_139_224 ();
 sg13g2_fill_8 FILLER_139_232 ();
 sg13g2_fill_8 FILLER_139_240 ();
 sg13g2_fill_8 FILLER_139_248 ();
 sg13g2_fill_8 FILLER_139_256 ();
 sg13g2_fill_8 FILLER_139_264 ();
 sg13g2_fill_8 FILLER_139_272 ();
 sg13g2_fill_8 FILLER_139_280 ();
 sg13g2_fill_8 FILLER_139_288 ();
 sg13g2_fill_8 FILLER_139_296 ();
 sg13g2_fill_8 FILLER_139_304 ();
 sg13g2_fill_8 FILLER_139_312 ();
 sg13g2_fill_8 FILLER_139_320 ();
 sg13g2_fill_8 FILLER_139_328 ();
 sg13g2_fill_8 FILLER_139_336 ();
 sg13g2_fill_8 FILLER_139_344 ();
 sg13g2_fill_8 FILLER_139_352 ();
 sg13g2_fill_8 FILLER_139_360 ();
 sg13g2_fill_8 FILLER_139_368 ();
 sg13g2_fill_8 FILLER_139_376 ();
 sg13g2_fill_8 FILLER_139_384 ();
 sg13g2_fill_8 FILLER_139_392 ();
 sg13g2_fill_8 FILLER_139_400 ();
 sg13g2_fill_8 FILLER_139_408 ();
 sg13g2_fill_8 FILLER_139_416 ();
 sg13g2_fill_8 FILLER_139_424 ();
 sg13g2_fill_8 FILLER_139_432 ();
 sg13g2_fill_8 FILLER_139_440 ();
 sg13g2_fill_8 FILLER_139_448 ();
 sg13g2_fill_8 FILLER_139_456 ();
 sg13g2_fill_8 FILLER_139_464 ();
 sg13g2_fill_8 FILLER_139_472 ();
 sg13g2_fill_8 FILLER_139_480 ();
 sg13g2_fill_8 FILLER_139_488 ();
 sg13g2_fill_8 FILLER_139_496 ();
 sg13g2_fill_8 FILLER_139_504 ();
 sg13g2_fill_8 FILLER_139_512 ();
 sg13g2_fill_8 FILLER_139_520 ();
 sg13g2_fill_8 FILLER_139_528 ();
 sg13g2_fill_8 FILLER_139_536 ();
 sg13g2_fill_8 FILLER_139_544 ();
 sg13g2_fill_8 FILLER_139_552 ();
 sg13g2_fill_8 FILLER_139_560 ();
 sg13g2_fill_8 FILLER_139_568 ();
 sg13g2_fill_8 FILLER_139_576 ();
 sg13g2_fill_8 FILLER_139_584 ();
 sg13g2_fill_8 FILLER_139_592 ();
 sg13g2_fill_8 FILLER_139_600 ();
 sg13g2_fill_8 FILLER_139_608 ();
 sg13g2_fill_8 FILLER_139_616 ();
 sg13g2_fill_8 FILLER_139_624 ();
 sg13g2_fill_8 FILLER_139_632 ();
 sg13g2_fill_8 FILLER_139_640 ();
 sg13g2_fill_8 FILLER_139_648 ();
 sg13g2_fill_8 FILLER_139_656 ();
 sg13g2_fill_8 FILLER_139_664 ();
 sg13g2_fill_8 FILLER_139_672 ();
 sg13g2_fill_8 FILLER_139_680 ();
 sg13g2_fill_8 FILLER_139_688 ();
 sg13g2_fill_8 FILLER_139_696 ();
 sg13g2_fill_8 FILLER_139_704 ();
 sg13g2_fill_8 FILLER_139_712 ();
 sg13g2_fill_8 FILLER_139_720 ();
 sg13g2_fill_8 FILLER_139_728 ();
 sg13g2_fill_8 FILLER_139_736 ();
 sg13g2_fill_8 FILLER_139_744 ();
 sg13g2_fill_8 FILLER_139_752 ();
 sg13g2_fill_8 FILLER_139_760 ();
 sg13g2_fill_8 FILLER_139_768 ();
 sg13g2_fill_8 FILLER_139_776 ();
 sg13g2_fill_8 FILLER_139_784 ();
 sg13g2_fill_8 FILLER_139_792 ();
 sg13g2_fill_8 FILLER_139_800 ();
 sg13g2_fill_8 FILLER_139_808 ();
 sg13g2_fill_8 FILLER_139_816 ();
 sg13g2_fill_8 FILLER_139_824 ();
 sg13g2_fill_8 FILLER_139_832 ();
 sg13g2_fill_8 FILLER_139_840 ();
 sg13g2_fill_8 FILLER_139_848 ();
 sg13g2_fill_8 FILLER_139_856 ();
 sg13g2_fill_8 FILLER_139_864 ();
 sg13g2_fill_8 FILLER_139_872 ();
 sg13g2_fill_8 FILLER_139_880 ();
 sg13g2_fill_8 FILLER_139_888 ();
 sg13g2_fill_8 FILLER_139_896 ();
 sg13g2_fill_8 FILLER_139_904 ();
 sg13g2_fill_8 FILLER_139_912 ();
 sg13g2_fill_8 FILLER_139_920 ();
 sg13g2_fill_8 FILLER_139_928 ();
 sg13g2_fill_8 FILLER_139_936 ();
 sg13g2_fill_8 FILLER_139_944 ();
 sg13g2_fill_8 FILLER_139_952 ();
 sg13g2_fill_8 FILLER_139_960 ();
 sg13g2_fill_8 FILLER_139_968 ();
 sg13g2_fill_8 FILLER_139_976 ();
 sg13g2_fill_8 FILLER_139_984 ();
 sg13g2_fill_8 FILLER_139_992 ();
 sg13g2_fill_8 FILLER_139_1000 ();
 sg13g2_fill_8 FILLER_139_1008 ();
 sg13g2_fill_8 FILLER_139_1016 ();
 sg13g2_fill_8 FILLER_139_1024 ();
 sg13g2_fill_8 FILLER_139_1032 ();
 sg13g2_fill_8 FILLER_139_1040 ();
 sg13g2_fill_8 FILLER_139_1048 ();
 sg13g2_fill_8 FILLER_139_1056 ();
 sg13g2_fill_8 FILLER_139_1064 ();
 sg13g2_fill_8 FILLER_139_1072 ();
 sg13g2_fill_8 FILLER_139_1080 ();
 sg13g2_fill_8 FILLER_139_1088 ();
 sg13g2_fill_8 FILLER_139_1096 ();
 sg13g2_fill_8 FILLER_139_1104 ();
 sg13g2_fill_8 FILLER_139_1112 ();
 sg13g2_fill_8 FILLER_139_1120 ();
 sg13g2_fill_8 FILLER_139_1128 ();
 sg13g2_fill_8 FILLER_139_1136 ();
 sg13g2_fill_8 FILLER_140_0 ();
 sg13g2_fill_8 FILLER_140_8 ();
 sg13g2_fill_8 FILLER_140_16 ();
 sg13g2_fill_8 FILLER_140_24 ();
 sg13g2_fill_8 FILLER_140_32 ();
 sg13g2_fill_8 FILLER_140_40 ();
 sg13g2_fill_8 FILLER_140_48 ();
 sg13g2_fill_8 FILLER_140_56 ();
 sg13g2_fill_8 FILLER_140_64 ();
 sg13g2_fill_8 FILLER_140_72 ();
 sg13g2_fill_8 FILLER_140_80 ();
 sg13g2_fill_8 FILLER_140_88 ();
 sg13g2_fill_8 FILLER_140_96 ();
 sg13g2_fill_8 FILLER_140_104 ();
 sg13g2_fill_8 FILLER_140_112 ();
 sg13g2_fill_8 FILLER_140_120 ();
 sg13g2_fill_8 FILLER_140_128 ();
 sg13g2_fill_8 FILLER_140_136 ();
 sg13g2_fill_8 FILLER_140_144 ();
 sg13g2_fill_8 FILLER_140_152 ();
 sg13g2_fill_8 FILLER_140_160 ();
 sg13g2_fill_8 FILLER_140_168 ();
 sg13g2_fill_8 FILLER_140_176 ();
 sg13g2_fill_8 FILLER_140_184 ();
 sg13g2_fill_8 FILLER_140_192 ();
 sg13g2_fill_8 FILLER_140_200 ();
 sg13g2_fill_8 FILLER_140_208 ();
 sg13g2_fill_8 FILLER_140_216 ();
 sg13g2_fill_8 FILLER_140_224 ();
 sg13g2_fill_8 FILLER_140_232 ();
 sg13g2_fill_8 FILLER_140_240 ();
 sg13g2_fill_8 FILLER_140_248 ();
 sg13g2_fill_8 FILLER_140_256 ();
 sg13g2_fill_8 FILLER_140_264 ();
 sg13g2_fill_8 FILLER_140_272 ();
 sg13g2_fill_8 FILLER_140_280 ();
 sg13g2_fill_8 FILLER_140_288 ();
 sg13g2_fill_8 FILLER_140_296 ();
 sg13g2_fill_8 FILLER_140_304 ();
 sg13g2_fill_8 FILLER_140_312 ();
 sg13g2_fill_8 FILLER_140_320 ();
 sg13g2_fill_8 FILLER_140_328 ();
 sg13g2_fill_8 FILLER_140_336 ();
 sg13g2_fill_8 FILLER_140_344 ();
 sg13g2_fill_8 FILLER_140_352 ();
 sg13g2_fill_8 FILLER_140_360 ();
 sg13g2_fill_8 FILLER_140_368 ();
 sg13g2_fill_8 FILLER_140_376 ();
 sg13g2_fill_8 FILLER_140_384 ();
 sg13g2_fill_8 FILLER_140_392 ();
 sg13g2_fill_8 FILLER_140_400 ();
 sg13g2_fill_8 FILLER_140_408 ();
 sg13g2_fill_8 FILLER_140_416 ();
 sg13g2_fill_8 FILLER_140_424 ();
 sg13g2_fill_8 FILLER_140_432 ();
 sg13g2_fill_8 FILLER_140_440 ();
 sg13g2_fill_8 FILLER_140_448 ();
 sg13g2_fill_8 FILLER_140_456 ();
 sg13g2_fill_8 FILLER_140_464 ();
 sg13g2_fill_8 FILLER_140_472 ();
 sg13g2_fill_8 FILLER_140_480 ();
 sg13g2_fill_8 FILLER_140_488 ();
 sg13g2_fill_8 FILLER_140_496 ();
 sg13g2_fill_8 FILLER_140_504 ();
 sg13g2_fill_8 FILLER_140_512 ();
 sg13g2_fill_8 FILLER_140_520 ();
 sg13g2_fill_8 FILLER_140_528 ();
 sg13g2_fill_8 FILLER_140_536 ();
 sg13g2_fill_8 FILLER_140_544 ();
 sg13g2_fill_8 FILLER_140_552 ();
 sg13g2_fill_8 FILLER_140_560 ();
 sg13g2_fill_8 FILLER_140_568 ();
 sg13g2_fill_8 FILLER_140_576 ();
 sg13g2_fill_8 FILLER_140_584 ();
 sg13g2_fill_8 FILLER_140_592 ();
 sg13g2_fill_8 FILLER_140_600 ();
 sg13g2_fill_8 FILLER_140_608 ();
 sg13g2_fill_8 FILLER_140_616 ();
 sg13g2_fill_8 FILLER_140_624 ();
 sg13g2_fill_8 FILLER_140_632 ();
 sg13g2_fill_8 FILLER_140_640 ();
 sg13g2_fill_8 FILLER_140_648 ();
 sg13g2_fill_8 FILLER_140_656 ();
 sg13g2_fill_8 FILLER_140_664 ();
 sg13g2_fill_8 FILLER_140_672 ();
 sg13g2_fill_8 FILLER_140_680 ();
 sg13g2_fill_8 FILLER_140_688 ();
 sg13g2_fill_8 FILLER_140_696 ();
 sg13g2_fill_8 FILLER_140_704 ();
 sg13g2_fill_8 FILLER_140_712 ();
 sg13g2_fill_8 FILLER_140_720 ();
 sg13g2_fill_8 FILLER_140_728 ();
 sg13g2_fill_8 FILLER_140_736 ();
 sg13g2_fill_8 FILLER_140_744 ();
 sg13g2_fill_8 FILLER_140_752 ();
 sg13g2_fill_8 FILLER_140_760 ();
 sg13g2_fill_8 FILLER_140_768 ();
 sg13g2_fill_8 FILLER_140_776 ();
 sg13g2_fill_8 FILLER_140_784 ();
 sg13g2_fill_8 FILLER_140_792 ();
 sg13g2_fill_8 FILLER_140_800 ();
 sg13g2_fill_8 FILLER_140_808 ();
 sg13g2_fill_8 FILLER_140_816 ();
 sg13g2_fill_8 FILLER_140_824 ();
 sg13g2_fill_8 FILLER_140_832 ();
 sg13g2_fill_8 FILLER_140_840 ();
 sg13g2_fill_8 FILLER_140_848 ();
 sg13g2_fill_8 FILLER_140_856 ();
 sg13g2_fill_8 FILLER_140_864 ();
 sg13g2_fill_8 FILLER_140_872 ();
 sg13g2_fill_8 FILLER_140_880 ();
 sg13g2_fill_8 FILLER_140_888 ();
 sg13g2_fill_8 FILLER_140_896 ();
 sg13g2_fill_8 FILLER_140_904 ();
 sg13g2_fill_8 FILLER_140_912 ();
 sg13g2_fill_8 FILLER_140_920 ();
 sg13g2_fill_8 FILLER_140_928 ();
 sg13g2_fill_8 FILLER_140_936 ();
 sg13g2_fill_8 FILLER_140_944 ();
 sg13g2_fill_8 FILLER_140_952 ();
 sg13g2_fill_8 FILLER_140_960 ();
 sg13g2_fill_8 FILLER_140_968 ();
 sg13g2_fill_8 FILLER_140_976 ();
 sg13g2_fill_8 FILLER_140_984 ();
 sg13g2_fill_8 FILLER_140_992 ();
 sg13g2_fill_8 FILLER_140_1000 ();
 sg13g2_fill_8 FILLER_140_1008 ();
 sg13g2_fill_8 FILLER_140_1016 ();
 sg13g2_fill_8 FILLER_140_1024 ();
 sg13g2_fill_8 FILLER_140_1032 ();
 sg13g2_fill_8 FILLER_140_1040 ();
 sg13g2_fill_8 FILLER_140_1048 ();
 sg13g2_fill_8 FILLER_140_1056 ();
 sg13g2_fill_8 FILLER_140_1064 ();
 sg13g2_fill_8 FILLER_140_1072 ();
 sg13g2_fill_8 FILLER_140_1080 ();
 sg13g2_fill_8 FILLER_140_1088 ();
 sg13g2_fill_8 FILLER_140_1096 ();
 sg13g2_fill_8 FILLER_140_1104 ();
 sg13g2_fill_8 FILLER_140_1112 ();
 sg13g2_fill_8 FILLER_140_1120 ();
 sg13g2_fill_8 FILLER_140_1128 ();
 sg13g2_fill_8 FILLER_140_1136 ();
 sg13g2_fill_8 FILLER_141_0 ();
 sg13g2_fill_8 FILLER_141_8 ();
 sg13g2_fill_8 FILLER_141_16 ();
 sg13g2_fill_8 FILLER_141_24 ();
 sg13g2_fill_8 FILLER_141_32 ();
 sg13g2_fill_8 FILLER_141_40 ();
 sg13g2_fill_8 FILLER_141_48 ();
 sg13g2_fill_8 FILLER_141_56 ();
 sg13g2_fill_8 FILLER_141_64 ();
 sg13g2_fill_8 FILLER_141_72 ();
 sg13g2_fill_8 FILLER_141_80 ();
 sg13g2_fill_8 FILLER_141_88 ();
 sg13g2_fill_8 FILLER_141_96 ();
 sg13g2_fill_8 FILLER_141_104 ();
 sg13g2_fill_8 FILLER_141_112 ();
 sg13g2_fill_8 FILLER_141_120 ();
 sg13g2_fill_8 FILLER_141_128 ();
 sg13g2_fill_8 FILLER_141_136 ();
 sg13g2_fill_8 FILLER_141_144 ();
 sg13g2_fill_8 FILLER_141_152 ();
 sg13g2_fill_8 FILLER_141_160 ();
 sg13g2_fill_8 FILLER_141_168 ();
 sg13g2_fill_8 FILLER_141_176 ();
 sg13g2_fill_8 FILLER_141_184 ();
 sg13g2_fill_8 FILLER_141_192 ();
 sg13g2_fill_8 FILLER_141_200 ();
 sg13g2_fill_8 FILLER_141_208 ();
 sg13g2_fill_8 FILLER_141_216 ();
 sg13g2_fill_8 FILLER_141_224 ();
 sg13g2_fill_8 FILLER_141_232 ();
 sg13g2_fill_8 FILLER_141_240 ();
 sg13g2_fill_8 FILLER_141_248 ();
 sg13g2_fill_8 FILLER_141_256 ();
 sg13g2_fill_8 FILLER_141_264 ();
 sg13g2_fill_8 FILLER_141_272 ();
 sg13g2_fill_8 FILLER_141_280 ();
 sg13g2_fill_8 FILLER_141_288 ();
 sg13g2_fill_8 FILLER_141_296 ();
 sg13g2_fill_8 FILLER_141_304 ();
 sg13g2_fill_8 FILLER_141_312 ();
 sg13g2_fill_8 FILLER_141_320 ();
 sg13g2_fill_8 FILLER_141_328 ();
 sg13g2_fill_8 FILLER_141_336 ();
 sg13g2_fill_8 FILLER_141_344 ();
 sg13g2_fill_8 FILLER_141_352 ();
 sg13g2_fill_8 FILLER_141_360 ();
 sg13g2_fill_8 FILLER_141_368 ();
 sg13g2_fill_8 FILLER_141_376 ();
 sg13g2_fill_8 FILLER_141_384 ();
 sg13g2_fill_8 FILLER_141_392 ();
 sg13g2_fill_8 FILLER_141_400 ();
 sg13g2_fill_8 FILLER_141_408 ();
 sg13g2_fill_8 FILLER_141_416 ();
 sg13g2_fill_8 FILLER_141_424 ();
 sg13g2_fill_8 FILLER_141_432 ();
 sg13g2_fill_8 FILLER_141_440 ();
 sg13g2_fill_8 FILLER_141_448 ();
 sg13g2_fill_8 FILLER_141_456 ();
 sg13g2_fill_8 FILLER_141_464 ();
 sg13g2_fill_8 FILLER_141_472 ();
 sg13g2_fill_8 FILLER_141_480 ();
 sg13g2_fill_8 FILLER_141_488 ();
 sg13g2_fill_8 FILLER_141_496 ();
 sg13g2_fill_8 FILLER_141_504 ();
 sg13g2_fill_8 FILLER_141_512 ();
 sg13g2_fill_8 FILLER_141_520 ();
 sg13g2_fill_8 FILLER_141_528 ();
 sg13g2_fill_8 FILLER_141_536 ();
 sg13g2_fill_8 FILLER_141_544 ();
 sg13g2_fill_8 FILLER_141_552 ();
 sg13g2_fill_8 FILLER_141_560 ();
 sg13g2_fill_8 FILLER_141_568 ();
 sg13g2_fill_8 FILLER_141_576 ();
 sg13g2_fill_8 FILLER_141_584 ();
 sg13g2_fill_8 FILLER_141_592 ();
 sg13g2_fill_8 FILLER_141_600 ();
 sg13g2_fill_8 FILLER_141_608 ();
 sg13g2_fill_8 FILLER_141_616 ();
 sg13g2_fill_8 FILLER_141_624 ();
 sg13g2_fill_8 FILLER_141_632 ();
 sg13g2_fill_8 FILLER_141_640 ();
 sg13g2_fill_8 FILLER_141_648 ();
 sg13g2_fill_8 FILLER_141_656 ();
 sg13g2_fill_8 FILLER_141_664 ();
 sg13g2_fill_8 FILLER_141_672 ();
 sg13g2_fill_8 FILLER_141_680 ();
 sg13g2_fill_8 FILLER_141_688 ();
 sg13g2_fill_8 FILLER_141_696 ();
 sg13g2_fill_8 FILLER_141_704 ();
 sg13g2_fill_8 FILLER_141_712 ();
 sg13g2_fill_8 FILLER_141_720 ();
 sg13g2_fill_8 FILLER_141_728 ();
 sg13g2_fill_8 FILLER_141_736 ();
 sg13g2_fill_8 FILLER_141_744 ();
 sg13g2_fill_8 FILLER_141_752 ();
 sg13g2_fill_8 FILLER_141_760 ();
 sg13g2_fill_8 FILLER_141_768 ();
 sg13g2_fill_8 FILLER_141_776 ();
 sg13g2_fill_8 FILLER_141_784 ();
 sg13g2_fill_8 FILLER_141_792 ();
 sg13g2_fill_8 FILLER_141_800 ();
 sg13g2_fill_8 FILLER_141_808 ();
 sg13g2_fill_8 FILLER_141_816 ();
 sg13g2_fill_8 FILLER_141_824 ();
 sg13g2_fill_8 FILLER_141_832 ();
 sg13g2_fill_8 FILLER_141_840 ();
 sg13g2_fill_8 FILLER_141_848 ();
 sg13g2_fill_8 FILLER_141_856 ();
 sg13g2_fill_8 FILLER_141_864 ();
 sg13g2_fill_8 FILLER_141_872 ();
 sg13g2_fill_8 FILLER_141_880 ();
 sg13g2_fill_8 FILLER_141_888 ();
 sg13g2_fill_8 FILLER_141_896 ();
 sg13g2_fill_8 FILLER_141_904 ();
 sg13g2_fill_8 FILLER_141_912 ();
 sg13g2_fill_8 FILLER_141_920 ();
 sg13g2_fill_8 FILLER_141_928 ();
 sg13g2_fill_8 FILLER_141_936 ();
 sg13g2_fill_8 FILLER_141_944 ();
 sg13g2_fill_8 FILLER_141_952 ();
 sg13g2_fill_8 FILLER_141_960 ();
 sg13g2_fill_8 FILLER_141_968 ();
 sg13g2_fill_8 FILLER_141_976 ();
 sg13g2_fill_8 FILLER_141_984 ();
 sg13g2_fill_8 FILLER_141_992 ();
 sg13g2_fill_8 FILLER_141_1000 ();
 sg13g2_fill_8 FILLER_141_1008 ();
 sg13g2_fill_8 FILLER_141_1016 ();
 sg13g2_fill_8 FILLER_141_1024 ();
 sg13g2_fill_8 FILLER_141_1032 ();
 sg13g2_fill_8 FILLER_141_1040 ();
 sg13g2_fill_8 FILLER_141_1048 ();
 sg13g2_fill_8 FILLER_141_1056 ();
 sg13g2_fill_8 FILLER_141_1064 ();
 sg13g2_fill_8 FILLER_141_1072 ();
 sg13g2_fill_8 FILLER_141_1080 ();
 sg13g2_fill_8 FILLER_141_1088 ();
 sg13g2_fill_8 FILLER_141_1096 ();
 sg13g2_fill_8 FILLER_141_1104 ();
 sg13g2_fill_8 FILLER_141_1112 ();
 sg13g2_fill_8 FILLER_141_1120 ();
 sg13g2_fill_8 FILLER_141_1128 ();
 sg13g2_fill_8 FILLER_141_1136 ();
 sg13g2_fill_8 FILLER_142_0 ();
 sg13g2_fill_8 FILLER_142_8 ();
 sg13g2_fill_8 FILLER_142_16 ();
 sg13g2_fill_8 FILLER_142_24 ();
 sg13g2_fill_8 FILLER_142_32 ();
 sg13g2_fill_8 FILLER_142_40 ();
 sg13g2_fill_8 FILLER_142_48 ();
 sg13g2_fill_8 FILLER_142_56 ();
 sg13g2_fill_8 FILLER_142_64 ();
 sg13g2_fill_8 FILLER_142_72 ();
 sg13g2_fill_8 FILLER_142_80 ();
 sg13g2_fill_8 FILLER_142_88 ();
 sg13g2_fill_8 FILLER_142_96 ();
 sg13g2_fill_8 FILLER_142_104 ();
 sg13g2_fill_8 FILLER_142_112 ();
 sg13g2_fill_8 FILLER_142_120 ();
 sg13g2_fill_8 FILLER_142_128 ();
 sg13g2_fill_8 FILLER_142_136 ();
 sg13g2_fill_8 FILLER_142_144 ();
 sg13g2_fill_8 FILLER_142_152 ();
 sg13g2_fill_8 FILLER_142_160 ();
 sg13g2_fill_8 FILLER_142_168 ();
 sg13g2_fill_8 FILLER_142_176 ();
 sg13g2_fill_8 FILLER_142_184 ();
 sg13g2_fill_8 FILLER_142_192 ();
 sg13g2_fill_8 FILLER_142_200 ();
 sg13g2_fill_8 FILLER_142_208 ();
 sg13g2_fill_8 FILLER_142_216 ();
 sg13g2_fill_8 FILLER_142_224 ();
 sg13g2_fill_8 FILLER_142_232 ();
 sg13g2_fill_8 FILLER_142_240 ();
 sg13g2_fill_8 FILLER_142_248 ();
 sg13g2_fill_8 FILLER_142_256 ();
 sg13g2_fill_8 FILLER_142_264 ();
 sg13g2_fill_8 FILLER_142_272 ();
 sg13g2_fill_8 FILLER_142_280 ();
 sg13g2_fill_8 FILLER_142_288 ();
 sg13g2_fill_8 FILLER_142_296 ();
 sg13g2_fill_8 FILLER_142_304 ();
 sg13g2_fill_8 FILLER_142_312 ();
 sg13g2_fill_8 FILLER_142_320 ();
 sg13g2_fill_8 FILLER_142_328 ();
 sg13g2_fill_8 FILLER_142_336 ();
 sg13g2_fill_8 FILLER_142_344 ();
 sg13g2_fill_8 FILLER_142_352 ();
 sg13g2_fill_8 FILLER_142_360 ();
 sg13g2_fill_8 FILLER_142_368 ();
 sg13g2_fill_8 FILLER_142_376 ();
 sg13g2_fill_8 FILLER_142_384 ();
 sg13g2_fill_8 FILLER_142_392 ();
 sg13g2_fill_8 FILLER_142_400 ();
 sg13g2_fill_8 FILLER_142_408 ();
 sg13g2_fill_8 FILLER_142_416 ();
 sg13g2_fill_8 FILLER_142_424 ();
 sg13g2_fill_8 FILLER_142_432 ();
 sg13g2_fill_8 FILLER_142_440 ();
 sg13g2_fill_8 FILLER_142_448 ();
 sg13g2_fill_8 FILLER_142_456 ();
 sg13g2_fill_8 FILLER_142_464 ();
 sg13g2_fill_8 FILLER_142_472 ();
 sg13g2_fill_8 FILLER_142_480 ();
 sg13g2_fill_8 FILLER_142_488 ();
 sg13g2_fill_8 FILLER_142_496 ();
 sg13g2_fill_8 FILLER_142_504 ();
 sg13g2_fill_8 FILLER_142_512 ();
 sg13g2_fill_8 FILLER_142_520 ();
 sg13g2_fill_8 FILLER_142_528 ();
 sg13g2_fill_8 FILLER_142_536 ();
 sg13g2_fill_8 FILLER_142_544 ();
 sg13g2_fill_8 FILLER_142_552 ();
 sg13g2_fill_8 FILLER_142_560 ();
 sg13g2_fill_8 FILLER_142_568 ();
 sg13g2_fill_8 FILLER_142_576 ();
 sg13g2_fill_8 FILLER_142_584 ();
 sg13g2_fill_8 FILLER_142_592 ();
 sg13g2_fill_8 FILLER_142_600 ();
 sg13g2_fill_8 FILLER_142_608 ();
 sg13g2_fill_8 FILLER_142_616 ();
 sg13g2_fill_8 FILLER_142_624 ();
 sg13g2_fill_8 FILLER_142_632 ();
 sg13g2_fill_8 FILLER_142_640 ();
 sg13g2_fill_8 FILLER_142_648 ();
 sg13g2_fill_8 FILLER_142_656 ();
 sg13g2_fill_8 FILLER_142_664 ();
 sg13g2_fill_8 FILLER_142_672 ();
 sg13g2_fill_8 FILLER_142_680 ();
 sg13g2_fill_8 FILLER_142_688 ();
 sg13g2_fill_8 FILLER_142_696 ();
 sg13g2_fill_8 FILLER_142_704 ();
 sg13g2_fill_8 FILLER_142_712 ();
 sg13g2_fill_8 FILLER_142_720 ();
 sg13g2_fill_8 FILLER_142_728 ();
 sg13g2_fill_8 FILLER_142_736 ();
 sg13g2_fill_8 FILLER_142_744 ();
 sg13g2_fill_8 FILLER_142_752 ();
 sg13g2_fill_8 FILLER_142_760 ();
 sg13g2_fill_8 FILLER_142_768 ();
 sg13g2_fill_8 FILLER_142_776 ();
 sg13g2_fill_8 FILLER_142_784 ();
 sg13g2_fill_8 FILLER_142_792 ();
 sg13g2_fill_8 FILLER_142_800 ();
 sg13g2_fill_8 FILLER_142_808 ();
 sg13g2_fill_8 FILLER_142_816 ();
 sg13g2_fill_8 FILLER_142_824 ();
 sg13g2_fill_8 FILLER_142_832 ();
 sg13g2_fill_8 FILLER_142_840 ();
 sg13g2_fill_8 FILLER_142_848 ();
 sg13g2_fill_8 FILLER_142_856 ();
 sg13g2_fill_8 FILLER_142_864 ();
 sg13g2_fill_8 FILLER_142_872 ();
 sg13g2_fill_8 FILLER_142_880 ();
 sg13g2_fill_8 FILLER_142_888 ();
 sg13g2_fill_8 FILLER_142_896 ();
 sg13g2_fill_8 FILLER_142_904 ();
 sg13g2_fill_8 FILLER_142_912 ();
 sg13g2_fill_8 FILLER_142_920 ();
 sg13g2_fill_8 FILLER_142_928 ();
 sg13g2_fill_8 FILLER_142_936 ();
 sg13g2_fill_8 FILLER_142_944 ();
 sg13g2_fill_8 FILLER_142_952 ();
 sg13g2_fill_8 FILLER_142_960 ();
 sg13g2_fill_8 FILLER_142_968 ();
 sg13g2_fill_8 FILLER_142_976 ();
 sg13g2_fill_8 FILLER_142_984 ();
 sg13g2_fill_8 FILLER_142_992 ();
 sg13g2_fill_8 FILLER_142_1000 ();
 sg13g2_fill_8 FILLER_142_1008 ();
 sg13g2_fill_8 FILLER_142_1016 ();
 sg13g2_fill_8 FILLER_142_1024 ();
 sg13g2_fill_8 FILLER_142_1032 ();
 sg13g2_fill_8 FILLER_142_1040 ();
 sg13g2_fill_8 FILLER_142_1048 ();
 sg13g2_fill_8 FILLER_142_1056 ();
 sg13g2_fill_8 FILLER_142_1064 ();
 sg13g2_fill_8 FILLER_142_1072 ();
 sg13g2_fill_8 FILLER_142_1080 ();
 sg13g2_fill_8 FILLER_142_1088 ();
 sg13g2_fill_8 FILLER_142_1096 ();
 sg13g2_fill_8 FILLER_142_1104 ();
 sg13g2_fill_8 FILLER_142_1112 ();
 sg13g2_fill_8 FILLER_142_1120 ();
 sg13g2_fill_8 FILLER_142_1128 ();
 sg13g2_fill_8 FILLER_142_1136 ();
 sg13g2_fill_8 FILLER_143_0 ();
 sg13g2_fill_8 FILLER_143_8 ();
 sg13g2_fill_8 FILLER_143_16 ();
 sg13g2_fill_8 FILLER_143_24 ();
 sg13g2_fill_8 FILLER_143_32 ();
 sg13g2_fill_8 FILLER_143_40 ();
 sg13g2_fill_8 FILLER_143_48 ();
 sg13g2_fill_8 FILLER_143_56 ();
 sg13g2_fill_8 FILLER_143_64 ();
 sg13g2_fill_8 FILLER_143_72 ();
 sg13g2_fill_8 FILLER_143_80 ();
 sg13g2_fill_8 FILLER_143_88 ();
 sg13g2_fill_8 FILLER_143_96 ();
 sg13g2_fill_8 FILLER_143_104 ();
 sg13g2_fill_8 FILLER_143_112 ();
 sg13g2_fill_8 FILLER_143_120 ();
 sg13g2_fill_8 FILLER_143_128 ();
 sg13g2_fill_8 FILLER_143_136 ();
 sg13g2_fill_8 FILLER_143_144 ();
 sg13g2_fill_8 FILLER_143_152 ();
 sg13g2_fill_8 FILLER_143_160 ();
 sg13g2_fill_8 FILLER_143_168 ();
 sg13g2_fill_8 FILLER_143_176 ();
 sg13g2_fill_8 FILLER_143_184 ();
 sg13g2_fill_8 FILLER_143_192 ();
 sg13g2_fill_8 FILLER_143_200 ();
 sg13g2_fill_8 FILLER_143_208 ();
 sg13g2_fill_8 FILLER_143_216 ();
 sg13g2_fill_8 FILLER_143_224 ();
 sg13g2_fill_8 FILLER_143_232 ();
 sg13g2_fill_8 FILLER_143_240 ();
 sg13g2_fill_8 FILLER_143_248 ();
 sg13g2_fill_8 FILLER_143_256 ();
 sg13g2_fill_8 FILLER_143_264 ();
 sg13g2_fill_8 FILLER_143_272 ();
 sg13g2_fill_8 FILLER_143_280 ();
 sg13g2_fill_8 FILLER_143_288 ();
 sg13g2_fill_8 FILLER_143_296 ();
 sg13g2_fill_8 FILLER_143_304 ();
 sg13g2_fill_8 FILLER_143_312 ();
 sg13g2_fill_8 FILLER_143_320 ();
 sg13g2_fill_8 FILLER_143_328 ();
 sg13g2_fill_8 FILLER_143_336 ();
 sg13g2_fill_8 FILLER_143_344 ();
 sg13g2_fill_8 FILLER_143_352 ();
 sg13g2_fill_8 FILLER_143_360 ();
 sg13g2_fill_8 FILLER_143_368 ();
 sg13g2_fill_8 FILLER_143_376 ();
 sg13g2_fill_8 FILLER_143_384 ();
 sg13g2_fill_8 FILLER_143_392 ();
 sg13g2_fill_8 FILLER_143_400 ();
 sg13g2_fill_8 FILLER_143_408 ();
 sg13g2_fill_8 FILLER_143_416 ();
 sg13g2_fill_8 FILLER_143_424 ();
 sg13g2_fill_8 FILLER_143_432 ();
 sg13g2_fill_8 FILLER_143_440 ();
 sg13g2_fill_8 FILLER_143_448 ();
 sg13g2_fill_8 FILLER_143_456 ();
 sg13g2_fill_8 FILLER_143_464 ();
 sg13g2_fill_8 FILLER_143_472 ();
 sg13g2_fill_8 FILLER_143_480 ();
 sg13g2_fill_8 FILLER_143_488 ();
 sg13g2_fill_8 FILLER_143_496 ();
 sg13g2_fill_8 FILLER_143_504 ();
 sg13g2_fill_8 FILLER_143_512 ();
 sg13g2_fill_8 FILLER_143_520 ();
 sg13g2_fill_8 FILLER_143_528 ();
 sg13g2_fill_8 FILLER_143_536 ();
 sg13g2_fill_8 FILLER_143_544 ();
 sg13g2_fill_8 FILLER_143_552 ();
 sg13g2_fill_8 FILLER_143_560 ();
 sg13g2_fill_8 FILLER_143_568 ();
 sg13g2_fill_8 FILLER_143_576 ();
 sg13g2_fill_8 FILLER_143_584 ();
 sg13g2_fill_8 FILLER_143_592 ();
 sg13g2_fill_8 FILLER_143_600 ();
 sg13g2_fill_8 FILLER_143_608 ();
 sg13g2_fill_8 FILLER_143_616 ();
 sg13g2_fill_8 FILLER_143_624 ();
 sg13g2_fill_8 FILLER_143_632 ();
 sg13g2_fill_8 FILLER_143_640 ();
 sg13g2_fill_8 FILLER_143_648 ();
 sg13g2_fill_8 FILLER_143_656 ();
 sg13g2_fill_8 FILLER_143_664 ();
 sg13g2_fill_8 FILLER_143_672 ();
 sg13g2_fill_8 FILLER_143_680 ();
 sg13g2_fill_8 FILLER_143_688 ();
 sg13g2_fill_8 FILLER_143_696 ();
 sg13g2_fill_8 FILLER_143_704 ();
 sg13g2_fill_8 FILLER_143_712 ();
 sg13g2_fill_8 FILLER_143_720 ();
 sg13g2_fill_8 FILLER_143_728 ();
 sg13g2_fill_8 FILLER_143_736 ();
 sg13g2_fill_8 FILLER_143_744 ();
 sg13g2_fill_8 FILLER_143_752 ();
 sg13g2_fill_8 FILLER_143_760 ();
 sg13g2_fill_8 FILLER_143_768 ();
 sg13g2_fill_8 FILLER_143_776 ();
 sg13g2_fill_8 FILLER_143_784 ();
 sg13g2_fill_8 FILLER_143_792 ();
 sg13g2_fill_8 FILLER_143_800 ();
 sg13g2_fill_8 FILLER_143_808 ();
 sg13g2_fill_8 FILLER_143_816 ();
 sg13g2_fill_8 FILLER_143_824 ();
 sg13g2_fill_8 FILLER_143_832 ();
 sg13g2_fill_8 FILLER_143_840 ();
 sg13g2_fill_8 FILLER_143_848 ();
 sg13g2_fill_8 FILLER_143_856 ();
 sg13g2_fill_8 FILLER_143_864 ();
 sg13g2_fill_8 FILLER_143_872 ();
 sg13g2_fill_8 FILLER_143_880 ();
 sg13g2_fill_8 FILLER_143_888 ();
 sg13g2_fill_8 FILLER_143_896 ();
 sg13g2_fill_8 FILLER_143_904 ();
 sg13g2_fill_8 FILLER_143_912 ();
 sg13g2_fill_8 FILLER_143_920 ();
 sg13g2_fill_8 FILLER_143_928 ();
 sg13g2_fill_8 FILLER_143_936 ();
 sg13g2_fill_8 FILLER_143_944 ();
 sg13g2_fill_8 FILLER_143_952 ();
 sg13g2_fill_8 FILLER_143_960 ();
 sg13g2_fill_8 FILLER_143_968 ();
 sg13g2_fill_8 FILLER_143_976 ();
 sg13g2_fill_8 FILLER_143_984 ();
 sg13g2_fill_8 FILLER_143_992 ();
 sg13g2_fill_8 FILLER_143_1000 ();
 sg13g2_fill_8 FILLER_143_1008 ();
 sg13g2_fill_8 FILLER_143_1016 ();
 sg13g2_fill_8 FILLER_143_1024 ();
 sg13g2_fill_8 FILLER_143_1032 ();
 sg13g2_fill_8 FILLER_143_1040 ();
 sg13g2_fill_8 FILLER_143_1048 ();
 sg13g2_fill_8 FILLER_143_1056 ();
 sg13g2_fill_8 FILLER_143_1064 ();
 sg13g2_fill_8 FILLER_143_1072 ();
 sg13g2_fill_8 FILLER_143_1080 ();
 sg13g2_fill_8 FILLER_143_1088 ();
 sg13g2_fill_8 FILLER_143_1096 ();
 sg13g2_fill_8 FILLER_143_1104 ();
 sg13g2_fill_8 FILLER_143_1112 ();
 sg13g2_fill_8 FILLER_143_1120 ();
 sg13g2_fill_8 FILLER_143_1128 ();
 sg13g2_fill_8 FILLER_143_1136 ();
 sg13g2_fill_8 FILLER_144_0 ();
 sg13g2_fill_8 FILLER_144_8 ();
 sg13g2_fill_8 FILLER_144_16 ();
 sg13g2_fill_8 FILLER_144_24 ();
 sg13g2_fill_8 FILLER_144_32 ();
 sg13g2_fill_8 FILLER_144_40 ();
 sg13g2_fill_8 FILLER_144_48 ();
 sg13g2_fill_8 FILLER_144_56 ();
 sg13g2_fill_8 FILLER_144_64 ();
 sg13g2_fill_8 FILLER_144_72 ();
 sg13g2_fill_8 FILLER_144_80 ();
 sg13g2_fill_8 FILLER_144_88 ();
 sg13g2_fill_8 FILLER_144_96 ();
 sg13g2_fill_8 FILLER_144_104 ();
 sg13g2_fill_8 FILLER_144_112 ();
 sg13g2_fill_8 FILLER_144_120 ();
 sg13g2_fill_8 FILLER_144_128 ();
 sg13g2_fill_8 FILLER_144_136 ();
 sg13g2_fill_8 FILLER_144_144 ();
 sg13g2_fill_8 FILLER_144_152 ();
 sg13g2_fill_8 FILLER_144_160 ();
 sg13g2_fill_8 FILLER_144_168 ();
 sg13g2_fill_8 FILLER_144_176 ();
 sg13g2_fill_8 FILLER_144_184 ();
 sg13g2_fill_8 FILLER_144_192 ();
 sg13g2_fill_8 FILLER_144_200 ();
 sg13g2_fill_8 FILLER_144_208 ();
 sg13g2_fill_8 FILLER_144_216 ();
 sg13g2_fill_8 FILLER_144_224 ();
 sg13g2_fill_8 FILLER_144_232 ();
 sg13g2_fill_8 FILLER_144_240 ();
 sg13g2_fill_8 FILLER_144_248 ();
 sg13g2_fill_8 FILLER_144_256 ();
 sg13g2_fill_8 FILLER_144_264 ();
 sg13g2_fill_8 FILLER_144_272 ();
 sg13g2_fill_8 FILLER_144_280 ();
 sg13g2_fill_8 FILLER_144_288 ();
 sg13g2_fill_8 FILLER_144_296 ();
 sg13g2_fill_8 FILLER_144_304 ();
 sg13g2_fill_8 FILLER_144_312 ();
 sg13g2_fill_8 FILLER_144_320 ();
 sg13g2_fill_8 FILLER_144_328 ();
 sg13g2_fill_8 FILLER_144_336 ();
 sg13g2_fill_8 FILLER_144_344 ();
 sg13g2_fill_8 FILLER_144_352 ();
 sg13g2_fill_8 FILLER_144_360 ();
 sg13g2_fill_8 FILLER_144_368 ();
 sg13g2_fill_8 FILLER_144_376 ();
 sg13g2_fill_8 FILLER_144_384 ();
 sg13g2_fill_8 FILLER_144_392 ();
 sg13g2_fill_8 FILLER_144_400 ();
 sg13g2_fill_8 FILLER_144_408 ();
 sg13g2_fill_8 FILLER_144_416 ();
 sg13g2_fill_8 FILLER_144_424 ();
 sg13g2_fill_8 FILLER_144_432 ();
 sg13g2_fill_8 FILLER_144_440 ();
 sg13g2_fill_8 FILLER_144_448 ();
 sg13g2_fill_8 FILLER_144_456 ();
 sg13g2_fill_8 FILLER_144_464 ();
 sg13g2_fill_8 FILLER_144_472 ();
 sg13g2_fill_8 FILLER_144_480 ();
 sg13g2_fill_8 FILLER_144_488 ();
 sg13g2_fill_8 FILLER_144_496 ();
 sg13g2_fill_8 FILLER_144_504 ();
 sg13g2_fill_8 FILLER_144_512 ();
 sg13g2_fill_8 FILLER_144_520 ();
 sg13g2_fill_8 FILLER_144_528 ();
 sg13g2_fill_8 FILLER_144_536 ();
 sg13g2_fill_8 FILLER_144_544 ();
 sg13g2_fill_8 FILLER_144_552 ();
 sg13g2_fill_8 FILLER_144_560 ();
 sg13g2_fill_8 FILLER_144_568 ();
 sg13g2_fill_8 FILLER_144_576 ();
 sg13g2_fill_8 FILLER_144_584 ();
 sg13g2_fill_8 FILLER_144_592 ();
 sg13g2_fill_8 FILLER_144_600 ();
 sg13g2_fill_8 FILLER_144_608 ();
 sg13g2_fill_8 FILLER_144_616 ();
 sg13g2_fill_8 FILLER_144_624 ();
 sg13g2_fill_8 FILLER_144_632 ();
 sg13g2_fill_8 FILLER_144_640 ();
 sg13g2_fill_8 FILLER_144_648 ();
 sg13g2_fill_8 FILLER_144_656 ();
 sg13g2_fill_8 FILLER_144_664 ();
 sg13g2_fill_8 FILLER_144_672 ();
 sg13g2_fill_8 FILLER_144_680 ();
 sg13g2_fill_8 FILLER_144_688 ();
 sg13g2_fill_8 FILLER_144_696 ();
 sg13g2_fill_8 FILLER_144_704 ();
 sg13g2_fill_8 FILLER_144_712 ();
 sg13g2_fill_8 FILLER_144_720 ();
 sg13g2_fill_8 FILLER_144_728 ();
 sg13g2_fill_8 FILLER_144_736 ();
 sg13g2_fill_8 FILLER_144_744 ();
 sg13g2_fill_8 FILLER_144_752 ();
 sg13g2_fill_8 FILLER_144_760 ();
 sg13g2_fill_8 FILLER_144_768 ();
 sg13g2_fill_8 FILLER_144_776 ();
 sg13g2_fill_8 FILLER_144_784 ();
 sg13g2_fill_8 FILLER_144_792 ();
 sg13g2_fill_8 FILLER_144_800 ();
 sg13g2_fill_8 FILLER_144_808 ();
 sg13g2_fill_8 FILLER_144_816 ();
 sg13g2_fill_8 FILLER_144_824 ();
 sg13g2_fill_8 FILLER_144_832 ();
 sg13g2_fill_8 FILLER_144_840 ();
 sg13g2_fill_8 FILLER_144_848 ();
 sg13g2_fill_8 FILLER_144_856 ();
 sg13g2_fill_8 FILLER_144_864 ();
 sg13g2_fill_8 FILLER_144_872 ();
 sg13g2_fill_8 FILLER_144_880 ();
 sg13g2_fill_8 FILLER_144_888 ();
 sg13g2_fill_8 FILLER_144_896 ();
 sg13g2_fill_8 FILLER_144_904 ();
 sg13g2_fill_8 FILLER_144_912 ();
 sg13g2_fill_8 FILLER_144_920 ();
 sg13g2_fill_8 FILLER_144_928 ();
 sg13g2_fill_8 FILLER_144_936 ();
 sg13g2_fill_8 FILLER_144_944 ();
 sg13g2_fill_8 FILLER_144_952 ();
 sg13g2_fill_8 FILLER_144_960 ();
 sg13g2_fill_8 FILLER_144_968 ();
 sg13g2_fill_8 FILLER_144_976 ();
 sg13g2_fill_8 FILLER_144_984 ();
 sg13g2_fill_8 FILLER_144_992 ();
 sg13g2_fill_8 FILLER_144_1000 ();
 sg13g2_fill_8 FILLER_144_1008 ();
 sg13g2_fill_8 FILLER_144_1016 ();
 sg13g2_fill_8 FILLER_144_1024 ();
 sg13g2_fill_8 FILLER_144_1032 ();
 sg13g2_fill_8 FILLER_144_1040 ();
 sg13g2_fill_8 FILLER_144_1048 ();
 sg13g2_fill_8 FILLER_144_1056 ();
 sg13g2_fill_8 FILLER_144_1064 ();
 sg13g2_fill_8 FILLER_144_1072 ();
 sg13g2_fill_8 FILLER_144_1080 ();
 sg13g2_fill_8 FILLER_144_1088 ();
 sg13g2_fill_8 FILLER_144_1096 ();
 sg13g2_fill_8 FILLER_144_1104 ();
 sg13g2_fill_8 FILLER_144_1112 ();
 sg13g2_fill_8 FILLER_144_1120 ();
 sg13g2_fill_8 FILLER_144_1128 ();
 sg13g2_fill_8 FILLER_144_1136 ();
endmodule
