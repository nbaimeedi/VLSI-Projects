//Latest Update Date: 11th Nov, 2025
//Owner: B Nithin Reddy


//Interface

interface mul_if;
  
  logic [3:0] a,b;
  logic [7:0] y;
  
endinterface
