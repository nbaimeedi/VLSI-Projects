VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MACRO cve2_core
  FOREIGN cve2_core 0 0 ;
  CLASS BLOCK ;
  SIZE 1300 BY 1273.86 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
  END VDD
  PIN VDDIO
    USE POWER ;
    DIRECTION INOUT ;
  END VDDIO
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
  END VSS
  PIN VSSIO
    USE GROUND ;
    DIRECTION INOUT ;
  END VSSIO
  PIN boot_addr_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1250.24 0.72 1250.44 ;
    END
  END boot_addr_i_0_
  PIN boot_addr_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 370.76 0.72 370.96 ;
    END
  END boot_addr_i_10_
  PIN boot_addr_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 650.48 0.72 650.68 ;
    END
  END boot_addr_i_11_
  PIN boot_addr_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 554.72 0.72 554.92 ;
    END
  END boot_addr_i_12_
  PIN boot_addr_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 647.96 0.72 648.16 ;
    END
  END boot_addr_i_13_
  PIN boot_addr_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 453.92 0.72 454.12 ;
    END
  END boot_addr_i_14_
  PIN boot_addr_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 607.64 0.72 607.84 ;
    END
  END boot_addr_i_15_
  PIN boot_addr_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 660.56 0.72 660.76 ;
    END
  END boot_addr_i_16_
  PIN boot_addr_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 552.2 0.72 552.4 ;
    END
  END boot_addr_i_17_
  PIN boot_addr_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 451.4 0.72 451.6 ;
    END
  END boot_addr_i_18_
  PIN boot_addr_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 605.12 0.72 605.32 ;
    END
  END boot_addr_i_19_
  PIN boot_addr_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1247.72 0.72 1247.92 ;
    END
  END boot_addr_i_1_
  PIN boot_addr_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 398.48 0.72 398.68 ;
    END
  END boot_addr_i_20_
  PIN boot_addr_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 642.92 0.72 643.12 ;
    END
  END boot_addr_i_21_
  PIN boot_addr_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 380.84 0.72 381.04 ;
    END
  END boot_addr_i_22_
  PIN boot_addr_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 511.88 0.72 512.08 ;
    END
  END boot_addr_i_23_
  PIN boot_addr_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 602.6 0.72 602.8 ;
    END
  END boot_addr_i_24_
  PIN boot_addr_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 640.4 0.72 640.6 ;
    END
  END boot_addr_i_25_
  PIN boot_addr_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 446.36 0.72 446.56 ;
    END
  END boot_addr_i_26_
  PIN boot_addr_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 663.08 0.72 663.28 ;
    END
  END boot_addr_i_27_
  PIN boot_addr_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 600.08 0.72 600.28 ;
    END
  END boot_addr_i_28_
  PIN boot_addr_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 481.64 0.72 481.84 ;
    END
  END boot_addr_i_29_
  PIN boot_addr_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1245.2 0.72 1245.4 ;
    END
  END boot_addr_i_2_
  PIN boot_addr_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 685.76 0.72 685.96 ;
    END
  END boot_addr_i_30_
  PIN boot_addr_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 443.84 0.72 444.04 ;
    END
  END boot_addr_i_31_
  PIN boot_addr_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1242.68 0.72 1242.88 ;
    END
  END boot_addr_i_3_
  PIN boot_addr_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1240.16 0.72 1240.36 ;
    END
  END boot_addr_i_4_
  PIN boot_addr_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1237.64 0.72 1237.84 ;
    END
  END boot_addr_i_5_
  PIN boot_addr_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1235.12 0.72 1235.32 ;
    END
  END boot_addr_i_6_
  PIN boot_addr_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1232.6 0.72 1232.8 ;
    END
  END boot_addr_i_7_
  PIN boot_addr_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 539.6 0.72 539.8 ;
    END
  END boot_addr_i_8_
  PIN boot_addr_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 597.56 0.72 597.76 ;
    END
  END boot_addr_i_9_
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 395.96 0.72 396.16 ;
    END
  END clk_i
  PIN core_busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 564.8 1300 565 ;
    END
  END core_busy_o
  PIN crash_dump_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 567.32 1300 567.52 ;
    END
  END crash_dump_o_0_
  PIN crash_dump_o_100_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 569.84 1300 570.04 ;
    END
  END crash_dump_o_100_
  PIN crash_dump_o_101_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 572.36 1300 572.56 ;
    END
  END crash_dump_o_101_
  PIN crash_dump_o_102_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 574.88 1300 575.08 ;
    END
  END crash_dump_o_102_
  PIN crash_dump_o_103_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 577.4 1300 577.6 ;
    END
  END crash_dump_o_103_
  PIN crash_dump_o_104_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 579.92 1300 580.12 ;
    END
  END crash_dump_o_104_
  PIN crash_dump_o_105_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 582.44 1300 582.64 ;
    END
  END crash_dump_o_105_
  PIN crash_dump_o_106_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 584.96 1300 585.16 ;
    END
  END crash_dump_o_106_
  PIN crash_dump_o_107_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 587.48 1300 587.68 ;
    END
  END crash_dump_o_107_
  PIN crash_dump_o_108_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 590 1300 590.2 ;
    END
  END crash_dump_o_108_
  PIN crash_dump_o_109_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 592.52 1300 592.72 ;
    END
  END crash_dump_o_109_
  PIN crash_dump_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 595.04 1300 595.24 ;
    END
  END crash_dump_o_10_
  PIN crash_dump_o_110_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 597.56 1300 597.76 ;
    END
  END crash_dump_o_110_
  PIN crash_dump_o_111_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 600.08 1300 600.28 ;
    END
  END crash_dump_o_111_
  PIN crash_dump_o_112_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 602.6 1300 602.8 ;
    END
  END crash_dump_o_112_
  PIN crash_dump_o_113_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 605.12 1300 605.32 ;
    END
  END crash_dump_o_113_
  PIN crash_dump_o_114_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 607.64 1300 607.84 ;
    END
  END crash_dump_o_114_
  PIN crash_dump_o_115_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 610.16 1300 610.36 ;
    END
  END crash_dump_o_115_
  PIN crash_dump_o_116_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 612.68 1300 612.88 ;
    END
  END crash_dump_o_116_
  PIN crash_dump_o_117_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 615.2 1300 615.4 ;
    END
  END crash_dump_o_117_
  PIN crash_dump_o_118_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 617.72 1300 617.92 ;
    END
  END crash_dump_o_118_
  PIN crash_dump_o_119_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 620.24 1300 620.44 ;
    END
  END crash_dump_o_119_
  PIN crash_dump_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 622.76 1300 622.96 ;
    END
  END crash_dump_o_11_
  PIN crash_dump_o_120_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 625.28 1300 625.48 ;
    END
  END crash_dump_o_120_
  PIN crash_dump_o_121_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 627.8 1300 628 ;
    END
  END crash_dump_o_121_
  PIN crash_dump_o_122_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 630.32 1300 630.52 ;
    END
  END crash_dump_o_122_
  PIN crash_dump_o_123_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 632.84 1300 633.04 ;
    END
  END crash_dump_o_123_
  PIN crash_dump_o_124_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 635.36 1300 635.56 ;
    END
  END crash_dump_o_124_
  PIN crash_dump_o_125_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 637.88 1300 638.08 ;
    END
  END crash_dump_o_125_
  PIN crash_dump_o_126_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 640.4 1300 640.6 ;
    END
  END crash_dump_o_126_
  PIN crash_dump_o_127_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 642.92 1300 643.12 ;
    END
  END crash_dump_o_127_
  PIN crash_dump_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 645.44 1300 645.64 ;
    END
  END crash_dump_o_12_
  PIN crash_dump_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 647.96 1300 648.16 ;
    END
  END crash_dump_o_13_
  PIN crash_dump_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 650.48 1300 650.68 ;
    END
  END crash_dump_o_14_
  PIN crash_dump_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 653 1300 653.2 ;
    END
  END crash_dump_o_15_
  PIN crash_dump_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 655.52 1300 655.72 ;
    END
  END crash_dump_o_16_
  PIN crash_dump_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 658.04 1300 658.24 ;
    END
  END crash_dump_o_17_
  PIN crash_dump_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 660.56 1300 660.76 ;
    END
  END crash_dump_o_18_
  PIN crash_dump_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 663.08 1300 663.28 ;
    END
  END crash_dump_o_19_
  PIN crash_dump_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 665.6 1300 665.8 ;
    END
  END crash_dump_o_1_
  PIN crash_dump_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 668.12 1300 668.32 ;
    END
  END crash_dump_o_20_
  PIN crash_dump_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 670.64 1300 670.84 ;
    END
  END crash_dump_o_21_
  PIN crash_dump_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 673.16 1300 673.36 ;
    END
  END crash_dump_o_22_
  PIN crash_dump_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 675.68 1300 675.88 ;
    END
  END crash_dump_o_23_
  PIN crash_dump_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 678.2 1300 678.4 ;
    END
  END crash_dump_o_24_
  PIN crash_dump_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 680.72 1300 680.92 ;
    END
  END crash_dump_o_25_
  PIN crash_dump_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 683.24 1300 683.44 ;
    END
  END crash_dump_o_26_
  PIN crash_dump_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 685.76 1300 685.96 ;
    END
  END crash_dump_o_27_
  PIN crash_dump_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 688.28 1300 688.48 ;
    END
  END crash_dump_o_28_
  PIN crash_dump_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 690.8 1300 691 ;
    END
  END crash_dump_o_29_
  PIN crash_dump_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 693.32 1300 693.52 ;
    END
  END crash_dump_o_2_
  PIN crash_dump_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 695.84 1300 696.04 ;
    END
  END crash_dump_o_30_
  PIN crash_dump_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 698.36 1300 698.56 ;
    END
  END crash_dump_o_31_
  PIN crash_dump_o_32_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 700.88 1300 701.08 ;
    END
  END crash_dump_o_32_
  PIN crash_dump_o_33_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 703.4 1300 703.6 ;
    END
  END crash_dump_o_33_
  PIN crash_dump_o_34_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 705.92 1300 706.12 ;
    END
  END crash_dump_o_34_
  PIN crash_dump_o_35_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 708.44 1300 708.64 ;
    END
  END crash_dump_o_35_
  PIN crash_dump_o_36_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 710.96 1300 711.16 ;
    END
  END crash_dump_o_36_
  PIN crash_dump_o_37_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 713.48 1300 713.68 ;
    END
  END crash_dump_o_37_
  PIN crash_dump_o_38_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 716 1300 716.2 ;
    END
  END crash_dump_o_38_
  PIN crash_dump_o_39_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 718.52 1300 718.72 ;
    END
  END crash_dump_o_39_
  PIN crash_dump_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 721.04 1300 721.24 ;
    END
  END crash_dump_o_3_
  PIN crash_dump_o_40_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 723.56 1300 723.76 ;
    END
  END crash_dump_o_40_
  PIN crash_dump_o_41_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 726.08 1300 726.28 ;
    END
  END crash_dump_o_41_
  PIN crash_dump_o_42_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 728.6 1300 728.8 ;
    END
  END crash_dump_o_42_
  PIN crash_dump_o_43_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 731.12 1300 731.32 ;
    END
  END crash_dump_o_43_
  PIN crash_dump_o_44_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 733.64 1300 733.84 ;
    END
  END crash_dump_o_44_
  PIN crash_dump_o_45_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 736.16 1300 736.36 ;
    END
  END crash_dump_o_45_
  PIN crash_dump_o_46_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 738.68 1300 738.88 ;
    END
  END crash_dump_o_46_
  PIN crash_dump_o_47_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 741.2 1300 741.4 ;
    END
  END crash_dump_o_47_
  PIN crash_dump_o_48_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 743.72 1300 743.92 ;
    END
  END crash_dump_o_48_
  PIN crash_dump_o_49_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 746.24 1300 746.44 ;
    END
  END crash_dump_o_49_
  PIN crash_dump_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 748.76 1300 748.96 ;
    END
  END crash_dump_o_4_
  PIN crash_dump_o_50_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 751.28 1300 751.48 ;
    END
  END crash_dump_o_50_
  PIN crash_dump_o_51_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 753.8 1300 754 ;
    END
  END crash_dump_o_51_
  PIN crash_dump_o_52_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 756.32 1300 756.52 ;
    END
  END crash_dump_o_52_
  PIN crash_dump_o_53_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 758.84 1300 759.04 ;
    END
  END crash_dump_o_53_
  PIN crash_dump_o_54_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 761.36 1300 761.56 ;
    END
  END crash_dump_o_54_
  PIN crash_dump_o_55_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 763.88 1300 764.08 ;
    END
  END crash_dump_o_55_
  PIN crash_dump_o_56_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 766.4 1300 766.6 ;
    END
  END crash_dump_o_56_
  PIN crash_dump_o_57_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 768.92 1300 769.12 ;
    END
  END crash_dump_o_57_
  PIN crash_dump_o_58_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 771.44 1300 771.64 ;
    END
  END crash_dump_o_58_
  PIN crash_dump_o_59_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 773.96 1300 774.16 ;
    END
  END crash_dump_o_59_
  PIN crash_dump_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 776.48 1300 776.68 ;
    END
  END crash_dump_o_5_
  PIN crash_dump_o_60_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 779 1300 779.2 ;
    END
  END crash_dump_o_60_
  PIN crash_dump_o_61_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 781.52 1300 781.72 ;
    END
  END crash_dump_o_61_
  PIN crash_dump_o_62_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 784.04 1300 784.24 ;
    END
  END crash_dump_o_62_
  PIN crash_dump_o_63_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 786.56 1300 786.76 ;
    END
  END crash_dump_o_63_
  PIN crash_dump_o_64_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 552.2 1300 552.4 ;
    END
  END crash_dump_o_64_
  PIN crash_dump_o_65_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 789.08 1300 789.28 ;
    END
  END crash_dump_o_65_
  PIN crash_dump_o_66_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 791.6 1300 791.8 ;
    END
  END crash_dump_o_66_
  PIN crash_dump_o_67_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 794.12 1300 794.32 ;
    END
  END crash_dump_o_67_
  PIN crash_dump_o_68_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 796.64 1300 796.84 ;
    END
  END crash_dump_o_68_
  PIN crash_dump_o_69_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 799.16 1300 799.36 ;
    END
  END crash_dump_o_69_
  PIN crash_dump_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 801.68 1300 801.88 ;
    END
  END crash_dump_o_6_
  PIN crash_dump_o_70_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 804.2 1300 804.4 ;
    END
  END crash_dump_o_70_
  PIN crash_dump_o_71_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 806.72 1300 806.92 ;
    END
  END crash_dump_o_71_
  PIN crash_dump_o_72_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 809.24 1300 809.44 ;
    END
  END crash_dump_o_72_
  PIN crash_dump_o_73_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 811.76 1300 811.96 ;
    END
  END crash_dump_o_73_
  PIN crash_dump_o_74_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 814.28 1300 814.48 ;
    END
  END crash_dump_o_74_
  PIN crash_dump_o_75_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 816.8 1300 817 ;
    END
  END crash_dump_o_75_
  PIN crash_dump_o_76_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 819.32 1300 819.52 ;
    END
  END crash_dump_o_76_
  PIN crash_dump_o_77_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 821.84 1300 822.04 ;
    END
  END crash_dump_o_77_
  PIN crash_dump_o_78_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 824.36 1300 824.56 ;
    END
  END crash_dump_o_78_
  PIN crash_dump_o_79_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 826.88 1300 827.08 ;
    END
  END crash_dump_o_79_
  PIN crash_dump_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 829.4 1300 829.6 ;
    END
  END crash_dump_o_7_
  PIN crash_dump_o_80_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 831.92 1300 832.12 ;
    END
  END crash_dump_o_80_
  PIN crash_dump_o_81_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 834.44 1300 834.64 ;
    END
  END crash_dump_o_81_
  PIN crash_dump_o_82_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 836.96 1300 837.16 ;
    END
  END crash_dump_o_82_
  PIN crash_dump_o_83_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 839.48 1300 839.68 ;
    END
  END crash_dump_o_83_
  PIN crash_dump_o_84_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 842 1300 842.2 ;
    END
  END crash_dump_o_84_
  PIN crash_dump_o_85_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 844.52 1300 844.72 ;
    END
  END crash_dump_o_85_
  PIN crash_dump_o_86_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 847.04 1300 847.24 ;
    END
  END crash_dump_o_86_
  PIN crash_dump_o_87_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 849.56 1300 849.76 ;
    END
  END crash_dump_o_87_
  PIN crash_dump_o_88_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 852.08 1300 852.28 ;
    END
  END crash_dump_o_88_
  PIN crash_dump_o_89_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 854.6 1300 854.8 ;
    END
  END crash_dump_o_89_
  PIN crash_dump_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 857.12 1300 857.32 ;
    END
  END crash_dump_o_8_
  PIN crash_dump_o_90_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 859.64 1300 859.84 ;
    END
  END crash_dump_o_90_
  PIN crash_dump_o_91_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 862.16 1300 862.36 ;
    END
  END crash_dump_o_91_
  PIN crash_dump_o_92_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 864.68 1300 864.88 ;
    END
  END crash_dump_o_92_
  PIN crash_dump_o_93_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 867.2 1300 867.4 ;
    END
  END crash_dump_o_93_
  PIN crash_dump_o_94_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 869.72 1300 869.92 ;
    END
  END crash_dump_o_94_
  PIN crash_dump_o_95_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 872.24 1300 872.44 ;
    END
  END crash_dump_o_95_
  PIN crash_dump_o_96_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 874.76 1300 874.96 ;
    END
  END crash_dump_o_96_
  PIN crash_dump_o_97_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 877.28 1300 877.48 ;
    END
  END crash_dump_o_97_
  PIN crash_dump_o_98_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 879.8 1300 880 ;
    END
  END crash_dump_o_98_
  PIN crash_dump_o_99_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 882.32 1300 882.52 ;
    END
  END crash_dump_o_99_
  PIN crash_dump_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 884.84 1300 885.04 ;
    END
  END crash_dump_o_9_
  PIN data_addr_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 554.72 1300 554.92 ;
    END
  END data_addr_o_0_
  PIN data_addr_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 887.36 1300 887.56 ;
    END
  END data_addr_o_10_
  PIN data_addr_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 889.88 1300 890.08 ;
    END
  END data_addr_o_11_
  PIN data_addr_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 892.4 1300 892.6 ;
    END
  END data_addr_o_12_
  PIN data_addr_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 894.92 1300 895.12 ;
    END
  END data_addr_o_13_
  PIN data_addr_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 897.44 1300 897.64 ;
    END
  END data_addr_o_14_
  PIN data_addr_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 899.96 1300 900.16 ;
    END
  END data_addr_o_15_
  PIN data_addr_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 902.48 1300 902.68 ;
    END
  END data_addr_o_16_
  PIN data_addr_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 905 1300 905.2 ;
    END
  END data_addr_o_17_
  PIN data_addr_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 907.52 1300 907.72 ;
    END
  END data_addr_o_18_
  PIN data_addr_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 910.04 1300 910.24 ;
    END
  END data_addr_o_19_
  PIN data_addr_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 557.24 1300 557.44 ;
    END
  END data_addr_o_1_
  PIN data_addr_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 912.56 1300 912.76 ;
    END
  END data_addr_o_20_
  PIN data_addr_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 915.08 1300 915.28 ;
    END
  END data_addr_o_21_
  PIN data_addr_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 917.6 1300 917.8 ;
    END
  END data_addr_o_22_
  PIN data_addr_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 920.12 1300 920.32 ;
    END
  END data_addr_o_23_
  PIN data_addr_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 922.64 1300 922.84 ;
    END
  END data_addr_o_24_
  PIN data_addr_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 925.16 1300 925.36 ;
    END
  END data_addr_o_25_
  PIN data_addr_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 927.68 1300 927.88 ;
    END
  END data_addr_o_26_
  PIN data_addr_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 930.2 1300 930.4 ;
    END
  END data_addr_o_27_
  PIN data_addr_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 932.72 1300 932.92 ;
    END
  END data_addr_o_28_
  PIN data_addr_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 935.24 1300 935.44 ;
    END
  END data_addr_o_29_
  PIN data_addr_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 937.76 1300 937.96 ;
    END
  END data_addr_o_2_
  PIN data_addr_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 940.28 1300 940.48 ;
    END
  END data_addr_o_30_
  PIN data_addr_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 942.8 1300 943 ;
    END
  END data_addr_o_31_
  PIN data_addr_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 945.32 1300 945.52 ;
    END
  END data_addr_o_3_
  PIN data_addr_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 947.84 1300 948.04 ;
    END
  END data_addr_o_4_
  PIN data_addr_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 950.36 1300 950.56 ;
    END
  END data_addr_o_5_
  PIN data_addr_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 952.88 1300 953.08 ;
    END
  END data_addr_o_6_
  PIN data_addr_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 955.4 1300 955.6 ;
    END
  END data_addr_o_7_
  PIN data_addr_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 957.92 1300 958.12 ;
    END
  END data_addr_o_8_
  PIN data_addr_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 960.44 1300 960.64 ;
    END
  END data_addr_o_9_
  PIN data_be_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 962.96 1300 963.16 ;
    END
  END data_be_o_0_
  PIN data_be_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 965.48 1300 965.68 ;
    END
  END data_be_o_1_
  PIN data_be_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 968 1300 968.2 ;
    END
  END data_be_o_2_
  PIN data_be_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 970.52 1300 970.72 ;
    END
  END data_be_o_3_
  PIN data_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 441.32 0.72 441.52 ;
    END
  END data_err_i
  PIN data_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 698.36 0.72 698.56 ;
    END
  END data_gnt_i
  PIN data_rdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 544.64 0.72 544.84 ;
    END
  END data_rdata_i_0_
  PIN data_rdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 534.56 0.72 534.76 ;
    END
  END data_rdata_i_10_
  PIN data_rdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 612.68 0.72 612.88 ;
    END
  END data_rdata_i_11_
  PIN data_rdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 438.8 0.72 439 ;
    END
  END data_rdata_i_12_
  PIN data_rdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 532.04 0.72 532.24 ;
    END
  END data_rdata_i_13_
  PIN data_rdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 592.52 0.72 592.72 ;
    END
  END data_rdata_i_14_
  PIN data_rdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 635.36 0.72 635.56 ;
    END
  END data_rdata_i_15_
  PIN data_rdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 436.28 0.72 436.48 ;
    END
  END data_rdata_i_16_
  PIN data_rdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 499.28 0.72 499.48 ;
    END
  END data_rdata_i_17_
  PIN data_rdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 590 0.72 590.2 ;
    END
  END data_rdata_i_18_
  PIN data_rdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 527 0.72 527.2 ;
    END
  END data_rdata_i_19_
  PIN data_rdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 721.04 0.72 721.24 ;
    END
  END data_rdata_i_1_
  PIN data_rdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 433.76 0.72 433.96 ;
    END
  END data_rdata_i_20_
  PIN data_rdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 524.48 0.72 524.68 ;
    END
  END data_rdata_i_21_
  PIN data_rdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 587.48 0.72 587.68 ;
    END
  END data_rdata_i_22_
  PIN data_rdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 700.88 0.72 701.08 ;
    END
  END data_rdata_i_23_
  PIN data_rdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 393.44 0.72 393.64 ;
    END
  END data_rdata_i_24_
  PIN data_rdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 675.68 0.72 675.88 ;
    END
  END data_rdata_i_25_
  PIN data_rdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 431.24 0.72 431.44 ;
    END
  END data_rdata_i_26_
  PIN data_rdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 519.44 0.72 519.64 ;
    END
  END data_rdata_i_27_
  PIN data_rdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 620.24 0.72 620.44 ;
    END
  END data_rdata_i_28_
  PIN data_rdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 655.52 0.72 655.72 ;
    END
  END data_rdata_i_29_
  PIN data_rdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 516.92 0.72 517.12 ;
    END
  END data_rdata_i_2_
  PIN data_rdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 582.44 0.72 582.64 ;
    END
  END data_rdata_i_30_
  PIN data_rdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 428.72 0.72 428.92 ;
    END
  END data_rdata_i_31_
  PIN data_rdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 390.92 0.72 391.12 ;
    END
  END data_rdata_i_3_
  PIN data_rdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 736.16 0.72 736.36 ;
    END
  END data_rdata_i_4_
  PIN data_rdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 489.2 0.72 489.4 ;
    END
  END data_rdata_i_5_
  PIN data_rdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 426.2 0.72 426.4 ;
    END
  END data_rdata_i_6_
  PIN data_rdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 537.08 0.72 537.28 ;
    END
  END data_rdata_i_7_
  PIN data_rdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 741.2 0.72 741.4 ;
    END
  END data_rdata_i_8_
  PIN data_rdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 509.36 0.72 509.56 ;
    END
  END data_rdata_i_9_
  PIN data_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 973.04 1300 973.24 ;
    END
  END data_req_o
  PIN data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 577.4 0.72 577.6 ;
    END
  END data_rvalid_i
  PIN data_wdata_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 975.56 1300 975.76 ;
    END
  END data_wdata_o_0_
  PIN data_wdata_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 978.08 1300 978.28 ;
    END
  END data_wdata_o_10_
  PIN data_wdata_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 980.6 1300 980.8 ;
    END
  END data_wdata_o_11_
  PIN data_wdata_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 983.12 1300 983.32 ;
    END
  END data_wdata_o_12_
  PIN data_wdata_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 985.64 1300 985.84 ;
    END
  END data_wdata_o_13_
  PIN data_wdata_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 988.16 1300 988.36 ;
    END
  END data_wdata_o_14_
  PIN data_wdata_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 990.68 1300 990.88 ;
    END
  END data_wdata_o_15_
  PIN data_wdata_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 993.2 1300 993.4 ;
    END
  END data_wdata_o_16_
  PIN data_wdata_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 995.72 1300 995.92 ;
    END
  END data_wdata_o_17_
  PIN data_wdata_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 998.24 1300 998.44 ;
    END
  END data_wdata_o_18_
  PIN data_wdata_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1000.76 1300 1000.96 ;
    END
  END data_wdata_o_19_
  PIN data_wdata_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1003.28 1300 1003.48 ;
    END
  END data_wdata_o_1_
  PIN data_wdata_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1005.8 1300 1006 ;
    END
  END data_wdata_o_20_
  PIN data_wdata_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1008.32 1300 1008.52 ;
    END
  END data_wdata_o_21_
  PIN data_wdata_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1010.84 1300 1011.04 ;
    END
  END data_wdata_o_22_
  PIN data_wdata_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1013.36 1300 1013.56 ;
    END
  END data_wdata_o_23_
  PIN data_wdata_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1015.88 1300 1016.08 ;
    END
  END data_wdata_o_24_
  PIN data_wdata_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1018.4 1300 1018.6 ;
    END
  END data_wdata_o_25_
  PIN data_wdata_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1020.92 1300 1021.12 ;
    END
  END data_wdata_o_26_
  PIN data_wdata_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1023.44 1300 1023.64 ;
    END
  END data_wdata_o_27_
  PIN data_wdata_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1025.96 1300 1026.16 ;
    END
  END data_wdata_o_28_
  PIN data_wdata_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1028.48 1300 1028.68 ;
    END
  END data_wdata_o_29_
  PIN data_wdata_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1031 1300 1031.2 ;
    END
  END data_wdata_o_2_
  PIN data_wdata_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1033.52 1300 1033.72 ;
    END
  END data_wdata_o_30_
  PIN data_wdata_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1036.04 1300 1036.24 ;
    END
  END data_wdata_o_31_
  PIN data_wdata_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1038.56 1300 1038.76 ;
    END
  END data_wdata_o_3_
  PIN data_wdata_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1041.08 1300 1041.28 ;
    END
  END data_wdata_o_4_
  PIN data_wdata_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1043.6 1300 1043.8 ;
    END
  END data_wdata_o_5_
  PIN data_wdata_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1046.12 1300 1046.32 ;
    END
  END data_wdata_o_6_
  PIN data_wdata_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1048.64 1300 1048.84 ;
    END
  END data_wdata_o_7_
  PIN data_wdata_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1051.16 1300 1051.36 ;
    END
  END data_wdata_o_8_
  PIN data_wdata_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 1053.68 1300 1053.88 ;
    END
  END data_wdata_o_9_
  PIN data_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 469.04 1300 469.24 ;
    END
  END data_we_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 743.72 0.72 743.92 ;
    END
  END debug_req_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 506.84 0.72 507.04 ;
    END
  END fetch_enable_i
  PIN hart_id_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 728.6 0.72 728.8 ;
    END
  END hart_id_i_0_
  PIN hart_id_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 610.16 0.72 610.36 ;
    END
  END hart_id_i_10_
  PIN hart_id_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 504.32 0.72 504.52 ;
    END
  END hart_id_i_11_
  PIN hart_id_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 637.88 0.72 638.08 ;
    END
  END hart_id_i_12_
  PIN hart_id_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 423.68 0.72 423.88 ;
    END
  END hart_id_i_13_
  PIN hart_id_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 501.8 0.72 502 ;
    END
  END hart_id_i_14_
  PIN hart_id_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 665.6 0.72 665.8 ;
    END
  END hart_id_i_15_
  PIN hart_id_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 378.32 0.72 378.52 ;
    END
  END hart_id_i_16_
  PIN hart_id_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 658.04 0.72 658.24 ;
    END
  END hart_id_i_17_
  PIN hart_id_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 421.16 0.72 421.36 ;
    END
  END hart_id_i_18_
  PIN hart_id_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 716 0.72 716.2 ;
    END
  END hart_id_i_19_
  PIN hart_id_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 713.48 0.72 713.68 ;
    END
  END hart_id_i_1_
  PIN hart_id_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 569.84 0.72 570.04 ;
    END
  END hart_id_i_20_
  PIN hart_id_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 496.76 0.72 496.96 ;
    END
  END hart_id_i_21_
  PIN hart_id_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 388.4 0.72 388.6 ;
    END
  END hart_id_i_22_
  PIN hart_id_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 680.72 0.72 680.92 ;
    END
  END hart_id_i_23_
  PIN hart_id_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 567.32 0.72 567.52 ;
    END
  END hart_id_i_24_
  PIN hart_id_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 494.24 0.72 494.44 ;
    END
  END hart_id_i_25_
  PIN hart_id_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 373.28 0.72 373.48 ;
    END
  END hart_id_i_26_
  PIN hart_id_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 418.64 0.72 418.84 ;
    END
  END hart_id_i_27_
  PIN hart_id_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 549.68 0.72 549.88 ;
    END
  END hart_id_i_28_
  PIN hart_id_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 491.72 0.72 491.92 ;
    END
  END hart_id_i_29_
  PIN hart_id_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 690.8 0.72 691 ;
    END
  END hart_id_i_2_
  PIN hart_id_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 630.32 0.72 630.52 ;
    END
  END hart_id_i_30_
  PIN hart_id_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 622.76 0.72 622.96 ;
    END
  END hart_id_i_31_
  PIN hart_id_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 416.12 0.72 416.32 ;
    END
  END hart_id_i_3_
  PIN hart_id_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 471.56 0.72 471.76 ;
    END
  END hart_id_i_4_
  PIN hart_id_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 678.2 0.72 678.4 ;
    END
  END hart_id_i_5_
  PIN hart_id_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 708.44 0.72 708.64 ;
    END
  END hart_id_i_6_
  PIN hart_id_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 486.68 0.72 486.88 ;
    END
  END hart_id_i_7_
  PIN hart_id_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 673.16 0.72 673.36 ;
    END
  END hart_id_i_8_
  PIN hart_id_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 718.52 0.72 718.72 ;
    END
  END hart_id_i_9_
  PIN instr_addr_o_0_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 559.76 1300 559.96 ;
    END
  END instr_addr_o_0_
  PIN instr_addr_o_10_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 549.68 1300 549.88 ;
    END
  END instr_addr_o_10_
  PIN instr_addr_o_11_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 547.16 1300 547.36 ;
    END
  END instr_addr_o_11_
  PIN instr_addr_o_12_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 544.64 1300 544.84 ;
    END
  END instr_addr_o_12_
  PIN instr_addr_o_13_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 542.12 1300 542.32 ;
    END
  END instr_addr_o_13_
  PIN instr_addr_o_14_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 539.6 1300 539.8 ;
    END
  END instr_addr_o_14_
  PIN instr_addr_o_15_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 537.08 1300 537.28 ;
    END
  END instr_addr_o_15_
  PIN instr_addr_o_16_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 534.56 1300 534.76 ;
    END
  END instr_addr_o_16_
  PIN instr_addr_o_17_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 532.04 1300 532.24 ;
    END
  END instr_addr_o_17_
  PIN instr_addr_o_18_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 529.52 1300 529.72 ;
    END
  END instr_addr_o_18_
  PIN instr_addr_o_19_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 527 1300 527.2 ;
    END
  END instr_addr_o_19_
  PIN instr_addr_o_1_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 562.28 1300 562.48 ;
    END
  END instr_addr_o_1_
  PIN instr_addr_o_20_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 524.48 1300 524.68 ;
    END
  END instr_addr_o_20_
  PIN instr_addr_o_21_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 521.96 1300 522.16 ;
    END
  END instr_addr_o_21_
  PIN instr_addr_o_22_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 519.44 1300 519.64 ;
    END
  END instr_addr_o_22_
  PIN instr_addr_o_23_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 516.92 1300 517.12 ;
    END
  END instr_addr_o_23_
  PIN instr_addr_o_24_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 514.4 1300 514.6 ;
    END
  END instr_addr_o_24_
  PIN instr_addr_o_25_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 511.88 1300 512.08 ;
    END
  END instr_addr_o_25_
  PIN instr_addr_o_26_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 509.36 1300 509.56 ;
    END
  END instr_addr_o_26_
  PIN instr_addr_o_27_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 506.84 1300 507.04 ;
    END
  END instr_addr_o_27_
  PIN instr_addr_o_28_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 504.32 1300 504.52 ;
    END
  END instr_addr_o_28_
  PIN instr_addr_o_29_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 501.8 1300 502 ;
    END
  END instr_addr_o_29_
  PIN instr_addr_o_2_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 499.28 1300 499.48 ;
    END
  END instr_addr_o_2_
  PIN instr_addr_o_30_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 496.76 1300 496.96 ;
    END
  END instr_addr_o_30_
  PIN instr_addr_o_31_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 494.24 1300 494.44 ;
    END
  END instr_addr_o_31_
  PIN instr_addr_o_3_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 491.72 1300 491.92 ;
    END
  END instr_addr_o_3_
  PIN instr_addr_o_4_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 489.2 1300 489.4 ;
    END
  END instr_addr_o_4_
  PIN instr_addr_o_5_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 486.68 1300 486.88 ;
    END
  END instr_addr_o_5_
  PIN instr_addr_o_6_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 484.16 1300 484.36 ;
    END
  END instr_addr_o_6_
  PIN instr_addr_o_7_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 481.64 1300 481.84 ;
    END
  END instr_addr_o_7_
  PIN instr_addr_o_8_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 479.12 1300 479.32 ;
    END
  END instr_addr_o_8_
  PIN instr_addr_o_9_
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 476.6 1300 476.8 ;
    END
  END instr_addr_o_9_
  PIN instr_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 668.12 0.72 668.32 ;
    END
  END instr_err_i
  PIN instr_gnt_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 484.16 0.72 484.36 ;
    END
  END instr_gnt_i
  PIN instr_rdata_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 693.32 0.72 693.52 ;
    END
  END instr_rdata_i_0_
  PIN instr_rdata_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 695.84 0.72 696.04 ;
    END
  END instr_rdata_i_10_
  PIN instr_rdata_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 617.72 0.72 617.92 ;
    END
  END instr_rdata_i_11_
  PIN instr_rdata_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 413.6 0.72 413.8 ;
    END
  END instr_rdata_i_12_
  PIN instr_rdata_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 653 0.72 653.2 ;
    END
  END instr_rdata_i_13_
  PIN instr_rdata_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 731.12 0.72 731.32 ;
    END
  END instr_rdata_i_14_
  PIN instr_rdata_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 627.8 0.72 628 ;
    END
  END instr_rdata_i_15_
  PIN instr_rdata_i_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 479.12 0.72 479.32 ;
    END
  END instr_rdata_i_16_
  PIN instr_rdata_i_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 710.96 0.72 711.16 ;
    END
  END instr_rdata_i_17_
  PIN instr_rdata_i_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 703.4 0.72 703.6 ;
    END
  END instr_rdata_i_18_
  PIN instr_rdata_i_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 411.08 0.72 411.28 ;
    END
  END instr_rdata_i_19_
  PIN instr_rdata_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 476.6 0.72 476.8 ;
    END
  END instr_rdata_i_1_
  PIN instr_rdata_i_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 645.44 0.72 645.64 ;
    END
  END instr_rdata_i_20_
  PIN instr_rdata_i_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 683.24 0.72 683.44 ;
    END
  END instr_rdata_i_21_
  PIN instr_rdata_i_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 746.24 0.72 746.44 ;
    END
  END instr_rdata_i_22_
  PIN instr_rdata_i_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 474.08 0.72 474.28 ;
    END
  END instr_rdata_i_23_
  PIN instr_rdata_i_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 733.64 0.72 733.84 ;
    END
  END instr_rdata_i_24_
  PIN instr_rdata_i_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 584.96 0.72 585.16 ;
    END
  END instr_rdata_i_25_
  PIN instr_rdata_i_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 726.08 0.72 726.28 ;
    END
  END instr_rdata_i_26_
  PIN instr_rdata_i_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 408.56 0.72 408.76 ;
    END
  END instr_rdata_i_27_
  PIN instr_rdata_i_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 615.2 0.72 615.4 ;
    END
  END instr_rdata_i_28_
  PIN instr_rdata_i_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 375.8 0.72 376 ;
    END
  END instr_rdata_i_29_
  PIN instr_rdata_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 385.88 0.72 386.08 ;
    END
  END instr_rdata_i_2_
  PIN instr_rdata_i_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 574.88 0.72 575.08 ;
    END
  END instr_rdata_i_30_
  PIN instr_rdata_i_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 469.04 0.72 469.24 ;
    END
  END instr_rdata_i_31_
  PIN instr_rdata_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 406.04 0.72 406.24 ;
    END
  END instr_rdata_i_3_
  PIN instr_rdata_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 738.68 0.72 738.88 ;
    END
  END instr_rdata_i_4_
  PIN instr_rdata_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 572.36 0.72 572.56 ;
    END
  END instr_rdata_i_5_
  PIN instr_rdata_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 595.04 0.72 595.24 ;
    END
  END instr_rdata_i_6_
  PIN instr_rdata_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 625.28 0.72 625.48 ;
    END
  END instr_rdata_i_7_
  PIN instr_rdata_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 403.52 0.72 403.72 ;
    END
  END instr_rdata_i_8_
  PIN instr_rdata_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 466.52 0.72 466.72 ;
    END
  END instr_rdata_i_9_
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 474.08 1300 474.28 ;
    END
  END instr_req_o
  PIN instr_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 688.28 0.72 688.48 ;
    END
  END instr_rvalid_i
  PIN irq_external_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 521.96 0.72 522.16 ;
    END
  END irq_external_i
  PIN irq_fast_i_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 542.12 0.72 542.32 ;
    END
  END irq_fast_i_0_
  PIN irq_fast_i_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 464 0.72 464.2 ;
    END
  END irq_fast_i_10_
  PIN irq_fast_i_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 383.36 0.72 383.56 ;
    END
  END irq_fast_i_11_
  PIN irq_fast_i_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 448.88 0.72 449.08 ;
    END
  END irq_fast_i_12_
  PIN irq_fast_i_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 632.84 0.72 633.04 ;
    END
  END irq_fast_i_13_
  PIN irq_fast_i_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 564.8 0.72 565 ;
    END
  END irq_fast_i_14_
  PIN irq_fast_i_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 529.52 0.72 529.72 ;
    END
  END irq_fast_i_15_
  PIN irq_fast_i_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 559.76 0.72 559.96 ;
    END
  END irq_fast_i_1_
  PIN irq_fast_i_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 514.4 0.72 514.6 ;
    END
  END irq_fast_i_2_
  PIN irq_fast_i_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 562.28 0.72 562.48 ;
    END
  END irq_fast_i_3_
  PIN irq_fast_i_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 461.48 0.72 461.68 ;
    END
  END irq_fast_i_4_
  PIN irq_fast_i_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 705.92 0.72 706.12 ;
    END
  END irq_fast_i_5_
  PIN irq_fast_i_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 723.56 0.72 723.76 ;
    END
  END irq_fast_i_6_
  PIN irq_fast_i_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 547.16 0.72 547.36 ;
    END
  END irq_fast_i_7_
  PIN irq_fast_i_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 458.96 0.72 459.16 ;
    END
  END irq_fast_i_8_
  PIN irq_fast_i_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 579.92 0.72 580.12 ;
    END
  END irq_fast_i_9_
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 670.64 0.72 670.84 ;
    END
  END irq_nm_i
  PIN irq_pending_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  1299.28 471.56 1300 471.76 ;
    END
  END irq_pending_o
  PIN irq_software_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 557.24 0.72 557.44 ;
    END
  END irq_software_i
  PIN irq_timer_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 401 0.72 401.2 ;
    END
  END irq_timer_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 456.44 0.72 456.64 ;
    END
  END rst_ni
  PIN test_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT  0 1230.08 0.72 1230.28 ;
    END
  END test_en_i
  OBS
    LAYER Metal1 ;
     RECT  25.44 26.24 1274.88 498.04 ;
     RECT  25.44 498.04 1275.44 499.88 ;
     RECT  1288.72 494.26 1288.88 500.3 ;
     RECT  1288.72 521.98 1288.88 528.44 ;
     RECT  25.44 499.88 1274.88 529.54 ;
     RECT  25.44 529.54 1275.44 537.1 ;
     RECT  25.44 537.1 1281.2 539.78 ;
     RECT  1298.8 474.1 1298.96 544.4 ;
     RECT  1297.36 574.9 1297.52 577.42 ;
     RECT  25.44 539.78 1274.88 577.715 ;
     RECT  25.44 577.715 1274.96 587.5 ;
     RECT  1296.4 577.42 1297.52 600.1 ;
     RECT  1289.68 600.1 1297.52 615.22 ;
     RECT  1289.68 615.22 1298 631.18 ;
     RECT  0.88 566.08 1.04 634.96 ;
     RECT  0.88 634.96 3.92 645.88 ;
     RECT  25.44 587.5 1277.84 646.46 ;
     RECT  1288.72 631.18 1298 649.24 ;
     RECT  1288.72 649.24 1298.48 655.96 ;
     RECT  0.88 645.88 5.36 678.38 ;
     RECT  1288.72 655.96 1298.96 678.38 ;
     RECT  0.88 678.38 1.04 680.9 ;
     RECT  1289.2 678.38 1298.96 681.16 ;
     RECT  1289.2 681.16 1299.44 691.24 ;
     RECT  1284.88 691.24 1299.44 710.72 ;
     RECT  25.44 646.46 1274.88 728.62 ;
     RECT  1284.88 710.72 1298.96 728.62 ;
     RECT  25.44 728.62 1298.96 773.3 ;
     RECT  1284.88 773.3 1298.96 784.48 ;
     RECT  1284.88 784.48 1299.44 793.04 ;
     RECT  1284.88 793.04 1298.96 804.38 ;
     RECT  1288.72 804.38 1298.96 833.78 ;
     RECT  25.44 773.3 1274.88 867.64 ;
     RECT  25.44 867.64 1277.84 920.3 ;
     RECT  1291.6 833.78 1298.96 921.4 ;
     RECT  1288.72 921.4 1298.96 940.46 ;
     RECT  1291.6 940.46 1298.96 942.98 ;
     RECT  1291.6 942.98 1291.76 945.5 ;
     RECT  25.44 920.3 1274.88 992.8 ;
     RECT  25.44 992.8 1275.92 1019.68 ;
     RECT  1288.72 996.58 1288.88 1019.68 ;
     RECT  25.44 1019.68 1288.88 1027.24 ;
     RECT  1298.8 1007.08 1298.96 1027.24 ;
     RECT  25.44 1027.24 1298.96 1041.26 ;
     RECT  1297.36 1041.26 1298.96 1048.82 ;
     RECT  1298.8 1048.82 1298.96 1051.34 ;
     RECT  25.44 1041.26 1284.08 1053.86 ;
     RECT  25.44 1053.86 1274.88 1274.08 ;
    LAYER Metal2 ;
     RECT  0.38 378.74 0.48 378.94 ;
     RECT  0.38 421.58 0.48 423.04 ;
     RECT  0.38 444.26 0.48 445.3 ;
     RECT  0.38 542.54 0.48 558.7 ;
     RECT  0.38 580.34 0.48 581.38 ;
     RECT  0.38 610.58 0.48 611.62 ;
     RECT  0.38 631.58 0.48 632.62 ;
     RECT  0.38 729.86 0.48 730.9 ;
     RECT  0.48 370.76 3.46 746.44 ;
     RECT  3.46 663.08 3.94 746.44 ;
     RECT  3.46 611.42 7.3 653.2 ;
     RECT  3.94 668.12 7.3 746.44 ;
     RECT  3.46 558.5 35.9 600.28 ;
     RECT  7.3 721.04 36.1 746.44 ;
     RECT  534.62 904.58 535.1 913.18 ;
     RECT  534.62 928.52 535.1 928.72 ;
     RECT  534.62 892.82 535.58 893.02 ;
     RECT  535.1 904.58 535.58 928.72 ;
     RECT  535.58 892.82 537.02 928.72 ;
     RECT  537.02 886.94 537.98 928.72 ;
     RECT  7.3 645.44 540.1 653.2 ;
     RECT  7.3 668.12 540.1 683.44 ;
     RECT  36.1 721.04 540.1 745.6 ;
     RECT  537.98 879.8 540.38 928.72 ;
     RECT  540.38 945.74 540.86 947.2 ;
     RECT  540.38 965.48 540.86 965.68 ;
     RECT  540.38 856.7 541.34 863.62 ;
     RECT  540.38 878.96 541.34 935.86 ;
     RECT  540.86 945.74 541.34 955.18 ;
     RECT  540.86 965.48 541.34 966.52 ;
     RECT  541.34 856.7 542.24 866.98 ;
     RECT  543.26 822.26 545.12 830.44 ;
     RECT  543.74 1139.36 545.18 1139.56 ;
     RECT  545.12 822.225 546.14 830.44 ;
     RECT  546.14 821.84 547.1 830.44 ;
     RECT  542.24 856.7 547.1 867.99 ;
     RECT  545.18 1139.36 547.1 1139.98 ;
     RECT  547.1 821.84 547.58 833.8 ;
     RECT  547.1 849.56 547.58 867.99 ;
     RECT  547.1 1138.52 547.58 1142.5 ;
     RECT  541.34 878.96 548.54 966.52 ;
     RECT  543.74 1080.14 548.54 1086.64 ;
     RECT  547.58 1101.56 548.54 1101.76 ;
     RECT  547.58 1130.54 548.54 1142.5 ;
     RECT  548.54 878.96 549.02 969.46 ;
     RECT  547.1 1181.36 549.02 1181.56 ;
     RECT  547.58 821.84 549.5 867.99 ;
     RECT  548.54 1064.18 549.5 1064.38 ;
     RECT  548.54 1074.26 549.5 1086.64 ;
     RECT  548.54 1101.56 549.5 1142.5 ;
     RECT  549.5 821.84 549.98 868.66 ;
     RECT  549.02 878.96 549.98 969.88 ;
     RECT  549.5 1064.18 549.98 1086.64 ;
     RECT  549.5 1101.56 549.98 1144.18 ;
     RECT  549.98 1101.14 550.46 1163.08 ;
     RECT  549.98 1059.56 550.88 1086.64 ;
     RECT  549.02 1174.22 550.94 1182.4 ;
     RECT  550.88 1059.56 551.42 1090.455 ;
     RECT  549.98 821.84 551.9 969.88 ;
     RECT  550.94 1172.54 552.38 1182.4 ;
     RECT  551.42 1059.56 552.86 1090.84 ;
     RECT  550.46 1100.72 552.86 1163.08 ;
     RECT  552.38 1172.54 554.3 1183.66 ;
     RECT  552.86 1059.56 554.78 1163.08 ;
     RECT  554.3 1172.54 554.78 1184.08 ;
     RECT  551.9 814.28 555.16 969.88 ;
     RECT  555.16 814.28 555.5 969.89 ;
     RECT  555.5 813.44 555.74 969.89 ;
     RECT  554.78 980.6 555.74 982.48 ;
     RECT  555.74 811.34 556.22 982.48 ;
     RECT  556.22 811.34 556.7 986.68 ;
     RECT  556.7 811.34 557.12 987.52 ;
     RECT  557.66 1019.66 558.14 1025.74 ;
     RECT  554.78 1059.56 558.325 1184.08 ;
     RECT  558.14 1012.1 558.62 1025.74 ;
     RECT  558.325 1097.78 558.62 1184.08 ;
     RECT  558.62 1044.02 559.1 1048.42 ;
     RECT  558.325 1059.56 559.1 1086.64 ;
     RECT  558.62 1004.54 559.52 1025.74 ;
     RECT  559.52 1004.54 560.54 1026.75 ;
     RECT  560.54 1002.02 561.02 1026.75 ;
     RECT  561.02 999.5 561.5 1026.75 ;
     RECT  558.62 1097.78 561.5 1193.32 ;
     RECT  557.12 810.33 562.46 987.52 ;
     RECT  561.5 1097.78 562.46 1204.66 ;
     RECT  554.78 1214.96 562.46 1215.16 ;
     RECT  562.46 810.33 562.94 988.36 ;
     RECT  561.5 998.24 562.94 1026.75 ;
     RECT  562.94 998.24 563.9 1029.1 ;
     RECT  562.46 1097.78 564.38 1218.1 ;
     RECT  563.42 1226.72 564.38 1226.92 ;
     RECT  563.9 998.24 565.34 1030.36 ;
     RECT  564.38 1097.78 565.82 1226.92 ;
     RECT  565.34 998.24 566.3 1032.88 ;
     RECT  565.82 1097.78 566.78 1234.06 ;
     RECT  562.46 1248.14 566.78 1248.34 ;
     RECT  562.94 810.33 568.7 989.62 ;
     RECT  566.3 998.24 568.7 1033.3 ;
     RECT  568.7 810.33 569.66 1034.14 ;
     RECT  559.1 1044.02 569.66 1086.64 ;
     RECT  569.66 807.14 570.56 1086.64 ;
     RECT  570.56 802.77 570.62 1086.64 ;
     RECT  566.78 1097.78 571.58 1248.34 ;
     RECT  570.62 802.77 572.06 1087.06 ;
     RECT  571.58 1097.36 572.54 1248.34 ;
     RECT  572.06 802.77 573.02 1087.48 ;
     RECT  572.54 1097.36 573.02 1249.6 ;
     RECT  573.02 802.77 573.22 1249.6 ;
     RECT  573.22 802.77 578.005 1248.34 ;
     RECT  578.005 802.94 582.14 1248.34 ;
     RECT  582.14 802.94 585.5 1249.6 ;
     RECT  585.5 802.94 589.82 1250.02 ;
     RECT  589.82 802.94 592.22 1252.54 ;
     RECT  592.22 800.42 593.18 1252.54 ;
     RECT  593.18 799.16 595.58 1252.54 ;
     RECT  595.58 799.16 599.9 1253.38 ;
     RECT  599.9 799.16 601.82 1257.58 ;
     RECT  601.82 796.22 602.02 1257.58 ;
     RECT  602.02 806.3 602.98 1257.58 ;
     RECT  602.02 796.22 603.46 796.42 ;
     RECT  540.1 723.56 604.62 745.6 ;
     RECT  604.22 776.48 604.7 776.68 ;
     RECT  604.62 723.56 605.395 753.58 ;
     RECT  602.78 762.62 605.395 765.76 ;
     RECT  605.395 723.56 605.66 765.76 ;
     RECT  604.7 776.48 605.66 777.52 ;
     RECT  7.3 611.42 606.34 635.56 ;
     RECT  540.1 668.54 607.78 683.44 ;
     RECT  602.98 806.3 608.26 1256.32 ;
     RECT  605.66 723.56 609.02 777.52 ;
     RECT  609.02 723.56 609.5 781.3 ;
     RECT  609.5 723.56 611.9 781.72 ;
     RECT  605.18 795.8 611.9 796 ;
     RECT  611.9 723.56 612.38 796 ;
     RECT  608.26 806.3 612.38 1254.22 ;
     RECT  3.46 489.2 615.94 548.62 ;
     RECT  612.38 723.56 618.14 1254.22 ;
     RECT  618.14 723.56 619.04 1256.74 ;
     RECT  607.78 668.54 619.1 668.74 ;
     RECT  619.1 668.54 619.3 669.16 ;
     RECT  619.04 723.56 619.33 1256.775 ;
     RECT  606.34 611.42 620.06 635.14 ;
     RECT  540.1 645.44 620.06 652.78 ;
     RECT  620.06 611.42 620.54 652.78 ;
     RECT  35.9 558.5 620.74 600.7 ;
     RECT  619.3 668.96 621.5 669.16 ;
     RECT  607.78 683.24 621.5 683.44 ;
     RECT  615.94 489.2 621.7 507.04 ;
     RECT  7.3 695.84 622.46 711.16 ;
     RECT  619.33 723.56 622.46 1256.74 ;
     RECT  622.46 695.84 623.9 1256.74 ;
     RECT  621.5 668.96 624.86 683.44 ;
     RECT  623.9 693.32 624.86 1256.74 ;
     RECT  624.86 668.96 626.485 1256.74 ;
     RECT  620.54 611.42 634.94 659.92 ;
     RECT  626.485 668.96 634.94 1255.9 ;
     RECT  634.94 611.42 637.76 1255.9 ;
     RECT  637.76 611.42 638.3 1256.775 ;
     RECT  620.74 590 639.94 600.7 ;
     RECT  3.46 370.76 644.26 479.32 ;
     RECT  638.3 611.42 650.78 1257.58 ;
     RECT  650.78 611.42 651.26 1260.1 ;
     RECT  651.26 611.42 651.74 1260.52 ;
     RECT  639.94 590 652.9 590.2 ;
     RECT  651.74 611.42 656.74 1261.36 ;
     RECT  615.94 516.92 660.1 548.62 ;
     RECT  656.74 611.42 661.06 1256.32 ;
     RECT  660.1 516.92 661.54 534.76 ;
     RECT  661.06 611.42 662.98 1254.22 ;
     RECT  662.98 624.44 664.9 1254.22 ;
     RECT  661.54 519.44 666.82 534.76 ;
     RECT  664.9 624.44 668.26 1250.44 ;
     RECT  668.26 624.44 671.14 1249.18 ;
     RECT  671.14 625.28 672.1 1249.18 ;
     RECT  666.82 519.44 677.86 532.24 ;
     RECT  644.26 436.28 682.18 479.32 ;
     RECT  662.98 611.42 687.94 612.88 ;
     RECT  644.26 370.76 689.86 423.88 ;
     RECT  689.86 370.76 691.78 406.24 ;
     RECT  621.7 489.2 692.74 494.44 ;
     RECT  672.1 625.28 693.22 1248.76 ;
     RECT  693.22 625.28 693.7 1237.42 ;
     RECT  677.86 522.8 696.58 532.24 ;
     RECT  693.7 625.28 702.62 1234.48 ;
     RECT  693.22 1248.56 702.82 1248.76 ;
     RECT  702.62 625.28 707.42 1235.32 ;
     RECT  707.42 625.28 712.7 1237 ;
     RECT  712.7 625.28 720.38 1242.04 ;
     RECT  720.38 625.28 722.78 1242.46 ;
     RECT  682.18 441.32 725.86 479.32 ;
     RECT  722.78 625.28 733.82 1242.88 ;
     RECT  733.82 621.08 739.945 1242.88 ;
     RECT  725.86 474.08 741.22 479.32 ;
     RECT  620.74 558.5 741.5 581.38 ;
     RECT  741.02 590.42 741.7 590.62 ;
     RECT  687.94 611.42 742.825 611.62 ;
     RECT  739.945 621.065 742.825 1242.88 ;
     RECT  742.825 611.42 750.08 1242.88 ;
     RECT  750.08 611.42 752.54 1245.99 ;
     RECT  752.54 611.42 753.7 1249.6 ;
     RECT  741.22 476.6 754.66 479.32 ;
     RECT  754.66 479.12 760.42 479.32 ;
     RECT  753.7 621.92 767.14 1249.6 ;
     RECT  767.14 621.92 767.65 1249.215 ;
     RECT  767.65 621.92 779.14 1249.18 ;
     RECT  779.14 643.745 780.035 1249.18 ;
     RECT  780.035 644.58 780.485 1249.18 ;
     RECT  780.485 645.44 780.86 1249.18 ;
     RECT  779.14 621.92 781.06 635.14 ;
     RECT  780.86 645.44 783.26 1252.96 ;
     RECT  783.26 645.44 785.86 1253.8 ;
     RECT  785.86 645.44 787.78 1249.18 ;
     RECT  787.78 645.86 790.18 1249.18 ;
     RECT  790.18 660.56 791.605 1249.18 ;
     RECT  791.605 660.56 794.02 1248.34 ;
     RECT  794.02 663.08 794.5 1248.34 ;
     RECT  781.06 629.9 798.505 635.14 ;
     RECT  794.5 663.5 800.06 1248.34 ;
     RECT  800.06 663.5 800.74 1249.6 ;
     RECT  790.18 645.86 801.02 647.74 ;
     RECT  800.74 664.34 801.22 1249.215 ;
     RECT  801.22 668.12 801.25 1249.215 ;
     RECT  801.02 645.86 801.7 649.42 ;
     RECT  639.94 600.5 802.46 600.7 ;
     RECT  725.86 441.32 802.66 464.2 ;
     RECT  801.7 645.86 803.14 648.16 ;
     RECT  801.25 668.12 804.1 1249.18 ;
     RECT  798.505 628.625 805.955 635.14 ;
     RECT  804.1 669.8 806.02 1249.18 ;
     RECT  803.14 645.86 806.3 647.74 ;
     RECT  805.955 629.46 806.405 635.14 ;
     RECT  806.3 644.18 806.5 647.74 ;
     RECT  802.46 592.52 808.7 600.7 ;
     RECT  753.7 611.42 808.7 611.62 ;
     RECT  806.405 629.48 810.34 635.14 ;
     RECT  808.7 592.52 810.62 611.62 ;
     RECT  810.34 630.32 810.62 635.14 ;
     RECT  806.5 644.18 810.62 646.06 ;
     RECT  810.62 630.32 810.82 646.06 ;
     RECT  806.02 669.8 810.82 1047.16 ;
     RECT  810.62 591.68 811.3 611.62 ;
     RECT  806.02 1055.78 813.02 1249.18 ;
     RECT  810.82 644.18 814.18 646.06 ;
     RECT  810.82 670.64 814.46 1047.16 ;
     RECT  813.02 1055.78 814.46 1249.6 ;
     RECT  814.46 670.64 815.42 1249.6 ;
     RECT  815.42 670.64 817.06 1250.02 ;
     RECT  817.06 670.64 819.94 1244.98 ;
     RECT  621.7 506.84 820.7 507.04 ;
     RECT  660.1 543.8 820.7 548.62 ;
     RECT  741.5 558.5 820.7 581.8 ;
     RECT  814.18 645.86 820.7 646.06 ;
     RECT  692.74 491.72 820.9 494.44 ;
     RECT  820.7 506.42 820.9 507.04 ;
     RECT  696.58 522.8 820.9 529.72 ;
     RECT  811.3 597.14 820.9 611.62 ;
     RECT  819.94 675.26 827.14 1244.98 ;
     RECT  820.7 645.86 827.9 646.9 ;
     RECT  827.9 643.76 828.38 652.78 ;
     RECT  827.14 675.26 829.34 1234.49 ;
     RECT  810.82 630.32 830.3 635.14 ;
     RECT  828.38 643.76 830.3 656.98 ;
     RECT  820.9 597.14 830.78 609.52 ;
     RECT  830.78 597.14 831.26 618.76 ;
     RECT  830.3 629.9 831.26 656.98 ;
     RECT  820.7 543.8 837.02 581.8 ;
     RECT  820.9 506.42 837.5 506.62 ;
     RECT  837.02 543.8 837.5 583.48 ;
     RECT  837.5 543.8 838.94 584.32 ;
     RECT  831.26 597.14 838.94 656.98 ;
     RECT  837.5 506.42 839.42 512.08 ;
     RECT  829.34 674.42 840.005 1234.49 ;
     RECT  802.66 441.32 840.1 449.08 ;
     RECT  838.94 543.8 840.265 659.92 ;
     RECT  840.005 674.42 840.565 1231.12 ;
     RECT  820.9 491.72 840.86 494.02 ;
     RECT  839.42 504.74 840.86 512.08 ;
     RECT  820.9 522.8 840.86 528.04 ;
     RECT  840.265 543.8 840.86 660.34 ;
     RECT  840.86 543.8 841.34 661.18 ;
     RECT  840.565 674.42 841.34 727.12 ;
     RECT  840.86 487.94 841.82 494.02 ;
     RECT  841.82 485 842.3 494.02 ;
     RECT  840.86 504.74 842.3 528.04 ;
     RECT  840.1 445.1 842.5 449.08 ;
     RECT  840.565 735.74 842.5 1231.12 ;
     RECT  842.3 485 842.725 528.04 ;
     RECT  842.725 481.64 843.26 528.04 ;
     RECT  843.26 481.22 844.22 528.04 ;
     RECT  841.34 543.8 846.06 727.12 ;
     RECT  846.06 539.18 846.835 727.12 ;
     RECT  844.22 475.34 847.1 528.04 ;
     RECT  847.1 474.08 847.58 528.04 ;
     RECT  846.835 538.34 847.58 727.12 ;
     RECT  847.58 474.08 850.46 727.12 ;
     RECT  842.5 735.74 850.46 1230.28 ;
     RECT  850.46 474.08 855.2 1230.28 ;
     RECT  855.2 474.08 857.18 1230.87 ;
     RECT  857.18 474.08 857.86 1234.48 ;
     RECT  842.5 445.52 858.34 449.08 ;
     RECT  857.86 474.08 858.37 1234.095 ;
     RECT  802.66 458.96 858.62 464.2 ;
     RECT  858.37 474.08 858.62 1234.06 ;
     RECT  858.62 458.96 865.525 1234.06 ;
     RECT  865.525 458.96 868.7 1229.86 ;
     RECT  858.34 445.52 872.06 446.56 ;
     RECT  868.7 456.02 872.06 1229.86 ;
     RECT  691.78 370.76 872.74 401.2 ;
     RECT  872.06 444.26 873.92 1229.86 ;
     RECT  873.92 444.225 874.94 1229.86 ;
     RECT  874.94 443.84 877.82 1229.86 ;
     RECT  877.82 443.84 881.66 1231.12 ;
     RECT  881.66 436.28 881.86 1231.12 ;
     RECT  881.86 436.28 883.1 1230.7 ;
     RECT  883.1 435.86 883.98 1230.7 ;
     RECT  883.98 433.34 884.755 1230.7 ;
     RECT  689.86 416.12 885.98 423.88 ;
     RECT  884.755 432.5 885.98 1230.7 ;
     RECT  872.74 370.76 893.86 398.68 ;
     RECT  885.98 416.12 898.18 1230.7 ;
     RECT  898.18 418.64 901.54 1230.7 ;
     RECT  893.86 380.84 905.86 398.68 ;
     RECT  901.54 422.84 914.78 1230.7 ;
     RECT  914.78 421.16 921.7 1230.7 ;
     RECT  921.7 421.545 921.92 1230.7 ;
     RECT  905.86 380.84 924.1 388.6 ;
     RECT  921.92 421.545 926.05 1230.87 ;
     RECT  926.05 421.58 935.62 1230.87 ;
     RECT  935.62 421.58 935.9 993.4 ;
     RECT  935.62 1003.7 936.38 1230.87 ;
     RECT  936.38 1003.7 937.82 1231.12 ;
     RECT  937.82 1003.7 938.3 1233.22 ;
     RECT  935.9 414.02 939.46 993.4 ;
     RECT  939.46 414.02 940.22 978.28 ;
     RECT  938.3 1003.7 940.42 1234.48 ;
     RECT  940.22 413.6 941.18 978.28 ;
     RECT  939.46 988.16 944.06 993.4 ;
     RECT  940.42 1003.7 944.06 1234.06 ;
     RECT  941.18 413.18 945.5 978.28 ;
     RECT  945.5 412.76 945.7 978.28 ;
     RECT  944.06 988.16 947.9 1234.06 ;
     RECT  945.7 413.18 948.38 978.28 ;
     RECT  947.9 987.74 948.38 1234.06 ;
     RECT  948.38 413.18 950.5 1234.06 ;
     RECT  950.5 413.18 957.7 1230.28 ;
     RECT  957.7 413.18 958.94 1218.94 ;
     RECT  958.94 412.76 959.14 1218.94 ;
     RECT  959.14 413.18 960.085 1218.94 ;
     RECT  960.085 413.18 963.46 1218.1 ;
     RECT  963.46 413.18 963.94 1211.8 ;
     RECT  963.94 413.6 964.9 1211.8 ;
     RECT  964.9 1191.44 965.38 1211.8 ;
     RECT  964.9 413.6 967.78 1182.4 ;
     RECT  967.78 1175.9 969.22 1182.4 ;
     RECT  965.38 1195.22 969.22 1211.8 ;
     RECT  969.22 1195.22 969.7 1210.54 ;
     RECT  969.7 1195.22 970.66 1201.3 ;
     RECT  969.22 1175.9 972.1 1177.95 ;
     RECT  967.78 413.6 973.06 1167.28 ;
     RECT  973.06 413.6 973.54 1166.45 ;
     RECT  973.54 413.6 974.81 1155.94 ;
     RECT  974.81 413.26 974.88 1155.94 ;
     RECT  973.54 1165.385 974.915 1166.45 ;
     RECT  974.915 1166.22 975.365 1166.45 ;
     RECT  972.1 1176.32 975.445 1177.95 ;
     RECT  970.66 1195.22 976.42 1200.895 ;
     RECT  975.445 1176.32 978.82 1176.52 ;
     RECT  974.88 413.18 979.1 1155.94 ;
     RECT  976.42 1197.32 979.1 1200.895 ;
     RECT  975.365 1166.24 979.3 1166.44 ;
     RECT  979.1 1197.32 979.3 1202.98 ;
     RECT  957.7 1230.08 979.3 1230.28 ;
     RECT  979.3 1199.42 980.26 1202.14 ;
     RECT  979.1 409.82 982.18 1155.94 ;
     RECT  982.18 412.76 983.42 1155.94 ;
     RECT  983.42 412.76 985.06 1157.2 ;
     RECT  985.06 413.26 985.82 1157.2 ;
     RECT  985.82 413.26 987.74 1158.88 ;
     RECT  987.74 413.26 989.66 1163.08 ;
     RECT  989.66 413.26 989.68 1169.8 ;
     RECT  989.68 413.6 991.1 1169.8 ;
     RECT  991.1 413.6 994.94 1173.16 ;
     RECT  994.94 413.6 995.9 1174 ;
     RECT  995.9 413.6 996.1 1176.94 ;
     RECT  996.1 421.16 996.38 1176.94 ;
     RECT  996.38 421.16 996.58 1184.08 ;
     RECT  996.58 421.58 999.74 1184.08 ;
     RECT  999.74 421.58 1002.325 1185.34 ;
     RECT  1002.325 425.15 1004.5 1185.34 ;
     RECT  1004.5 425.36 1005.02 1185.34 ;
     RECT  1005.02 425.36 1009.54 1192.06 ;
     RECT  1009.54 427.88 1010.78 1192.06 ;
     RECT  1010.78 427.88 1015.1 1192.9 ;
     RECT  1015.1 427.88 1015.58 1195 ;
     RECT  1015.58 427.88 1015.78 1196.68 ;
     RECT  1015.78 427.88 1021.06 1196.26 ;
     RECT  1021.06 427.88 1023.46 1193.32 ;
     RECT  1023.46 429.56 1030.66 1193.32 ;
     RECT  1030.66 438.38 1032.58 1193.32 ;
     RECT  1032.58 439.64 1035.46 1193.32 ;
     RECT  1030.66 429.56 1036.42 429.76 ;
     RECT  1035.46 440.48 1040.26 1193.32 ;
     RECT  1040.26 440.48 1041.22 1189.54 ;
     RECT  905.86 398.48 1041.7 398.68 ;
     RECT  1041.22 440.48 1047.46 1186.18 ;
     RECT  1047.46 458.96 1048.42 1186.18 ;
     RECT  1048.42 462.57 1052.26 1186.18 ;
     RECT  1052.26 462.57 1052.725 1185.76 ;
     RECT  1052.725 462.74 1054.66 1185.76 ;
     RECT  924.1 380.84 1057.06 381.04 ;
     RECT  1047.46 440.48 1058.02 449.5 ;
     RECT  1054.66 465.68 1058.02 1185.76 ;
     RECT  1058.02 465.68 1060.42 533.92 ;
     RECT  1060.42 466.94 1066.94 533.92 ;
     RECT  1058.02 542.54 1066.94 1185.76 ;
     RECT  1066.94 466.94 1071.46 1185.76 ;
     RECT  1058.02 445.1 1072.9 449.5 ;
     RECT  1071.46 486.26 1072.9 1185.76 ;
     RECT  1072.9 486.68 1081.06 1183.66 ;
     RECT  1071.46 466.94 1082.5 473.44 ;
     RECT  1081.06 486.68 1089.7 1183.24 ;
     RECT  1089.7 496.76 1090.66 1183.24 ;
     RECT  893.86 370.76 1092.1 370.96 ;
     RECT  1090.66 499.7 1092.58 1183.24 ;
     RECT  1082.5 466.94 1094.3 467.14 ;
     RECT  1094.3 466.94 1094.5 467.98 ;
     RECT  1092.58 503.48 1097.86 1183.24 ;
     RECT  1094.5 467.78 1103.14 467.98 ;
     RECT  1097.86 503.9 1108.42 1183.24 ;
     RECT  1089.7 486.68 1112.26 486.88 ;
     RECT  1072.9 445.1 1120.42 445.3 ;
     RECT  1108.42 504.32 1123.3 1183.24 ;
     RECT  1123.3 504.32 1130.5 1182.4 ;
     RECT  1130.5 1182.2 1141.06 1182.4 ;
     RECT  1130.5 504.32 1142.02 1171.48 ;
     RECT  1142.02 522.785 1143.94 1171.48 ;
     RECT  1142.02 504.32 1146.34 513.34 ;
     RECT  1143.94 522.785 1153.285 1168.12 ;
     RECT  1153.285 522.785 1153.475 1169.38 ;
     RECT  1153.475 523.62 1153.925 1169.38 ;
     RECT  1153.925 523.64 1154.5 1169.38 ;
     RECT  1154.5 526.58 1154.78 1169.38 ;
     RECT  1154.78 526.58 1155.94 1169.8 ;
     RECT  1155.94 530.78 1160.26 1169.38 ;
     RECT  1160.26 1153.64 1161.22 1168.54 ;
     RECT  1161.22 1154.06 1163.62 1168.54 ;
     RECT  1163.62 1154.48 1165.54 1159.72 ;
     RECT  1165.54 1155.74 1166.02 1159.72 ;
     RECT  1160.26 530.78 1166.5 1144.6 ;
     RECT  1166.02 1158.68 1167.22 1159.72 ;
     RECT  1167.22 1158.68 1167.94 1158.88 ;
     RECT  1163.62 1168.34 1167.94 1168.54 ;
     RECT  1146.34 504.32 1168.42 511.66 ;
     RECT  1166.5 532.46 1168.9 1144.6 ;
     RECT  1168.9 1144.4 1170.82 1144.6 ;
     RECT  1168.9 532.46 1171.3 1125.28 ;
     RECT  1168.42 507.26 1174.18 511.66 ;
     RECT  1171.3 532.46 1176.38 1124.86 ;
     RECT  1176.38 532.04 1176.58 1124.86 ;
     RECT  1176.58 532.04 1180.9 1123.6 ;
     RECT  1180.9 532.04 1181.14 1120.66 ;
     RECT  1181.14 532.04 1181.86 1117.72 ;
     RECT  1181.86 532.04 1183.3 1116.04 ;
     RECT  1183.3 532.04 1184.74 1113.94 ;
     RECT  1184.74 532.04 1186.66 1112.68 ;
     RECT  1186.66 532.04 1188.1 1111 ;
     RECT  1188.1 532.04 1189.54 1110.58 ;
     RECT  1189.54 1081.82 1190.02 1109.32 ;
     RECT  1190.02 1081.82 1190.74 1108.48 ;
     RECT  1189.54 532.04 1190.98 1072.78 ;
     RECT  1190.98 532.04 1191.46 1072.36 ;
     RECT  1191.46 532.04 1192.7 1071.94 ;
     RECT  1190.74 1081.82 1194.82 1107.22 ;
     RECT  1192.7 527.42 1195.3 1071.94 ;
     RECT  1195.3 527.42 1196.06 1066.06 ;
     RECT  1194.82 1083.08 1196.26 1107.22 ;
     RECT  1196.06 526.58 1197.02 1066.06 ;
     RECT  1174.18 507.26 1197.5 507.46 ;
     RECT  1197.02 524.06 1197.92 1066.06 ;
     RECT  1197.5 504.74 1197.98 507.46 ;
     RECT  1197.98 504.74 1198.4 508.3 ;
     RECT  1197.02 495.92 1199.42 496.12 ;
     RECT  1198.4 504.705 1199.42 508.3 ;
     RECT  1199.42 495.92 1199.9 512.5 ;
     RECT  1197.92 523.05 1199.9 1066.06 ;
     RECT  1196.26 1091.9 1200.58 1107.22 ;
     RECT  1200.58 1094 1201.06 1097.56 ;
     RECT  1200.58 1107.02 1201.54 1107.22 ;
     RECT  1201.06 1094.21 1202.02 1097.56 ;
     RECT  1199.9 495.92 1203.46 1066.06 ;
     RECT  1203.46 495.92 1203.94 1062.28 ;
     RECT  1203.94 495.92 1204.9 1058.92 ;
     RECT  1204.9 495.92 1207.3 1055.98 ;
     RECT  1207.3 496.76 1216.7 1049.43 ;
     RECT  1216.7 496.76 1217.66 1049.68 ;
     RECT  1217.66 492.98 1221.02 1049.68 ;
     RECT  1221.02 492.14 1223.14 1049.68 ;
     RECT  1223.14 492.14 1223.9 1046.74 ;
     RECT  1223.9 491.72 1226.5 1046.74 ;
     RECT  1226.5 491.72 1226.98 1045.48 ;
     RECT  1226.98 1036.88 1229.38 1045.48 ;
     RECT  1229.38 1037.72 1231.3 1045.48 ;
     RECT  1231.3 1037.72 1234.18 1037.92 ;
     RECT  1226.98 491.72 1245.98 1027.84 ;
     RECT  1240.7 476.6 1255.58 476.8 ;
     RECT  1245.98 487.94 1260.38 1027.84 ;
     RECT  1260.38 487.94 1262.3 1029.1 ;
     RECT  1260.38 1046.12 1263.74 1046.32 ;
     RECT  1255.58 476.6 1264.22 479.32 ;
     RECT  1262.3 487.94 1264.22 1030.36 ;
     RECT  1264.22 476.6 1265.18 1030.36 ;
     RECT  1265.18 476.6 1265.66 1031.2 ;
     RECT  1265.66 476.6 1268.5 1033.72 ;
     RECT  1268.5 621.5 1268.73 1033.72 ;
     RECT  1268.73 621.5 1270.41 852.7 ;
     RECT  1268.5 476.6 1271.62 611.62 ;
     RECT  1268.73 863 1272.1 1033.72 ;
     RECT  1271.62 611.42 1273.06 611.62 ;
     RECT  1272.1 863 1273.06 889.66 ;
     RECT  1272.1 898.7 1273.06 1033.72 ;
     RECT  1271.62 476.6 1273.54 601.96 ;
     RECT  1270.41 621.92 1273.54 852.7 ;
     RECT  1273.06 863 1273.54 877.48 ;
     RECT  1273.06 898.7 1273.54 937.96 ;
     RECT  1273.06 947.84 1273.54 961.06 ;
     RECT  1273.06 970.52 1273.82 1033.72 ;
     RECT  1263.74 1043.6 1273.82 1046.32 ;
     RECT  1273.54 621.92 1274.02 670.84 ;
     RECT  1273.54 679.88 1274.02 852.7 ;
     RECT  1273.54 476.6 1274.5 595.24 ;
     RECT  1273.54 863 1274.5 876.64 ;
     RECT  1273.06 886.52 1274.5 889.66 ;
     RECT  1274.5 579.08 1274.98 595.24 ;
     RECT  1274.5 886.52 1274.98 888.82 ;
     RECT  1273.82 970.52 1283.9 1046.32 ;
     RECT  1274.5 476.6 1288.7 570.04 ;
     RECT  1274.98 582.44 1288.7 595.24 ;
     RECT  1274.02 623.18 1288.7 670.84 ;
     RECT  1274.02 679.88 1288.7 833.8 ;
     RECT  1274.5 863.42 1288.7 876.64 ;
     RECT  1273.54 899.96 1288.7 937.96 ;
     RECT  1273.54 947.84 1288.7 960.64 ;
     RECT  1283.9 970.52 1288.7 1053.88 ;
     RECT  1274.98 887.36 1289.18 888.82 ;
     RECT  1288.7 897.44 1289.18 1053.88 ;
     RECT  1288.7 582.44 1290.14 602.8 ;
     RECT  1290.14 582.44 1292.54 607.84 ;
     RECT  1274.02 849.56 1293.02 852.7 ;
     RECT  1288.7 862.16 1293.02 876.64 ;
     RECT  1293.02 849.56 1293.5 876.64 ;
     RECT  1289.18 887.36 1293.5 1053.88 ;
     RECT  1292.54 582.44 1294.46 612.88 ;
     RECT  1288.7 622.76 1294.46 833.8 ;
     RECT  1293.5 849.56 1294.46 1053.88 ;
     RECT  1288.7 469.04 1295.9 570.04 ;
     RECT  1295.9 469.04 1296.38 572.56 ;
     RECT  1294.46 582.44 1296.38 1053.88 ;
     RECT  1296.38 469.04 1299.36 1053.88 ;
     RECT  1299.36 487.94 1299.46 518.38 ;
     RECT  1299.36 533.3 1299.46 564.16 ;
     RECT  1299.36 661.82 1299.46 662.86 ;
     RECT  1299.36 681.14 1299.46 681.34 ;
     RECT  1299.36 708.86 1299.46 718.3 ;
     RECT  1299.36 731.54 1299.46 738.46 ;
     RECT  1299.36 755.9 1299.46 763.24 ;
     RECT  1299.36 784.46 1299.46 801.04 ;
     RECT  1299.36 867.62 1299.46 869.08 ;
     RECT  1299.36 888.62 1299.46 889.66 ;
     RECT  1299.36 933.56 1299.46 935.02 ;
     RECT  1299.36 988.58 1299.46 1014.82 ;
     RECT  1299.36 1024.28 1299.46 1025.74 ;
    LAYER Metal3 ;
     RECT  694.94 375.8 695.14 390.92 ;
     RECT  690.14 390.92 695.14 393.44 ;
     RECT  866.78 383.36 866.98 401 ;
     RECT  979.1 409.82 979.3 410.24 ;
     RECT  979.1 410.24 982.66 410.66 ;
     RECT  979.1 410.66 983.14 412.76 ;
     RECT  979.1 412.76 985.06 413.6 ;
     RECT  940.22 413.6 963.94 414.02 ;
     RECT  979.1 413.6 995.62 414.02 ;
     RECT  893.66 373.28 893.86 416.12 ;
     RECT  905.66 395.96 905.86 416.12 ;
     RECT  940.22 414.02 995.62 417.38 ;
     RECT  893.66 416.12 905.86 417.5 ;
     RECT  938.3 417.38 996.1 420.74 ;
     RECT  893.66 417.5 906.34 421.16 ;
     RECT  923.9 388.4 924.1 421.16 ;
     RECT  937.82 420.74 996.1 421.16 ;
     RECT  893.66 421.16 926.98 421.58 ;
     RECT  937.82 421.16 996.58 421.58 ;
     RECT  893.66 421.58 996.58 422 ;
     RECT  893.66 422 1003.3 422.42 ;
     RECT  893.66 422.42 1005.7 424.94 ;
     RECT  893.66 424.94 1009.06 426.2 ;
     RECT  893.66 426.2 1010.02 428.72 ;
     RECT  1041.5 398.48 1041.7 429.56 ;
     RECT  641.66 426.2 641.86 431.24 ;
     RECT  893.66 428.72 1016.74 432.08 ;
     RECT  885.98 432.08 1016.74 432.92 ;
     RECT  626.78 385.88 626.98 433.76 ;
     RECT  641.66 431.24 644.26 433.76 ;
     RECT  885.98 432.92 1024.42 435.86 ;
     RECT  1036.22 429.56 1041.7 435.86 ;
     RECT  0.38 378.74 0.58 436.06 ;
     RECT  885.98 435.86 1041.7 436.28 ;
     RECT  626.78 433.76 644.26 438.8 ;
     RECT  884.06 436.28 1044.58 439.1 ;
     RECT  866.78 401 872.74 444.26 ;
     RECT  884.06 439.1 1045.06 444.26 ;
     RECT  866.78 444.26 1045.06 448.88 ;
     RECT  1091.9 370.76 1092.1 453.92 ;
     RECT  858.14 448.88 1045.06 459.38 ;
     RECT  1056.86 380.84 1057.06 459.38 ;
     RECT  858.14 459.38 1057.06 464 ;
     RECT  858.14 464 1058.02 466.1 ;
     RECT  858.14 466.1 1058.5 467.9 ;
     RECT  858.14 467.9 1058.98 471.14 ;
     RECT  1288.7 471.56 1288.9 472.18 ;
     RECT  1089.5 453.92 1092.1 473.24 ;
     RECT  839.9 441.32 840.1 474.08 ;
     RECT  858.14 471.14 1068.1 474.08 ;
     RECT  839.9 474.08 1068.1 486.26 ;
     RECT  1104.38 451.4 1104.58 486.68 ;
     RECT  1120.22 445.1 1120.42 486.68 ;
     RECT  1255.58 486.68 1255.78 487.94 ;
     RECT  839.9 486.26 1068.58 488.78 ;
     RECT  1082.3 473.24 1092.1 488.78 ;
     RECT  1255.58 487.94 1260.1 488.78 ;
     RECT  1255.58 488.78 1263.46 489.2 ;
     RECT  1253.18 489.2 1263.46 492.56 ;
     RECT  1253.18 492.56 1273.06 492.98 ;
     RECT  1247.9 492.98 1273.06 493.4 ;
     RECT  1218.14 492.98 1228.9 496.34 ;
     RECT  1197.02 495.92 1197.22 496.76 ;
     RECT  1218.14 496.34 1230.34 496.76 ;
     RECT  1244.06 493.4 1273.06 497.18 ;
     RECT  1197.02 496.76 1230.34 498.02 ;
     RECT  1240.7 497.18 1273.06 498.02 ;
     RECT  7.1 496.76 7.3 498.22 ;
     RECT  839.9 488.78 1092.1 500.96 ;
     RECT  1197.02 498.02 1273.06 501.8 ;
     RECT  839.9 500.96 1094.5 503.48 ;
     RECT  1104.38 486.68 1120.42 503.48 ;
     RECT  1197.02 501.8 1281.7 504.94 ;
     RECT  1255.58 504.94 1281.7 505.36 ;
     RECT  839.9 503.48 1120.42 508.94 ;
     RECT  1131.26 508.52 1131.46 508.94 ;
     RECT  1197.02 504.94 1245.22 508.94 ;
     RECT  608.54 428.72 608.74 509.36 ;
     RECT  619.58 438.8 644.26 509.36 ;
     RECT  839.9 508.94 1138.18 513.14 ;
     RECT  660.86 403.52 661.06 516.92 ;
     RECT  1195.58 508.94 1245.22 518.6 ;
     RECT  1255.58 505.36 1272.1 518.6 ;
     RECT  680.54 393.44 695.14 519.44 ;
     RECT  1195.58 518.6 1272.1 523.84 ;
     RECT  677.66 519.44 695.14 524.48 ;
     RECT  839.9 513.14 1146.34 526.58 ;
     RECT  1195.58 523.84 1245.22 527.42 ;
     RECT  839.9 526.58 1155.94 528.26 ;
     RECT  839.9 528.26 1159.3 530.78 ;
     RECT  1169.66 484.16 1169.86 530.78 ;
     RECT  839.9 530.78 1169.86 532.04 ;
     RECT  660.86 516.92 661.54 534.56 ;
     RECT  1184.06 534.14 1184.26 534.56 ;
     RECT  1195.1 527.42 1245.22 534.56 ;
     RECT  1256.06 523.84 1272.1 534.56 ;
     RECT  660.86 534.56 666.82 537.08 ;
     RECT  754.46 476.6 754.66 539.9 ;
     RECT  754.46 539.9 755.14 540.1 ;
     RECT  839.9 532.04 1174.18 541.7 ;
     RECT  1184.06 534.56 1272.1 541.7 ;
     RECT  838.94 541.7 1272.1 542.32 ;
     RECT  659.9 537.08 666.82 544.64 ;
     RECT  677.66 524.48 700.9 544.64 ;
     RECT  838.94 542.32 1266.82 546.94 ;
     RECT  1186.46 546.94 1266.82 550.3 ;
     RECT  838.94 546.94 1175.14 561.02 ;
     RECT  838.94 561.02 1179.46 562.28 ;
     RECT  1191.74 550.3 1266.82 562.28 ;
     RECT  838.94 562.28 1266.82 564.38 ;
     RECT  1.34 569.42 1.54 569.84 ;
     RECT  838.94 564.38 1271.14 574.04 ;
     RECT  838.94 574.04 1272.58 574.46 ;
     RECT  838.94 574.46 1273.54 577.4 ;
     RECT  1295.9 572.36 1296.1 579.92 ;
     RECT  838.46 577.4 1273.54 580.12 ;
     RECT  838.46 580.12 1271.62 580.54 ;
     RECT  608.54 509.36 644.26 582.44 ;
     RECT  606.62 582.44 644.26 590 ;
     RECT  659.9 544.64 700.9 590 ;
     RECT  802.46 456.44 802.66 592.1 ;
     RECT  802.46 592.1 809.38 592.72 ;
     RECT  838.46 580.54 1267.3 597.14 ;
     RECT  835.1 597.14 1267.3 598.4 ;
     RECT  835.1 598.4 1269.22 599.44 ;
     RECT  1281.5 592.52 1281.7 602.6 ;
     RECT  1295.9 579.92 1298.98 602.6 ;
     RECT  754.94 540.1 755.14 604.7 ;
     RECT  809.18 592.72 809.38 607.64 ;
     RECT  835.1 599.44 1268.26 610.16 ;
     RECT  833.66 610.16 1268.26 613.3 ;
     RECT  833.66 613.3 1264.9 614.56 ;
     RECT  754.94 604.7 760.42 617.72 ;
     RECT  835.1 614.56 1264.9 617.92 ;
     RECT  808.7 607.64 809.38 620.66 ;
     RECT  1281.5 602.6 1298.98 622.96 ;
     RECT  741.02 590.42 741.22 624.44 ;
     RECT  753.5 617.72 760.42 624.44 ;
     RECT  741.02 624.44 760.42 625.28 ;
     RECT  1.34 569.84 5.38 626.12 ;
     RECT  734.78 625.28 760.42 627.8 ;
     RECT  730.94 627.8 760.42 629.06 ;
     RECT  606.62 590 700.9 629.48 ;
     RECT  716.54 629.06 760.42 629.48 ;
     RECT  1281.5 622.96 1281.7 630.1 ;
     RECT  606.62 629.48 760.42 632.42 ;
     RECT  836.54 617.92 1264.9 632.42 ;
     RECT  798.62 632.42 798.82 632.84 ;
     RECT  808.7 620.66 812.26 632.84 ;
     RECT  798.62 632.84 812.26 634.72 ;
     RECT  606.62 632.42 762.34 635.36 ;
     RECT  836.54 632.42 1266.82 636.82 ;
     RECT  606.14 635.36 762.34 637.46 ;
     RECT  837.98 636.82 1266.82 637.88 ;
     RECT  0.86 626.12 5.38 638.3 ;
     RECT  606.14 637.46 768.58 640.4 ;
     RECT  0.86 638.3 7.3 640.6 ;
     RECT  606.14 640.4 769.54 640.82 ;
     RECT  780.86 621.92 781.06 640.82 ;
     RECT  1295.9 622.96 1298.98 642.92 ;
     RECT  606.14 640.82 781.06 645.44 ;
     RECT  837.98 637.88 1270.66 647.96 ;
     RECT  806.78 634.72 812.26 649.22 ;
     RECT  1290.62 642.92 1298.98 650.48 ;
     RECT  837.98 647.96 1272.1 651.74 ;
     RECT  829.82 651.74 1272.1 652.36 ;
     RECT  606.14 645.44 787.78 653 ;
     RECT  1288.7 650.48 1298.98 658.24 ;
     RECT  1289.18 658.24 1298.98 659.5 ;
     RECT  606.14 653 790.18 663.08 ;
     RECT  801.5 649.22 812.26 663.08 ;
     RECT  829.82 652.36 1270.66 667.28 ;
     RECT  606.14 663.08 812.26 669.8 ;
     RECT  1289.66 659.5 1298.98 670.64 ;
     RECT  1281.5 670.64 1298.98 671.26 ;
     RECT  606.14 669.8 813.22 674.42 ;
     RECT  829.82 667.28 1271.14 674.84 ;
     RECT  606.14 674.42 814.66 675.68 ;
     RECT  827.42 674.84 1271.62 675.68 ;
     RECT  1281.5 671.26 1298.5 676.72 ;
     RECT  606.14 675.68 1271.62 693.32 ;
     RECT  1288.7 676.72 1298.5 698.56 ;
     RECT  606.14 693.32 1272.1 700.88 ;
     RECT  0.86 640.6 5.38 715.58 ;
     RECT  606.14 700.88 1281.7 717.04 ;
     RECT  606.14 717.04 1274.02 720.4 ;
     RECT  1293.5 698.56 1298.5 723.56 ;
     RECT  0.86 715.58 7.3 723.76 ;
     RECT  1288.7 723.56 1298.5 726.92 ;
     RECT  606.14 720.4 1143.94 727.12 ;
     RECT  0.86 723.76 1.06 728.8 ;
     RECT  851.9 727.12 1143.94 730.7 ;
     RECT  1153.82 720.4 1274.02 730.7 ;
     RECT  1288.7 726.92 1298.98 731.54 ;
     RECT  1288.7 731.54 1299.46 738.04 ;
     RECT  606.14 727.12 840.58 739.1 ;
     RECT  606.14 739.1 842.02 739.94 ;
     RECT  851.9 730.7 1274.02 739.94 ;
     RECT  4.22 736.16 4.42 743.92 ;
     RECT  606.14 739.94 1274.02 751.48 ;
     RECT  606.14 751.48 802.18 755.06 ;
     RECT  1293.5 738.04 1299.46 756.1 ;
     RECT  605.66 755.06 802.18 763.04 ;
     RECT  605.66 763.04 803.14 764.3 ;
     RECT  813.5 751.48 1274.02 764.3 ;
     RECT  605.66 764.3 1274.02 776.26 ;
     RECT  606.14 776.26 1274.02 777.52 ;
     RECT  606.62 777.52 1274.02 779.62 ;
     RECT  608.54 779.62 1274.02 780.88 ;
     RECT  609.02 780.88 1274.02 781.3 ;
     RECT  609.5 781.3 1274.02 781.72 ;
     RECT  614.78 781.72 1274.02 791.8 ;
     RECT  614.78 791.8 623.14 792.02 ;
     RECT  633.5 791.8 738.34 798.52 ;
     RECT  614.3 792.02 623.14 799.36 ;
     RECT  662.78 798.52 738.34 802.94 ;
     RECT  751.58 791.8 1274.02 803.56 ;
     RECT  572.06 803.36 572.26 803.78 ;
     RECT  569.66 803.78 572.26 804.2 ;
     RECT  614.3 799.36 614.5 806.72 ;
     RECT  633.5 798.52 652.42 806.72 ;
     RECT  569.66 804.2 581.38 807.98 ;
     RECT  595.58 806.72 597.22 807.98 ;
     RECT  610.94 806.72 614.5 807.98 ;
     RECT  662.78 802.94 740.74 807.98 ;
     RECT  751.58 803.56 1273.54 807.98 ;
     RECT  569.66 807.98 583.3 810.5 ;
     RECT  595.58 807.98 614.5 810.5 ;
     RECT  569.66 810.5 614.5 810.92 ;
     RECT  561.5 810.92 614.5 811.34 ;
     RECT  625.34 806.72 652.42 811.34 ;
     RECT  662.78 807.98 1273.54 811.34 ;
     RECT  558.14 811.34 614.5 813.86 ;
     RECT  625.34 811.34 1273.54 814.06 ;
     RECT  553.82 813.86 615.46 814.28 ;
     RECT  625.34 814.06 722.02 814.28 ;
     RECT  733.34 814.06 1273.54 821.62 ;
     RECT  553.82 814.28 722.02 821.84 ;
     RECT  548.06 821.84 722.02 825.2 ;
     RECT  733.34 821.62 777.22 825.2 ;
     RECT  788.06 821.62 1273.54 826.66 ;
     RECT  548.06 825.2 777.22 833.6 ;
     RECT  788.54 826.66 1273.54 837.38 ;
     RECT  547.1 833.6 777.22 841.16 ;
     RECT  788.54 837.38 1274.02 841.16 ;
     RECT  547.1 841.16 1274.02 844.72 ;
     RECT  1293.5 756.1 1298.98 857.32 ;
     RECT  547.1 844.72 1267.78 860.06 ;
     RECT  543.74 860.06 1267.78 863.62 ;
     RECT  1293.5 857.32 1298.5 874.34 ;
     RECT  543.74 863.62 1265.86 878.96 ;
     RECT  543.26 878.96 1265.86 882.32 ;
     RECT  1289.18 874.34 1298.5 882.74 ;
     RECT  539.9 882.32 1267.3 885.46 ;
     RECT  539.9 885.46 1265.38 886.72 ;
     RECT  1288.7 882.74 1298.5 897.64 ;
     RECT  541.82 886.72 1262.98 902.48 ;
     RECT  541.82 902.48 1272.1 904.78 ;
     RECT  541.82 904.78 1267.3 905 ;
     RECT  1298.3 897.64 1298.5 912.76 ;
     RECT  537.98 905 1267.3 919.48 ;
     RECT  541.82 919.48 1267.3 947.2 ;
     RECT  547.1 947.2 1267.3 962.32 ;
     RECT  1289.18 961.28 1289.38 963.8 ;
     RECT  569.18 962.32 1267.3 964.22 ;
     RECT  1288.7 963.8 1289.38 965.68 ;
     RECT  1288.7 965.68 1288.9 968.2 ;
     RECT  548.54 962.32 559.3 969.46 ;
     RECT  549.02 969.46 559.3 969.88 ;
     RECT  569.18 964.22 1269.22 972.4 ;
     RECT  556.22 969.88 559.3 974.3 ;
     RECT  569.18 972.4 1268.26 974.3 ;
     RECT  556.22 974.3 1268.26 983.74 ;
     RECT  557.66 983.74 1268.26 984.8 ;
     RECT  557.66 984.8 1268.74 985 ;
     RECT  1288.7 983.12 1288.9 989.2 ;
     RECT  562.46 985 1268.74 992.78 ;
     RECT  562.46 992.78 1274.02 1000.12 ;
     RECT  1256.54 1000.12 1274.02 1003.06 ;
     RECT  562.46 1000.12 1246.66 1003.28 ;
     RECT  561.98 1003.28 1246.66 1003.48 ;
     RECT  1257.5 1003.06 1274.02 1005.8 ;
     RECT  561.98 1003.48 1246.18 1006 ;
     RECT  1257.5 1005.8 1274.5 1006 ;
     RECT  1257.5 1006 1273.06 1013.36 ;
     RECT  563.42 1006 1246.18 1014.2 ;
     RECT  1256.06 1013.36 1273.06 1014.2 ;
     RECT  563.42 1014.2 1273.06 1018.6 ;
     RECT  564.38 1018.6 1273.06 1022.5 ;
     RECT  1244.06 1022.5 1273.06 1022.8 ;
     RECT  1247.9 1022.8 1273.06 1026.16 ;
     RECT  1257.02 1026.16 1273.06 1026.58 ;
     RECT  1262.3 1026.58 1273.06 1029.94 ;
     RECT  564.38 1022.5 1234.18 1030.36 ;
     RECT  1262.3 1029.94 1272.58 1030.36 ;
     RECT  1298.78 989.42 1298.98 1031.2 ;
     RECT  566.3 1030.36 588.1 1033.3 ;
     RECT  1265.66 1030.36 1265.86 1033.72 ;
     RECT  597.98 1030.36 1234.18 1037.92 ;
     RECT  567.74 1033.3 588.1 1041.08 ;
     RECT  597.98 1037.92 1231.3 1041.08 ;
     RECT  567.74 1041.08 1231.3 1044.86 ;
     RECT  561.5 1044.86 1231.3 1045.06 ;
     RECT  561.5 1045.06 1217.86 1045.48 ;
     RECT  1229.66 1045.06 1231.3 1045.48 ;
     RECT  1229.66 1045.48 1229.86 1046.32 ;
     RECT  562.46 1045.48 1217.86 1049.26 ;
     RECT  1216.7 1049.26 1216.9 1049.68 ;
     RECT  562.46 1049.26 1205.38 1055.98 ;
     RECT  562.46 1055.98 1204.9 1058.5 ;
     RECT  557.66 1059.98 558.34 1060.4 ;
     RECT  569.18 1058.5 1203.94 1060.6 ;
     RECT  1175.9 1060.6 1203.94 1062.28 ;
     RECT  1175.9 1062.28 1200.58 1063.54 ;
     RECT  556.7 1060.4 558.34 1063.76 ;
     RECT  1175.9 1063.54 1199.14 1063.96 ;
     RECT  1175.9 1063.96 1196.26 1065.64 ;
     RECT  553.82 1063.76 558.34 1067.54 ;
     RECT  552.86 1067.54 558.34 1070.9 ;
     RECT  569.18 1060.6 1165.54 1070.9 ;
     RECT  552.86 1070.9 1165.54 1071.32 ;
     RECT  1175.9 1065.64 1195.3 1071.32 ;
     RECT  551.42 1071.32 1195.3 1079.72 ;
     RECT  549.98 1079.72 1195.3 1083.5 ;
     RECT  549.02 1083.5 1195.3 1087.48 ;
     RECT  549.98 1087.48 1195.3 1090.42 ;
     RECT  551.42 1090.42 1195.3 1090.84 ;
     RECT  552.38 1090.84 1195.3 1093.58 ;
     RECT  552.38 1093.58 1196.74 1098.2 ;
     RECT  552.38 1098.2 1197.7 1101.56 ;
     RECT  552.38 1101.56 1200.58 1102.6 ;
     RECT  552.38 1102.6 1192.42 1104.7 ;
     RECT  552.38 1104.7 1190.5 1105.76 ;
     RECT  550.46 1105.76 1190.5 1108.48 ;
     RECT  550.46 1108.48 1188.1 1109.32 ;
     RECT  552.38 1109.32 1188.1 1109.74 ;
     RECT  552.86 1109.74 1188.1 1111 ;
     RECT  552.86 1111 1186.66 1112.68 ;
     RECT  552.86 1112.68 1184.74 1113.94 ;
     RECT  552.86 1113.94 1184.26 1114.36 ;
     RECT  552.86 1114.36 1180.9 1114.78 ;
     RECT  552.86 1114.78 962.5 1116.88 ;
     RECT  972.38 1114.78 1180.9 1123.6 ;
     RECT  552.86 1116.88 957.22 1124.24 ;
     RECT  972.38 1123.6 1176.1 1124.44 ;
     RECT  972.86 1124.44 1171.3 1125.28 ;
     RECT  550.46 1124.24 957.22 1127.6 ;
     RECT  549.5 1127.6 957.22 1136.42 ;
     RECT  972.86 1125.28 1170.82 1136.42 ;
     RECT  548.54 1136.42 957.22 1140.4 ;
     RECT  970.94 1136.42 1170.82 1141.24 ;
     RECT  970.94 1141.24 1160.26 1143.34 ;
     RECT  551.42 1140.4 957.22 1143.76 ;
     RECT  1170.62 1141.24 1170.82 1144.6 ;
     RECT  554.3 1143.76 957.22 1146.92 ;
     RECT  554.3 1146.92 958.18 1150.7 ;
     RECT  970.94 1143.34 1159.78 1150.7 ;
     RECT  554.3 1150.7 1159.78 1154.48 ;
     RECT  552.86 1154.48 1160.74 1154.9 ;
     RECT  552.86 1154.9 1163.14 1157.84 ;
     RECT  552.86 1157.84 1163.62 1158.88 ;
     RECT  1114.46 1158.88 1163.62 1159.3 ;
     RECT  1023.26 1158.88 1102.18 1160.98 ;
     RECT  989.18 1158.88 1010.98 1162.24 ;
     RECT  1114.46 1159.3 1163.14 1162.24 ;
     RECT  1114.94 1162.24 1163.14 1163.08 ;
     RECT  1119.26 1163.08 1163.14 1163.92 ;
     RECT  1126.94 1163.92 1163.14 1166.02 ;
     RECT  554.3 1158.88 975.94 1166.44 ;
     RECT  1023.26 1160.98 1101.22 1166.44 ;
     RECT  1127.9 1166.02 1163.14 1166.44 ;
     RECT  1127.9 1166.44 1160.26 1166.86 ;
     RECT  554.3 1166.44 973.06 1167.28 ;
     RECT  1127.9 1166.86 1141.06 1167.28 ;
     RECT  1127.9 1167.28 1139.62 1168.96 ;
     RECT  991.1 1162.24 1010.98 1169.18 ;
     RECT  1023.26 1166.44 1098.82 1169.18 ;
     RECT  1150.94 1166.86 1160.26 1169.38 ;
     RECT  1130.3 1168.96 1139.62 1169.8 ;
     RECT  1150.94 1169.38 1156.9 1169.8 ;
     RECT  1130.3 1169.8 1138.18 1170.22 ;
     RECT  1130.3 1170.22 1133.38 1171.48 ;
     RECT  991.1 1169.18 1098.82 1173.16 ;
     RECT  995.9 1173.16 1098.82 1176.74 ;
     RECT  995.9 1176.74 1099.78 1176.94 ;
     RECT  1130.3 1171.48 1130.5 1176.94 ;
     RECT  554.3 1167.28 967.3 1177.16 ;
     RECT  997.34 1176.94 1099.78 1177.16 ;
     RECT  997.34 1177.16 1101.7 1177.78 ;
     RECT  997.34 1177.78 1096.42 1181.14 ;
     RECT  554.3 1177.16 969.22 1181.56 ;
     RECT  1067.42 1181.14 1095.94 1181.56 ;
     RECT  1068.38 1181.56 1074.34 1181.98 ;
     RECT  1074.14 1181.98 1074.34 1182.4 ;
     RECT  1087.1 1181.56 1094.5 1182.4 ;
     RECT  554.3 1181.56 741.7 1184.08 ;
     RECT  997.34 1181.14 1056.58 1184.08 ;
     RECT  1000.22 1184.08 1056.58 1184.5 ;
     RECT  561.5 1184.08 741.7 1184.92 ;
     RECT  1051.1 1184.5 1056.58 1184.92 ;
     RECT  1005.98 1184.5 1040.26 1189.12 ;
     RECT  1012.7 1189.12 1040.26 1192.48 ;
     RECT  561.98 1184.92 741.7 1192.9 ;
     RECT  1012.7 1192.48 1027.3 1192.9 ;
     RECT  1040.06 1192.48 1040.26 1193.32 ;
     RECT  1015.1 1192.9 1021.06 1195 ;
     RECT  1016.54 1195 1021.06 1196.26 ;
     RECT  751.58 1181.56 969.22 1196.48 ;
     RECT  561.98 1192.9 738.82 1196.68 ;
     RECT  1016.54 1196.26 1016.74 1196.68 ;
     RECT  748.7 1196.48 969.22 1199.2 ;
     RECT  910.94 1199.2 969.22 1204.24 ;
     RECT  748.7 1199.2 901.06 1206.76 ;
     RECT  562.46 1196.68 738.82 1207.82 ;
     RECT  748.7 1206.76 896.74 1207.82 ;
     RECT  910.94 1204.24 960.1 1211.38 ;
     RECT  910.94 1211.38 959.14 1214.32 ;
     RECT  910.94 1214.32 957.7 1214.96 ;
     RECT  562.46 1207.82 896.74 1217.9 ;
     RECT  562.46 1217.9 897.22 1220 ;
     RECT  907.1 1214.96 957.7 1220 ;
     RECT  562.46 1220 957.7 1221.88 ;
     RECT  921.02 1221.88 957.7 1223.56 ;
     RECT  904.22 1221.88 911.14 1223.98 ;
     RECT  921.02 1223.56 950.98 1225.24 ;
     RECT  562.46 1221.88 893.38 1225.66 ;
     RECT  904.22 1223.98 909.22 1225.66 ;
     RECT  562.46 1225.66 823.78 1226.5 ;
     RECT  835.1 1225.66 893.38 1226.5 ;
     RECT  836.06 1226.5 893.38 1226.92 ;
     RECT  905.18 1225.66 908.26 1226.92 ;
     RECT  950.78 1225.24 950.98 1227.34 ;
     RECT  836.54 1226.92 891.94 1227.76 ;
     RECT  908.06 1226.92 908.26 1227.76 ;
     RECT  836.54 1227.76 878.02 1228.18 ;
     RECT  840.38 1228.18 878.02 1229.86 ;
     RECT  891.74 1227.76 891.94 1229.86 ;
     RECT  921.02 1225.24 940.9 1229.86 ;
     RECT  928.7 1229.86 940.9 1230.7 ;
     RECT  840.38 1229.86 843.94 1231.12 ;
     RECT  857.66 1229.86 878.02 1231.12 ;
     RECT  857.66 1231.12 868.9 1233.22 ;
     RECT  937.82 1230.7 940.9 1233.22 ;
     RECT  562.46 1226.5 819.46 1234.06 ;
     RECT  562.46 1234.06 738.82 1234.48 ;
     RECT  840.38 1231.12 840.58 1234.48 ;
     RECT  857.66 1233.22 859.3 1234.48 ;
     RECT  938.3 1233.22 940.9 1234.48 ;
     RECT  940.7 1234.48 940.9 1234.9 ;
     RECT  719.42 1234.48 738.82 1237 ;
     RECT  719.42 1237 737.86 1237.42 ;
     RECT  732.86 1237.42 737.86 1237.84 ;
     RECT  719.42 1237.42 721.54 1238.26 ;
     RECT  562.46 1234.48 695.14 1238.68 ;
     RECT  562.46 1238.68 685.54 1240.78 ;
     RECT  719.42 1238.26 720.58 1240.78 ;
     RECT  749.18 1234.06 818.02 1240.78 ;
     RECT  573.02 1240.78 685.54 1241.62 ;
     RECT  573.02 1241.62 680.74 1242.04 ;
     RECT  749.18 1240.78 817.54 1242.04 ;
     RECT  720.38 1240.78 720.58 1242.46 ;
     RECT  573.02 1242.04 676.42 1244.56 ;
     RECT  584.54 1244.56 676.42 1244.98 ;
     RECT  749.18 1242.04 817.06 1244.98 ;
     RECT  750.14 1244.98 817.06 1245.4 ;
     RECT  750.14 1245.4 752.74 1245.82 ;
     RECT  562.46 1240.78 562.66 1248.34 ;
     RECT  584.54 1244.98 672.1 1249.18 ;
     RECT  764.06 1245.4 817.06 1249.18 ;
     RECT  573.02 1244.56 573.22 1249.6 ;
     RECT  585.5 1249.18 667.78 1249.6 ;
     RECT  752.54 1245.82 752.74 1249.6 ;
     RECT  764.06 1249.18 768.58 1249.6 ;
     RECT  800.54 1249.18 802.18 1249.6 ;
     RECT  813.02 1249.18 817.06 1249.6 ;
     RECT  764.06 1249.6 764.26 1250.02 ;
     RECT  816.86 1249.6 817.06 1250.02 ;
     RECT  587.9 1249.6 624.58 1252.96 ;
     RECT  780.86 1249.18 785.86 1252.96 ;
     RECT  591.26 1252.96 607.78 1253.8 ;
     RECT  783.26 1252.96 783.46 1253.8 ;
     RECT  599.9 1253.8 607.78 1254.22 ;
     RECT  636.86 1249.6 661.54 1254.22 ;
     RECT  620.06 1252.96 624.58 1255.9 ;
     RECT  636.86 1254.22 656.74 1255.9 ;
     RECT  655.58 1255.9 656.74 1256.32 ;
     RECT  620.06 1255.9 621.22 1256.74 ;
     RECT  636.86 1255.9 645.7 1256.74 ;
     RECT  599.9 1254.22 601.06 1257.16 ;
     RECT  620.06 1256.74 620.26 1257.16 ;
     RECT  638.3 1256.74 638.98 1257.16 ;
     RECT  599.9 1257.16 600.1 1257.58 ;
     RECT  638.3 1257.16 638.5 1257.58 ;
     RECT  655.58 1256.32 655.78 1257.58 ;
    LAYER Metal4 ;
     RECT  1.34 569.42 2.3 569.62 ;
     RECT  1.82 583.7 2.3 583.9 ;
     RECT  0.86 626.12 3.26 626.32 ;
     RECT  3.26 501.8 7.1 514.6 ;
     RECT  3.26 622.76 7.1 626.32 ;
     RECT  3.26 642.92 7.1 660.76 ;
     RECT  3.26 685.76 7.1 718.72 ;
     RECT  554.3 934.82 556.22 935.02 ;
     RECT  554.3 1116.68 556.7 1116.88 ;
     RECT  541.82 894.08 561.02 894.28 ;
     RECT  561.02 890.72 562.46 894.28 ;
     RECT  556.22 928.1 562.94 935.02 ;
     RECT  561.5 1044.86 562.94 1045.06 ;
     RECT  562.94 928.1 563.14 942.16 ;
     RECT  556.7 1116.68 565.54 1120.66 ;
     RECT  565.54 1120.46 566.78 1120.66 ;
     RECT  564.86 869.72 567.94 869.92 ;
     RECT  562.94 1044.86 567.94 1049.26 ;
     RECT  562.46 890.72 568.7 901.84 ;
     RECT  568.22 1082.66 568.7 1082.86 ;
     RECT  563.14 941.96 568.9 942.16 ;
     RECT  568.7 886.52 569.18 901.84 ;
     RECT  566.78 1120.46 569.18 1124.44 ;
     RECT  569.18 1120.46 570.62 1127.8 ;
     RECT  561.98 841.16 571.1 841.36 ;
     RECT  563.14 928.1 571.1 932.5 ;
     RECT  564.38 855.86 571.58 860.26 ;
     RECT  571.1 924.74 571.58 932.5 ;
     RECT  567.26 981.02 571.58 981.22 ;
     RECT  570.62 1120.46 571.78 1128.64 ;
     RECT  566.3 950.78 572.54 950.98 ;
     RECT  571.58 922.22 573.02 932.5 ;
     RECT  568.7 1078.88 573.7 1086.22 ;
     RECT  573.7 1086.02 573.98 1086.22 ;
     RECT  569.66 965.48 574.46 965.68 ;
     RECT  571.58 981.02 574.46 985.42 ;
     RECT  573.98 1086.02 575.42 1088.32 ;
     RECT  571.78 1123.82 575.42 1128.64 ;
     RECT  575.42 1086.02 575.9 1091.68 ;
     RECT  554.3 1101.98 575.9 1102.18 ;
     RECT  569.18 885.68 576.38 901.84 ;
     RECT  575.9 1101.98 576.38 1109.32 ;
     RECT  575.42 1123.82 576.38 1129.06 ;
     RECT  564.38 818.9 576.86 819.1 ;
     RECT  562.94 829.4 576.86 829.6 ;
     RECT  571.1 841.16 576.86 841.78 ;
     RECT  573.02 921.8 576.86 932.5 ;
     RECT  574.46 965.48 577.06 985.42 ;
     RECT  576.86 818.48 577.34 819.1 ;
     RECT  576.38 1101.98 577.34 1110.16 ;
     RECT  577.34 1101.98 577.54 1110.58 ;
     RECT  576.86 921.8 578.78 935.44 ;
     RECT  558.14 1060.4 578.78 1060.6 ;
     RECT  577.82 1071.32 578.78 1071.52 ;
     RECT  575.9 1086.02 578.78 1092.52 ;
     RECT  567.94 1044.86 578.98 1045.48 ;
     RECT  572.54 948.68 579.46 950.98 ;
     RECT  577.54 1101.98 579.94 1110.16 ;
     RECT  576.38 1123.82 580.22 1129.9 ;
     RECT  578.78 1060.4 581.38 1071.52 ;
     RECT  580.22 1123.4 582.14 1129.9 ;
     RECT  582.14 1120.88 582.34 1129.9 ;
     RECT  570.14 1188.5 582.34 1188.7 ;
     RECT  581.38 1060.4 582.62 1064.38 ;
     RECT  582.34 1120.88 583.3 1129.06 ;
     RECT  577.34 814.28 584.06 819.1 ;
     RECT  576.86 829.4 584.06 841.78 ;
     RECT  570.14 1177.16 584.06 1177.36 ;
     RECT  584.06 814.28 584.26 841.78 ;
     RECT  574.94 1233.86 584.74 1234.06 ;
     RECT  578.78 916.76 585.02 935.44 ;
     RECT  578.3 1150.7 585.02 1150.9 ;
     RECT  571.58 852.5 585.22 860.26 ;
     RECT  574.94 870.98 585.5 871.18 ;
     RECT  582.62 1056.62 586.46 1064.38 ;
     RECT  576.38 881.9 586.66 901.84 ;
     RECT  585.5 870.98 587.42 871.6 ;
     RECT  586.66 881.9 587.42 899.32 ;
     RECT  579.94 1101.98 589.54 1102.18 ;
     RECT  578.98 1045.28 590.02 1045.48 ;
     RECT  585.22 852.5 590.98 856.48 ;
     RECT  587.42 870.98 591.94 899.32 ;
     RECT  583.3 1120.88 591.94 1128.64 ;
     RECT  586.46 1056.2 592.42 1064.38 ;
     RECT  589.34 1075.1 592.42 1075.3 ;
     RECT  592.42 1056.2 592.7 1058.5 ;
     RECT  591.94 871.4 593.38 899.32 ;
     RECT  591.94 1122.98 596.26 1128.64 ;
     RECT  585.02 912.98 596.54 939.64 ;
     RECT  590.98 855.86 597.5 856.48 ;
     RECT  577.06 984.38 599.14 985.42 ;
     RECT  584.26 837.8 599.9 841.78 ;
     RECT  577.06 973.04 599.9 973.24 ;
     RECT  599.14 984.38 599.9 985 ;
     RECT  578.3 1007.48 600.1 1007.68 ;
     RECT  584.26 814.28 600.86 822.04 ;
     RECT  579.46 948.68 601.82 948.88 ;
     RECT  599.9 973.04 602.02 985 ;
     RECT  596.54 912.56 604.42 939.64 ;
     RECT  601.82 948.68 604.7 951.4 ;
     RECT  602.02 973.04 604.7 976.18 ;
     RECT  585.02 1150.7 604.7 1158.88 ;
     RECT  590.78 1192.28 604.7 1192.48 ;
     RECT  567.74 1201.94 604.7 1202.14 ;
     RECT  602.3 1214.54 604.7 1214.74 ;
     RECT  593.38 873.92 604.9 899.32 ;
     RECT  604.7 948.68 604.9 976.18 ;
     RECT  604.7 1150.7 604.9 1159.3 ;
     RECT  592.7 1052.84 605.18 1058.5 ;
     RECT  604.9 950.36 605.38 976.18 ;
     RECT  604.7 1030.58 605.66 1030.78 ;
     RECT  604.7 1192.28 606.14 1193.32 ;
     RECT  604.7 1201.94 606.14 1214.74 ;
     RECT  605.38 965.48 606.34 976.18 ;
     RECT  605.66 1030.16 606.82 1030.78 ;
     RECT  599.9 835.28 607.78 841.78 ;
     RECT  602.02 984.8 608.06 985 ;
     RECT  578.78 1086.02 608.06 1093.36 ;
     RECT  606.82 1030.16 608.26 1030.36 ;
     RECT  7.1 685.76 608.54 723.34 ;
     RECT  4.22 736.16 608.54 736.36 ;
     RECT  605.18 1050.32 608.54 1058.5 ;
     RECT  608.06 984.8 609.02 992.56 ;
     RECT  608.06 1086.02 609.5 1098.4 ;
     RECT  584.06 1177.16 609.5 1181.98 ;
     RECT  606.14 1192.28 609.5 1219.36 ;
     RECT  608.54 685.76 609.7 736.36 ;
     RECT  608.54 1044.02 609.98 1058.5 ;
     RECT  609.98 1044.02 611.62 1063.96 ;
     RECT  605.38 950.36 612.1 954.76 ;
     RECT  609.5 1177.16 612.38 1219.36 ;
     RECT  600.86 814.28 613.34 826.24 ;
     RECT  607.78 835.28 613.34 840.1 ;
     RECT  609.02 984.8 613.34 1000.12 ;
     RECT  604.9 1150.7 615.26 1150.9 ;
     RECT  612.86 1162.04 615.26 1162.24 ;
     RECT  596.26 1122.98 615.46 1124.44 ;
     RECT  597.5 855.86 616.22 859 ;
     RECT  612.38 1173.8 616.22 1219.36 ;
     RECT  607.1 1234.28 616.22 1234.48 ;
     RECT  604.42 916.76 616.7 939.64 ;
     RECT  616.22 855.02 617.18 859 ;
     RECT  615.26 1150.7 617.18 1162.24 ;
     RECT  616.7 914.66 618.14 939.64 ;
     RECT  618.14 913.82 618.34 939.64 ;
     RECT  613.34 814.28 618.62 840.1 ;
     RECT  618.62 814.28 619.1 840.94 ;
     RECT  604.9 873.92 619.1 894.28 ;
     RECT  616.22 1173.8 620.54 1234.48 ;
     RECT  618.34 916.76 621.5 939.64 ;
     RECT  612.1 950.78 621.5 954.76 ;
     RECT  617.18 1143.56 623.9 1162.24 ;
     RECT  619.1 873.92 624.1 897.64 ;
     RECT  609.5 1084.76 624.1 1098.4 ;
     RECT  617.18 854.6 624.38 859 ;
     RECT  624.38 854.6 624.58 863.62 ;
     RECT  609.7 685.76 624.86 723.34 ;
     RECT  623.9 1142.3 624.86 1162.24 ;
     RECT  606.34 965.48 625.34 973.24 ;
     RECT  613.34 981.86 625.34 1000.12 ;
     RECT  619.1 814.28 625.82 841.36 ;
     RECT  615.46 1124.24 625.82 1124.44 ;
     RECT  606.62 750.44 626.3 750.64 ;
     RECT  621.5 916.76 626.98 954.76 ;
     RECT  619.58 784.04 627.74 784.24 ;
     RECT  611.62 1044.02 629.18 1057.66 ;
     RECT  624.86 685.76 629.38 727.54 ;
     RECT  607.58 765.98 629.66 766.18 ;
     RECT  7.1 670.64 630.14 670.84 ;
     RECT  629.38 685.76 630.14 723.34 ;
     RECT  628.22 1033.52 630.14 1033.72 ;
     RECT  626.3 746.24 631.1 750.64 ;
     RECT  624.1 1084.76 631.1 1097.98 ;
     RECT  619.58 1010.84 631.3 1011.04 ;
     RECT  627.74 784.04 631.58 791.8 ;
     RECT  626.98 916.76 632.26 939.64 ;
     RECT  631.1 746.24 632.54 752.32 ;
     RECT  629.66 765.14 632.54 766.18 ;
     RECT  625.34 965.48 632.54 1000.12 ;
     RECT  631.1 1072.58 632.54 1072.78 ;
     RECT  631.1 1082.66 632.54 1097.98 ;
     RECT  624.1 873.92 632.74 894.28 ;
     RECT  632.54 746.24 633.02 766.18 ;
     RECT  633.02 746.24 633.5 769.12 ;
     RECT  631.58 783.62 633.5 791.8 ;
     RECT  633.5 746.24 633.98 791.8 ;
     RECT  626.98 950.78 634.18 954.76 ;
     RECT  624.86 1138.52 634.18 1162.24 ;
     RECT  624.58 855.44 634.46 863.62 ;
     RECT  632.74 873.92 634.46 890.08 ;
     RECT  625.82 813.86 634.94 841.36 ;
     RECT  634.46 855.44 634.94 890.08 ;
     RECT  630.14 1029.74 635.42 1033.72 ;
     RECT  633.98 746.24 636.86 796 ;
     RECT  620.54 1173.8 638.5 1242.04 ;
     RECT  635.42 1023.02 638.78 1033.72 ;
     RECT  630.14 670.64 639.94 723.34 ;
     RECT  634.94 813.86 640.42 890.08 ;
     RECT  638.78 1018.4 640.42 1033.72 ;
     RECT  636.86 746.24 640.7 796.42 ;
     RECT  632.54 965.06 641.18 1000.12 ;
     RECT  632.26 916.76 641.66 934.6 ;
     RECT  638.5 1173.8 642.62 1237.84 ;
     RECT  632.54 1072.58 643.58 1097.98 ;
     RECT  642.14 1106.6 643.58 1106.8 ;
     RECT  642.62 1166.66 643.78 1237.84 ;
     RECT  643.58 1072.58 644.06 1106.8 ;
     RECT  644.06 1072.16 645.22 1106.8 ;
     RECT  639.26 1249.4 645.22 1249.6 ;
     RECT  639.94 670.64 646.18 671.26 ;
     RECT  640.7 746.24 646.46 798.1 ;
     RECT  646.46 746.24 646.66 803.56 ;
     RECT  641.66 916.76 647.42 935.86 ;
     RECT  634.18 950.78 647.42 951.4 ;
     RECT  643.78 1173.8 647.62 1237.84 ;
     RECT  647.42 916.76 648.86 951.4 ;
     RECT  641.18 965.06 648.86 1007.26 ;
     RECT  648.86 916.76 649.06 1007.26 ;
     RECT  649.06 994.88 649.34 1007.26 ;
     RECT  640.42 1018.4 649.34 1018.6 ;
     RECT  647.62 1173.8 649.54 1211.8 ;
     RECT  646.66 759.68 650.02 803.56 ;
     RECT  625.82 1115.84 650.3 1124.44 ;
     RECT  634.18 1138.52 650.3 1157.62 ;
     RECT  649.34 994.88 650.98 1018.6 ;
     RECT  639.94 685.76 651.26 723.34 ;
     RECT  609.7 736.16 651.26 736.36 ;
     RECT  649.06 916.76 653.38 985 ;
     RECT  645.22 1072.16 653.86 1102.18 ;
     RECT  650.3 1138.52 654.14 1158.46 ;
     RECT  654.14 1138.52 654.62 1158.88 ;
     RECT  629.18 1044.02 654.82 1058.5 ;
     RECT  647.62 1222.52 654.82 1237.84 ;
     RECT  7.1 638.3 655.1 660.76 ;
     RECT  646.18 670.64 655.1 670.84 ;
     RECT  654.82 1044.02 655.1 1058.08 ;
     RECT  651.26 685.76 655.3 736.36 ;
     RECT  654.62 1138.52 655.3 1159.72 ;
     RECT  649.54 1177.16 655.3 1211.8 ;
     RECT  654.82 1229.24 655.3 1237.84 ;
     RECT  650.02 759.68 655.58 793.48 ;
     RECT  655.58 758 657.02 793.48 ;
     RECT  655.3 1201.94 657.5 1211.8 ;
     RECT  657.02 757.58 658.94 793.48 ;
     RECT  650.02 803.36 658.94 803.56 ;
     RECT  655.3 1234.28 658.94 1237.84 ;
     RECT  650.98 1010 660.86 1018.6 ;
     RECT  650.3 1115.84 661.34 1128.22 ;
     RECT  655.3 1138.52 661.34 1158.88 ;
     RECT  653.38 965.06 661.82 985 ;
     RECT  650.98 994.88 661.82 1000.12 ;
     RECT  658.94 757.58 663.74 803.56 ;
     RECT  653.38 916.76 663.74 951.4 ;
     RECT  658.94 1234.28 663.94 1241.62 ;
     RECT  640.42 814.28 665.86 890.08 ;
     RECT  661.82 965.06 666.14 1000.12 ;
     RECT  655.3 736.16 667.1 736.36 ;
     RECT  662.78 1105.76 667.1 1105.96 ;
     RECT  661.34 1115.84 667.1 1158.88 ;
     RECT  660.86 1009.58 667.58 1018.6 ;
     RECT  653.86 1072.16 667.78 1093.78 ;
     RECT  663.74 757.58 668.26 803.98 ;
     RECT  655.3 685.76 668.54 723.76 ;
     RECT  667.1 736.16 668.54 743.08 ;
     RECT  667.58 1009.58 668.74 1019.02 ;
     RECT  667.1 1105.76 669.7 1158.88 ;
     RECT  663.94 1237.64 669.7 1241.62 ;
     RECT  668.54 685.76 670.18 743.08 ;
     RECT  666.14 962.54 670.46 1000.12 ;
     RECT  665.86 818.48 671.14 890.08 ;
     RECT  670.46 962.12 674.5 1000.12 ;
     RECT  672.86 907.1 674.78 907.3 ;
     RECT  663.74 916.76 674.78 951.82 ;
     RECT  670.18 685.76 674.98 736.36 ;
     RECT  640.42 1029.74 675.74 1033.72 ;
     RECT  674.78 907.1 675.94 951.82 ;
     RECT  671.14 818.48 676.42 864.46 ;
     RECT  674.98 685.76 677.38 723.76 ;
     RECT  668.74 1009.58 679.3 1018.6 ;
     RECT  675.74 1029.74 681.98 1034.14 ;
     RECT  655.1 1043.6 681.98 1058.08 ;
     RECT  667.78 1072.58 682.46 1093.78 ;
     RECT  668.26 760.52 684.58 803.98 ;
     RECT  676.42 825.62 685.06 864.46 ;
     RECT  655.1 638.3 685.34 670.84 ;
     RECT  669.7 1241.42 685.54 1241.62 ;
     RECT  675.94 909.2 686.78 951.82 ;
     RECT  674.5 962.12 686.78 983.74 ;
     RECT  669.7 1113.32 687.26 1158.88 ;
     RECT  684.58 760.52 687.74 803.56 ;
     RECT  674.5 994.88 687.74 1000.12 ;
     RECT  677.38 685.76 689.18 723.34 ;
     RECT  687.26 1113.32 689.86 1159.72 ;
     RECT  687.74 758 691.3 803.56 ;
     RECT  686.78 909.2 691.78 983.74 ;
     RECT  655.3 1177.16 692.06 1192.48 ;
     RECT  657.5 1201.94 692.06 1218.94 ;
     RECT  679.1 899.12 692.26 899.32 ;
     RECT  689.18 681.56 693.22 723.34 ;
     RECT  687.74 994.04 693.5 1000.12 ;
     RECT  681.98 1029.74 695.14 1058.08 ;
     RECT  685.34 638.3 696.1 671.68 ;
     RECT  682.46 1071.32 696.58 1093.78 ;
     RECT  685.06 825.62 698.3 829.6 ;
     RECT  685.06 844.52 698.3 864.46 ;
     RECT  689.86 1113.32 698.3 1124.44 ;
     RECT  698.3 1113.32 698.5 1126.96 ;
     RECT  696.1 660.56 699.46 671.68 ;
     RECT  671.14 873.92 700.22 890.08 ;
     RECT  692.06 1177.16 700.7 1218.94 ;
     RECT  691.3 760.52 701.66 803.56 ;
     RECT  693.98 813.44 701.66 813.64 ;
     RECT  700.22 873.92 701.86 896.38 ;
     RECT  691.78 909.2 702.34 951.4 ;
     RECT  702.34 924.32 702.62 951.4 ;
     RECT  691.78 961.28 702.62 983.74 ;
     RECT  702.62 924.32 702.82 983.74 ;
     RECT  700.7 1173.8 703.3 1218.94 ;
     RECT  689.86 1138.52 704.54 1159.72 ;
     RECT  696.58 1072.58 705.02 1093.78 ;
     RECT  693.22 685.76 705.5 723.34 ;
     RECT  695.14 1041.08 705.5 1058.08 ;
     RECT  698.5 1113.32 705.5 1116.04 ;
     RECT  698.5 1126.76 705.5 1126.96 ;
     RECT  704.54 1136 705.5 1159.72 ;
     RECT  702.82 934.4 705.7 983.74 ;
     RECT  695.14 1029.74 705.7 1031.62 ;
     RECT  698.3 825.62 705.98 864.46 ;
     RECT  701.86 873.92 705.98 890.08 ;
     RECT  705.5 1041.08 706.46 1058.92 ;
     RECT  705.02 1072.58 706.46 1094.2 ;
     RECT  705.5 1126.76 707.14 1159.72 ;
     RECT  701.66 760.52 708.38 813.64 ;
     RECT  708.38 755.06 709.06 813.64 ;
     RECT  707.14 1136 709.82 1159.72 ;
     RECT  709.06 764.72 710.3 813.64 ;
     RECT  705.98 825.62 710.3 890.08 ;
     RECT  705.7 960.02 712.7 983.74 ;
     RECT  693.5 992.36 712.7 1000.12 ;
     RECT  705.5 1109.12 713.18 1116.04 ;
     RECT  702.34 909.2 715.1 915.7 ;
     RECT  702.82 924.32 715.1 924.52 ;
     RECT  696.1 638.3 716.06 650.68 ;
     RECT  699.46 660.56 716.06 660.76 ;
     RECT  710.3 764.72 716.06 890.08 ;
     RECT  715.1 908.36 716.06 924.52 ;
     RECT  705.7 934.4 716.06 950.56 ;
     RECT  716.06 764.72 716.54 897.22 ;
     RECT  706.46 1041.08 717.02 1094.2 ;
     RECT  713.18 1105.76 717.98 1116.04 ;
     RECT  707.14 1126.76 717.98 1126.96 ;
     RECT  709.82 1136 717.98 1161.82 ;
     RECT  716.06 908.36 718.18 950.56 ;
     RECT  705.7 1029.74 718.66 1030.36 ;
     RECT  717.02 1041.08 718.66 1094.62 ;
     RECT  709.06 755.06 718.94 755.26 ;
     RECT  716.54 764.72 718.94 897.64 ;
     RECT  717.98 1105.76 719.14 1126.96 ;
     RECT  703.3 1173.8 719.14 1216.42 ;
     RECT  705.5 685.76 719.9 727.54 ;
     RECT  674.98 736.16 719.9 736.36 ;
     RECT  712.7 960.02 719.9 1000.12 ;
     RECT  719.9 960.02 720.86 1000.54 ;
     RECT  718.18 934.4 721.34 950.56 ;
     RECT  720.86 959.18 721.34 1000.54 ;
     RECT  718.94 755.06 721.82 897.64 ;
     RECT  719.9 685.76 722.3 743.08 ;
     RECT  721.82 753.8 722.3 897.64 ;
     RECT  718.18 908.36 722.3 924.52 ;
     RECT  722.3 685.76 722.5 924.52 ;
     RECT  721.34 934.4 724.42 1000.54 ;
     RECT  719.14 1105.76 724.9 1116.04 ;
     RECT  722.5 873.92 727.1 924.52 ;
     RECT  724.42 934.4 727.1 951.4 ;
     RECT  719.14 1173.8 727.3 1214.74 ;
     RECT  719.14 1126.76 728.06 1126.96 ;
     RECT  717.98 1136 728.06 1162.24 ;
     RECT  7.1 622.76 731.14 628 ;
     RECT  718.66 1029.74 733.82 1029.94 ;
     RECT  718.66 1041.08 733.82 1058.92 ;
     RECT  724.9 1105.76 734.3 1105.96 ;
     RECT  724.9 1115.84 734.3 1116.04 ;
     RECT  679.3 1009.58 734.98 1010.2 ;
     RECT  734.3 1105.76 735.46 1116.04 ;
     RECT  718.66 1070.48 736.22 1094.62 ;
     RECT  735.46 1105.76 736.22 1105.96 ;
     RECT  736.22 1070.48 737.18 1105.96 ;
     RECT  733.82 1022.6 737.38 1058.92 ;
     RECT  734.98 1010 739.3 1010.2 ;
     RECT  737.18 1068.8 739.3 1105.96 ;
     RECT  739.3 1102.82 739.78 1105.96 ;
     RECT  739.3 1068.8 741.7 1093.78 ;
     RECT  727.1 873.92 742.18 951.4 ;
     RECT  737.38 1031.84 742.66 1058.92 ;
     RECT  724.42 960.02 743.62 1000.54 ;
     RECT  743.62 961.28 744.1 1000.54 ;
     RECT  722.5 685.76 744.86 864.46 ;
     RECT  737.38 1022.6 745.54 1022.8 ;
     RECT  716.06 638.3 746.02 660.76 ;
     RECT  727.3 1173.8 746.5 1212.64 ;
     RECT  739.58 1230.5 746.78 1230.7 ;
     RECT  746.02 660.56 747.26 660.76 ;
     RECT  699.46 670.64 747.26 671.68 ;
     RECT  742.66 1031.84 747.26 1058.08 ;
     RECT  742.18 873.92 747.46 903.1 ;
     RECT  731.14 622.76 747.74 626.32 ;
     RECT  746.02 638.3 747.74 650.68 ;
     RECT  744.86 685.34 748.22 864.46 ;
     RECT  747.46 873.92 748.22 889.66 ;
     RECT  728.06 1126.76 748.22 1162.24 ;
     RECT  746.5 1173.8 748.22 1204.24 ;
     RECT  742.18 912.98 748.7 951.4 ;
     RECT  747.26 660.56 749.38 671.68 ;
     RECT  747.26 1031 749.38 1058.08 ;
     RECT  746.78 1230.5 750.34 1234.48 ;
     RECT  739.78 1105.76 750.62 1105.96 ;
     RECT  735.46 1115.84 750.62 1116.04 ;
     RECT  744.1 961.28 753.22 1000.12 ;
     RECT  750.34 1234.28 753.5 1234.48 ;
     RECT  747.74 622.76 754.18 650.68 ;
     RECT  748.22 685.34 755.14 889.66 ;
     RECT  747.46 902.9 755.9 903.1 ;
     RECT  748.7 912.98 755.9 951.82 ;
     RECT  752.06 1224.2 755.9 1224.4 ;
     RECT  748.22 1126.76 756.1 1204.24 ;
     RECT  754.46 1011.26 756.38 1011.46 ;
     RECT  755.14 685.34 757.34 864.46 ;
     RECT  755.14 873.92 759.26 889.66 ;
     RECT  756.38 1011.26 760.22 1011.88 ;
     RECT  755.9 1223.36 760.42 1224.4 ;
     RECT  757.34 682.4 760.9 864.46 ;
     RECT  759.26 873.92 761.18 890.92 ;
     RECT  755.9 902.9 761.18 952.24 ;
     RECT  760.22 1011.26 763.1 1013.98 ;
     RECT  749.38 1031.84 763.1 1058.08 ;
     RECT  753.22 961.28 763.58 998.44 ;
     RECT  763.1 1008.32 763.58 1013.98 ;
     RECT  753.5 1234.28 763.58 1237.42 ;
     RECT  763.58 961.28 764.06 1013.98 ;
     RECT  763.1 1026.38 764.06 1058.08 ;
     RECT  760.42 1223.36 764.06 1223.56 ;
     RECT  750.62 1105.76 766.94 1116.04 ;
     RECT  756.1 1126.76 766.94 1158.46 ;
     RECT  760.9 685.76 768.38 864.46 ;
     RECT  761.18 873.92 768.38 952.24 ;
     RECT  764.06 1219.16 768.38 1223.56 ;
     RECT  764.06 961.28 768.58 1058.08 ;
     RECT  766.94 1105.76 769.54 1158.46 ;
     RECT  768.38 685.76 771.94 952.24 ;
     RECT  741.7 1071.32 773.18 1093.78 ;
     RECT  769.54 1105.76 773.18 1116.04 ;
     RECT  768.58 1026.38 777.02 1058.08 ;
     RECT  773.18 1071.32 777.02 1116.04 ;
     RECT  768.38 1218.74 777.22 1223.56 ;
     RECT  769.54 1126.76 777.98 1158.46 ;
     RECT  749.38 670.64 778.18 671.68 ;
     RECT  768.58 961.28 778.94 1014.82 ;
     RECT  777.02 1026.38 778.94 1116.04 ;
     RECT  763.58 1234.28 779.9 1242.04 ;
     RECT  777.22 1218.74 784.42 1219.36 ;
     RECT  779.9 1230.5 784.42 1242.04 ;
     RECT  756.1 1173.8 784.9 1204.24 ;
     RECT  778.18 670.64 787.1 671.26 ;
     RECT  771.94 685.76 787.1 897.64 ;
     RECT  771.94 907.94 789.7 952.24 ;
     RECT  787.1 670.64 790.18 897.64 ;
     RECT  784.42 1219.16 791.9 1219.36 ;
     RECT  784.42 1230.5 791.9 1238.26 ;
     RECT  784.9 1177.58 793.34 1204.24 ;
     RECT  793.34 1177.58 793.54 1207.18 ;
     RECT  791.9 1219.16 795.94 1238.26 ;
     RECT  790.18 679.46 796.9 897.64 ;
     RECT  778.94 961.28 797.86 1116.04 ;
     RECT  796.9 679.46 798.34 864.46 ;
     RECT  793.54 1180.52 798.34 1207.18 ;
     RECT  795.94 1222.52 798.82 1238.26 ;
     RECT  798.34 679.46 799.3 751.48 ;
     RECT  799.3 679.46 800.26 748.96 ;
     RECT  797.86 961.28 800.26 1058.92 ;
     RECT  790.18 670.64 800.54 670.84 ;
     RECT  777.98 1126.76 800.74 1161.82 ;
     RECT  798.34 760.94 801.7 864.46 ;
     RECT  800.26 685.76 802.66 748.96 ;
     RECT  789.7 907.94 802.94 951.82 ;
     RECT  800.26 961.28 802.94 998.44 ;
     RECT  800.26 1010 803.62 1058.92 ;
     RECT  796.9 873.92 804.38 897.64 ;
     RECT  802.94 907.94 804.38 998.44 ;
     RECT  797.86 1071.32 804.58 1116.04 ;
     RECT  798.82 1232.18 806.5 1238.26 ;
     RECT  804.58 1071.32 808.22 1097.14 ;
     RECT  804.38 873.92 808.42 998.44 ;
     RECT  808.42 873.92 809.38 951.82 ;
     RECT  800.74 1126.76 809.66 1158.46 ;
     RECT  809.38 950.78 810.82 951.82 ;
     RECT  806.5 1234.28 811.78 1238.26 ;
     RECT  754.18 622.76 812.06 626.32 ;
     RECT  801.7 761.78 812.06 864.46 ;
     RECT  809.38 873.92 812.06 942.16 ;
     RECT  804.58 1105.76 812.26 1116.04 ;
     RECT  811.78 1235.54 812.26 1238.26 ;
     RECT  800.54 669.8 813.22 670.84 ;
     RECT  798.34 1180.52 813.22 1205.08 ;
     RECT  812.06 761.78 813.5 942.16 ;
     RECT  812.26 1235.54 814.18 1237 ;
     RECT  813.22 1180.52 814.46 1181.14 ;
     RECT  803.62 1029.74 815.42 1058.92 ;
     RECT  814.18 1236.8 815.62 1237 ;
     RECT  803.62 1010 816.38 1016.92 ;
     RECT  814.46 1179.26 816.86 1181.14 ;
     RECT  813.5 756.32 817.54 942.16 ;
     RECT  813.22 670.64 818.3 670.84 ;
     RECT  802.66 685.76 818.3 746.44 ;
     RECT  816.38 1010 818.5 1019.02 ;
     RECT  816.86 1175.9 818.5 1181.14 ;
     RECT  813.22 1191.44 819.26 1205.08 ;
     RECT  818.5 1179.26 819.46 1181.14 ;
     RECT  819.46 1179.68 819.94 1181.14 ;
     RECT  810.82 950.78 820.22 950.98 ;
     RECT  808.42 961.28 820.22 998.44 ;
     RECT  818.3 670.64 820.42 746.44 ;
     RECT  812.26 1108.7 820.7 1116.04 ;
     RECT  818.5 1010 823.58 1016.92 ;
     RECT  819.94 1180.52 823.58 1181.14 ;
     RECT  817.54 873.92 824.74 942.16 ;
     RECT  815.42 1029.74 828.1 1060.6 ;
     RECT  749.38 660.56 830.78 660.76 ;
     RECT  820.42 670.64 830.78 743.08 ;
     RECT  817.54 756.32 830.78 864.46 ;
     RECT  824.74 873.92 830.78 938.8 ;
     RECT  820.7 1106.18 831.74 1116.04 ;
     RECT  809.66 1126.76 831.74 1162.66 ;
     RECT  830.78 756.32 832.22 938.8 ;
     RECT  831.74 1106.18 833.38 1162.66 ;
     RECT  823.58 1008.74 834.14 1016.92 ;
     RECT  832.22 754.22 834.62 938.8 ;
     RECT  828.1 1029.74 834.82 1058.08 ;
     RECT  819.26 1191.44 834.82 1211.38 ;
     RECT  834.62 754.22 835.1 939.22 ;
     RECT  833.38 1109.12 835.3 1162.66 ;
     RECT  830.78 660.56 836.06 743.08 ;
     RECT  835.1 751.7 836.06 939.22 ;
     RECT  834.82 1033.1 837.98 1058.08 ;
     RECT  3.26 539.6 838.94 539.8 ;
     RECT  836.06 660.56 838.94 939.22 ;
     RECT  838.94 660.56 840.1 940.48 ;
     RECT  838.94 539.6 840.38 541.9 ;
     RECT  3.26 552.2 840.38 554.92 ;
     RECT  834.14 1008.32 841.34 1016.92 ;
     RECT  823.58 1180.52 841.34 1181.56 ;
     RECT  834.82 1191.44 841.34 1204.24 ;
     RECT  820.22 950.78 842.02 998.44 ;
     RECT  837.98 1033.1 842.98 1060.6 ;
     RECT  812.06 620.66 843.74 626.32 ;
     RECT  754.18 638.3 843.74 650.68 ;
     RECT  843.74 620.66 844.22 650.68 ;
     RECT  840.1 660.56 844.22 938.38 ;
     RECT  844.22 620.66 844.42 938.38 ;
     RECT  808.22 1070.9 845.86 1097.14 ;
     RECT  835.3 1126.76 845.86 1162.66 ;
     RECT  842.98 1036.46 846.14 1060.6 ;
     RECT  835.3 1109.12 846.62 1116.04 ;
     RECT  844.42 620.66 849.5 889.66 ;
     RECT  849.5 618.56 849.7 889.66 ;
     RECT  846.14 1036.46 849.7 1061.02 ;
     RECT  845.86 1071.32 850.46 1097.14 ;
     RECT  846.62 1105.76 850.46 1116.04 ;
     RECT  849.7 1040.24 850.66 1061.02 ;
     RECT  840.38 539.6 856.7 554.92 ;
     RECT  3.26 597.56 856.7 607.84 ;
     RECT  849.7 618.56 856.7 889.24 ;
     RECT  844.42 901.64 856.7 938.38 ;
     RECT  841.34 1008.32 856.7 1022.8 ;
     RECT  2.3 569.42 857.18 583.9 ;
     RECT  856.7 597.56 857.18 889.24 ;
     RECT  856.7 901.64 857.38 945.1 ;
     RECT  7.1 498.02 857.66 514.6 ;
     RECT  842.02 954.56 858.62 998.44 ;
     RECT  856.7 539.6 859.1 557.02 ;
     RECT  856.7 1007.9 859.3 1022.8 ;
     RECT  859.1 534.56 860.06 557.44 ;
     RECT  857.18 569 860.06 583.9 ;
     RECT  857.18 593.78 860.26 889.24 ;
     RECT  850.66 1040.24 860.54 1060.6 ;
     RECT  850.46 1071.32 860.54 1116.04 ;
     RECT  845.86 1126.76 860.54 1158.46 ;
     RECT  857.66 498.02 861.02 515.86 ;
     RECT  860.06 534.56 861.02 583.9 ;
     RECT  860.26 593.78 861.02 691 ;
     RECT  860.26 701.3 861.7 889.24 ;
     RECT  861.7 851.24 861.98 889.24 ;
     RECT  857.38 901.64 861.98 928.72 ;
     RECT  860.54 1040.24 863.9 1116.04 ;
     RECT  861.02 534.56 864.1 691 ;
     RECT  864.1 534.56 865.34 583.9 ;
     RECT  859.3 1007.9 866.98 1015.66 ;
     RECT  861.02 498.02 869.18 520.9 ;
     RECT  865.34 531.62 869.18 583.9 ;
     RECT  857.38 938.18 869.18 945.1 ;
     RECT  858.62 954.14 869.18 998.44 ;
     RECT  869.18 938.18 870.14 998.44 ;
     RECT  866.98 1007.9 870.14 1014.82 ;
     RECT  861.98 851.24 871.58 928.72 ;
     RECT  863.9 1033.52 872.54 1116.04 ;
     RECT  860.54 1125.08 872.54 1158.88 ;
     RECT  861.7 701.3 873.02 841.78 ;
     RECT  871.58 850.82 873.02 928.72 ;
     RECT  3.26 471.56 873.5 471.76 ;
     RECT  798.82 1222.52 875.62 1222.72 ;
     RECT  864.1 593.78 878.3 691 ;
     RECT  873.02 701.3 878.3 928.72 ;
     RECT  869.18 498.02 878.78 583.9 ;
     RECT  878.3 593.78 878.78 928.72 ;
     RECT  878.78 498.02 878.98 928.72 ;
     RECT  873.5 471.56 879.74 472.18 ;
     RECT  870.14 938.18 879.74 1014.82 ;
     RECT  879.74 938.18 881.18 1021.54 ;
     RECT  872.54 1033.52 881.18 1158.88 ;
     RECT  879.74 466.52 881.66 472.18 ;
     RECT  881.18 938.18 883.3 1158.88 ;
     RECT  3.26 481.64 883.58 486.88 ;
     RECT  878.98 498.02 883.58 527.2 ;
     RECT  881.66 464 884.54 472.18 ;
     RECT  883.58 481.64 884.54 527.2 ;
     RECT  883.3 951.2 884.74 1158.88 ;
     RECT  841.34 1180.52 885.7 1204.24 ;
     RECT  0.38 435.86 885.98 436.06 ;
     RECT  878.98 539.6 886.94 928.72 ;
     RECT  883.3 938.18 886.94 938.38 ;
     RECT  3.26 451.4 887.42 454.12 ;
     RECT  884.54 464 887.42 527.2 ;
     RECT  886.94 539.6 887.62 938.38 ;
     RECT  884.74 954.14 890.98 1158.88 ;
     RECT  885.7 1196.9 890.98 1204.24 ;
     RECT  887.42 451.4 891.26 527.2 ;
     RECT  873.98 1169.6 891.46 1169.8 ;
     RECT  887.62 539.6 892.22 928.72 ;
     RECT  890.98 954.14 893.38 981.64 ;
     RECT  890.78 1214.96 893.38 1215.16 ;
     RECT  891.26 451.4 896.26 528.88 ;
     RECT  890.98 991.94 897.7 1158.88 ;
     RECT  896.26 471.56 899.62 528.88 ;
     RECT  897.7 991.94 901.06 1158.46 ;
     RECT  896.26 451.4 902.02 462.94 ;
     RECT  892.22 537.92 902.02 928.72 ;
     RECT  885.98 435.86 902.5 440.68 ;
     RECT  885.7 1180.52 902.78 1184.92 ;
     RECT  902.02 537.92 903.94 890.08 ;
     RECT  887.62 938.18 904.7 938.38 ;
     RECT  893.38 954.14 906.62 980.8 ;
     RECT  902.02 451.4 907.1 454.12 ;
     RECT  902.78 1176.74 907.1 1184.92 ;
     RECT  890.98 1196.9 907.1 1197.1 ;
     RECT  901.06 1115.84 907.3 1158.46 ;
     RECT  907.1 1176.74 907.3 1197.1 ;
     RECT  904.7 938.18 908.54 939.64 ;
     RECT  902.02 462.74 909.02 462.94 ;
     RECT  899.62 471.56 909.02 527.2 ;
     RECT  907.3 1180.52 911.62 1197.1 ;
     RECT  907.1 448.04 915.26 454.12 ;
     RECT  909.02 462.74 915.26 527.2 ;
     RECT  906.62 949.94 915.46 980.8 ;
     RECT  907.3 1127.18 915.74 1158.46 ;
     RECT  902.5 435.86 916.22 436.06 ;
     RECT  916.22 428.72 918.14 436.06 ;
     RECT  911.62 1180.52 918.14 1181.56 ;
     RECT  908.54 938.18 918.62 941.32 ;
     RECT  902.02 901.64 919.3 928.72 ;
     RECT  915.74 1126.76 920.74 1158.46 ;
     RECT  915.46 957.08 921.5 980.8 ;
     RECT  920.74 1127.18 921.5 1158.46 ;
     RECT  920.54 1210.76 921.5 1210.96 ;
     RECT  921.5 1210.76 921.7 1211.38 ;
     RECT  901.06 991.94 923.42 1105.96 ;
     RECT  921.5 957.08 923.62 981.64 ;
     RECT  918.62 938.18 923.9 948.46 ;
     RECT  918.14 1180.1 925.06 1181.56 ;
     RECT  923.9 938.18 925.54 950.14 ;
     RECT  923.42 991.52 925.82 1105.96 ;
     RECT  907.3 1115.84 925.82 1118.14 ;
     RECT  925.82 991.52 927.46 1118.14 ;
     RECT  911.62 1192.28 928.22 1197.1 ;
     RECT  925.54 938.18 929.38 948.46 ;
     RECT  929.38 938.18 929.86 941.32 ;
     RECT  927.46 991.94 930.34 1118.14 ;
     RECT  918.14 428.72 930.62 437.74 ;
     RECT  915.26 448.04 930.62 527.2 ;
     RECT  930.34 1115.84 930.62 1118.14 ;
     RECT  921.5 1127.18 930.62 1158.88 ;
     RECT  930.62 428.72 931.58 527.2 ;
     RECT  929.86 938.18 931.78 939.64 ;
     RECT  928.22 1192.28 932.06 1200.04 ;
     RECT  925.06 1180.52 932.26 1181.56 ;
     RECT  930.34 991.94 933.22 1105.96 ;
     RECT  931.58 428.72 933.5 527.62 ;
     RECT  919.3 902.06 933.7 928.72 ;
     RECT  932.06 1190.18 933.7 1200.04 ;
     RECT  933.5 425.36 934.66 527.62 ;
     RECT  934.66 451.4 935.14 527.62 ;
     RECT  933.22 1061.24 935.62 1105.96 ;
     RECT  903.94 537.92 935.9 889.66 ;
     RECT  932.26 1180.52 935.9 1181.14 ;
     RECT  930.62 1115.84 936.1 1158.88 ;
     RECT  933.7 1193.12 937.06 1200.04 ;
     RECT  934.66 425.36 938.3 437.74 ;
     RECT  937.06 1199.84 938.5 1200.04 ;
     RECT  935.14 462.74 938.78 527.62 ;
     RECT  935.9 537.5 938.78 889.66 ;
     RECT  938.78 462.74 939.46 889.66 ;
     RECT  936.1 1122.56 939.94 1158.88 ;
     RECT  935.62 1081.82 940.7 1105.96 ;
     RECT  939.94 1143.56 942.14 1158.88 ;
     RECT  942.14 1143.56 942.34 1162.66 ;
     RECT  939.94 1122.56 944.26 1134.94 ;
     RECT  938.3 417.38 944.54 437.74 ;
     RECT  939.46 467.36 944.74 889.66 ;
     RECT  944.26 1127.18 950.3 1134.94 ;
     RECT  942.34 1143.56 950.3 1149.64 ;
     RECT  935.9 1178.42 950.3 1181.14 ;
     RECT  942.34 1158.26 950.98 1162.66 ;
     RECT  950.3 1173.8 951.94 1181.14 ;
     RECT  923.62 960.86 952.22 981.64 ;
     RECT  933.22 991.94 952.22 1051.78 ;
     RECT  944.54 417.38 952.9 440.68 ;
     RECT  935.14 451.4 953.18 454.12 ;
     RECT  950.3 1127.18 953.38 1149.64 ;
     RECT  950.98 1158.26 953.86 1158.88 ;
     RECT  951.94 1173.8 953.86 1174 ;
     RECT  952.22 960.86 954.14 1051.78 ;
     RECT  953.18 451.4 954.62 455.8 ;
     RECT  952.9 432.5 954.82 440.68 ;
     RECT  948.86 1196.9 955.3 1197.1 ;
     RECT  944.74 467.78 956.06 889.66 ;
     RECT  954.14 954.56 956.06 1051.78 ;
     RECT  953.86 1158.26 956.26 1158.46 ;
     RECT  956.06 467.78 957.98 893.02 ;
     RECT  933.7 903.32 957.98 928.72 ;
     RECT  931.78 938.18 957.98 938.38 ;
     RECT  952.9 417.38 958.46 421.36 ;
     RECT  956.06 950.36 958.46 1051.78 ;
     RECT  954.62 451.4 958.94 456.22 ;
     RECT  957.98 467.78 958.94 938.38 ;
     RECT  958.46 950.36 958.94 1052.62 ;
     RECT  958.94 451.4 960.1 1052.62 ;
     RECT  960.1 451.4 960.38 488.98 ;
     RECT  958.46 413.6 962.5 421.36 ;
     RECT  960.1 497.6 963.26 1052.62 ;
     RECT  935.62 1063.34 963.26 1070.68 ;
     RECT  940.7 1081.82 964.7 1112.26 ;
     RECT  953.38 1127.18 964.7 1134.94 ;
     RECT  953.38 1143.56 964.7 1149.64 ;
     RECT  963.26 497.6 966.82 1070.68 ;
     RECT  954.82 432.5 968.54 436.9 ;
     RECT  964.7 1081.82 968.74 1113.1 ;
     RECT  966.82 497.6 969.7 981.64 ;
     RECT  960.38 450.98 971.42 488.98 ;
     RECT  969.7 497.6 971.42 944.68 ;
     RECT  964.7 1127.18 972.38 1149.64 ;
     RECT  962.5 421.16 973.34 421.36 ;
     RECT  966.82 992.36 974.78 1070.68 ;
     RECT  971.42 450.98 974.98 944.68 ;
     RECT  974.78 992.36 975.74 1071.52 ;
     RECT  968.74 1111.64 975.74 1113.1 ;
     RECT  972.38 1123.4 975.74 1149.64 ;
     RECT  968.54 432.5 975.94 440.68 ;
     RECT  969.7 955.4 978.62 981.64 ;
     RECT  975.74 1111.64 978.82 1149.64 ;
     RECT  978.82 1123.4 980.74 1149.64 ;
     RECT  973.34 421.16 981.02 422.2 ;
     RECT  975.94 432.5 981.02 436.9 ;
     RECT  978.62 953.3 981.02 981.64 ;
     RECT  975.74 992.36 981.02 1072.36 ;
     RECT  981.02 953.3 981.22 1072.36 ;
     RECT  981.02 421.16 981.5 436.9 ;
     RECT  981.22 1070.48 981.5 1072.36 ;
     RECT  968.74 1081.82 981.5 1101.76 ;
     RECT  974.98 941.54 982.94 944.68 ;
     RECT  981.22 953.3 982.94 1058.08 ;
     RECT  978.82 1111.64 983.62 1113.52 ;
     RECT  980.74 1127.18 987.26 1149.64 ;
     RECT  981.5 420.74 988.22 436.9 ;
     RECT  974.98 450.98 988.22 930.82 ;
     RECT  981.5 1070.48 988.9 1101.76 ;
     RECT  988.22 420.74 991.58 930.82 ;
     RECT  982.94 941.54 991.58 1058.08 ;
     RECT  987.26 1127.18 993.7 1153.84 ;
     RECT  991.58 420.74 994.18 1058.08 ;
     RECT  994.18 420.74 995.14 985 ;
     RECT  995.14 420.74 995.62 436.9 ;
     RECT  994.18 995.3 997.82 1058.08 ;
     RECT  988.9 1070.48 997.82 1073.2 ;
     RECT  996.38 1174.22 997.82 1174.42 ;
     RECT  995.62 422 1002.34 436.9 ;
     RECT  1002.34 422 1003.3 436.48 ;
     RECT  995.14 451.4 1003.58 981.64 ;
     RECT  997.82 1173.8 1003.58 1174.42 ;
     RECT  997.34 1183.88 1003.58 1184.08 ;
     RECT  1003.58 1173.8 1006.66 1184.08 ;
     RECT  1003.3 429.14 1007.14 436.48 ;
     RECT  1006.66 1173.8 1007.14 1174 ;
     RECT  983.62 1111.64 1007.9 1111.84 ;
     RECT  1003.58 451.4 1008.38 986.68 ;
     RECT  997.82 995.3 1008.38 1073.2 ;
     RECT  1008.38 451.4 1009.34 1073.2 ;
     RECT  988.9 1081.82 1009.34 1101.76 ;
     RECT  1007.14 429.98 1009.54 436.48 ;
     RECT  1009.34 451.4 1011.74 1101.76 ;
     RECT  1007.9 1111.64 1011.74 1116.88 ;
     RECT  1011.74 451.4 1013.38 1116.88 ;
     RECT  1009.82 1166.24 1013.86 1166.44 ;
     RECT  1013.38 466.1 1014.14 1116.88 ;
     RECT  993.7 1127.18 1014.62 1149.64 ;
     RECT  1008.38 1184.72 1014.62 1184.92 ;
     RECT  1014.62 1184.72 1015.58 1188.7 ;
     RECT  1014.14 466.1 1015.78 1118.14 ;
     RECT  1015.78 466.94 1016.26 1118.14 ;
     RECT  1009.54 433.34 1018.66 436.48 ;
     RECT  1015.58 1177.16 1018.66 1188.7 ;
     RECT  1016.26 467.78 1019.9 1118.14 ;
     RECT  1014.62 1126.76 1019.9 1149.64 ;
     RECT  1019.9 467.78 1020.86 1149.64 ;
     RECT  1018.66 1177.16 1021.54 1177.36 ;
     RECT  1018.66 1188.5 1022.78 1188.7 ;
     RECT  1022.78 1188.5 1022.98 1189.54 ;
     RECT  1020.86 467.78 1023.46 1154.68 ;
     RECT  1023.46 467.78 1023.94 1150.06 ;
     RECT  1022.98 1188.5 1027.1 1189.12 ;
     RECT  1023.94 467.78 1028.06 472.18 ;
     RECT  1024.7 1169.6 1028.74 1169.8 ;
     RECT  1013.38 451.4 1031.9 454.12 ;
     RECT  1027.1 1184.3 1033.06 1189.12 ;
     RECT  1031.9 451.4 1034.02 455.8 ;
     RECT  1033.06 1188.92 1035.94 1189.12 ;
     RECT  1023.94 481.22 1036.9 1150.06 ;
     RECT  1033.82 1163.72 1039.58 1163.92 ;
     RECT  1018.66 435.44 1039.78 436.48 ;
     RECT  1028.06 465.68 1041.22 472.18 ;
     RECT  1036.9 481.64 1043.14 1150.06 ;
     RECT  1043.14 481.64 1044.1 1129.48 ;
     RECT  1043.14 1142.3 1044.38 1150.06 ;
     RECT  1039.58 1158.68 1044.38 1163.92 ;
     RECT  1039.78 436.28 1044.58 436.48 ;
     RECT  1039.1 1173.8 1046.02 1174 ;
     RECT  1044.1 484.16 1055.62 1129.48 ;
     RECT  1041.22 468.2 1057.54 472.18 ;
     RECT  1055.62 484.16 1057.54 492.34 ;
     RECT  1055.62 505.16 1057.54 1129.48 ;
     RECT  1044.38 1142.3 1057.54 1163.92 ;
     RECT  1057.54 1142.3 1058.02 1158.88 ;
     RECT  1058.02 1142.3 1058.5 1154.26 ;
     RECT  1057.54 507.68 1058.78 1129.48 ;
     RECT  1058.5 1142.3 1058.78 1150.06 ;
     RECT  1048.22 1174.64 1059.26 1177.36 ;
     RECT  1059.26 1172.54 1059.74 1177.36 ;
     RECT  1058.78 507.68 1060.42 1150.06 ;
     RECT  1057.54 484.16 1064.74 489.4 ;
     RECT  1059.74 1169.6 1064.74 1177.36 ;
     RECT  1064.74 1172.54 1065.02 1177.36 ;
     RECT  1060.42 1142.72 1065.22 1150.06 ;
     RECT  1060.42 507.68 1065.98 1129.48 ;
     RECT  1065.02 1172.54 1068.1 1181.14 ;
     RECT  1065.98 500.96 1070.78 1129.48 ;
     RECT  1070.78 493.4 1070.98 1129.48 ;
     RECT  1068.1 1172.54 1071.94 1175.26 ;
     RECT  1070.98 511.46 1072.22 1129.48 ;
     RECT  1071.94 1172.54 1072.9 1172.74 ;
     RECT  1071.26 1158.68 1073.38 1158.88 ;
     RECT  1070.98 493.4 1073.86 501.16 ;
     RECT  1072.22 511.46 1075.3 1131.58 ;
     RECT  1075.3 511.88 1077.7 1131.58 ;
     RECT  1077.7 511.88 1079.62 1053.88 ;
     RECT  1081.82 1168.76 1083.26 1168.96 ;
     RECT  1065.22 1143.56 1083.74 1150.06 ;
     RECT  1083.26 1168.76 1084.22 1177.36 ;
     RECT  1083.74 1143.56 1084.7 1153.84 ;
     RECT  1079.62 511.88 1085.38 1053.04 ;
     RECT  1073.86 500.96 1086.82 501.16 ;
     RECT  1034.02 451.4 1089.7 454.12 ;
     RECT  1085.38 511.88 1091.14 1048.84 ;
     RECT  1084.7 1143.56 1091.9 1158.88 ;
     RECT  1084.22 1168.76 1091.9 1177.78 ;
     RECT  1077.7 1063.76 1100.26 1131.58 ;
     RECT  1091.9 1143.56 1101.22 1177.78 ;
     RECT  1101.22 1143.56 1101.7 1162.24 ;
     RECT  1101.22 1174.64 1101.7 1177.78 ;
     RECT  1091.14 516.08 1103.14 1048.84 ;
     RECT  1103.14 516.08 1103.62 1045.9 ;
     RECT  1101.7 1174.64 1104.1 1174.84 ;
     RECT  1089.7 451.4 1104.58 451.6 ;
     RECT  1103.62 516.08 1105.06 1045.48 ;
     RECT  1100.26 1063.76 1105.54 1129.06 ;
     RECT  1105.06 516.08 1113.7 1041.7 ;
     RECT  1113.7 533.72 1114.46 1041.7 ;
     RECT  1101.7 1143.56 1114.46 1153.84 ;
     RECT  1105.54 1083.5 1115.42 1129.06 ;
     RECT  1114.46 533.72 1115.9 1048 ;
     RECT  1105.54 1063.76 1115.9 1074.46 ;
     RECT  1115.42 1083.5 1116.58 1133.68 ;
     RECT  1115.9 533.72 1116.86 1074.46 ;
     RECT  1116.58 1083.5 1116.86 1101.76 ;
     RECT  1116.86 533.72 1119.46 1101.76 ;
     RECT  1114.46 1143.56 1119.94 1159.72 ;
     RECT  1116.58 1112.48 1122.34 1133.68 ;
     RECT  1119.46 533.72 1125.7 1098.4 ;
     RECT  1119.94 1149.86 1127.9 1159.72 ;
     RECT  1125.7 1065.86 1128.1 1098.4 ;
     RECT  1127.9 1149.86 1131.26 1166.44 ;
     RECT  1125.7 533.72 1131.46 1056.82 ;
     RECT  1122.34 1112.48 1131.94 1129.48 ;
     RECT  1131.26 1143.56 1132.22 1166.44 ;
     RECT  1131.46 536.66 1134.34 1056.82 ;
     RECT  1132.22 1142.72 1134.82 1166.44 ;
     RECT  1134.82 1142.72 1135.1 1162.24 ;
     RECT  1113.7 516.08 1135.3 524.68 ;
     RECT  1134.34 563.96 1136.54 1056.82 ;
     RECT  1128.1 1070.48 1136.74 1098.4 ;
     RECT  1136.54 563.96 1137.02 1060.18 ;
     RECT  1136.74 1070.48 1137.02 1075.3 ;
     RECT  1131.94 1112.48 1137.22 1124.44 ;
     RECT  1135.1 1136 1137.7 1162.24 ;
     RECT  1137.22 1116.68 1138.66 1124.44 ;
     RECT  1137.7 1136.84 1139.62 1162.24 ;
     RECT  1135.3 524.48 1144.42 524.68 ;
     RECT  1137.02 563.96 1144.42 1075.3 ;
     RECT  1139.62 1142.3 1144.7 1162.24 ;
     RECT  1144.7 1142.3 1147.58 1165.18 ;
     RECT  1147.58 1142.3 1147.78 1166.44 ;
     RECT  1136.74 1086.02 1149.7 1098.4 ;
     RECT  1138.66 1124.24 1149.7 1124.44 ;
     RECT  1134.34 536.66 1151.14 554.08 ;
     RECT  1144.42 1070.48 1151.62 1075.3 ;
     RECT  1151.62 1071.32 1152.1 1075.3 ;
     RECT  1149.7 1090.64 1152.1 1091.26 ;
     RECT  1144.42 563.96 1154.98 1060.6 ;
     RECT  1147.78 1149.86 1155.46 1166.44 ;
     RECT  1152.86 1122.56 1155.94 1122.76 ;
     RECT  1154.98 583.7 1156.42 1060.6 ;
     RECT  1156.42 1052.42 1156.9 1060.6 ;
     RECT  1156.9 1052.84 1157.38 1060.6 ;
     RECT  1157.38 1053.68 1158.34 1060.6 ;
     RECT  1155.46 1154.48 1158.82 1166.44 ;
     RECT  1151.14 541.7 1159.1 554.08 ;
     RECT  1159.1 541.7 1159.3 554.5 ;
     RECT  1159.1 1136 1159.58 1136.2 ;
     RECT  1158.82 1155.74 1159.78 1166.44 ;
     RECT  1154.98 563.96 1160.26 567.52 ;
     RECT  1159.78 1155.74 1161.22 1165.18 ;
     RECT  1152.1 1071.32 1162.66 1071.52 ;
     RECT  1161.22 1155.74 1162.66 1162.66 ;
     RECT  1159.58 1135.58 1163.14 1136.2 ;
     RECT  1162.66 1158.68 1163.14 1161.82 ;
     RECT  1163.14 1135.58 1164.58 1135.78 ;
     RECT  1163.14 1158.68 1164.58 1159.72 ;
     RECT  1152.1 1090.64 1165.06 1090.84 ;
     RECT  1164.58 1159.52 1165.06 1159.72 ;
     RECT  1158.34 1053.68 1166.02 1056.82 ;
     RECT  1166.02 1053.68 1166.98 1053.88 ;
     RECT  1166.78 1120.46 1167.74 1120.66 ;
     RECT  1167.74 1120.04 1169.18 1120.66 ;
     RECT  1064.74 484.16 1169.86 484.36 ;
     RECT  1156.42 583.7 1170.34 1041.28 ;
     RECT  1170.34 983.54 1171.78 1041.28 ;
     RECT  1170.34 583.7 1173.7 973.24 ;
     RECT  1171.78 983.96 1174.46 1041.28 ;
     RECT  1159.3 541.7 1174.66 549.04 ;
     RECT  1169.18 1120.04 1176.1 1124.44 ;
     RECT  1172.54 1078.88 1177.34 1079.08 ;
     RECT  1177.34 1070.48 1177.54 1079.08 ;
     RECT  1177.54 1070.48 1178.3 1072.36 ;
     RECT  1176.1 1120.04 1178.5 1123.6 ;
     RECT  1174.46 983.96 1179.94 1042.12 ;
     RECT  1178.5 1120.04 1179.94 1121.08 ;
     RECT  1174.66 541.7 1180.42 541.9 ;
     RECT  1180.7 1105.76 1181.18 1105.96 ;
     RECT  1175.9 1090.22 1181.38 1090.42 ;
     RECT  1181.18 1105.76 1183.78 1113.1 ;
     RECT  1183.78 1105.76 1184.06 1106.38 ;
     RECT  1178.3 1063.76 1186.94 1072.36 ;
     RECT  1184.06 1102.4 1186.94 1106.38 ;
     RECT  1186.94 1056.2 1187.14 1072.36 ;
     RECT  1187.14 1056.2 1187.9 1057.24 ;
     RECT  1186.94 1094 1192.42 1106.38 ;
     RECT  1173.7 583.7 1192.7 641.44 ;
     RECT  1179.94 983.96 1192.9 1041.28 ;
     RECT  1187.14 1071.32 1193.38 1071.52 ;
     RECT  1192.7 579.92 1193.66 641.44 ;
     RECT  1187.9 1052.84 1193.86 1057.24 ;
     RECT  1192.9 1037.3 1194.82 1041.28 ;
     RECT  1160.26 565.64 1195.1 567.52 ;
     RECT  1193.66 576.56 1195.1 641.44 ;
     RECT  1194.82 1038.56 1196.26 1041.28 ;
     RECT  1195.1 557.66 1196.74 641.44 ;
     RECT  1193.86 1053.26 1197.98 1057.24 ;
     RECT  1192.42 1094 1198.66 1102.6 ;
     RECT  1196.74 564.8 1198.94 641.44 ;
     RECT  1173.7 650.48 1198.94 973.24 ;
     RECT  1198.94 564.8 1200.1 973.24 ;
     RECT  1196.26 1041.08 1200.58 1041.28 ;
     RECT  1198.66 1102.4 1200.58 1102.6 ;
     RECT  1200.1 564.8 1201.54 748.96 ;
     RECT  1200.1 758.42 1201.54 973.24 ;
     RECT  1201.54 761.36 1202.5 973.24 ;
     RECT  1197.98 1053.26 1202.98 1060.6 ;
     RECT  1202.98 1053.26 1203.74 1055.98 ;
     RECT  1201.54 579.92 1204.42 748.96 ;
     RECT  1203.74 1045.28 1204.42 1055.98 ;
     RECT  1204.42 1055.78 1205.38 1055.98 ;
     RECT  1202.5 765.56 1205.66 973.24 ;
     RECT  1192.9 983.96 1205.66 1026.58 ;
     RECT  1195.58 508.94 1206.34 509.14 ;
     RECT  1204.42 1045.28 1206.34 1045.48 ;
     RECT  1205.66 765.56 1207.3 1026.58 ;
     RECT  1201.54 564.8 1207.78 567.52 ;
     RECT  1207.3 765.56 1208.74 1022.8 ;
     RECT  1204.42 579.92 1209.7 635.98 ;
     RECT  1208.74 765.56 1209.7 964 ;
     RECT  1208.74 973.04 1209.7 1022.8 ;
     RECT  1207.58 504.32 1213.82 504.52 ;
     RECT  1204.42 647.54 1214.78 706.12 ;
     RECT  1213.34 538.34 1215.74 538.54 ;
     RECT  1209.7 983.96 1216.42 1022.8 ;
     RECT  1215.74 538.34 1217.38 539.8 ;
     RECT  1214.78 647.12 1217.66 706.12 ;
     RECT  1204.42 716.42 1217.66 748.96 ;
     RECT  1209.7 765.56 1222.66 887.14 ;
     RECT  1209.7 579.92 1223.9 633.88 ;
     RECT  1222.66 765.56 1224.1 886.3 ;
     RECT  1217.66 647.12 1225.54 748.96 ;
     RECT  1213.82 496.76 1226.98 504.52 ;
     RECT  1207.78 565.64 1229.66 567.52 ;
     RECT  1225.54 647.12 1230.14 727.12 ;
     RECT  1229.66 565.64 1231.58 568.78 ;
     RECT  1209.7 896.18 1232.06 964 ;
     RECT  1209.7 973.04 1232.06 973.24 ;
     RECT  1216.42 983.96 1232.54 1018.6 ;
     RECT  1223.9 578.66 1233.5 633.88 ;
     RECT  1230.14 646.28 1233.5 727.12 ;
     RECT  1231.58 565.64 1233.98 569.2 ;
     RECT  1233.5 578.66 1233.98 727.12 ;
     RECT  1232.06 896.18 1234.66 973.24 ;
     RECT  1225.54 739.1 1237.06 748.96 ;
     RECT  1224.1 765.56 1238.98 885.88 ;
     RECT  1217.38 538.34 1239.46 538.54 ;
     RECT  1233.98 565.64 1240.42 727.12 ;
     RECT  1238.98 822.68 1240.9 885.88 ;
     RECT  1232.54 983.54 1240.9 1018.6 ;
     RECT  1238.98 765.56 1241.38 812.38 ;
     RECT  1240.9 836.96 1241.38 885.88 ;
     RECT  1241.38 840.74 1242.34 885.88 ;
     RECT  1242.34 854.6 1245.02 885.88 ;
     RECT  1245.02 854.6 1245.22 886.72 ;
     RECT  1241.38 765.56 1245.7 802.72 ;
     RECT  1240.9 983.96 1246.18 1018.6 ;
     RECT  1246.18 983.96 1246.66 1015.66 ;
     RECT  1245.22 870.98 1248.58 886.72 ;
     RECT  1240.9 822.68 1249.06 825.82 ;
     RECT  1240.42 565.64 1249.82 580.12 ;
     RECT  1240.42 592.94 1250.02 727.12 ;
     RECT  1250.02 592.94 1250.3 633.88 ;
     RECT  1237.06 742.88 1250.3 748.96 ;
     RECT  1242.34 840.74 1250.98 845.98 ;
     RECT  1248.58 870.98 1250.98 885.88 ;
     RECT  1249.82 565.64 1251.26 581.38 ;
     RECT  1250.3 591.68 1251.26 633.88 ;
     RECT  1234.66 896.18 1251.46 964 ;
     RECT  1250.3 736.58 1252.9 748.96 ;
     RECT  1251.26 565.64 1253.38 633.88 ;
     RECT  1252.9 736.58 1253.38 746.02 ;
     RECT  1250.98 870.98 1253.86 882.94 ;
     RECT  1253.38 565.64 1254.82 633.04 ;
     RECT  1250.02 647.54 1255.3 727.12 ;
     RECT  1245.7 765.98 1256.26 802.72 ;
     RECT  1251.46 897.86 1256.54 964 ;
     RECT  1234.66 973.04 1256.54 973.24 ;
     RECT  1255.3 647.96 1256.74 727.12 ;
     RECT  1256.54 897.86 1256.74 973.24 ;
     RECT  1253.38 736.58 1257.22 743.08 ;
     RECT  1254.82 565.64 1257.7 577.18 ;
     RECT  1254.82 585.8 1257.7 633.04 ;
     RECT  1256.74 938.18 1257.7 973.24 ;
     RECT  1257.7 586.64 1258.18 633.04 ;
     RECT  1257.22 736.58 1258.18 742.24 ;
     RECT  1257.7 565.64 1258.66 574.24 ;
     RECT  1256.74 897.86 1258.66 923.68 ;
     RECT  1257.7 942.8 1258.66 973.24 ;
     RECT  1258.66 565.64 1259.14 573.82 ;
     RECT  1241.38 812.18 1259.14 812.38 ;
     RECT  1259.14 565.64 1259.62 570.46 ;
     RECT  1258.18 613.52 1259.62 633.04 ;
     RECT  1258.66 903.32 1259.62 923.68 ;
     RECT  1259.62 615.62 1260.1 633.04 ;
     RECT  1256.74 647.96 1260.1 705.7 ;
     RECT  1245.22 854.6 1260.1 862.36 ;
     RECT  1259.62 903.32 1260.1 911.5 ;
     RECT  1259.62 920.12 1261.06 923.68 ;
     RECT  1250.98 845.78 1261.54 845.98 ;
     RECT  1260.86 534.98 1263.46 535.18 ;
     RECT  1258.18 586.64 1263.46 597.76 ;
     RECT  1263.46 587.48 1263.94 597.76 ;
     RECT  1256.26 765.98 1265.86 797.26 ;
     RECT  1263.94 587.9 1266.34 588.1 ;
     RECT  1261.06 923.48 1266.34 923.68 ;
     RECT  1246.66 983.96 1266.34 1014.82 ;
     RECT  1258.18 742.04 1266.82 742.24 ;
     RECT  1260.1 903.32 1267.3 907.72 ;
     RECT  1266.34 1009.58 1267.3 1014.82 ;
     RECT  1249.06 822.68 1267.78 822.88 ;
     RECT  1266.34 983.96 1267.78 999.28 ;
     RECT  1267.3 1010 1267.78 1014.82 ;
     RECT  1259.62 565.64 1268.26 567.52 ;
     RECT  1267.78 983.96 1268.26 985 ;
     RECT  1268.26 984.8 1268.74 985 ;
     RECT  1260.1 647.96 1272.1 703.6 ;
     RECT  1267.78 993.62 1272.1 999.28 ;
     RECT  1272.1 999.08 1272.58 999.28 ;
     RECT  1267.78 1014.62 1273.06 1014.82 ;
     RECT  1260.1 615.62 1281.7 631.36 ;
     RECT  1272.1 652.58 1281.7 703.6 ;
     RECT  1057.54 469.04 1288.9 472.18 ;
     RECT  1226.98 504.32 1288.9 504.52 ;
     RECT  1268.26 567.32 1288.9 567.52 ;
     RECT  1263.94 597.56 1288.9 597.76 ;
     RECT  1281.7 615.62 1288.9 621.7 ;
     RECT  1281.7 652.58 1288.9 673.36 ;
     RECT  1281.7 683.24 1288.9 703.6 ;
     RECT  1260.1 862.16 1288.9 862.36 ;
     RECT  1253.86 874.34 1288.9 882.94 ;
     RECT  1267.3 907.52 1288.9 907.72 ;
     RECT  1258.66 950.36 1288.9 964 ;
     RECT  1258.66 973.04 1288.9 973.24 ;
     RECT  1288.9 656.78 1289.38 671.26 ;
     RECT  1288.9 874.34 1289.38 874.54 ;
     RECT  1288.9 961.28 1289.38 961.48 ;
     RECT  1289.38 666.44 1289.86 671.26 ;
     RECT  1289.38 656.78 1290.34 656.98 ;
     RECT  1256.74 716.42 1294.18 727.12 ;
     RECT  1265.86 789.08 1294.18 797.26 ;
     RECT  1265.86 765.98 1294.66 777.1 ;
     RECT  1294.66 773.12 1295.14 777.1 ;
     RECT  1294.18 789.08 1295.62 789.28 ;
     RECT  1294.18 723.14 1297.06 727.12 ;
     RECT  1281.7 631.16 1298.02 631.36 ;
     RECT  1288.9 685.76 1298.02 702.34 ;
     RECT  1298.02 685.76 1298.5 694.36 ;
     RECT  1295.14 776.9 1298.5 777.1 ;
     RECT  1289.86 671.06 1298.98 671.26 ;
     RECT  1297.06 726.92 1298.98 727.12 ;
    LAYER Metal5 ;
     RECT  933.5 453.5 933.7 462.74 ;
     RECT  933.5 462.74 939.46 491.92 ;
     RECT  974.78 463.16 974.98 495.5 ;
     RECT  974.78 495.5 977.86 502.84 ;
     RECT  887.9 472.4 888.1 504.1 ;
     RECT  977.18 502.84 977.86 504.74 ;
     RECT  935.9 491.92 939.46 508.1 ;
     RECT  951.26 511.46 951.46 518.6 ;
     RECT  931.58 508.1 939.46 520.28 ;
     RECT  977.18 504.74 978.82 520.9 ;
     RECT  977.18 520.9 978.34 522.16 ;
     RECT  951.26 518.6 959.62 524.9 ;
     RECT  931.1 520.28 939.46 528.46 ;
     RECT  989.66 521.54 989.86 535.6 ;
     RECT  977.18 522.16 977.38 537.28 ;
     RECT  935.9 528.46 939.46 538.96 ;
     RECT  935.9 538.96 937.06 541.48 ;
     RECT  951.26 524.9 960.58 558.08 ;
     RECT  936.38 541.48 937.06 561.64 ;
     RECT  1029.98 540.02 1030.18 565 ;
     RECT  918.62 549.68 918.82 567.1 ;
     RECT  951.26 558.08 968.26 569.2 ;
     RECT  936.86 561.64 937.06 572.78 ;
     RECT  994.46 563.12 994.66 577.82 ;
     RECT  967.58 569.2 968.26 578.24 ;
     RECT  859.1 554.3 859.3 579.7 ;
     RECT  936.86 572.78 939.94 579.92 ;
     RECT  934.94 579.92 939.94 580.34 ;
     RECT  951.26 569.2 956.74 580.34 ;
     RECT  967.58 578.24 969.22 580.34 ;
     RECT  979.1 562.28 979.3 580.34 ;
     RECT  1107.74 576.98 1107.94 580.54 ;
     RECT  934.94 580.34 956.74 581.18 ;
     RECT  967.58 580.34 979.3 581.18 ;
     RECT  934.94 581.18 979.3 583.28 ;
     RECT  994.46 577.82 998.5 583.7 ;
     RECT  906.62 583.28 906.82 584.12 ;
     RECT  906.62 584.12 916.42 584.54 ;
     RECT  933.02 583.28 979.3 584.54 ;
     RECT  906.62 584.54 979.3 588.1 ;
     RECT  994.46 583.7 998.98 591.68 ;
     RECT  1198.94 553.88 1199.14 597.56 ;
     RECT  906.62 588.1 953.38 597.98 ;
     RECT  906.62 597.98 953.86 599.02 ;
     RECT  989.66 591.68 998.98 599.02 ;
     RECT  964.7 588.1 979.3 600.08 ;
     RECT  989.66 599.02 998.5 600.08 ;
     RECT  1250.78 582.02 1250.98 600.28 ;
     RECT  1098.14 600.08 1098.34 600.5 ;
     RECT  916.22 599.02 953.86 600.7 ;
     RECT  964.7 600.08 998.5 601.12 ;
     RECT  1098.14 600.5 1099.3 601.2 ;
     RECT  1109.18 602.18 1109.38 604.28 ;
     RECT  916.22 600.7 940.42 604.9 ;
     RECT  1151.9 602.18 1152.1 604.9 ;
     RECT  964.7 601.12 985.54 608.26 ;
     RECT  953.18 600.7 953.86 611 ;
     RECT  1109.18 604.28 1117.54 611.62 ;
     RECT  1109.18 611.62 1114.18 612.04 ;
     RECT  1137.5 600.92 1137.7 612.26 ;
     RECT  964.7 608.26 980.74 614.56 ;
     RECT  1129.82 612.26 1137.7 614.56 ;
     RECT  924.86 604.9 940.42 615.62 ;
     RECT  952.22 611 953.86 615.62 ;
     RECT  1081.34 602.18 1081.54 620.02 ;
     RECT  1110.14 612.04 1114.18 620.02 ;
     RECT  924.86 615.62 954.82 621.28 ;
     RECT  1039.1 614.36 1039.3 621.5 ;
     RECT  926.3 621.28 954.82 623.6 ;
     RECT  998.3 601.12 998.5 623.6 ;
     RECT  926.3 623.6 955.3 624.44 ;
     RECT  967.58 614.56 980.74 624.44 ;
     RECT  1110.14 620.02 1112.74 625.48 ;
     RECT  926.3 624.44 980.74 626.12 ;
     RECT  992.06 623.6 998.5 626.12 ;
     RECT  926.3 626.12 998.5 627.58 ;
     RECT  967.1 627.58 998.5 628.42 ;
     RECT  1158.62 625.7 1158.82 632.62 ;
     RECT  1034.78 621.5 1039.3 632.84 ;
     RECT  967.1 628.42 967.78 637.66 ;
     RECT  926.3 627.58 953.86 638.08 ;
     RECT  1245.98 631.16 1246.18 640.4 ;
     RECT  1110.14 625.48 1110.34 640.6 ;
     RECT  1033.82 632.84 1039.3 643.54 ;
     RECT  1198.94 597.56 1202.02 643.54 ;
     RECT  1034.3 643.54 1039.3 644.38 ;
     RECT  979.1 628.42 998.5 646.06 ;
     RECT  1034.3 644.38 1038.34 646.06 ;
     RECT  1034.78 646.06 1038.34 648.16 ;
     RECT  926.3 638.08 934.18 650.68 ;
     RECT  926.3 650.68 929.86 651.94 ;
     RECT  1201.82 643.54 1202.02 652.36 ;
     RECT  926.3 651.94 926.5 654.04 ;
     RECT  945.02 638.08 953.86 655.3 ;
     RECT  1244.06 640.4 1246.18 655.3 ;
     RECT  1129.82 614.56 1130.02 655.94 ;
     RECT  1034.78 648.16 1034.98 656.56 ;
     RECT  1112.06 657.2 1112.26 657.62 ;
     RECT  1129.82 655.94 1134.34 659.72 ;
     RECT  1084.22 654.68 1084.42 660.76 ;
     RECT  979.1 646.06 993.22 666.44 ;
     RECT  1129.82 659.72 1136.74 669.16 ;
     RECT  979.1 666.44 999.94 670 ;
     RECT  1129.82 669.16 1134.34 670 ;
     RECT  1250.78 656.36 1250.98 670 ;
     RECT  949.82 655.3 953.86 670.42 ;
     RECT  1212.38 669.38 1216.42 672.74 ;
     RECT  1031.42 660.98 1031.62 673.16 ;
     RECT  1112.06 657.62 1115.14 676.52 ;
     RECT  1112.06 676.52 1122.82 679.88 ;
     RECT  1031.42 673.16 1035.94 682.18 ;
     RECT  1211.9 672.74 1216.42 685.96 ;
     RECT  979.1 670 993.22 687.02 ;
     RECT  1035.74 682.18 1035.94 688.48 ;
     RECT  979.1 687.02 999.46 690.16 ;
     RECT  979.1 690.16 993.22 692.68 ;
     RECT  1110.62 679.88 1122.82 693.32 ;
     RECT  1134.14 670 1134.34 694.36 ;
     RECT  1109.18 693.32 1122.82 696.04 ;
     RECT  967.58 637.66 967.78 696.68 ;
     RECT  979.1 692.68 990.34 696.68 ;
     RECT  953.18 670.42 953.86 698.14 ;
     RECT  967.58 696.68 990.34 698.14 ;
     RECT  979.1 698.14 990.34 705.7 ;
     RECT  1008.38 702.14 1008.58 705.7 ;
     RECT  1074.62 679.88 1074.82 705.7 ;
     RECT  1110.62 696.04 1122.82 705.7 ;
     RECT  1211.9 685.96 1212.1 705.7 ;
     RECT  921.02 692.9 921.22 708.64 ;
     RECT  1114.46 705.7 1122.82 710.54 ;
     RECT  1114.46 710.54 1127.62 711.8 ;
     RECT  907.58 683.66 907.78 712.22 ;
     RECT  967.58 698.14 967.78 713.26 ;
     RECT  979.1 705.7 984.1 715.78 ;
     RECT  907.58 712.22 908.26 719.14 ;
     RECT  983.9 715.78 984.1 719.36 ;
     RECT  983.9 719.36 984.58 719.98 ;
     RECT  856.22 717.26 856.42 720.82 ;
     RECT  984.38 719.98 984.58 720.82 ;
     RECT  1245.02 719.78 1245.22 720.82 ;
     RECT  1114.46 711.8 1129.06 722.5 ;
     RECT  784.22 728.18 784.42 729.02 ;
     RECT  870.62 722.3 870.82 730.9 ;
     RECT  730.94 733.64 731.14 734.06 ;
     RECT  1114.46 722.5 1128.1 734.26 ;
     RECT  728.54 734.06 731.14 734.48 ;
     RECT  728.54 734.48 731.62 734.9 ;
     RECT  781.34 729.02 784.42 738.68 ;
     RECT  728.54 734.9 732.58 739.52 ;
     RECT  975.26 739.1 975.46 741.62 ;
     RECT  1142.78 728.18 1142.98 741.62 ;
     RECT  1142.78 741.62 1143.46 745.4 ;
     RECT  728.54 739.52 737.38 745.82 ;
     RECT  973.34 741.62 975.46 748.54 ;
     RECT  990.62 746.24 990.82 750.44 ;
     RECT  1122.62 734.26 1128.1 750.44 ;
     RECT  728.54 745.82 743.14 750.64 ;
     RECT  907.58 719.14 907.78 751.28 ;
     RECT  1142.78 745.4 1147.3 755.26 ;
     RECT  781.34 738.68 789.22 755.9 ;
     RECT  990.62 750.44 991.3 755.9 ;
     RECT  1101.98 753.38 1102.18 755.9 ;
     RECT  1122.62 750.44 1132.42 756.1 ;
     RECT  772.7 755.9 789.22 756.32 ;
     RECT  953.18 698.14 953.38 757.36 ;
     RECT  728.54 750.64 741.22 758 ;
     RECT  1127.9 756.1 1132.42 758 ;
     RECT  1147.1 755.26 1147.3 758 ;
     RECT  905.18 751.28 907.78 760.94 ;
     RECT  905.18 760.94 912.1 761.36 ;
     RECT  1147.1 758 1149.22 761.36 ;
     RECT  1147.1 761.36 1154.98 761.56 ;
     RECT  905.18 761.36 913.06 761.78 ;
     RECT  727.58 758 741.22 761.98 ;
     RECT  1127.9 758 1135.78 764.08 ;
     RECT  990.62 755.9 1009.06 765.34 ;
     RECT  974.3 748.54 975.46 765.56 ;
     RECT  990.62 765.34 1005.22 765.56 ;
     RECT  772.7 756.32 790.66 765.76 ;
     RECT  1101.98 755.9 1105.06 766.4 ;
     RECT  761.66 753.8 761.86 766.6 ;
     RECT  772.7 765.76 772.9 767.02 ;
     RECT  937.34 765.98 937.54 768.08 ;
     RECT  1149.02 761.56 1154.98 769.34 ;
     RECT  785.66 765.76 790.66 769.76 ;
     RECT  729.98 761.98 741.22 770.18 ;
     RECT  785.66 769.76 792.1 770.18 ;
     RECT  1135.58 764.08 1135.78 770.38 ;
     RECT  729.98 770.18 744.1 770.8 ;
     RECT  737.66 770.8 744.1 771.22 ;
     RECT  785.66 770.18 793.06 771.22 ;
     RECT  937.34 768.08 939.94 771.22 ;
     RECT  960.86 769.76 961.06 772.7 ;
     RECT  1196.06 768.5 1196.26 773.54 ;
     RECT  737.66 771.22 741.22 774.16 ;
     RECT  789.02 771.22 793.06 775.84 ;
     RECT  937.34 771.22 937.54 775.84 ;
     RECT  636.86 765.98 637.06 776.26 ;
     RECT  789.02 775.84 792.1 778.78 ;
     RECT  957.98 772.7 961.06 780.68 ;
     RECT  974.3 765.56 1005.22 780.68 ;
     RECT  1074.14 755.9 1074.34 780.68 ;
     RECT  791.9 778.78 792.1 780.88 ;
     RECT  741.02 774.16 741.22 788.02 ;
     RECT  1101.98 766.4 1108.42 788.86 ;
     RECT  1074.14 780.68 1080.58 789.7 ;
     RECT  1051.58 782.78 1051.78 789.92 ;
     RECT  1149.02 769.34 1158.34 790.76 ;
     RECT  1196.06 773.54 1197.22 791.18 ;
     RECT  1196.06 791.18 1201.54 791.6 ;
     RECT  1149.02 790.76 1166.02 794.54 ;
     RECT  1080.38 789.7 1080.58 794.74 ;
     RECT  1120.7 794.54 1120.9 795.8 ;
     RECT  1186.46 791.6 1201.54 796.22 ;
     RECT  957.98 780.68 1005.22 797.48 ;
     RECT  1120.7 795.8 1128.58 797.9 ;
     RECT  957.98 797.48 1011.46 799.16 ;
     RECT  1101.98 788.86 1105.06 799.16 ;
     RECT  904.22 761.78 913.06 800.42 ;
     RECT  1186.46 796.22 1202.98 800.62 ;
     RECT  1098.62 799.16 1105.06 800.84 ;
     RECT  1117.34 797.9 1128.58 801.26 ;
     RECT  1148.06 794.54 1166.02 801.26 ;
     RECT  1045.82 789.92 1051.78 803.36 ;
     RECT  904.22 800.42 918.34 804.62 ;
     RECT  956.06 799.16 1011.46 804.82 ;
     RECT  1038.14 803.36 1051.78 805.88 ;
     RECT  1116.86 801.26 1128.58 805.88 ;
     RECT  956.06 804.82 962.5 806.3 ;
     RECT  976.7 804.82 1011.46 806.5 ;
     RECT  1095.74 800.84 1105.06 806.72 ;
     RECT  1116.86 805.88 1137.22 806.72 ;
     RECT  1148.06 801.26 1169.86 806.72 ;
     RECT  1023.26 803.36 1023.46 807.14 ;
     RECT  1038.14 805.88 1053.7 807.14 ;
     RECT  1116.86 806.72 1169.86 807.76 ;
     RECT  1023.26 807.14 1053.7 810.08 ;
     RECT  1116.86 807.76 1120.9 810.7 ;
     RECT  1195.58 800.62 1202.98 810.7 ;
     RECT  894.62 804.62 918.34 810.92 ;
     RECT  894.62 810.92 923.14 811.34 ;
     RECT  886.46 811.34 923.14 811.96 ;
     RECT  1023.26 810.08 1056.1 812.6 ;
     RECT  1066.46 810.5 1074.34 812.6 ;
     RECT  1131.74 807.76 1169.86 812.6 ;
     RECT  1089.02 806.72 1105.06 813.02 ;
     RECT  1131.74 812.6 1175.62 813.22 ;
     RECT  1023.26 812.6 1074.34 813.86 ;
     RECT  1133.18 813.22 1175.62 814.06 ;
     RECT  1196.06 810.7 1202.98 814.06 ;
     RECT  976.7 806.5 990.34 817.64 ;
     RECT  1002.14 806.5 1011.46 817.64 ;
     RECT  952.7 806.3 962.5 818.48 ;
     RECT  976.7 817.64 1011.46 818.48 ;
     RECT  1022.3 813.86 1074.34 818.48 ;
     RECT  886.46 811.96 894.82 819.52 ;
     RECT  976.7 818.48 1074.34 819.74 ;
     RECT  1137.02 814.06 1175.62 819.94 ;
     RECT  1137.02 819.94 1174.18 820.36 ;
     RECT  973.34 819.74 1074.34 820.78 ;
     RECT  1196.06 814.06 1201.54 820.78 ;
     RECT  1226.3 807.14 1226.5 820.78 ;
     RECT  1118.3 810.7 1120.9 821.84 ;
     RECT  1089.02 813.02 1106.98 822.04 ;
     RECT  1139.9 820.36 1174.18 822.46 ;
     RECT  1140.38 822.46 1174.18 823.3 ;
     RECT  952.7 818.48 962.98 825.62 ;
     RECT  1041.98 820.78 1074.34 826.24 ;
     RECT  1118.3 821.84 1122.34 826.46 ;
     RECT  1140.38 823.3 1172.26 827.5 ;
     RECT  894.62 819.52 894.82 828.34 ;
     RECT  944.06 825.62 962.98 828.34 ;
     RECT  1041.98 826.24 1042.66 829.18 ;
     RECT  952.7 828.34 962.98 830.02 ;
     RECT  1053.5 826.24 1074.34 830.66 ;
     RECT  1089.02 822.04 1103.14 830.66 ;
     RECT  973.34 820.78 1032.1 830.86 ;
     RECT  1114.94 826.46 1122.34 830.86 ;
     RECT  1031.9 830.86 1032.1 834.64 ;
     RECT  857.18 811.34 857.38 835.48 ;
     RECT  907.58 811.96 923.14 836.32 ;
     RECT  1041.98 829.18 1042.18 836.32 ;
     RECT  1053.5 830.66 1103.14 838.22 ;
     RECT  1114.94 830.86 1121.38 838.22 ;
     RECT  908.54 836.32 923.14 839.06 ;
     RECT  1140.38 827.5 1144.9 840.32 ;
     RECT  1154.78 827.5 1172.26 840.32 ;
     RECT  1140.38 840.32 1172.26 842 ;
     RECT  1053.5 838.22 1121.38 842.42 ;
     RECT  1140.38 842 1174.18 842.42 ;
     RECT  908.54 839.06 923.62 843.04 ;
     RECT  1140.38 842.42 1181.38 843.26 ;
     RECT  1052.06 842.42 1121.38 843.88 ;
     RECT  973.34 830.86 1021.54 845.14 ;
     RECT  1039.58 838.64 1040.26 848.92 ;
     RECT  1114.94 843.88 1121.38 848.92 ;
     RECT  1119.74 848.92 1121.38 849.34 ;
     RECT  952.7 830.02 962.5 851.02 ;
     RECT  1140.38 843.26 1185.22 851.02 ;
     RECT  908.54 843.04 914.02 851.86 ;
     RECT  908.54 851.86 912.1 853.12 ;
     RECT  1012.7 845.14 1021.54 853.12 ;
     RECT  956.06 851.02 962.5 853.34 ;
     RECT  973.34 845.14 1002.34 853.34 ;
     RECT  1140.38 851.02 1178.98 853.34 ;
     RECT  1119.74 849.34 1120.9 853.54 ;
     RECT  1240.7 806.72 1240.9 853.96 ;
     RECT  1052.06 843.88 1103.62 854.8 ;
     RECT  1120.7 853.54 1120.9 855.64 ;
     RECT  908.54 853.12 908.74 856.06 ;
     RECT  1137.5 853.34 1178.98 856.06 ;
     RECT  956.06 853.34 1002.34 856.28 ;
     RECT  1012.7 853.12 1012.9 856.28 ;
     RECT  1074.14 854.8 1103.62 856.28 ;
     RECT  956.06 856.28 1012.9 856.48 ;
     RECT  1052.06 854.8 1062.34 856.7 ;
     RECT  1074.14 856.28 1107.46 856.9 ;
     RECT  1143.74 856.06 1178.98 856.9 ;
     RECT  1074.14 856.9 1077.7 857.32 ;
     RECT  1168.7 856.9 1178.98 857.74 ;
     RECT  931.1 854.18 931.3 859.64 ;
     RECT  1093.34 856.9 1107.46 860.48 ;
     RECT  1209.02 856.7 1209.22 860.68 ;
     RECT  1093.34 860.48 1107.94 860.9 ;
     RECT  1093.34 860.9 1109.38 861.1 ;
     RECT  929.18 859.64 931.3 861.52 ;
     RECT  1045.82 856.7 1062.34 864.88 ;
     RECT  1024.22 863 1024.42 865.52 ;
     RECT  1100.54 861.1 1109.38 865.72 ;
     RECT  1143.74 856.9 1158.82 866.78 ;
     RECT  1133.66 866.78 1158.82 867.4 ;
     RECT  1023.26 865.52 1024.42 867.82 ;
     RECT  1045.82 864.88 1061.86 867.82 ;
     RECT  1045.82 867.82 1047.94 868.04 ;
     RECT  1023.26 867.82 1023.46 868.66 ;
     RECT  1143.74 867.4 1158.82 869.08 ;
     RECT  1101.02 865.72 1109.38 869.5 ;
     RECT  1059.74 867.82 1061.86 870.34 ;
     RECT  1173.98 857.74 1178.98 870.56 ;
     RECT  929.18 861.52 929.38 871.18 ;
     RECT  956.06 856.48 1007.62 871.18 ;
     RECT  1171.58 870.56 1178.98 871.4 ;
     RECT  1101.02 869.5 1107.46 871.6 ;
     RECT  1171.1 871.4 1178.98 871.6 ;
     RECT  1043.42 868.04 1047.94 873.28 ;
     RECT  956.06 871.18 964.42 874.12 ;
     RECT  1077.5 857.32 1077.7 874.12 ;
     RECT  1146.62 869.08 1158.82 874.54 ;
     RECT  1171.1 871.6 1178.5 874.54 ;
     RECT  1171.1 874.54 1173.22 875.38 ;
     RECT  713.66 863.42 713.86 875.8 ;
     RECT  1171.58 875.38 1173.22 876.22 ;
     RECT  1171.58 876.22 1171.78 880 ;
     RECT  976.7 871.18 1007.62 881.9 ;
     RECT  976.7 881.9 1012.9 882.52 ;
     RECT  1045.82 873.28 1047.94 883.36 ;
     RECT  1045.82 883.36 1046.02 884.2 ;
     RECT  1146.62 874.54 1158.34 886.1 ;
     RECT  981.5 882.52 1012.9 886.3 ;
     RECT  1196.06 820.78 1197.22 890.08 ;
     RECT  956.06 874.12 961.06 893.02 ;
     RECT  1143.26 886.1 1158.34 893.24 ;
     RECT  1059.74 870.34 1059.94 894.5 ;
     RECT  1056.86 894.5 1059.94 894.92 ;
     RECT  1101.98 871.6 1107.46 895.12 ;
     RECT  982.46 886.3 1012.9 896.38 ;
     RECT  1091.42 887.78 1091.62 897.44 ;
     RECT  1101.98 895.12 1102.18 897.44 ;
     RECT  572.06 856.7 572.26 898.48 ;
     RECT  1056.86 894.92 1061.86 899.32 ;
     RECT  991.1 896.38 1012.9 899.74 ;
     RECT  1057.82 899.32 1061.86 899.96 ;
     RECT  765.5 889.88 765.7 901.84 ;
     RECT  1140.38 893.24 1158.34 905.84 ;
     RECT  1178.3 893.66 1178.5 905.84 ;
     RECT  1140.38 905.84 1161.22 906.68 ;
     RECT  1091.42 897.44 1102.18 907.52 ;
     RECT  1140.38 906.68 1161.7 907.52 ;
     RECT  1177.34 905.84 1178.5 907.52 ;
     RECT  1091.42 907.52 1113.7 908.36 ;
     RECT  993.02 899.74 1012.9 909.2 ;
     RECT  1197.02 890.08 1197.22 909.2 ;
     RECT  1032.38 907.1 1040.74 909.62 ;
     RECT  1077.02 906.52 1078.66 909.62 ;
     RECT  1091.42 908.36 1119.46 909.62 ;
     RECT  1140.38 907.52 1178.5 910.88 ;
     RECT  1194.62 909.2 1197.22 910.88 ;
     RECT  1140.38 910.88 1197.22 911.3 ;
     RECT  1032.38 909.62 1047.46 911.72 ;
     RECT  1057.82 899.96 1067.14 911.72 ;
     RECT  1077.02 909.62 1119.46 912.98 ;
     RECT  1133.18 911.3 1197.22 912.98 ;
     RECT  1032.38 911.72 1067.14 914.66 ;
     RECT  1077.02 912.98 1197.22 914.66 ;
     RECT  993.02 909.2 1021.54 916.76 ;
     RECT  1032.38 914.66 1197.22 916.76 ;
     RECT  957.98 893.02 961.06 916.96 ;
     RECT  993.02 916.76 1197.22 921.16 ;
     RECT  899.9 912.56 900.1 924.52 ;
     RECT  717.02 907.1 717.22 925.16 ;
     RECT  654.14 923.06 654.34 927.88 ;
     RECT  1021.34 921.16 1197.22 927.88 ;
     RECT  957.98 916.96 958.66 930.82 ;
     RECT  993.02 921.16 1010.02 931.46 ;
     RECT  1021.34 927.88 1181.86 931.46 ;
     RECT  993.02 931.46 1181.86 931.66 ;
     RECT  957.98 930.82 958.18 932.08 ;
     RECT  993.02 931.66 993.22 935.86 ;
     RECT  1194.62 927.88 1197.22 935.86 ;
     RECT  1194.62 935.86 1194.82 936.28 ;
     RECT  829.82 932.3 830.02 937.34 ;
     RECT  1003.1 931.66 1181.86 939.22 ;
     RECT  1003.1 939.22 1081.54 939.64 ;
     RECT  829.82 937.34 831.94 939.86 ;
     RECT  717.02 925.16 720.1 940.48 ;
     RECT  820.22 939.86 831.94 940.48 ;
     RECT  1004.06 939.64 1081.54 942.16 ;
     RECT  1021.34 942.16 1081.54 942.58 ;
     RECT  1029.5 942.58 1081.54 943 ;
     RECT  1091.9 939.22 1181.86 943.64 ;
     RECT  1091.9 943.64 1187.62 943.84 ;
     RECT  1045.82 943 1081.54 944.26 ;
     RECT  1096.22 943.84 1187.62 944.26 ;
     RECT  1096.22 944.26 1119.94 945.52 ;
     RECT  1132.22 944.26 1187.62 946.16 ;
     RECT  1045.82 944.26 1080.58 946.78 ;
     RECT  1132.22 946.16 1188.1 948.26 ;
     RECT  1132.22 948.26 1194.82 948.88 ;
     RECT  1149.5 948.88 1194.82 949.72 ;
     RECT  1048.22 946.78 1080.58 950.14 ;
     RECT  1049.66 950.14 1080.58 950.56 ;
     RECT  719.9 940.48 720.1 950.98 ;
     RECT  1133.18 948.88 1133.38 951.82 ;
     RECT  1149.5 949.72 1181.86 953.08 ;
     RECT  1192.7 949.72 1194.82 953.92 ;
     RECT  820.22 940.48 830.02 954.76 ;
     RECT  1096.22 945.52 1116.58 955.6 ;
     RECT  1149.5 953.08 1161.22 955.6 ;
     RECT  1051.1 950.56 1080.58 956.02 ;
     RECT  1029.5 943 1031.14 956.44 ;
     RECT  1096.22 955.6 1098.82 956.86 ;
     RECT  1194.62 953.92 1194.82 956.86 ;
     RECT  829.82 954.76 830.02 957.7 ;
     RECT  1030.94 956.44 1031.14 957.7 ;
     RECT  1051.1 956.02 1068.58 957.7 ;
     RECT  1080.38 956.02 1080.58 957.7 ;
     RECT  1172.06 953.08 1181.86 957.7 ;
     RECT  1110.14 955.6 1116.58 959.8 ;
     RECT  1156.7 955.6 1161.22 959.8 ;
     RECT  1172.06 957.7 1172.26 965.26 ;
     RECT  605.18 957.92 605.38 965.68 ;
     RECT  1158.14 959.8 1161.22 965.68 ;
     RECT  691.58 949.1 691.78 968.42 ;
     RECT  766.46 957.5 766.66 969.68 ;
     RECT  1051.1 957.7 1061.86 973.88 ;
     RECT  766.46 969.68 772.9 974.5 ;
     RECT  1051.1 973.88 1065.22 974.92 ;
     RECT  1052.54 974.92 1065.22 975.76 ;
     RECT  957.98 969.26 958.18 976.4 ;
     RECT  691.58 968.42 694.66 979.54 ;
     RECT  694.46 979.54 694.66 980.8 ;
     RECT  1053.98 975.76 1065.22 980.8 ;
     RECT  1053.98 980.8 1057.54 982.06 ;
     RECT  1096.7 956.86 1098.82 983.32 ;
     RECT  1158.62 965.68 1161.22 983.32 ;
     RECT  1004.06 942.16 1006.18 986.68 ;
     RECT  957.98 976.4 959.62 988.36 ;
     RECT  957.98 988.36 958.18 992.56 ;
     RECT  1161.02 983.32 1161.22 992.98 ;
     RECT  1110.14 959.8 1110.34 995.92 ;
     RECT  880.22 961.7 880.42 996.34 ;
     RECT  1005.98 986.68 1006.18 996.76 ;
     RECT  1098.62 983.32 1098.82 998.86 ;
     RECT  1057.34 982.06 1057.54 1003.9 ;
     RECT  766.46 974.5 766.66 1004.32 ;
     RECT  1057.82 1008.32 1058.02 1018.82 ;
     RECT  1069.34 1016.72 1069.54 1018.82 ;
     RECT  968.06 1022.6 968.26 1027.84 ;
     RECT  893.66 999.92 893.86 1030.36 ;
     RECT  1024.22 992.36 1024.42 1036.88 ;
     RECT  1057.82 1018.82 1069.54 1045.48 ;
     RECT  1057.82 1045.48 1063.3 1050.52 ;
     RECT  1024.22 1036.88 1024.9 1052.42 ;
     RECT  832.22 1033.1 832.42 1052.62 ;
     RECT  1010.3 1007.9 1010.5 1058.5 ;
     RECT  1021.34 1052.42 1024.9 1060.82 ;
     RECT  1063.1 1050.52 1063.3 1060.82 ;
     RECT  896.06 1058.72 896.26 1061.44 ;
     RECT  1146.62 1052.84 1146.82 1063.96 ;
     RECT  1063.1 1060.82 1068.58 1064.18 ;
     RECT  1015.58 1060.82 1024.9 1067.12 ;
     RECT  1063.1 1064.18 1072.9 1067.12 ;
     RECT  1063.1 1067.12 1075.3 1067.96 ;
     RECT  1015.58 1067.12 1026.34 1068.16 ;
     RECT  1063.1 1067.96 1080.1 1068.38 ;
     RECT  918.62 1062.92 918.82 1072.78 ;
     RECT  705.98 1058.72 706.18 1073.84 ;
     RECT  1061.18 1068.38 1080.1 1077.82 ;
     RECT  703.1 1073.84 706.18 1079.08 ;
     RECT  1061.18 1077.82 1074.34 1084.12 ;
     RECT  1061.18 1084.12 1072.9 1085.18 ;
     RECT  858.14 1075.52 858.34 1089.58 ;
     RECT  705.98 1079.08 706.18 1090.42 ;
     RECT  1016.06 1068.16 1026.34 1102.18 ;
     RECT  1058.78 1085.18 1072.9 1104.7 ;
     RECT  1060.22 1104.7 1063.3 1108.9 ;
     RECT  1060.22 1108.9 1060.9 1115.84 ;
     RECT  1058.78 1115.84 1060.9 1122.34 ;
     RECT  640.22 1122.98 640.42 1124.02 ;
     RECT  578.78 1109.54 578.98 1124.66 ;
     RECT  578.78 1124.66 584.26 1124.86 ;
     RECT  1058.78 1122.34 1060.42 1128.86 ;
     RECT  1016.06 1102.18 1024.42 1129.06 ;
     RECT  1050.14 1128.86 1060.42 1136.2 ;
     RECT  806.78 1135.16 806.98 1136.84 ;
     RECT  806.78 1136.84 807.46 1139.14 ;
     RECT  807.26 1139.14 807.46 1139.56 ;
     RECT  918.62 1101.14 918.82 1143.34 ;
     RECT  1050.14 1136.2 1058.98 1147.12 ;
     RECT  1024.22 1129.06 1024.42 1150.06 ;
     RECT  584.06 1124.86 584.26 1156.78 ;
     RECT  652.7 1108.7 652.9 1159.3 ;
     RECT  1050.14 1147.12 1050.34 1159.3 ;
     RECT  654.62 1159.52 654.82 1181.56 ;
     RECT  805.82 1184.3 806.02 1200.88 ;
     RECT  811.1 1201.94 811.3 1212.22 ;
  END
END cve2_core
END LIBRARY
